/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 20:57:04 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2237795551 */

module carry_lookahead_adder_4bit__6_8(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   INV_X1 i_8 (.A(in0[0]), .ZN(sum[0]));
   XOR2_X1 i_0_0 (.A(in0[1]), .B(in0[0]), .Z(sum[1]));
   NOR2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(sum[2]));
   AOI21_X1 i_0_2 (.A(in0[2]), .B1(in0[1]), .B2(in0[0]), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[3]), .B(n_0_2), .ZN(sum[3]));
   AND2_X1 i_0_4 (.A1(in0[3]), .A2(n_0_1), .ZN(cout));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_0_1));
   NAND3_X1 i_0_6 (.A1(in0[2]), .A2(in0[1]), .A3(in0[0]), .ZN(n_0_2));
endmodule

module carry_lookahead_adder_4bit__6_17(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(cin), .Z(sum[0]));
   NOR2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum[1]));
   AOI21_X1 i_0_2 (.A(in0[1]), .B1(in0[0]), .B2(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[2]), .B(n_0_3), .ZN(sum[2]));
   XNOR2_X1 i_0_4 (.A(in0[3]), .B(n_0_1), .ZN(sum[3]));
   AND3_X1 i_0_5 (.A1(in0[3]), .A2(in0[2]), .A3(n_0_2), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in0[2]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_8 (.A1(in0[1]), .A2(in0[0]), .A3(cin), .ZN(n_0_3));
endmodule

module carry_lookahead_adder_4bit__6_26(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(cin), .Z(sum[0]));
   NOR2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum[1]));
   AOI21_X1 i_0_2 (.A(in0[1]), .B1(in0[0]), .B2(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[2]), .B(n_0_3), .ZN(sum[2]));
   XNOR2_X1 i_0_4 (.A(in0[3]), .B(n_0_1), .ZN(sum[3]));
   AND3_X1 i_0_5 (.A1(in0[3]), .A2(in0[2]), .A3(n_0_2), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in0[2]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_8 (.A1(in0[1]), .A2(in0[0]), .A3(cin), .ZN(n_0_3));
endmodule

module carry_lookahead_adder_4bit__6_35(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   XOR2_X1 i_0_0 (.A(in0[3]), .B(cin), .Z(sum[0]));
endmodule

module carry_lookahead_adder_20bit__0_1376(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [19:0]in0;
   input [19:0]in1;
   input cin;
   output [19:0]sum;
   output cout;
   output v;

   wire c1;
   wire c2;
   wire c3;

   carry_lookahead_adder_4bit__6_8 cla0 (.in0({in0[3], in0[2], in0[1], in0[0]}), 
      .in1(), .cin(), .sum({sum[3], sum[2], sum[1], sum[0]}), .cout(c1), .v());
   carry_lookahead_adder_4bit__6_17 cla1 (.in0({in0[7], in0[6], in0[5], in0[4]}), 
      .in1(), .cin(c1), .sum({sum[7], sum[6], sum[5], sum[4]}), .cout(c2), .v());
   carry_lookahead_adder_4bit__6_26 cla2 (.in0({in0[11], in0[10], in0[9], in0[8]}), 
      .in1(), .cin(c2), .sum({sum[11], sum[10], sum[9], sum[8]}), .cout(c3), 
      .v());
   carry_lookahead_adder_4bit__6_35 cla3 (.in0({in0[19], uc_0, uc_1, uc_2}), 
      .in1(), .cin(c3), .sum({uc_3, uc_4, uc_5, sum[12]}), .cout(), .v());
endmodule

module add_sub_cla__0_1377__GU(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   carry_lookahead_adder_20bit__0_1376 cs0 (.sub(), .in0({in1[12], uc_0, uc_1, 
      uc_2, uc_3, uc_4, uc_5, uc_6, in1[11], in1[10], in1[9], in1[8], in1[7], 
      in1[6], in1[5], in1[4], in1[3], in1[2], in1[1], in1[0]}), .in1(), .cin(), 
      .sum({uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, out[12], out[11], 
      out[10], out[9], out[8], out[7], out[6], out[5], out[4], out[3], out[2], 
      out[1], out[0]}), .cout(), .v());
endmodule

module carry_lookahead_adder_4bit__4_8(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   INV_X1 i_8 (.A(in0[0]), .ZN(sum[0]));
   XOR2_X1 i_0_0 (.A(in0[1]), .B(in0[0]), .Z(sum[1]));
   NOR2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(sum[2]));
   AOI21_X1 i_0_2 (.A(in0[2]), .B1(in0[1]), .B2(in0[0]), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[3]), .B(n_0_2), .ZN(sum[3]));
   AND2_X1 i_0_4 (.A1(in0[3]), .A2(n_0_1), .ZN(cout));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_0_1));
   NAND3_X1 i_0_6 (.A1(in0[2]), .A2(in0[1]), .A3(in0[0]), .ZN(n_0_2));
endmodule

module carry_lookahead_adder_4bit__4_17(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(cin), .Z(sum[0]));
   NOR2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum[1]));
   AOI21_X1 i_0_2 (.A(in0[1]), .B1(in0[0]), .B2(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[2]), .B(n_0_3), .ZN(sum[2]));
   XNOR2_X1 i_0_4 (.A(in0[3]), .B(n_0_1), .ZN(sum[3]));
   AND3_X1 i_0_5 (.A1(in0[3]), .A2(in0[2]), .A3(n_0_2), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in0[2]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_8 (.A1(in0[1]), .A2(in0[0]), .A3(cin), .ZN(n_0_3));
endmodule

module carry_lookahead_adder_4bit__4_26(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(cin), .Z(sum[0]));
   NOR2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum[1]));
   AOI21_X1 i_0_2 (.A(in0[1]), .B1(in0[0]), .B2(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[2]), .B(n_0_3), .ZN(sum[2]));
   XNOR2_X1 i_0_4 (.A(in0[3]), .B(n_0_1), .ZN(sum[3]));
   AND3_X1 i_0_5 (.A1(in0[3]), .A2(in0[2]), .A3(n_0_2), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in0[2]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_8 (.A1(in0[1]), .A2(in0[0]), .A3(cin), .ZN(n_0_3));
endmodule

module carry_lookahead_adder_4bit__4_35(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   XOR2_X1 i_0_0 (.A(in0[3]), .B(cin), .Z(sum[0]));
endmodule

module carry_lookahead_adder_20bit__0_1320(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [19:0]in0;
   input [19:0]in1;
   input cin;
   output [19:0]sum;
   output cout;
   output v;

   wire c1;
   wire c2;
   wire c3;

   carry_lookahead_adder_4bit__4_8 cla0 (.in0({in0[3], in0[2], in0[1], in0[0]}), 
      .in1(), .cin(), .sum({sum[3], sum[2], sum[1], sum[0]}), .cout(c1), .v());
   carry_lookahead_adder_4bit__4_17 cla1 (.in0({in0[7], in0[6], in0[5], in0[4]}), 
      .in1(), .cin(c1), .sum({sum[7], sum[6], sum[5], sum[4]}), .cout(c2), .v());
   carry_lookahead_adder_4bit__4_26 cla2 (.in0({in0[11], in0[10], in0[9], in0[8]}), 
      .in1(), .cin(c2), .sum({sum[11], sum[10], sum[9], sum[8]}), .cout(c3), 
      .v());
   carry_lookahead_adder_4bit__4_35 cla3 (.in0({in0[19], uc_0, uc_1, uc_2}), 
      .in1(), .cin(c3), .sum({uc_3, uc_4, uc_5, sum[12]}), .cout(), .v());
endmodule

module add_sub_cla__0_1321__GU(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   carry_lookahead_adder_20bit__0_1320 cs0 (.sub(), .in0({in1[12], uc_0, uc_1, 
      uc_2, uc_3, uc_4, uc_5, uc_6, in1[11], in1[10], in1[9], in1[8], in1[7], 
      in1[6], in1[5], in1[4], in1[3], in1[2], in1[1], in1[0]}), .in1(), .cin(), 
      .sum({uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, out[12], out[11], 
      out[10], out[9], out[8], out[7], out[6], out[5], out[4], out[3], out[2], 
      out[1], out[0]}), .cout(), .v());
endmodule

module carry_lookahead_adder_4bit__9_8(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   INV_X1 i_8 (.A(in0[0]), .ZN(sum[0]));
   XOR2_X1 i_0_0 (.A(in0[1]), .B(in0[0]), .Z(sum[1]));
   NOR2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(sum[2]));
   AOI21_X1 i_0_2 (.A(in0[2]), .B1(in0[1]), .B2(in0[0]), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[3]), .B(n_0_2), .ZN(sum[3]));
   AND2_X1 i_0_4 (.A1(in0[3]), .A2(n_0_1), .ZN(cout));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_0_1));
   NAND3_X1 i_0_6 (.A1(in0[2]), .A2(in0[1]), .A3(in0[0]), .ZN(n_0_2));
endmodule

module carry_lookahead_adder_4bit__9_17(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(cin), .Z(sum[0]));
   NOR2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum[1]));
   AOI21_X1 i_0_2 (.A(in0[1]), .B1(in0[0]), .B2(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[2]), .B(n_0_3), .ZN(sum[2]));
   XNOR2_X1 i_0_4 (.A(in0[3]), .B(n_0_1), .ZN(sum[3]));
   AND3_X1 i_0_5 (.A1(in0[3]), .A2(in0[2]), .A3(n_0_2), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in0[2]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_8 (.A1(in0[1]), .A2(in0[0]), .A3(cin), .ZN(n_0_3));
endmodule

module carry_lookahead_adder_4bit__9_26(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(cin), .Z(sum[0]));
   NOR2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum[1]));
   AOI21_X1 i_0_2 (.A(in0[1]), .B1(in0[0]), .B2(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[2]), .B(n_0_3), .ZN(sum[2]));
   XNOR2_X1 i_0_4 (.A(in0[3]), .B(n_0_1), .ZN(sum[3]));
   AND3_X1 i_0_5 (.A1(in0[3]), .A2(in0[2]), .A3(n_0_2), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in0[2]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_8 (.A1(in0[1]), .A2(in0[0]), .A3(cin), .ZN(n_0_3));
endmodule

module carry_lookahead_adder_4bit__9_35(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   XOR2_X1 i_0_0 (.A(in0[3]), .B(cin), .Z(sum[0]));
endmodule

module carry_lookahead_adder_20bit(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [19:0]in0;
   input [19:0]in1;
   input cin;
   output [19:0]sum;
   output cout;
   output v;

   wire c1;
   wire c2;
   wire c3;

   carry_lookahead_adder_4bit__9_8 cla0 (.in0({in0[3], in0[2], in0[1], in0[0]}), 
      .in1(), .cin(), .sum({sum[3], sum[2], sum[1], sum[0]}), .cout(c1), .v());
   carry_lookahead_adder_4bit__9_17 cla1 (.in0({in0[7], in0[6], in0[5], in0[4]}), 
      .in1(), .cin(c1), .sum({sum[7], sum[6], sum[5], sum[4]}), .cout(c2), .v());
   carry_lookahead_adder_4bit__9_26 cla2 (.in0({in0[11], in0[10], in0[9], in0[8]}), 
      .in1(), .cin(c2), .sum({sum[11], sum[10], sum[9], sum[8]}), .cout(c3), 
      .v());
   carry_lookahead_adder_4bit__9_35 cla3 (.in0({in0[19], uc_0, uc_1, uc_2}), 
      .in1(), .cin(c3), .sum({uc_3, uc_4, uc_5, sum[12]}), .cout(), .v());
endmodule

module add_sub_cla__GU(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   carry_lookahead_adder_20bit cs0 (.sub(), .in0({in1[12], uc_0, uc_1, uc_2, 
      uc_3, uc_4, uc_5, uc_6, in1[11], in1[10], in1[9], in1[8], in1[7], in1[6], 
      in1[5], in1[4], in1[3], in1[2], in1[1], in1[0]}), .in1(), .cin(), .sum({
      uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, out[12], out[11], out[10], 
      out[9], out[8], out[7], out[6], out[5], out[4], out[3], out[2], out[1], 
      out[0]}), .cout(), .v());
endmodule

module carry_lookahead_adder_4bit__8_8(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   INV_X1 i_8 (.A(in0[0]), .ZN(sum[0]));
   XOR2_X1 i_0_0 (.A(in0[1]), .B(in0[0]), .Z(sum[1]));
   NOR2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(sum[2]));
   AOI21_X1 i_0_2 (.A(in0[2]), .B1(in0[1]), .B2(in0[0]), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[3]), .B(n_0_2), .ZN(sum[3]));
   AND2_X1 i_0_4 (.A1(in0[3]), .A2(n_0_1), .ZN(cout));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_0_1));
   NAND3_X1 i_0_6 (.A1(in0[2]), .A2(in0[1]), .A3(in0[0]), .ZN(n_0_2));
endmodule

module carry_lookahead_adder_4bit__8_17(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(cin), .Z(sum[0]));
   NOR2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum[1]));
   AOI21_X1 i_0_2 (.A(in0[1]), .B1(in0[0]), .B2(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[2]), .B(n_0_3), .ZN(sum[2]));
   XNOR2_X1 i_0_4 (.A(in0[3]), .B(n_0_1), .ZN(sum[3]));
   AND3_X1 i_0_5 (.A1(in0[3]), .A2(in0[2]), .A3(n_0_2), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in0[2]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_8 (.A1(in0[1]), .A2(in0[0]), .A3(cin), .ZN(n_0_3));
endmodule

module carry_lookahead_adder_4bit__8_26(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(cin), .Z(sum[0]));
   NOR2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum[1]));
   AOI21_X1 i_0_2 (.A(in0[1]), .B1(in0[0]), .B2(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[2]), .B(n_0_3), .ZN(sum[2]));
   XNOR2_X1 i_0_4 (.A(in0[3]), .B(n_0_1), .ZN(sum[3]));
   AND3_X1 i_0_5 (.A1(in0[3]), .A2(in0[2]), .A3(n_0_2), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in0[2]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_8 (.A1(in0[1]), .A2(in0[0]), .A3(cin), .ZN(n_0_3));
endmodule

module carry_lookahead_adder_4bit__8_35(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   XOR2_X1 i_0_0 (.A(in0[3]), .B(cin), .Z(sum[0]));
endmodule

module carry_lookahead_adder_20bit__0_1432(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [19:0]in0;
   input [19:0]in1;
   input cin;
   output [19:0]sum;
   output cout;
   output v;

   wire c1;
   wire c2;
   wire c3;

   carry_lookahead_adder_4bit__8_8 cla0 (.in0({in0[3], in0[2], in0[1], in0[0]}), 
      .in1(), .cin(), .sum({sum[3], sum[2], sum[1], sum[0]}), .cout(c1), .v());
   carry_lookahead_adder_4bit__8_17 cla1 (.in0({in0[7], in0[6], in0[5], in0[4]}), 
      .in1(), .cin(c1), .sum({sum[7], sum[6], sum[5], sum[4]}), .cout(c2), .v());
   carry_lookahead_adder_4bit__8_26 cla2 (.in0({in0[11], in0[10], in0[9], in0[8]}), 
      .in1(), .cin(c2), .sum({sum[11], sum[10], sum[9], sum[8]}), .cout(c3), 
      .v());
   carry_lookahead_adder_4bit__8_35 cla3 (.in0({in0[19], uc_0, uc_1, uc_2}), 
      .in1(), .cin(c3), .sum({uc_3, uc_4, uc_5, sum[12]}), .cout(), .v());
endmodule

module add_sub_cla__0_1433__GU(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   carry_lookahead_adder_20bit__0_1432 cs0 (.sub(), .in0({in1[12], uc_0, uc_1, 
      uc_2, uc_3, uc_4, uc_5, uc_6, in1[11], in1[10], in1[9], in1[8], in1[7], 
      in1[6], in1[5], in1[4], in1[3], in1[2], in1[1], in1[0]}), .in1(), .cin(), 
      .sum({uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, out[12], out[11], 
      out[10], out[9], out[8], out[7], out[6], out[5], out[4], out[3], out[2], 
      out[1], out[0]}), .cout(), .v());
endmodule

module carry_lookahead_adder_4bit__7_8(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   INV_X1 i_8 (.A(in0[0]), .ZN(sum[0]));
   XOR2_X1 i_0_0 (.A(in0[1]), .B(in0[0]), .Z(sum[1]));
   NOR2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(sum[2]));
   AOI21_X1 i_0_2 (.A(in0[2]), .B1(in0[1]), .B2(in0[0]), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[3]), .B(n_0_2), .ZN(sum[3]));
   AND2_X1 i_0_4 (.A1(in0[3]), .A2(n_0_1), .ZN(cout));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_0_1));
   NAND3_X1 i_0_6 (.A1(in0[2]), .A2(in0[1]), .A3(in0[0]), .ZN(n_0_2));
endmodule

module carry_lookahead_adder_4bit__7_17(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(cin), .Z(sum[0]));
   NOR2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum[1]));
   AOI21_X1 i_0_2 (.A(in0[1]), .B1(in0[0]), .B2(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[2]), .B(n_0_3), .ZN(sum[2]));
   XNOR2_X1 i_0_4 (.A(in0[3]), .B(n_0_1), .ZN(sum[3]));
   AND3_X1 i_0_5 (.A1(in0[3]), .A2(in0[2]), .A3(n_0_2), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in0[2]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_8 (.A1(in0[1]), .A2(in0[0]), .A3(cin), .ZN(n_0_3));
endmodule

module carry_lookahead_adder_4bit__7_26(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(cin), .Z(sum[0]));
   NOR2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum[1]));
   AOI21_X1 i_0_2 (.A(in0[1]), .B1(in0[0]), .B2(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[2]), .B(n_0_3), .ZN(sum[2]));
   XNOR2_X1 i_0_4 (.A(in0[3]), .B(n_0_1), .ZN(sum[3]));
   AND3_X1 i_0_5 (.A1(in0[3]), .A2(in0[2]), .A3(n_0_2), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in0[2]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_8 (.A1(in0[1]), .A2(in0[0]), .A3(cin), .ZN(n_0_3));
endmodule

module carry_lookahead_adder_4bit__7_35(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   XOR2_X1 i_0_0 (.A(in0[3]), .B(cin), .Z(sum[0]));
endmodule

module carry_lookahead_adder_20bit__0_1404(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [19:0]in0;
   input [19:0]in1;
   input cin;
   output [19:0]sum;
   output cout;
   output v;

   wire c1;
   wire c2;
   wire c3;

   carry_lookahead_adder_4bit__7_8 cla0 (.in0({in0[3], in0[2], in0[1], in0[0]}), 
      .in1(), .cin(), .sum({sum[3], sum[2], sum[1], sum[0]}), .cout(c1), .v());
   carry_lookahead_adder_4bit__7_17 cla1 (.in0({in0[7], in0[6], in0[5], in0[4]}), 
      .in1(), .cin(c1), .sum({sum[7], sum[6], sum[5], sum[4]}), .cout(c2), .v());
   carry_lookahead_adder_4bit__7_26 cla2 (.in0({in0[11], in0[10], in0[9], in0[8]}), 
      .in1(), .cin(c2), .sum({sum[11], sum[10], sum[9], sum[8]}), .cout(c3), 
      .v());
   carry_lookahead_adder_4bit__7_35 cla3 (.in0({in0[19], uc_0, uc_1, uc_2}), 
      .in1(), .cin(c3), .sum({uc_3, uc_4, uc_5, sum[12]}), .cout(), .v());
endmodule

module add_sub_cla__0_1405__GU(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   carry_lookahead_adder_20bit__0_1404 cs0 (.sub(), .in0({in1[12], uc_0, uc_1, 
      uc_2, uc_3, uc_4, uc_5, uc_6, in1[11], in1[10], in1[9], in1[8], in1[7], 
      in1[6], in1[5], in1[4], in1[3], in1[2], in1[1], in1[0]}), .in1(), .cin(), 
      .sum({uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, out[12], out[11], 
      out[10], out[9], out[8], out[7], out[6], out[5], out[4], out[3], out[2], 
      out[1], out[0]}), .cout(), .v());
endmodule

module carry_lookahead_adder_4bit__5_8(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;

   INV_X1 i_8 (.A(in0[0]), .ZN(sum[0]));
   XOR2_X1 i_0_0 (.A(in0[1]), .B(in0[0]), .Z(sum[1]));
   NOR2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(sum[2]));
   AOI21_X1 i_0_2 (.A(in0[2]), .B1(in0[1]), .B2(in0[0]), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[3]), .B(n_0_2), .ZN(sum[3]));
   AND2_X1 i_0_4 (.A1(in0[3]), .A2(n_0_1), .ZN(cout));
   INV_X1 i_0_5 (.A(n_0_2), .ZN(n_0_1));
   NAND3_X1 i_0_6 (.A1(in0[2]), .A2(in0[1]), .A3(in0[0]), .ZN(n_0_2));
endmodule

module carry_lookahead_adder_4bit__5_17(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(cin), .Z(sum[0]));
   NOR2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum[1]));
   AOI21_X1 i_0_2 (.A(in0[1]), .B1(in0[0]), .B2(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[2]), .B(n_0_3), .ZN(sum[2]));
   XNOR2_X1 i_0_4 (.A(in0[3]), .B(n_0_1), .ZN(sum[3]));
   AND3_X1 i_0_5 (.A1(in0[3]), .A2(in0[2]), .A3(n_0_2), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in0[2]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_8 (.A1(in0[1]), .A2(in0[0]), .A3(cin), .ZN(n_0_3));
endmodule

module carry_lookahead_adder_4bit__5_26(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(cin), .Z(sum[0]));
   NOR2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_0), .ZN(sum[1]));
   AOI21_X1 i_0_2 (.A(in0[1]), .B1(in0[0]), .B2(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(in0[2]), .B(n_0_3), .ZN(sum[2]));
   XNOR2_X1 i_0_4 (.A(in0[3]), .B(n_0_1), .ZN(sum[3]));
   AND3_X1 i_0_5 (.A1(in0[3]), .A2(in0[2]), .A3(n_0_2), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in0[2]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_7 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_8 (.A1(in0[1]), .A2(in0[0]), .A3(cin), .ZN(n_0_3));
endmodule

module carry_lookahead_adder_4bit__5_35(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   XOR2_X1 i_0_0 (.A(in0[3]), .B(cin), .Z(sum[0]));
endmodule

module carry_lookahead_adder_20bit__0_1348(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [19:0]in0;
   input [19:0]in1;
   input cin;
   output [19:0]sum;
   output cout;
   output v;

   wire c1;
   wire c2;
   wire c3;

   carry_lookahead_adder_4bit__5_8 cla0 (.in0({in0[3], in0[2], in0[1], in0[0]}), 
      .in1(), .cin(), .sum({sum[3], sum[2], sum[1], sum[0]}), .cout(c1), .v());
   carry_lookahead_adder_4bit__5_17 cla1 (.in0({in0[7], in0[6], in0[5], in0[4]}), 
      .in1(), .cin(c1), .sum({sum[7], sum[6], sum[5], sum[4]}), .cout(c2), .v());
   carry_lookahead_adder_4bit__5_26 cla2 (.in0({in0[11], in0[10], in0[9], in0[8]}), 
      .in1(), .cin(c2), .sum({sum[11], sum[10], sum[9], sum[8]}), .cout(c3), 
      .v());
   carry_lookahead_adder_4bit__5_35 cla3 (.in0({in0[19], uc_0, uc_1, uc_2}), 
      .in1(), .cin(c3), .sum({uc_3, uc_4, uc_5, sum[12]}), .cout(), .v());
endmodule

module add_sub_cla__0_1349__GU(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   carry_lookahead_adder_20bit__0_1348 cs0 (.sub(), .in0({in1[12], uc_0, uc_1, 
      uc_2, uc_3, uc_4, uc_5, uc_6, in1[11], in1[10], in1[9], in1[8], in1[7], 
      in1[6], in1[5], in1[4], in1[3], in1[2], in1[1], in1[0]}), .in1(), .cin(), 
      .sum({uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, out[12], out[11], 
      out[10], out[9], out[8], out[7], out[6], out[5], out[4], out[3], out[2], 
      out[1], out[0]}), .cout(), .v());
endmodule

module datapath__0_1(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   INV_X1 i_0 (.A(n_0), .ZN(p_1[0]));
   OAI21_X1 i_1 (.A(n_65), .B1(B[0]), .B2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_65), .B(n_1), .Z(p_1[1]));
   OAI21_X1 i_3 (.A(n_64), .B1(B[1]), .B2(p_0[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_63), .B(n_2), .ZN(p_1[2]));
   OAI21_X1 i_5 (.A(n_67), .B1(B[2]), .B2(p_0[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_61), .B(n_3), .Z(p_1[3]));
   XOR2_X1 i_7 (.A(B[3]), .B(p_0[3]), .Z(n_3));
   XOR2_X1 i_8 (.A(n_60), .B(n_10), .Z(p_1[4]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_1[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_1[6]));
   NOR2_X1 i_11 (.A1(n_57), .A2(n_48), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_1[7]));
   OAI22_X1 i_13 (.A1(B[6]), .A2(p_0[6]), .B1(n_48), .B2(n_7), .ZN(n_5));
   AOI21_X1 i_14 (.A(n_58), .B1(B[5]), .B2(p_0[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_58), .B1(n_52), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_55), .B1(n_60), .B2(n_53), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_53), .B1(B[4]), .B2(p_0[4]), .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_59), .A2(n_50), .ZN(n_11));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_1[10]));
   NOR2_X1 i_23 (.A1(n_43), .A2(n_34), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_1[11]));
   OAI22_X1 i_25 (.A1(B[10]), .A2(p_0[10]), .B1(n_34), .B2(n_15), .ZN(n_13));
   AOI21_X1 i_27 (.A(n_44), .B1(n_38), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   NOR2_X1 i_31 (.A1(n_45), .A2(n_36), .ZN(n_19));
   XNOR2_X1 i_32 (.A(n_32), .B(n_31), .ZN(p_1[12]));
   XOR2_X1 i_33 (.A(n_29), .B(n_25), .Z(p_1[13]));
   XOR2_X1 i_34 (.A(n_21), .B(n_20), .Z(p_1[14]));
   OAI22_X1 i_35 (.A1(B[15]), .A2(p_0[13]), .B1(n_29), .B2(n_26), .ZN(n_20));
   AOI21_X1 i_36 (.A(n_28), .B1(p_0[14]), .B2(n_70), .ZN(n_21));
   XNOR2_X1 i_37 (.A(n_23), .B(n_22), .ZN(p_1[15]));
   XOR2_X1 i_38 (.A(p_0[15]), .B(p_0[14]), .Z(n_22));
   AOI222_X1 i_39 (.A1(p_0[14]), .A2(n_70), .B1(B[15]), .B2(p_0[14]), .C1(n_29), 
      .C2(n_24), .ZN(n_23));
   NOR2_X1 i_40 (.A1(n_28), .A2(n_25), .ZN(n_24));
   OAI21_X1 i_41 (.A(n_27), .B1(B[15]), .B2(p_0[13]), .ZN(n_25));
   INV_X1 i_42 (.A(n_27), .ZN(n_26));
   NAND2_X1 i_43 (.A1(B[15]), .A2(p_0[13]), .ZN(n_27));
   NOR2_X1 i_44 (.A1(p_0[14]), .A2(n_70), .ZN(n_28));
   INV_X1 i_45 (.A(n_30), .ZN(n_29));
   AOI21_X1 i_46 (.A(n_69), .B1(n_32), .B2(n_31), .ZN(n_30));
   AOI21_X1 i_47 (.A(n_69), .B1(B[15]), .B2(p_0[12]), .ZN(n_31));
   NOR4_X1 i_48 (.A1(n_36), .A2(n_33), .A3(n_37), .A4(n_40), .ZN(n_32));
   NOR2_X1 i_49 (.A1(n_45), .A2(n_35), .ZN(n_33));
   INV_X1 i_50 (.A(n_35), .ZN(n_34));
   NAND2_X1 i_51 (.A1(B[10]), .A2(p_0[10]), .ZN(n_35));
   AND2_X1 i_52 (.A1(B[11]), .A2(p_0[11]), .ZN(n_36));
   AOI21_X1 i_53 (.A(n_42), .B1(n_39), .B2(n_38), .ZN(n_37));
   NAND2_X1 i_54 (.A1(B[9]), .A2(p_0[9]), .ZN(n_38));
   NOR3_X1 i_56 (.A1(n_42), .A2(n_41), .A3(n_46), .ZN(n_40));
   OR3_X1 i_58 (.A1(n_45), .A2(n_43), .A3(n_44), .ZN(n_42));
   NOR2_X1 i_59 (.A1(B[10]), .A2(p_0[10]), .ZN(n_43));
   NOR2_X1 i_60 (.A1(B[9]), .A2(p_0[9]), .ZN(n_44));
   NOR2_X1 i_61 (.A1(B[11]), .A2(p_0[11]), .ZN(n_45));
   INV_X1 i_64 (.A(n_49), .ZN(n_48));
   NAND2_X1 i_77 (.A1(n_67), .A2(n_62), .ZN(n_61));
   OAI21_X1 i_78 (.A(n_63), .B1(B[2]), .B2(p_0[2]), .ZN(n_62));
   AOI21_X1 i_79 (.A(n_66), .B1(n_65), .B2(n_64), .ZN(n_63));
   NAND2_X1 i_80 (.A1(B[1]), .A2(p_0[1]), .ZN(n_64));
   NAND2_X1 i_81 (.A1(B[0]), .A2(p_0[0]), .ZN(n_65));
   NOR2_X1 i_82 (.A1(B[1]), .A2(p_0[1]), .ZN(n_66));
   NAND2_X1 i_83 (.A1(B[2]), .A2(p_0[2]), .ZN(n_67));
   AND2_X1 i_84 (.A1(B[3]), .A2(p_0[3]), .ZN(n_68));
   NOR2_X1 i_85 (.A1(B[15]), .A2(p_0[12]), .ZN(n_69));
   INV_X1 i_86 (.A(p_0[13]), .ZN(n_70));
   INV_X1 i_20 (.A(n_73), .ZN(n_50));
   XNOR2_X1 i_21 (.A(n_14), .B(n_71), .ZN(p_1[8]));
   NAND2_X1 i_26 (.A1(n_18), .A2(n_39), .ZN(n_14));
   INV_X1 i_29 (.A(n_41), .ZN(n_18));
   NAND2_X1 i_30 (.A1(n_47), .A2(n_54), .ZN(p_1[9]));
   OAI21_X1 i_55 (.A(n_17), .B1(n_44), .B2(n_51), .ZN(n_47));
   INV_X1 i_57 (.A(n_79), .ZN(n_51));
   NAND3_X1 i_62 (.A1(n_80), .A2(n_79), .A3(n_56), .ZN(n_54));
   INV_X1 i_63 (.A(n_17), .ZN(n_56));
   OAI21_X1 i_65 (.A(n_39), .B1(n_46), .B2(n_41), .ZN(n_17));
   INV_X1 i_66 (.A(n_71), .ZN(n_46));
   NAND4_X1 i_67 (.A1(n_72), .A2(n_76), .A3(n_74), .A4(n_73), .ZN(n_71));
   OR2_X1 i_68 (.A1(n_59), .A2(n_49), .ZN(n_72));
   NAND2_X1 i_69 (.A1(p_0[6]), .A2(B[6]), .ZN(n_49));
   NOR2_X1 i_70 (.A1(p_0[7]), .A2(B[7]), .ZN(n_59));
   NAND2_X1 i_71 (.A1(p_0[7]), .A2(B[7]), .ZN(n_73));
   OAI211_X1 i_72 (.A(n_78), .B(n_75), .C1(p_0[7]), .C2(B[7]), .ZN(n_74));
   NAND2_X1 i_73 (.A1(n_52), .A2(n_53), .ZN(n_75));
   NAND2_X1 i_74 (.A1(p_0[5]), .A2(B[5]), .ZN(n_52));
   NAND2_X1 i_75 (.A1(p_0[4]), .A2(B[4]), .ZN(n_53));
   OAI211_X1 i_76 (.A(n_78), .B(n_77), .C1(p_0[7]), .C2(B[7]), .ZN(n_76));
   NOR2_X1 i_87 (.A1(n_55), .A2(n_60), .ZN(n_77));
   NOR2_X1 i_88 (.A1(p_0[4]), .A2(B[4]), .ZN(n_55));
   OAI22_X1 i_89 (.A1(n_68), .A2(n_61), .B1(B[3]), .B2(p_0[3]), .ZN(n_60));
   NOR2_X1 i_90 (.A1(n_57), .A2(n_58), .ZN(n_78));
   NOR2_X1 i_91 (.A1(p_0[6]), .A2(B[6]), .ZN(n_57));
   NOR2_X1 i_92 (.A1(p_0[5]), .A2(B[5]), .ZN(n_58));
   NOR2_X1 i_93 (.A1(p_0[8]), .A2(B[8]), .ZN(n_41));
   NAND2_X1 i_94 (.A1(p_0[8]), .A2(B[8]), .ZN(n_39));
   NAND2_X1 i_95 (.A1(p_0[9]), .A2(B[9]), .ZN(n_79));
   INV_X1 i_96 (.A(n_44), .ZN(n_80));
endmodule

module datapath__0_6(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   INV_X1 i_0 (.A(n_0), .ZN(p_1[0]));
   OAI21_X1 i_1 (.A(n_60), .B1(B[0]), .B2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_60), .B(n_1), .Z(p_1[1]));
   OAI21_X1 i_3 (.A(n_59), .B1(B[1]), .B2(p_0[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_58), .B(n_2), .ZN(p_1[2]));
   OAI21_X1 i_5 (.A(n_62), .B1(B[2]), .B2(p_0[2]), .ZN(n_2));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_1[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_1[6]));
   NOR2_X1 i_11 (.A1(n_52), .A2(n_43), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_1[7]));
   OAI22_X1 i_13 (.A1(B[6]), .A2(p_0[6]), .B1(n_43), .B2(n_7), .ZN(n_5));
   AOI21_X1 i_14 (.A(n_53), .B1(B[5]), .B2(p_0[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_53), .B1(n_47), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_50), .B1(n_55), .B2(n_48), .ZN(n_9));
   NOR2_X1 i_19 (.A1(n_54), .A2(n_45), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_41), .B(n_18), .ZN(p_1[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_1[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_1[10]));
   NOR2_X1 i_23 (.A1(n_38), .A2(n_29), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_1[11]));
   OAI22_X1 i_25 (.A1(B[10]), .A2(p_0[10]), .B1(n_29), .B2(n_15), .ZN(n_13));
   AOI21_X1 i_26 (.A(n_39), .B1(B[9]), .B2(p_0[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_39), .B1(n_33), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_36), .B1(n_41), .B2(n_34), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_36), .B1(B[8]), .B2(p_0[8]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_40), .A2(n_31), .ZN(n_19));
   XNOR2_X1 i_32 (.A(n_27), .B(n_26), .ZN(p_1[12]));
   XNOR2_X1 i_33 (.A(n_25), .B(n_24), .ZN(p_1[13]));
   XNOR2_X1 i_34 (.A(p_0[14]), .B(n_20), .ZN(p_1[14]));
   AOI21_X1 i_35 (.A(n_21), .B1(n_65), .B2(n_25), .ZN(n_20));
   NOR3_X1 i_36 (.A1(n_68), .A2(p_0[13]), .A3(n_25), .ZN(n_21));
   OAI22_X1 i_37 (.A1(n_67), .A2(n_65), .B1(n_25), .B2(n_22), .ZN(p_1[15]));
   OAI21_X1 i_38 (.A(n_23), .B1(p_0[14]), .B2(n_66), .ZN(n_22));
   INV_X1 i_39 (.A(n_24), .ZN(n_23));
   AOI21_X1 i_40 (.A(n_65), .B1(B[15]), .B2(n_66), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_64), .B1(n_27), .B2(n_26), .ZN(n_25));
   AOI21_X1 i_42 (.A(n_64), .B1(B[15]), .B2(p_0[12]), .ZN(n_26));
   NOR4_X1 i_43 (.A1(n_31), .A2(n_28), .A3(n_32), .A4(n_35), .ZN(n_27));
   NOR2_X1 i_44 (.A1(n_40), .A2(n_30), .ZN(n_28));
   INV_X1 i_45 (.A(n_30), .ZN(n_29));
   NAND2_X1 i_46 (.A1(B[10]), .A2(p_0[10]), .ZN(n_30));
   AND2_X1 i_47 (.A1(B[11]), .A2(p_0[11]), .ZN(n_31));
   AOI21_X1 i_48 (.A(n_37), .B1(n_34), .B2(n_33), .ZN(n_32));
   NAND2_X1 i_49 (.A1(B[9]), .A2(p_0[9]), .ZN(n_33));
   NAND2_X1 i_50 (.A1(B[8]), .A2(p_0[8]), .ZN(n_34));
   NOR3_X1 i_51 (.A1(n_37), .A2(n_36), .A3(n_41), .ZN(n_35));
   NOR2_X1 i_52 (.A1(B[8]), .A2(p_0[8]), .ZN(n_36));
   OR3_X1 i_53 (.A1(n_40), .A2(n_38), .A3(n_39), .ZN(n_37));
   NOR2_X1 i_54 (.A1(B[10]), .A2(p_0[10]), .ZN(n_38));
   NOR2_X1 i_55 (.A1(B[9]), .A2(p_0[9]), .ZN(n_39));
   NOR2_X1 i_56 (.A1(B[11]), .A2(p_0[11]), .ZN(n_40));
   NOR4_X1 i_57 (.A1(n_45), .A2(n_42), .A3(n_46), .A4(n_49), .ZN(n_41));
   NOR2_X1 i_58 (.A1(n_54), .A2(n_44), .ZN(n_42));
   INV_X1 i_59 (.A(n_44), .ZN(n_43));
   NAND2_X1 i_60 (.A1(B[6]), .A2(p_0[6]), .ZN(n_44));
   AND2_X1 i_61 (.A1(B[7]), .A2(p_0[7]), .ZN(n_45));
   AOI21_X1 i_62 (.A(n_51), .B1(n_48), .B2(n_47), .ZN(n_46));
   NAND2_X1 i_63 (.A1(B[5]), .A2(p_0[5]), .ZN(n_47));
   NAND2_X1 i_64 (.A1(B[4]), .A2(p_0[4]), .ZN(n_48));
   NOR3_X1 i_65 (.A1(n_51), .A2(n_50), .A3(n_55), .ZN(n_49));
   NOR2_X1 i_66 (.A1(B[4]), .A2(p_0[4]), .ZN(n_50));
   OR3_X1 i_67 (.A1(n_54), .A2(n_52), .A3(n_53), .ZN(n_51));
   NOR2_X1 i_68 (.A1(B[6]), .A2(p_0[6]), .ZN(n_52));
   NOR2_X1 i_69 (.A1(B[5]), .A2(p_0[5]), .ZN(n_53));
   NOR2_X1 i_70 (.A1(B[7]), .A2(p_0[7]), .ZN(n_54));
   NOR2_X1 i_80 (.A1(B[15]), .A2(p_0[12]), .ZN(n_64));
   NOR2_X1 i_81 (.A1(B[15]), .A2(n_66), .ZN(n_65));
   INV_X1 i_82 (.A(p_0[13]), .ZN(n_66));
   INV_X1 i_83 (.A(p_0[14]), .ZN(n_67));
   INV_X1 i_84 (.A(B[15]), .ZN(n_68));
   NOR2_X1 i_6 (.A1(n_73), .A2(n_74), .ZN(n_58));
   NAND2_X1 i_7 (.A1(p_0[1]), .A2(B[1]), .ZN(n_59));
   NAND2_X1 i_8 (.A1(p_0[0]), .A2(B[0]), .ZN(n_60));
   OAI21_X1 i_18 (.A(n_3), .B1(n_10), .B2(n_57), .ZN(p_1[3]));
   NAND3_X1 i_71 (.A1(n_57), .A2(n_77), .A3(n_76), .ZN(n_3));
   INV_X1 i_72 (.A(n_56), .ZN(n_10));
   NAND2_X1 i_73 (.A1(n_77), .A2(n_76), .ZN(n_56));
   OAI21_X1 i_74 (.A(n_72), .B1(B[2]), .B2(p_0[2]), .ZN(n_57));
   NAND2_X1 i_75 (.A1(n_61), .A2(n_69), .ZN(p_1[4]));
   NAND2_X1 i_76 (.A1(n_55), .A2(n_63), .ZN(n_61));
   NAND2_X1 i_77 (.A1(n_70), .A2(n_77), .ZN(n_55));
   INV_X1 i_78 (.A(n_80), .ZN(n_63));
   NAND3_X1 i_79 (.A1(n_70), .A2(n_80), .A3(n_77), .ZN(n_69));
   OAI21_X1 i_85 (.A(n_76), .B1(n_71), .B2(n_75), .ZN(n_70));
   INV_X1 i_86 (.A(n_72), .ZN(n_71));
   OAI21_X1 i_87 (.A(n_62), .B1(n_73), .B2(n_74), .ZN(n_72));
   AOI22_X1 i_88 (.A1(p_0[1]), .A2(B[1]), .B1(p_0[0]), .B2(B[0]), .ZN(n_73));
   NOR2_X1 i_89 (.A1(p_0[1]), .A2(B[1]), .ZN(n_74));
   NAND2_X1 i_90 (.A1(p_0[2]), .A2(B[2]), .ZN(n_62));
   NOR2_X1 i_91 (.A1(p_0[2]), .A2(B[2]), .ZN(n_75));
   NAND2_X1 i_92 (.A1(p_0[3]), .A2(B[3]), .ZN(n_76));
   NAND2_X1 i_93 (.A1(n_78), .A2(n_79), .ZN(n_77));
   INV_X1 i_94 (.A(p_0[3]), .ZN(n_78));
   INV_X1 i_95 (.A(B[3]), .ZN(n_79));
   OAI21_X1 i_96 (.A(n_48), .B1(B[4]), .B2(p_0[4]), .ZN(n_80));
endmodule

module datapath__0_7(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   INV_X1 i_0 (.A(n_0), .ZN(p_2[0]));
   OAI21_X1 i_1 (.A(n_63), .B1(p_0[0]), .B2(p_1[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_63), .B(n_1), .Z(p_2[1]));
   OAI21_X1 i_3 (.A(n_62), .B1(p_0[1]), .B2(p_1[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_61), .B(n_2), .ZN(p_2[2]));
   OAI21_X1 i_5 (.A(n_66), .B1(p_0[2]), .B2(p_1[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_60), .B(n_3), .Z(p_2[3]));
   OAI21_X1 i_7 (.A(n_67), .B1(n_71), .B2(n_69), .ZN(n_3));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_2[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_2[6]));
   NOR2_X1 i_11 (.A1(n_55), .A2(n_46), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_2[7]));
   OAI22_X1 i_13 (.A1(p_0[6]), .A2(p_1[6]), .B1(n_46), .B2(n_7), .ZN(n_5));
   AOI21_X1 i_14 (.A(n_56), .B1(p_0[5]), .B2(p_1[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_56), .B1(n_50), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_53), .B1(n_58), .B2(n_51), .ZN(n_9));
   NOR2_X1 i_19 (.A1(n_57), .A2(n_48), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_44), .B(n_18), .ZN(p_2[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_2[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_2[10]));
   NOR2_X1 i_23 (.A1(n_41), .A2(n_32), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_2[11]));
   OAI22_X1 i_25 (.A1(p_0[10]), .A2(p_1[10]), .B1(n_32), .B2(n_15), .ZN(n_13));
   AOI21_X1 i_26 (.A(n_42), .B1(p_0[9]), .B2(p_1[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_42), .B1(n_36), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_39), .B1(n_44), .B2(n_37), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_39), .B1(p_0[8]), .B2(p_1[8]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_43), .A2(n_34), .ZN(n_19));
   XNOR2_X1 i_32 (.A(n_30), .B(n_29), .ZN(p_2[12]));
   XOR2_X1 i_33 (.A(n_28), .B(n_24), .Z(p_2[13]));
   XNOR2_X1 i_34 (.A(n_21), .B(n_20), .ZN(p_2[14]));
   OAI22_X1 i_35 (.A1(p_0[14]), .A2(p_1[14]), .B1(n_72), .B2(n_70), .ZN(n_20));
   NOR2_X1 i_36 (.A1(n_27), .A2(n_26), .ZN(n_21));
   XNOR2_X1 i_37 (.A(n_23), .B(n_22), .ZN(p_2[15]));
   XNOR2_X1 i_38 (.A(p_0[15]), .B(p_0[14]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_25), .B1(n_72), .B2(n_70), .ZN(n_23));
   AOI21_X1 i_40 (.A(n_26), .B1(p_0[13]), .B2(p_1[13]), .ZN(n_24));
   AOI211_X1 i_41 (.A(n_26), .B(n_27), .C1(p_0[14]), .C2(p_1[14]), .ZN(n_25));
   NOR2_X1 i_42 (.A1(p_0[13]), .A2(p_1[13]), .ZN(n_26));
   AOI21_X1 i_43 (.A(n_28), .B1(p_0[13]), .B2(p_1[13]), .ZN(n_27));
   AOI21_X1 i_44 (.A(n_68), .B1(n_30), .B2(n_29), .ZN(n_28));
   AOI21_X1 i_45 (.A(n_68), .B1(p_0[12]), .B2(p_1[12]), .ZN(n_29));
   NOR4_X1 i_46 (.A1(n_34), .A2(n_31), .A3(n_35), .A4(n_38), .ZN(n_30));
   NOR2_X1 i_47 (.A1(n_43), .A2(n_33), .ZN(n_31));
   INV_X1 i_48 (.A(n_33), .ZN(n_32));
   NAND2_X1 i_49 (.A1(p_0[10]), .A2(p_1[10]), .ZN(n_33));
   AND2_X1 i_50 (.A1(p_0[11]), .A2(p_1[11]), .ZN(n_34));
   AOI21_X1 i_51 (.A(n_40), .B1(n_37), .B2(n_36), .ZN(n_35));
   NAND2_X1 i_52 (.A1(p_0[9]), .A2(p_1[9]), .ZN(n_36));
   NAND2_X1 i_53 (.A1(p_0[8]), .A2(p_1[8]), .ZN(n_37));
   NOR3_X1 i_54 (.A1(n_40), .A2(n_39), .A3(n_44), .ZN(n_38));
   NOR2_X1 i_55 (.A1(p_0[8]), .A2(p_1[8]), .ZN(n_39));
   OR3_X1 i_56 (.A1(n_43), .A2(n_41), .A3(n_42), .ZN(n_40));
   NOR2_X1 i_57 (.A1(p_0[10]), .A2(p_1[10]), .ZN(n_41));
   NOR2_X1 i_58 (.A1(p_0[9]), .A2(p_1[9]), .ZN(n_42));
   NOR2_X1 i_59 (.A1(p_0[11]), .A2(p_1[11]), .ZN(n_43));
   NOR4_X1 i_60 (.A1(n_48), .A2(n_45), .A3(n_49), .A4(n_52), .ZN(n_44));
   NOR2_X1 i_61 (.A1(n_57), .A2(n_47), .ZN(n_45));
   INV_X1 i_62 (.A(n_47), .ZN(n_46));
   NAND2_X1 i_63 (.A1(p_0[6]), .A2(p_1[6]), .ZN(n_47));
   AND2_X1 i_64 (.A1(p_0[7]), .A2(p_1[7]), .ZN(n_48));
   AOI21_X1 i_65 (.A(n_54), .B1(n_51), .B2(n_50), .ZN(n_49));
   NAND2_X1 i_66 (.A1(p_0[5]), .A2(p_1[5]), .ZN(n_50));
   NAND2_X1 i_67 (.A1(p_0[4]), .A2(p_1[4]), .ZN(n_51));
   NOR3_X1 i_68 (.A1(n_54), .A2(n_53), .A3(n_58), .ZN(n_52));
   NOR2_X1 i_69 (.A1(p_0[4]), .A2(p_1[4]), .ZN(n_53));
   OR3_X1 i_70 (.A1(n_57), .A2(n_55), .A3(n_56), .ZN(n_54));
   NOR2_X1 i_71 (.A1(p_0[6]), .A2(p_1[6]), .ZN(n_55));
   NOR2_X1 i_72 (.A1(p_0[5]), .A2(p_1[5]), .ZN(n_56));
   NOR2_X1 i_73 (.A1(p_0[7]), .A2(p_1[7]), .ZN(n_57));
   NAND2_X1 i_78 (.A1(p_0[1]), .A2(p_1[1]), .ZN(n_62));
   NAND2_X1 i_79 (.A1(p_0[0]), .A2(p_1[0]), .ZN(n_63));
   NOR2_X1 i_80 (.A1(p_0[1]), .A2(p_1[1]), .ZN(n_64));
   NOR2_X1 i_84 (.A1(p_0[12]), .A2(p_1[12]), .ZN(n_68));
   INV_X1 i_86 (.A(p_1[14]), .ZN(n_70));
   INV_X1 i_88 (.A(p_0[14]), .ZN(n_72));
   NAND2_X1 i_8 (.A1(n_73), .A2(n_67), .ZN(n_58));
   NOR2_X1 i_18 (.A1(n_59), .A2(n_10), .ZN(p_2[4]));
   AOI21_X1 i_74 (.A(n_77), .B1(n_73), .B2(n_67), .ZN(n_10));
   INV_X1 i_75 (.A(n_65), .ZN(n_59));
   NAND3_X1 i_76 (.A1(n_73), .A2(n_77), .A3(n_67), .ZN(n_65));
   NAND2_X1 i_77 (.A1(n_60), .A2(n_76), .ZN(n_73));
   OAI21_X1 i_81 (.A(n_75), .B1(n_61), .B2(n_74), .ZN(n_60));
   AOI21_X1 i_82 (.A(n_64), .B1(n_62), .B2(n_63), .ZN(n_61));
   INV_X1 i_83 (.A(n_66), .ZN(n_74));
   NAND2_X1 i_85 (.A1(p_1[2]), .A2(p_0[2]), .ZN(n_66));
   OR2_X1 i_87 (.A1(p_1[2]), .A2(p_0[2]), .ZN(n_75));
   NAND2_X1 i_89 (.A1(p_1[3]), .A2(p_0[3]), .ZN(n_76));
   NAND2_X1 i_90 (.A1(n_69), .A2(n_71), .ZN(n_67));
   INV_X1 i_91 (.A(p_1[3]), .ZN(n_69));
   INV_X1 i_92 (.A(p_0[3]), .ZN(n_71));
   INV_X1 i_93 (.A(n_78), .ZN(n_77));
   OAI21_X1 i_94 (.A(n_51), .B1(p_0[4]), .B2(p_1[4]), .ZN(n_78));
endmodule

module datapath__0_12(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   INV_X1 i_0 (.A(n_0), .ZN(p_1[0]));
   OAI21_X1 i_1 (.A(n_60), .B1(B[0]), .B2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_60), .B(n_1), .Z(p_1[1]));
   OAI21_X1 i_3 (.A(n_59), .B1(B[1]), .B2(p_0[1]), .ZN(n_1));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_1[6]));
   NOR2_X1 i_11 (.A1(n_52), .A2(n_43), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_1[7]));
   OAI22_X1 i_13 (.A1(B[6]), .A2(p_0[6]), .B1(n_43), .B2(n_7), .ZN(n_5));
   AOI21_X1 i_15 (.A(n_53), .B1(n_47), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   NOR2_X1 i_19 (.A1(n_54), .A2(n_45), .ZN(n_11));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_1[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_1[10]));
   NOR2_X1 i_23 (.A1(n_38), .A2(n_29), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_1[11]));
   OAI22_X1 i_25 (.A1(B[10]), .A2(p_0[10]), .B1(n_29), .B2(n_15), .ZN(n_13));
   AOI21_X1 i_26 (.A(n_39), .B1(B[9]), .B2(p_0[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_39), .B1(n_33), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_36), .B1(n_41), .B2(n_34), .ZN(n_17));
   NOR2_X1 i_31 (.A1(n_40), .A2(n_31), .ZN(n_19));
   XNOR2_X1 i_32 (.A(n_27), .B(n_26), .ZN(p_1[12]));
   XNOR2_X1 i_33 (.A(n_25), .B(n_24), .ZN(p_1[13]));
   XNOR2_X1 i_34 (.A(p_0[14]), .B(n_20), .ZN(p_1[14]));
   AOI21_X1 i_35 (.A(n_21), .B1(n_65), .B2(n_25), .ZN(n_20));
   NOR3_X1 i_36 (.A1(n_68), .A2(p_0[13]), .A3(n_25), .ZN(n_21));
   OAI22_X1 i_37 (.A1(n_67), .A2(n_65), .B1(n_25), .B2(n_22), .ZN(p_1[15]));
   OAI21_X1 i_38 (.A(n_23), .B1(p_0[14]), .B2(n_66), .ZN(n_22));
   INV_X1 i_39 (.A(n_24), .ZN(n_23));
   AOI21_X1 i_40 (.A(n_65), .B1(B[15]), .B2(n_66), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_64), .B1(n_27), .B2(n_26), .ZN(n_25));
   AOI21_X1 i_42 (.A(n_64), .B1(B[15]), .B2(p_0[12]), .ZN(n_26));
   NOR4_X1 i_43 (.A1(n_31), .A2(n_28), .A3(n_32), .A4(n_35), .ZN(n_27));
   NOR2_X1 i_44 (.A1(n_40), .A2(n_30), .ZN(n_28));
   INV_X1 i_45 (.A(n_30), .ZN(n_29));
   NAND2_X1 i_46 (.A1(B[10]), .A2(p_0[10]), .ZN(n_30));
   AND2_X1 i_47 (.A1(B[11]), .A2(p_0[11]), .ZN(n_31));
   AOI21_X1 i_48 (.A(n_37), .B1(n_34), .B2(n_33), .ZN(n_32));
   NAND2_X1 i_49 (.A1(B[9]), .A2(p_0[9]), .ZN(n_33));
   NAND2_X1 i_50 (.A1(B[8]), .A2(p_0[8]), .ZN(n_34));
   NOR3_X1 i_51 (.A1(n_37), .A2(n_36), .A3(n_41), .ZN(n_35));
   NOR2_X1 i_52 (.A1(B[8]), .A2(p_0[8]), .ZN(n_36));
   OR3_X1 i_53 (.A1(n_40), .A2(n_38), .A3(n_39), .ZN(n_37));
   NOR2_X1 i_54 (.A1(B[10]), .A2(p_0[10]), .ZN(n_38));
   NOR2_X1 i_55 (.A1(B[9]), .A2(p_0[9]), .ZN(n_39));
   NOR2_X1 i_56 (.A1(B[11]), .A2(p_0[11]), .ZN(n_40));
   INV_X1 i_59 (.A(n_44), .ZN(n_43));
   NAND2_X1 i_60 (.A1(B[6]), .A2(p_0[6]), .ZN(n_44));
   NOR2_X1 i_80 (.A1(B[15]), .A2(p_0[12]), .ZN(n_64));
   NOR2_X1 i_81 (.A1(B[15]), .A2(n_66), .ZN(n_65));
   INV_X1 i_82 (.A(p_0[13]), .ZN(n_66));
   INV_X1 i_83 (.A(p_0[14]), .ZN(n_67));
   INV_X1 i_84 (.A(B[15]), .ZN(n_68));
   INV_X1 i_4 (.A(n_18), .ZN(n_45));
   NOR2_X1 i_5 (.A1(p_0[6]), .A2(B[6]), .ZN(n_52));
   NAND2_X1 i_6 (.A1(n_6), .A2(n_2), .ZN(p_1[8]));
   NAND3_X1 i_7 (.A1(n_3), .A2(n_61), .A3(n_41), .ZN(n_2));
   INV_X1 i_8 (.A(n_10), .ZN(n_41));
   INV_X1 i_9 (.A(n_36), .ZN(n_3));
   OAI21_X1 i_14 (.A(n_10), .B1(n_36), .B2(n_58), .ZN(n_6));
   NAND4_X1 i_17 (.A1(n_42), .A2(n_49), .A3(n_46), .A4(n_18), .ZN(n_10));
   NAND2_X1 i_18 (.A1(p_0[7]), .A2(B[7]), .ZN(n_18));
   OR2_X1 i_20 (.A1(n_54), .A2(n_44), .ZN(n_42));
   INV_X1 i_30 (.A(n_57), .ZN(n_54));
   NAND3_X1 i_57 (.A1(n_57), .A2(n_55), .A3(n_48), .ZN(n_46));
   NOR2_X1 i_58 (.A1(n_77), .A2(n_62), .ZN(n_48));
   NAND3_X1 i_61 (.A1(n_57), .A2(n_55), .A3(n_50), .ZN(n_49));
   NAND2_X1 i_62 (.A1(n_47), .A2(n_51), .ZN(n_50));
   NAND2_X1 i_63 (.A1(p_0[4]), .A2(B[4]), .ZN(n_51));
   INV_X1 i_64 (.A(n_56), .ZN(n_55));
   OAI21_X1 i_65 (.A(n_88), .B1(B[6]), .B2(p_0[6]), .ZN(n_56));
   OR2_X1 i_66 (.A1(p_0[7]), .A2(B[7]), .ZN(n_57));
   INV_X1 i_67 (.A(n_61), .ZN(n_58));
   NAND2_X1 i_68 (.A1(p_0[8]), .A2(B[8]), .ZN(n_61));
   INV_X1 i_69 (.A(n_78), .ZN(n_62));
   XOR2_X1 i_70 (.A(n_63), .B(n_83), .Z(p_1[2]));
   NAND2_X1 i_71 (.A1(n_85), .A2(n_82), .ZN(n_63));
   XOR2_X1 i_72 (.A(n_80), .B(n_69), .Z(p_1[3]));
   NAND2_X1 i_73 (.A1(n_70), .A2(n_86), .ZN(n_69));
   INV_X1 i_74 (.A(n_79), .ZN(n_70));
   XNOR2_X1 i_75 (.A(n_78), .B(n_71), .ZN(p_1[4]));
   NAND2_X1 i_76 (.A1(n_51), .A2(n_76), .ZN(n_71));
   NAND2_X1 i_77 (.A1(n_72), .A2(n_74), .ZN(p_1[5]));
   OAI21_X1 i_78 (.A(n_9), .B1(n_73), .B2(n_53), .ZN(n_72));
   INV_X1 i_79 (.A(n_75), .ZN(n_9));
   INV_X1 i_85 (.A(n_47), .ZN(n_73));
   NOR2_X1 i_86 (.A1(p_0[5]), .A2(B[5]), .ZN(n_53));
   NAND3_X1 i_87 (.A1(n_88), .A2(n_75), .A3(n_47), .ZN(n_74));
   OAI21_X1 i_88 (.A(n_76), .B1(n_78), .B2(n_87), .ZN(n_75));
   INV_X1 i_89 (.A(n_77), .ZN(n_76));
   NOR2_X1 i_90 (.A1(p_0[4]), .A2(B[4]), .ZN(n_77));
   AOI21_X1 i_91 (.A(n_79), .B1(n_80), .B2(n_86), .ZN(n_78));
   NOR2_X1 i_92 (.A1(p_0[3]), .A2(B[3]), .ZN(n_79));
   NAND2_X1 i_93 (.A1(n_81), .A2(n_85), .ZN(n_80));
   NAND2_X1 i_94 (.A1(n_83), .A2(n_82), .ZN(n_81));
   NAND2_X1 i_95 (.A1(p_0[2]), .A2(B[2]), .ZN(n_82));
   OAI21_X1 i_96 (.A(n_84), .B1(B[1]), .B2(p_0[1]), .ZN(n_83));
   NAND2_X1 i_97 (.A1(n_60), .A2(n_59), .ZN(n_84));
   NAND2_X1 i_98 (.A1(p_0[1]), .A2(B[1]), .ZN(n_59));
   NAND2_X1 i_99 (.A1(p_0[0]), .A2(B[0]), .ZN(n_60));
   OR2_X1 i_100 (.A1(p_0[2]), .A2(B[2]), .ZN(n_85));
   NAND2_X1 i_101 (.A1(p_0[3]), .A2(B[3]), .ZN(n_86));
   INV_X1 i_102 (.A(n_51), .ZN(n_87));
   NAND2_X1 i_103 (.A1(p_0[5]), .A2(B[5]), .ZN(n_47));
   NAND2_X1 i_104 (.A1(n_89), .A2(n_90), .ZN(n_88));
   INV_X1 i_105 (.A(p_0[5]), .ZN(n_89));
   INV_X1 i_106 (.A(B[5]), .ZN(n_90));
endmodule

module datapath__0_13(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   INV_X1 i_0 (.A(n_0), .ZN(p_2[0]));
   OAI21_X1 i_1 (.A(n_63), .B1(p_0[0]), .B2(p_1[0]), .ZN(n_0));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_2[7]));
   OAI22_X1 i_13 (.A1(p_0[6]), .A2(p_1[6]), .B1(n_46), .B2(n_7), .ZN(n_5));
   NOR2_X1 i_19 (.A1(n_57), .A2(n_48), .ZN(n_11));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_2[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_2[10]));
   NOR2_X1 i_23 (.A1(n_41), .A2(n_32), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_2[11]));
   OAI22_X1 i_25 (.A1(p_0[10]), .A2(p_1[10]), .B1(n_32), .B2(n_15), .ZN(n_13));
   AOI21_X1 i_26 (.A(n_42), .B1(p_0[9]), .B2(p_1[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_42), .B1(n_36), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_39), .B1(n_44), .B2(n_37), .ZN(n_17));
   NOR2_X1 i_31 (.A1(n_43), .A2(n_34), .ZN(n_19));
   XNOR2_X1 i_32 (.A(n_30), .B(n_29), .ZN(p_2[12]));
   XOR2_X1 i_33 (.A(n_28), .B(n_24), .Z(p_2[13]));
   XNOR2_X1 i_34 (.A(n_21), .B(n_20), .ZN(p_2[14]));
   OAI22_X1 i_35 (.A1(p_0[14]), .A2(p_1[14]), .B1(n_72), .B2(n_70), .ZN(n_20));
   NOR2_X1 i_36 (.A1(n_27), .A2(n_26), .ZN(n_21));
   XNOR2_X1 i_37 (.A(n_23), .B(n_22), .ZN(p_2[15]));
   XNOR2_X1 i_38 (.A(p_0[15]), .B(p_0[14]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_25), .B1(n_72), .B2(n_70), .ZN(n_23));
   AOI21_X1 i_40 (.A(n_26), .B1(p_0[13]), .B2(p_1[13]), .ZN(n_24));
   AOI211_X1 i_41 (.A(n_26), .B(n_27), .C1(p_0[14]), .C2(p_1[14]), .ZN(n_25));
   NOR2_X1 i_42 (.A1(p_0[13]), .A2(p_1[13]), .ZN(n_26));
   AOI21_X1 i_43 (.A(n_28), .B1(p_0[13]), .B2(p_1[13]), .ZN(n_27));
   AOI21_X1 i_44 (.A(n_68), .B1(n_30), .B2(n_29), .ZN(n_28));
   AOI21_X1 i_45 (.A(n_68), .B1(p_0[12]), .B2(p_1[12]), .ZN(n_29));
   NOR4_X1 i_46 (.A1(n_34), .A2(n_31), .A3(n_35), .A4(n_38), .ZN(n_30));
   NOR2_X1 i_47 (.A1(n_43), .A2(n_33), .ZN(n_31));
   INV_X1 i_48 (.A(n_33), .ZN(n_32));
   NAND2_X1 i_49 (.A1(p_0[10]), .A2(p_1[10]), .ZN(n_33));
   AND2_X1 i_50 (.A1(p_0[11]), .A2(p_1[11]), .ZN(n_34));
   AOI21_X1 i_51 (.A(n_40), .B1(n_37), .B2(n_36), .ZN(n_35));
   NAND2_X1 i_52 (.A1(p_0[9]), .A2(p_1[9]), .ZN(n_36));
   NAND2_X1 i_53 (.A1(p_0[8]), .A2(p_1[8]), .ZN(n_37));
   NOR3_X1 i_54 (.A1(n_40), .A2(n_39), .A3(n_44), .ZN(n_38));
   OR3_X1 i_56 (.A1(n_43), .A2(n_41), .A3(n_42), .ZN(n_40));
   NOR2_X1 i_57 (.A1(p_0[10]), .A2(p_1[10]), .ZN(n_41));
   NOR2_X1 i_58 (.A1(p_0[9]), .A2(p_1[9]), .ZN(n_42));
   NOR2_X1 i_59 (.A1(p_0[11]), .A2(p_1[11]), .ZN(n_43));
   INV_X1 i_62 (.A(n_47), .ZN(n_46));
   NAND2_X1 i_63 (.A1(p_0[6]), .A2(p_1[6]), .ZN(n_47));
   NOR2_X1 i_84 (.A1(p_0[12]), .A2(p_1[12]), .ZN(n_68));
   INV_X1 i_86 (.A(p_1[14]), .ZN(n_70));
   INV_X1 i_88 (.A(p_0[14]), .ZN(n_72));
   NOR2_X1 i_2 (.A1(p_1[8]), .A2(p_0[8]), .ZN(n_39));
   NAND2_X1 i_3 (.A1(p_1[7]), .A2(p_0[7]), .ZN(n_1));
   INV_X1 i_4 (.A(n_1), .ZN(n_48));
   NOR2_X1 i_5 (.A1(p_1[7]), .A2(p_0[7]), .ZN(n_2));
   NOR2_X1 i_6 (.A1(p_1[6]), .A2(p_0[6]), .ZN(n_3));
   NAND2_X1 i_7 (.A1(p_1[0]), .A2(p_0[0]), .ZN(n_4));
   NOR2_X1 i_8 (.A1(p_1[1]), .A2(p_0[1]), .ZN(n_6));
   INV_X1 i_9 (.A(n_6), .ZN(n_8));
   NAND2_X1 i_10 (.A1(p_1[1]), .A2(p_0[1]), .ZN(n_10));
   NAND2_X1 i_11 (.A1(n_8), .A2(n_10), .ZN(n_18));
   XOR2_X1 i_14 (.A(n_18), .B(n_4), .Z(p_2[1]));
   OR2_X1 i_15 (.A1(p_1[2]), .A2(p_0[2]), .ZN(n_45));
   NAND2_X1 i_16 (.A1(p_1[2]), .A2(p_0[2]), .ZN(n_49));
   NAND2_X1 i_17 (.A1(n_45), .A2(n_49), .ZN(n_50));
   AOI21_X1 i_18 (.A(n_6), .B1(n_4), .B2(n_10), .ZN(n_51));
   XNOR2_X1 i_20 (.A(n_50), .B(n_51), .ZN(p_2[2]));
   OR2_X1 i_30 (.A1(p_1[3]), .A2(p_0[3]), .ZN(n_52));
   NAND2_X1 i_55 (.A1(p_1[3]), .A2(p_0[3]), .ZN(n_53));
   NAND2_X1 i_60 (.A1(n_52), .A2(n_53), .ZN(n_54));
   INV_X1 i_61 (.A(n_49), .ZN(n_56));
   OAI21_X1 i_64 (.A(n_45), .B1(n_51), .B2(n_56), .ZN(n_58));
   XOR2_X1 i_65 (.A(n_54), .B(n_58), .Z(p_2[3]));
   NOR2_X1 i_66 (.A1(p_1[4]), .A2(p_0[4]), .ZN(n_59));
   INV_X1 i_67 (.A(n_59), .ZN(n_60));
   NAND2_X1 i_68 (.A1(p_1[4]), .A2(p_0[4]), .ZN(n_61));
   NAND2_X1 i_69 (.A1(n_60), .A2(n_61), .ZN(n_62));
   NAND2_X1 i_70 (.A1(n_58), .A2(n_53), .ZN(n_64));
   NAND2_X1 i_71 (.A1(n_64), .A2(n_52), .ZN(n_65));
   XOR2_X1 i_72 (.A(n_62), .B(n_65), .Z(p_2[4]));
   AOI21_X1 i_73 (.A(n_59), .B1(n_61), .B2(n_65), .ZN(n_66));
   NAND2_X1 i_74 (.A1(p_1[5]), .A2(p_0[5]), .ZN(n_67));
   INV_X1 i_75 (.A(n_86), .ZN(n_69));
   NAND2_X1 i_76 (.A1(n_69), .A2(n_67), .ZN(n_71));
   XNOR2_X1 i_77 (.A(n_71), .B(n_66), .ZN(p_2[5]));
   NAND3_X1 i_78 (.A1(n_60), .A2(n_52), .A3(n_64), .ZN(n_73));
   AND3_X1 i_79 (.A1(n_73), .A2(n_67), .A3(n_61), .ZN(n_74));
   OR3_X1 i_80 (.A1(n_74), .A2(n_86), .A3(n_3), .ZN(n_75));
   NAND3_X1 i_81 (.A1(n_1), .A2(n_47), .A3(n_75), .ZN(n_76));
   INV_X1 i_82 (.A(n_2), .ZN(n_77));
   NAND2_X1 i_83 (.A1(n_76), .A2(n_77), .ZN(n_78));
   XNOR2_X1 i_85 (.A(p_1[8]), .B(p_0[8]), .ZN(n_79));
   NAND3_X1 i_87 (.A1(n_79), .A2(n_77), .A3(n_76), .ZN(n_80));
   INV_X1 i_89 (.A(n_78), .ZN(n_81));
   OAI21_X1 i_90 (.A(n_80), .B1(n_79), .B2(n_81), .ZN(p_2[8]));
   BUF_X1 i_91 (.A(n_2), .Z(n_57));
   BUF_X1 i_92 (.A(n_3), .Z(n_55));
   BUF_X1 i_93 (.A(n_4), .Z(n_63));
   BUF_X1 i_94 (.A(n_66), .Z(n_9));
   BUF_X1 i_95 (.A(n_78), .Z(n_44));
   NAND2_X1 i_96 (.A1(n_88), .A2(n_82), .ZN(p_2[6]));
   NAND2_X1 i_97 (.A1(n_83), .A2(n_7), .ZN(n_82));
   NAND2_X1 i_98 (.A1(n_85), .A2(n_84), .ZN(n_83));
   INV_X1 i_99 (.A(n_46), .ZN(n_84));
   INV_X1 i_100 (.A(n_55), .ZN(n_85));
   AOI21_X1 i_101 (.A(n_86), .B1(n_87), .B2(n_67), .ZN(n_7));
   NOR2_X1 i_102 (.A1(p_1[5]), .A2(p_0[5]), .ZN(n_86));
   INV_X1 i_103 (.A(n_9), .ZN(n_87));
   NAND2_X1 i_104 (.A1(n_89), .A2(n_90), .ZN(n_88));
   NOR2_X1 i_105 (.A1(n_55), .A2(n_46), .ZN(n_89));
   OAI22_X1 i_106 (.A1(n_91), .A2(n_9), .B1(p_0[5]), .B2(p_1[5]), .ZN(n_90));
   INV_X1 i_107 (.A(n_67), .ZN(n_91));
endmodule

module datapath__0_18(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   INV_X1 i_0 (.A(n_0), .ZN(p_1[0]));
   OAI21_X1 i_1 (.A(n_60), .B1(B[0]), .B2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_1[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_1[6]));
   NOR2_X1 i_11 (.A1(n_52), .A2(n_43), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_1[7]));
   OAI22_X1 i_13 (.A1(B[6]), .A2(p_0[6]), .B1(n_43), .B2(n_7), .ZN(n_5));
   AOI21_X1 i_14 (.A(n_53), .B1(B[5]), .B2(p_0[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_53), .B1(n_47), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_50), .B1(n_55), .B2(n_48), .ZN(n_9));
   NOR2_X1 i_19 (.A1(n_54), .A2(n_45), .ZN(n_11));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_1[10]));
   NOR2_X1 i_23 (.A1(n_38), .A2(n_29), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_1[11]));
   OAI22_X1 i_25 (.A1(B[10]), .A2(p_0[10]), .B1(n_29), .B2(n_15), .ZN(n_13));
   AOI21_X1 i_27 (.A(n_39), .B1(n_33), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   NOR2_X1 i_31 (.A1(n_40), .A2(n_31), .ZN(n_19));
   XNOR2_X1 i_32 (.A(n_27), .B(n_26), .ZN(p_1[12]));
   XNOR2_X1 i_33 (.A(n_25), .B(n_24), .ZN(p_1[13]));
   XNOR2_X1 i_34 (.A(p_0[14]), .B(n_20), .ZN(p_1[14]));
   AOI21_X1 i_35 (.A(n_21), .B1(n_65), .B2(n_25), .ZN(n_20));
   NOR3_X1 i_36 (.A1(n_68), .A2(p_0[13]), .A3(n_25), .ZN(n_21));
   OAI22_X1 i_37 (.A1(n_67), .A2(n_65), .B1(n_25), .B2(n_22), .ZN(p_1[15]));
   OAI21_X1 i_38 (.A(n_23), .B1(p_0[14]), .B2(n_66), .ZN(n_22));
   INV_X1 i_39 (.A(n_24), .ZN(n_23));
   AOI21_X1 i_40 (.A(n_65), .B1(B[15]), .B2(n_66), .ZN(n_24));
   AOI21_X1 i_41 (.A(n_64), .B1(n_27), .B2(n_26), .ZN(n_25));
   AOI21_X1 i_42 (.A(n_64), .B1(B[15]), .B2(p_0[12]), .ZN(n_26));
   NOR4_X1 i_43 (.A1(n_31), .A2(n_28), .A3(n_32), .A4(n_35), .ZN(n_27));
   NOR2_X1 i_44 (.A1(n_40), .A2(n_30), .ZN(n_28));
   INV_X1 i_45 (.A(n_30), .ZN(n_29));
   NAND2_X1 i_46 (.A1(B[10]), .A2(p_0[10]), .ZN(n_30));
   AND2_X1 i_47 (.A1(B[11]), .A2(p_0[11]), .ZN(n_31));
   AOI21_X1 i_48 (.A(n_37), .B1(n_34), .B2(n_33), .ZN(n_32));
   NAND2_X1 i_49 (.A1(B[9]), .A2(p_0[9]), .ZN(n_33));
   NOR3_X1 i_51 (.A1(n_37), .A2(n_36), .A3(n_41), .ZN(n_35));
   OR3_X1 i_53 (.A1(n_40), .A2(n_38), .A3(n_39), .ZN(n_37));
   NOR2_X1 i_54 (.A1(B[10]), .A2(p_0[10]), .ZN(n_38));
   NOR2_X1 i_55 (.A1(B[9]), .A2(p_0[9]), .ZN(n_39));
   NOR2_X1 i_56 (.A1(B[11]), .A2(p_0[11]), .ZN(n_40));
   INV_X1 i_59 (.A(n_44), .ZN(n_43));
   NAND2_X1 i_60 (.A1(B[6]), .A2(p_0[6]), .ZN(n_44));
   OAI21_X1 i_73 (.A(n_58), .B1(B[2]), .B2(p_0[2]), .ZN(n_57));
   AND2_X1 i_79 (.A1(B[3]), .A2(p_0[3]), .ZN(n_63));
   NOR2_X1 i_80 (.A1(B[15]), .A2(p_0[12]), .ZN(n_64));
   NOR2_X1 i_81 (.A1(B[15]), .A2(n_66), .ZN(n_65));
   INV_X1 i_82 (.A(p_0[13]), .ZN(n_66));
   INV_X1 i_83 (.A(p_0[14]), .ZN(n_67));
   INV_X1 i_84 (.A(B[15]), .ZN(n_68));
   INV_X1 i_2 (.A(n_46), .ZN(n_45));
   NOR2_X1 i_3 (.A1(p_0[7]), .A2(B[7]), .ZN(n_54));
   XNOR2_X1 i_4 (.A(n_1), .B(n_42), .ZN(p_1[8]));
   NAND2_X1 i_5 (.A1(n_2), .A2(n_34), .ZN(n_1));
   INV_X1 i_6 (.A(n_36), .ZN(n_2));
   NAND2_X1 i_7 (.A1(n_3), .A2(n_14), .ZN(p_1[9]));
   OAI21_X1 i_8 (.A(n_17), .B1(n_39), .B2(n_10), .ZN(n_3));
   INV_X1 i_18 (.A(n_71), .ZN(n_10));
   NAND3_X1 i_20 (.A1(n_72), .A2(n_71), .A3(n_18), .ZN(n_14));
   INV_X1 i_21 (.A(n_17), .ZN(n_18));
   OAI21_X1 i_26 (.A(n_34), .B1(n_36), .B2(n_41), .ZN(n_17));
   INV_X1 i_29 (.A(n_42), .ZN(n_41));
   NAND4_X1 i_30 (.A1(n_61), .A2(n_56), .A3(n_49), .A4(n_46), .ZN(n_42));
   NAND2_X1 i_50 (.A1(p_0[7]), .A2(B[7]), .ZN(n_46));
   OAI21_X1 i_52 (.A(n_51), .B1(p_0[7]), .B2(B[7]), .ZN(n_49));
   INV_X1 i_57 (.A(n_44), .ZN(n_51));
   OAI211_X1 i_58 (.A(n_70), .B(n_59), .C1(p_0[7]), .C2(B[7]), .ZN(n_56));
   NAND2_X1 i_61 (.A1(n_47), .A2(n_48), .ZN(n_59));
   NAND2_X1 i_62 (.A1(p_0[5]), .A2(B[5]), .ZN(n_47));
   OAI211_X1 i_63 (.A(n_70), .B(n_62), .C1(p_0[7]), .C2(B[7]), .ZN(n_61));
   NOR2_X1 i_64 (.A1(n_50), .A2(n_55), .ZN(n_62));
   NAND2_X1 i_65 (.A1(p_0[2]), .A2(B[2]), .ZN(n_69));
   NOR2_X1 i_66 (.A1(n_52), .A2(n_53), .ZN(n_70));
   NOR2_X1 i_67 (.A1(p_0[5]), .A2(B[5]), .ZN(n_53));
   NOR2_X1 i_68 (.A1(p_0[6]), .A2(B[6]), .ZN(n_52));
   NOR2_X1 i_69 (.A1(p_0[8]), .A2(B[8]), .ZN(n_36));
   NAND2_X1 i_70 (.A1(p_0[8]), .A2(B[8]), .ZN(n_34));
   NAND2_X1 i_71 (.A1(p_0[9]), .A2(B[9]), .ZN(n_71));
   INV_X1 i_72 (.A(n_39), .ZN(n_72));
   XOR2_X1 i_74 (.A(n_60), .B(n_73), .Z(p_1[1]));
   NAND2_X1 i_75 (.A1(n_74), .A2(n_76), .ZN(n_73));
   INV_X1 i_76 (.A(n_77), .ZN(n_74));
   XOR2_X1 i_77 (.A(n_58), .B(n_75), .Z(p_1[2]));
   XOR2_X1 i_78 (.A(B[2]), .B(p_0[2]), .Z(n_75));
   AOI21_X1 i_85 (.A(n_77), .B1(n_76), .B2(n_60), .ZN(n_58));
   NAND2_X1 i_86 (.A1(p_0[0]), .A2(B[0]), .ZN(n_60));
   NAND2_X1 i_87 (.A1(p_0[1]), .A2(B[1]), .ZN(n_76));
   NOR2_X1 i_88 (.A1(p_0[1]), .A2(B[1]), .ZN(n_77));
   XNOR2_X1 i_89 (.A(n_78), .B(n_86), .ZN(p_1[3]));
   XNOR2_X1 i_90 (.A(p_0[3]), .B(B[3]), .ZN(n_78));
   NAND2_X1 i_91 (.A1(n_83), .A2(n_79), .ZN(p_1[4]));
   NAND3_X1 i_92 (.A1(n_80), .A2(n_55), .A3(n_48), .ZN(n_79));
   NAND2_X1 i_93 (.A1(n_81), .A2(n_82), .ZN(n_80));
   INV_X1 i_94 (.A(p_0[4]), .ZN(n_81));
   INV_X1 i_95 (.A(B[4]), .ZN(n_82));
   OAI21_X1 i_96 (.A(n_85), .B1(n_84), .B2(n_50), .ZN(n_83));
   INV_X1 i_97 (.A(n_48), .ZN(n_84));
   NAND2_X1 i_98 (.A1(p_0[4]), .A2(B[4]), .ZN(n_48));
   NOR2_X1 i_99 (.A1(p_0[4]), .A2(B[4]), .ZN(n_50));
   INV_X1 i_100 (.A(n_55), .ZN(n_85));
   OAI22_X1 i_101 (.A1(n_63), .A2(n_86), .B1(B[3]), .B2(p_0[3]), .ZN(n_55));
   NAND2_X1 i_102 (.A1(n_57), .A2(n_69), .ZN(n_86));
endmodule

module datapath__0_19(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   INV_X1 i_0 (.A(n_0), .ZN(p_2[0]));
   OAI21_X1 i_1 (.A(n_63), .B1(p_0[0]), .B2(p_1[0]), .ZN(n_0));
   XOR2_X1 i_8 (.A(n_58), .B(n_10), .Z(p_2[4]));
   XOR2_X1 i_9 (.A(n_9), .B(n_6), .Z(p_2[5]));
   XOR2_X1 i_10 (.A(n_7), .B(n_4), .Z(p_2[6]));
   NOR2_X1 i_11 (.A1(n_55), .A2(n_46), .ZN(n_4));
   XNOR2_X1 i_12 (.A(n_11), .B(n_5), .ZN(p_2[7]));
   OAI22_X1 i_13 (.A1(p_0[6]), .A2(p_1[6]), .B1(n_46), .B2(n_7), .ZN(n_5));
   AOI21_X1 i_14 (.A(n_56), .B1(p_0[5]), .B2(p_1[5]), .ZN(n_6));
   AOI21_X1 i_15 (.A(n_56), .B1(n_50), .B2(n_8), .ZN(n_7));
   INV_X1 i_16 (.A(n_9), .ZN(n_8));
   AOI21_X1 i_17 (.A(n_53), .B1(n_58), .B2(n_51), .ZN(n_9));
   OAI21_X1 i_18 (.A(n_51), .B1(p_0[4]), .B2(p_1[4]), .ZN(n_10));
   NOR2_X1 i_19 (.A1(n_57), .A2(n_48), .ZN(n_11));
   XNOR2_X1 i_20 (.A(n_44), .B(n_18), .ZN(p_2[8]));
   XOR2_X1 i_21 (.A(n_17), .B(n_14), .Z(p_2[9]));
   XOR2_X1 i_22 (.A(n_15), .B(n_12), .Z(p_2[10]));
   NOR2_X1 i_23 (.A1(n_41), .A2(n_32), .ZN(n_12));
   XNOR2_X1 i_24 (.A(n_19), .B(n_13), .ZN(p_2[11]));
   OAI22_X1 i_25 (.A1(p_0[10]), .A2(p_1[10]), .B1(n_32), .B2(n_15), .ZN(n_13));
   AOI21_X1 i_26 (.A(n_42), .B1(p_0[9]), .B2(p_1[9]), .ZN(n_14));
   AOI21_X1 i_27 (.A(n_42), .B1(n_36), .B2(n_16), .ZN(n_15));
   INV_X1 i_28 (.A(n_17), .ZN(n_16));
   AOI21_X1 i_29 (.A(n_39), .B1(n_44), .B2(n_37), .ZN(n_17));
   AOI21_X1 i_30 (.A(n_39), .B1(p_0[8]), .B2(p_1[8]), .ZN(n_18));
   NOR2_X1 i_31 (.A1(n_43), .A2(n_34), .ZN(n_19));
   XNOR2_X1 i_32 (.A(n_30), .B(n_29), .ZN(p_2[12]));
   XOR2_X1 i_33 (.A(n_28), .B(n_24), .Z(p_2[13]));
   XNOR2_X1 i_34 (.A(n_21), .B(n_20), .ZN(p_2[14]));
   OAI22_X1 i_35 (.A1(p_0[14]), .A2(p_1[14]), .B1(n_72), .B2(n_70), .ZN(n_20));
   NOR2_X1 i_36 (.A1(n_27), .A2(n_26), .ZN(n_21));
   XNOR2_X1 i_37 (.A(n_23), .B(n_22), .ZN(p_2[15]));
   XNOR2_X1 i_38 (.A(p_0[15]), .B(p_0[14]), .ZN(n_22));
   AOI21_X1 i_39 (.A(n_25), .B1(n_72), .B2(n_70), .ZN(n_23));
   AOI21_X1 i_40 (.A(n_26), .B1(p_0[13]), .B2(p_1[13]), .ZN(n_24));
   AOI211_X1 i_41 (.A(n_26), .B(n_27), .C1(p_0[14]), .C2(p_1[14]), .ZN(n_25));
   NOR2_X1 i_42 (.A1(p_0[13]), .A2(p_1[13]), .ZN(n_26));
   AOI21_X1 i_43 (.A(n_28), .B1(p_0[13]), .B2(p_1[13]), .ZN(n_27));
   AOI21_X1 i_44 (.A(n_68), .B1(n_30), .B2(n_29), .ZN(n_28));
   AOI21_X1 i_45 (.A(n_68), .B1(p_0[12]), .B2(p_1[12]), .ZN(n_29));
   NOR4_X1 i_46 (.A1(n_34), .A2(n_31), .A3(n_35), .A4(n_38), .ZN(n_30));
   NOR2_X1 i_47 (.A1(n_43), .A2(n_33), .ZN(n_31));
   INV_X1 i_48 (.A(n_33), .ZN(n_32));
   NAND2_X1 i_49 (.A1(p_0[10]), .A2(p_1[10]), .ZN(n_33));
   AND2_X1 i_50 (.A1(p_0[11]), .A2(p_1[11]), .ZN(n_34));
   AOI21_X1 i_51 (.A(n_40), .B1(n_37), .B2(n_36), .ZN(n_35));
   NAND2_X1 i_52 (.A1(p_0[9]), .A2(p_1[9]), .ZN(n_36));
   NAND2_X1 i_53 (.A1(p_0[8]), .A2(p_1[8]), .ZN(n_37));
   NOR3_X1 i_54 (.A1(n_40), .A2(n_39), .A3(n_44), .ZN(n_38));
   NOR2_X1 i_55 (.A1(p_0[8]), .A2(p_1[8]), .ZN(n_39));
   OR3_X1 i_56 (.A1(n_43), .A2(n_41), .A3(n_42), .ZN(n_40));
   NOR2_X1 i_57 (.A1(p_0[10]), .A2(p_1[10]), .ZN(n_41));
   NOR2_X1 i_58 (.A1(p_0[9]), .A2(p_1[9]), .ZN(n_42));
   NOR2_X1 i_59 (.A1(p_0[11]), .A2(p_1[11]), .ZN(n_43));
   NOR4_X1 i_60 (.A1(n_48), .A2(n_45), .A3(n_49), .A4(n_52), .ZN(n_44));
   NOR2_X1 i_61 (.A1(n_57), .A2(n_47), .ZN(n_45));
   INV_X1 i_62 (.A(n_47), .ZN(n_46));
   NAND2_X1 i_63 (.A1(p_0[6]), .A2(p_1[6]), .ZN(n_47));
   AND2_X1 i_64 (.A1(p_0[7]), .A2(p_1[7]), .ZN(n_48));
   AOI21_X1 i_65 (.A(n_54), .B1(n_51), .B2(n_50), .ZN(n_49));
   NAND2_X1 i_66 (.A1(p_0[5]), .A2(p_1[5]), .ZN(n_50));
   NAND2_X1 i_67 (.A1(p_0[4]), .A2(p_1[4]), .ZN(n_51));
   NOR3_X1 i_68 (.A1(n_54), .A2(n_53), .A3(n_58), .ZN(n_52));
   NOR2_X1 i_69 (.A1(p_0[4]), .A2(p_1[4]), .ZN(n_53));
   OR3_X1 i_70 (.A1(n_57), .A2(n_55), .A3(n_56), .ZN(n_54));
   NOR2_X1 i_71 (.A1(p_0[6]), .A2(p_1[6]), .ZN(n_55));
   NOR2_X1 i_72 (.A1(p_0[5]), .A2(p_1[5]), .ZN(n_56));
   NOR2_X1 i_73 (.A1(p_0[7]), .A2(p_1[7]), .ZN(n_57));
   NAND2_X1 i_74 (.A1(n_67), .A2(n_59), .ZN(n_58));
   OAI21_X1 i_75 (.A(n_60), .B1(n_71), .B2(n_69), .ZN(n_59));
   NOR2_X1 i_80 (.A1(p_0[1]), .A2(p_1[1]), .ZN(n_64));
   INV_X1 i_81 (.A(n_66), .ZN(n_65));
   NOR2_X1 i_84 (.A1(p_0[12]), .A2(p_1[12]), .ZN(n_68));
   INV_X1 i_86 (.A(p_1[14]), .ZN(n_70));
   INV_X1 i_88 (.A(p_0[14]), .ZN(n_72));
   NAND2_X1 i_2 (.A1(p_1[2]), .A2(p_0[2]), .ZN(n_66));
   NAND2_X1 i_3 (.A1(p_1[0]), .A2(p_0[0]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(p_1[1]), .B(p_0[1]), .ZN(n_2));
   XOR2_X1 i_5 (.A(n_2), .B(n_1), .Z(p_2[1]));
   XNOR2_X1 i_6 (.A(p_1[2]), .B(p_0[2]), .ZN(n_3));
   NAND2_X1 i_7 (.A1(p_1[1]), .A2(p_0[1]), .ZN(n_61));
   AOI21_X1 i_76 (.A(n_64), .B1(n_1), .B2(n_61), .ZN(n_62));
   XNOR2_X1 i_77 (.A(n_3), .B(n_62), .ZN(p_2[2]));
   OAI22_X1 i_78 (.A1(n_62), .A2(n_65), .B1(p_1[2]), .B2(p_0[2]), .ZN(n_73));
   INV_X1 i_79 (.A(p_1[3]), .ZN(n_69));
   INV_X1 i_82 (.A(p_0[3]), .ZN(n_71));
   NOR2_X1 i_83 (.A1(p_1[3]), .A2(p_0[3]), .ZN(n_74));
   INV_X1 i_85 (.A(n_74), .ZN(n_75));
   INV_X1 i_87 (.A(n_73), .ZN(n_76));
   NAND2_X1 i_89 (.A1(p_1[3]), .A2(p_0[3]), .ZN(n_77));
   INV_X1 i_90 (.A(n_77), .ZN(n_78));
   OAI21_X1 i_91 (.A(n_76), .B1(n_78), .B2(n_74), .ZN(n_79));
   NAND3_X1 i_92 (.A1(n_75), .A2(n_73), .A3(n_77), .ZN(n_80));
   NAND2_X1 i_93 (.A1(n_79), .A2(n_80), .ZN(p_2[3]));
   BUF_X1 i_94 (.A(n_1), .Z(n_63));
   BUF_X1 i_95 (.A(n_73), .Z(n_60));
   BUF_X1 i_96 (.A(n_75), .Z(n_67));
endmodule

module booth_16bit_multiplier__1(A, B, product);
   input [15:0]A;
   input [15:0]B;
   output [31:0]product;

   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_80;
   wire n_0_100;
   wire n_0_120;
   wire n_0_140;
   wire n_0_160;
   wire n_0_180;
   wire n_0_200;
   wire n_0_214;
   wire n_0_216;
   wire n_0_220;
   wire n_0_230;
   wire n_0_231;
   wire n_0_234;
   wire n_0_235;
   wire n_0_0;
   wire n_0_4;
   wire n_0_5;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_24;
   wire n_0_25;
   wire n_0_34;
   wire n_0_35;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_44;
   wire n_0_50;
   wire n_0_55;
   wire n_0_57;
   wire n_0_58;
   wire n_0_69;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_215;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_16;
   wire n_0_26;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_36;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_56;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_76;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_75;
   wire n_0_105;
   wire n_0_27;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_77;
   wire n_0_79;
   wire n_0_113;
   wire n_0_78;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_98;
   wire n_0_97;
   wire n_0_141;
   wire n_0_99;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_117;
   wire n_0_118;
   wire n_0_166;
   wire n_0_119;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_137;
   wire n_0_138;
   wire n_0_193;
   wire n_0_139;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_157;
   wire n_0_158;
   wire n_0_229;
   wire n_0_159;
   wire n_0_232;
   wire n_0_233;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_178;
   wire n_0_177;
   wire n_0_257;
   wire n_0_179;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_197;
   wire n_0_198;
   wire n_0_283;
   wire n_0_199;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_217;
   wire n_0_310;
   wire n_0_311;
   wire n_0_218;
   wire n_0_312;
   wire n_0_219;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_2;
   wire n_0_1;
   wire n_0_332;
   wire n_0_3;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_21;
   wire n_0_345;
   wire n_0_346;
   wire n_0_22;
   wire n_0_347;
   wire n_0_23;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_41;
   wire n_0_43;
   wire n_0_363;
   wire n_0_42;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_59;
   wire n_0_68;
   wire n_0_377;
   wire n_0_70;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_132;
   wire n_0_404;
   wire n_0_134;
   wire n_0_133;
   wire n_0_136;
   wire n_0_135;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_0;
   wire n_1_1;
   wire n_1_15;
   wire n_1_16;
   wire n_1_17;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;
   wire n_1_28;
   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire n_1_60;
   wire n_1_61;
   wire n_1_62;
   wire n_1_63;
   wire n_1_64;
   wire n_1_65;
   wire n_1_66;
   wire n_1_67;
   wire n_1_68;
   wire n_1_69;
   wire n_1_70;
   wire n_1_71;
   wire n_1_72;
   wire n_1_73;
   wire n_1_74;
   wire n_1_75;
   wire n_1_76;
   wire n_1_77;
   wire n_1_78;
   wire n_1_79;
   wire n_1_80;
   wire n_1_81;
   wire n_1_82;
   wire n_1_83;
   wire n_1_84;
   wire n_1_85;
   wire n_1_86;
   wire n_1_87;
   wire n_1_88;
   wire n_1_89;
   wire n_1_90;
   wire n_1_91;
   wire n_1_92;
   wire n_1_93;
   wire n_1_94;
   wire n_1_95;
   wire n_1_96;
   wire n_1_97;
   wire n_1_98;
   wire n_1_99;
   wire n_1_100;
   wire n_1_101;
   wire n_1_102;
   wire n_1_103;
   wire n_1_104;
   wire n_1_105;
   wire n_1_106;
   wire n_1_107;
   wire n_1_108;
   wire n_1_109;
   wire n_1_110;
   wire n_1_111;
   wire n_1_112;
   wire n_1_113;
   wire n_1_114;
   wire n_1_115;
   wire n_1_116;
   wire n_1_117;
   wire n_1_118;
   wire n_1_119;
   wire n_1_120;
   wire n_1_121;
   wire n_1_122;
   wire n_1_123;
   wire n_1_124;
   wire n_1_125;
   wire n_1_126;
   wire n_1_127;
   wire n_1_128;
   wire n_1_129;
   wire n_1_130;
   wire n_1_131;
   wire n_1_132;
   wire n_1_133;
   wire n_1_134;
   wire n_1_135;
   wire n_1_136;
   wire n_1_137;
   wire n_1_138;
   wire n_1_139;
   wire n_1_140;
   wire n_1_141;
   wire n_1_142;
   wire n_1_143;
   wire n_1_144;
   wire n_1_145;
   wire n_1_146;
   wire n_1_147;
   wire n_1_148;
   wire n_1_149;
   wire n_1_150;
   wire n_1_151;
   wire n_1_152;
   wire n_1_153;
   wire n_1_154;
   wire n_1_155;
   wire n_1_156;
   wire n_1_157;
   wire n_1_158;
   wire n_1_159;
   wire n_1_160;
   wire n_1_161;
   wire n_1_162;
   wire n_1_163;
   wire n_1_164;
   wire n_1_165;
   wire n_1_166;
   wire n_1_167;
   wire n_1_168;
   wire n_1_169;
   wire n_1_170;
   wire n_1_171;
   wire n_1_172;
   wire n_1_173;
   wire n_1_174;
   wire n_1_175;
   wire n_1_176;
   wire n_1_177;

   datapath__0_1 i_2 (.B({B[15], uc_0, uc_1, uc_2, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({n_124, n_126, 
      n_125, n_264, n_263, n_262, n_261, n_260, n_259, n_258, n_257, n_256, 
      n_255, n_148, n_147, n_146}), .p_1({n_15, n_14, n_13, n_12, n_11, n_10, 
      n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0}));
   datapath__0_6 i_5 (.B({B[15], uc_3, uc_4, uc_5, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_6, n_123, n_122, 
      n_254, n_253, n_121, n_252, n_251, n_250, n_249, n_145, n_248, n_247, 
      n_144, n_143, n_142}), .p_1({n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
      n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16}));
   datapath__0_7 i_6 (.p_0({n_126, n_125, n_264, n_263, n_262, n_261, n_260, 
      n_259, n_258, n_257, n_256, n_255, n_148, n_147, n_146, B[0]}), .p_1({uc_7, 
      n_123, n_122, n_254, n_253, n_121, n_252, n_251, n_250, n_249, n_145, 
      n_248, n_247, n_144, n_143, n_142}), .p_2({n_47, n_46, n_45, n_44, n_43, 
      n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32}));
   datapath__0_12 i_9 (.B({B[15], uc_8, uc_9, uc_10, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_11, n_120, 
      n_119, n_246, n_245, n_118, n_117, n_244, n_243, n_242, n_241, n_141, 
      n_240, n_239, n_140, n_116}), .p_1({n_63, n_62, n_61, n_60, n_59, n_58, 
      n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48}));
   datapath__0_13 i_10 (.p_0({n_126, n_125, n_264, n_263, n_262, n_261, n_260, 
      n_259, n_258, n_257, n_256, n_255, n_148, n_147, n_146, B[0]}), .p_1({
      uc_12, n_120, n_119, n_246, n_245, n_118, n_117, n_244, n_243, n_242, 
      n_241, n_141, n_240, n_239, n_140, n_116}), .p_2({n_79, n_78, n_77, n_76, 
      n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64}));
   datapath__0_18 i_13 (.B({B[15], uc_13, uc_14, uc_15, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_16, n_115, 
      n_238, n_237, n_236, n_114, n_235, n_234, n_233, n_232, n_231, n_230, 
      n_139, n_229, n_138, n_113}), .p_1({n_95, n_94, n_93, n_92, n_91, n_90, 
      n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80}));
   datapath__0_19 i_14 (.p_0({n_126, n_125, n_264, n_263, n_262, n_261, n_260, 
      n_259, n_258, n_257, n_256, n_255, n_148, n_147, n_146, B[0]}), .p_1({
      uc_17, n_115, n_238, n_237, n_236, n_114, n_235, n_234, n_233, n_232, 
      n_231, n_230, n_139, n_229, n_138, n_113}), .p_2({n_111, n_110, n_109, 
      n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
      n_97, n_96}));
   INV_X1 i_0_108 (.A(n_0_60), .ZN(product[12]));
   AOI222_X1 i_0_109 (.A1(n_438), .A2(n_0_79), .B1(n_438), .B2(n_0_78), .C1(
      n_149), .C2(n_0_77), .ZN(n_0_60));
   INV_X1 i_0_110 (.A(n_0_61), .ZN(product[13]));
   AOI222_X1 i_0_111 (.A1(n_424), .A2(n_0_79), .B1(n_417), .B2(n_0_78), .C1(
      n_150), .C2(n_0_77), .ZN(n_0_61));
   INV_X1 i_0_112 (.A(n_0_62), .ZN(product[14]));
   AOI222_X1 i_0_113 (.A1(n_425), .A2(n_0_79), .B1(n_418), .B2(n_0_78), .C1(
      n_151), .C2(n_0_77), .ZN(n_0_62));
   INV_X1 i_0_144 (.A(n_0_80), .ZN(product[11]));
   AOI222_X1 i_0_145 (.A1(n_437), .A2(n_0_98), .B1(n_437), .B2(n_0_99), .C1(
      n_156), .C2(n_0_97), .ZN(n_0_80));
   INV_X1 i_0_180 (.A(n_0_100), .ZN(product[10]));
   AOI222_X1 i_0_181 (.A1(n_436), .A2(n_0_118), .B1(n_436), .B2(n_0_119), 
      .C1(n_164), .C2(n_0_117), .ZN(n_0_100));
   INV_X1 i_0_216 (.A(n_0_120), .ZN(product[9]));
   AOI222_X1 i_0_217 (.A1(n_435), .A2(n_0_138), .B1(n_435), .B2(n_0_139), 
      .C1(n_173), .C2(n_0_137), .ZN(n_0_120));
   INV_X1 i_0_252 (.A(n_0_140), .ZN(product[8]));
   AOI222_X1 i_0_253 (.A1(n_434), .A2(n_0_158), .B1(n_434), .B2(n_0_159), 
      .C1(n_183), .C2(n_0_157), .ZN(n_0_140));
   INV_X1 i_0_288 (.A(n_0_160), .ZN(product[7]));
   AOI222_X1 i_0_289 (.A1(n_433), .A2(n_0_178), .B1(n_433), .B2(n_0_179), 
      .C1(n_194), .C2(n_0_177), .ZN(n_0_160));
   INV_X1 i_0_324 (.A(n_0_180), .ZN(product[6]));
   AOI222_X1 i_0_325 (.A1(n_432), .A2(n_0_198), .B1(n_432), .B2(n_0_199), 
      .C1(n_206), .C2(n_0_197), .ZN(n_0_180));
   INV_X1 i_0_360 (.A(n_0_200), .ZN(product[5]));
   AOI222_X1 i_0_361 (.A1(n_431), .A2(n_0_218), .B1(n_431), .B2(n_0_219), 
      .C1(n_134), .C2(n_0_217), .ZN(n_0_200));
   AOI221_X1 i_0_389 (.A(n_0_216), .B1(n_440), .B2(n_0_218), .C1(n_439), 
      .C2(n_0_219), .ZN(n_0_214));
   AND2_X1 i_0_392 (.A1(n_112), .A2(n_0_217), .ZN(n_0_216));
   INV_X1 i_0_396 (.A(n_0_220), .ZN(product[4]));
   AOI222_X1 i_0_397 (.A1(n_80), .A2(n_0_2), .B1(n_96), .B2(n_0_3), .C1(n_113), 
      .C2(n_0_1), .ZN(n_0_220));
   AOI222_X1 i_0_417 (.A1(n_90), .A2(n_0_2), .B1(n_106), .B2(n_0_3), .C1(n_114), 
      .C2(n_0_1), .ZN(n_0_230));
   AOI222_X1 i_0_419 (.A1(n_107), .A2(n_0_3), .B1(n_91), .B2(n_0_2), .C1(n_236), 
      .C2(n_0_1), .ZN(n_0_231));
   AOI221_X1 i_0_425 (.A(n_0_0), .B1(n_94), .B2(n_0_2), .C1(n_110), .C2(n_0_3), 
      .ZN(n_0_234));
   INV_X1 i_0_426 (.A(n_0_235), .ZN(n_112));
   AOI221_X1 i_0_427 (.A(n_0_0), .B1(n_95), .B2(n_0_2), .C1(n_111), .C2(n_0_3), 
      .ZN(n_0_235));
   AND2_X1 i_0_428 (.A1(n_115), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_432 (.A(n_0_4), .ZN(product[3]));
   AOI222_X1 i_0_433 (.A1(n_48), .A2(n_0_22), .B1(n_64), .B2(n_0_23), .C1(n_116), 
      .C2(n_0_21), .ZN(n_0_4));
   INV_X1 i_0_434 (.A(n_0_5), .ZN(n_113));
   AOI222_X1 i_0_435 (.A1(n_49), .A2(n_0_22), .B1(n_65), .B2(n_0_23), .C1(n_140), 
      .C2(n_0_21), .ZN(n_0_5));
   AOI222_X1 i_0_451 (.A1(n_57), .A2(n_0_22), .B1(n_73), .B2(n_0_23), .C1(n_117), 
      .C2(n_0_21), .ZN(n_0_13));
   AOI222_X1 i_0_453 (.A1(n_58), .A2(n_0_22), .B1(n_74), .B2(n_0_23), .C1(n_118), 
      .C2(n_0_21), .ZN(n_0_14));
   INV_X1 i_0_454 (.A(n_0_15), .ZN(n_114));
   AOI222_X1 i_0_455 (.A1(n_59), .A2(n_0_22), .B1(n_75), .B2(n_0_23), .C1(n_245), 
      .C2(n_0_21), .ZN(n_0_15));
   AOI222_X1 i_0_459 (.A1(n_77), .A2(n_0_23), .B1(n_61), .B2(n_0_22), .C1(n_119), 
      .C2(n_0_21), .ZN(n_0_17));
   AOI221_X1 i_0_461 (.A(n_0_20), .B1(n_62), .B2(n_0_22), .C1(n_78), .C2(n_0_23), 
      .ZN(n_0_18));
   INV_X1 i_0_462 (.A(n_0_19), .ZN(n_115));
   AOI221_X1 i_0_463 (.A(n_0_20), .B1(n_63), .B2(n_0_22), .C1(n_79), .C2(n_0_23), 
      .ZN(n_0_19));
   AND2_X1 i_0_464 (.A1(n_120), .A2(n_0_21), .ZN(n_0_20));
   INV_X1 i_0_468 (.A(n_0_24), .ZN(product[2]));
   AOI222_X1 i_0_469 (.A1(n_16), .A2(n_0_42), .B1(n_32), .B2(n_0_43), .C1(n_142), 
      .C2(n_0_41), .ZN(n_0_24));
   INV_X1 i_0_470 (.A(n_0_25), .ZN(n_116));
   AOI222_X1 i_0_471 (.A1(n_17), .A2(n_0_42), .B1(n_33), .B2(n_0_43), .C1(n_143), 
      .C2(n_0_41), .ZN(n_0_25));
   INV_X1 i_0_488 (.A(n_0_34), .ZN(n_117));
   AOI222_X1 i_0_489 (.A1(n_26), .A2(n_0_42), .B1(n_42), .B2(n_0_43), .C1(n_121), 
      .C2(n_0_41), .ZN(n_0_34));
   INV_X1 i_0_490 (.A(n_0_35), .ZN(n_118));
   AOI222_X1 i_0_491 (.A1(n_27), .A2(n_0_42), .B1(n_43), .B2(n_0_43), .C1(n_253), 
      .C2(n_0_41), .ZN(n_0_35));
   AOI222_X1 i_0_495 (.A1(n_45), .A2(n_0_43), .B1(n_29), .B2(n_0_42), .C1(n_122), 
      .C2(n_0_41), .ZN(n_0_37));
   INV_X1 i_0_496 (.A(n_0_38), .ZN(n_119));
   AOI221_X1 i_0_497 (.A(n_0_40), .B1(n_30), .B2(n_0_42), .C1(n_46), .C2(n_0_43), 
      .ZN(n_0_38));
   INV_X1 i_0_498 (.A(n_0_39), .ZN(n_120));
   AOI221_X1 i_0_499 (.A(n_0_40), .B1(n_31), .B2(n_0_42), .C1(n_47), .C2(n_0_43), 
      .ZN(n_0_39));
   AND2_X1 i_0_500 (.A1(n_123), .A2(n_0_41), .ZN(n_0_40));
   INV_X1 i_0_504 (.A(n_0_44), .ZN(product[1]));
   AOI222_X1 i_0_505 (.A1(n_0), .A2(n_0_70), .B1(B[0]), .B2(n_0_59), .C1(n_146), 
      .C2(n_0_68), .ZN(n_0_44));
   AOI222_X1 i_0_517 (.A1(n_6), .A2(n_0_70), .B1(n_257), .B2(n_0_59), .C1(n_258), 
      .C2(n_0_68), .ZN(n_0_50));
   INV_X1 i_0_526 (.A(n_0_55), .ZN(n_121));
   AOI222_X1 i_0_527 (.A1(n_262), .A2(n_0_59), .B1(n_11), .B2(n_0_70), .C1(n_263), 
      .C2(n_0_68), .ZN(n_0_55));
   AOI222_X1 i_0_531 (.A1(n_13), .A2(n_0_70), .B1(n_264), .B2(n_0_59), .C1(n_125), 
      .C2(n_0_68), .ZN(n_0_57));
   INV_X1 i_0_532 (.A(n_0_58), .ZN(n_122));
   AOI222_X1 i_0_533 (.A1(n_125), .A2(n_0_59), .B1(n_14), .B2(n_0_70), .C1(n_126), 
      .C2(n_0_68), .ZN(n_0_58));
   INV_X1 i_0_536 (.A(n_0_69), .ZN(n_123));
   AOI22_X1 i_0_537 (.A1(n_15), .A2(n_0_70), .B1(A[1]), .B2(n_126), .ZN(n_0_69));
   AND2_X1 i_0_539 (.A1(B[0]), .A2(A[0]), .ZN(product[0]));
   AND2_X1 i_0_540 (.A1(A[0]), .A2(n_126), .ZN(n_124));
   AOI21_X1 i_0_554 (.A(n_0_71), .B1(B[15]), .B2(n_0_72), .ZN(n_125));
   XNOR2_X1 i_0_555 (.A(B[15]), .B(n_0_71), .ZN(n_126));
   NOR2_X1 i_0_556 (.A1(B[15]), .A2(n_0_72), .ZN(n_0_71));
   INV_X1 i_0_557 (.A(n_0_73), .ZN(n_0_72));
   NOR2_X1 i_0_558 (.A1(B[15]), .A2(n_0_74), .ZN(n_0_73));
   INV_X1 i_0_559 (.A(n_0_75), .ZN(n_0_74));
   INV_X1 i_0_584 (.A(A[1]), .ZN(n_0_153));
   INV_X1 i_0_585 (.A(A[2]), .ZN(n_0_154));
   INV_X1 i_0_586 (.A(A[3]), .ZN(n_0_155));
   INV_X1 i_0_587 (.A(A[4]), .ZN(n_0_156));
   INV_X1 i_0_588 (.A(A[5]), .ZN(n_0_173));
   INV_X1 i_0_589 (.A(A[6]), .ZN(n_0_174));
   INV_X1 i_0_590 (.A(A[7]), .ZN(n_0_175));
   INV_X1 i_0_591 (.A(A[8]), .ZN(n_0_176));
   INV_X1 i_0_592 (.A(A[9]), .ZN(n_0_194));
   INV_X1 i_0_593 (.A(A[10]), .ZN(n_0_195));
   INV_X1 i_0_594 (.A(A[11]), .ZN(n_0_196));
   INV_X1 i_0_595 (.A(A[15]), .ZN(n_0_215));
   NAND3_X1 i_0_0 (.A1(n_0_6), .A2(n_0_8), .A3(n_0_7), .ZN(product[19]));
   NAND2_X1 i_0_1 (.A1(n_430), .A2(n_0_79), .ZN(n_0_6));
   NAND2_X1 i_0_2 (.A1(n_127), .A2(n_0_77), .ZN(n_0_7));
   NAND2_X1 i_0_3 (.A1(n_423), .A2(n_0_78), .ZN(n_0_8));
   OAI21_X1 i_0_4 (.A(n_0_9), .B1(n_0_11), .B2(n_0_141), .ZN(n_127));
   AOI22_X1 i_0_5 (.A1(n_408), .A2(n_0_98), .B1(n_128), .B2(n_0_97), .ZN(n_0_9));
   OR2_X1 i_0_6 (.A1(n_0_99), .A2(n_0_98), .ZN(n_0_10));
   INV_X1 i_0_7 (.A(n_416), .ZN(n_0_11));
   OAI21_X1 i_0_8 (.A(n_0_12), .B1(n_0_16), .B2(n_0_166), .ZN(n_128));
   AOI22_X1 i_0_9 (.A1(n_391), .A2(n_0_118), .B1(n_129), .B2(n_0_117), .ZN(
      n_0_12));
   INV_X1 i_0_10 (.A(n_400), .ZN(n_0_16));
   OAI21_X1 i_0_11 (.A(n_0_26), .B1(n_0_28), .B2(n_0_193), .ZN(n_129));
   AOI22_X1 i_0_12 (.A1(n_372), .A2(n_0_138), .B1(n_130), .B2(n_0_137), .ZN(
      n_0_26));
   INV_X1 i_0_13 (.A(n_382), .ZN(n_0_28));
   OAI21_X1 i_0_14 (.A(n_0_29), .B1(n_0_30), .B2(n_0_229), .ZN(n_130));
   AOI22_X1 i_0_15 (.A1(n_351), .A2(n_0_158), .B1(n_131), .B2(n_0_157), .ZN(
      n_0_29));
   INV_X1 i_0_16 (.A(n_362), .ZN(n_0_30));
   OAI21_X1 i_0_17 (.A(n_0_31), .B1(n_0_33), .B2(n_0_257), .ZN(n_131));
   AOI22_X1 i_0_18 (.A1(n_328), .A2(n_0_178), .B1(n_132), .B2(n_0_177), .ZN(
      n_0_31));
   NAND2_X1 i_0_19 (.A1(n_0_257), .A2(n_0_246), .ZN(n_0_32));
   INV_X1 i_0_20 (.A(n_340), .ZN(n_0_33));
   OAI21_X1 i_0_21 (.A(n_0_36), .B1(n_0_45), .B2(n_0_283), .ZN(n_132));
   AOI22_X1 i_0_22 (.A1(n_303), .A2(n_0_198), .B1(n_133), .B2(n_0_197), .ZN(
      n_0_36));
   INV_X1 i_0_23 (.A(n_316), .ZN(n_0_45));
   INV_X1 i_0_24 (.A(n_0_214), .ZN(n_133));
   NAND2_X1 i_0_25 (.A1(n_0_47), .A2(n_0_46), .ZN(n_134));
   NAND2_X1 i_0_26 (.A1(n_97), .A2(n_0_3), .ZN(n_0_46));
   AOI22_X1 i_0_27 (.A1(n_81), .A2(n_0_2), .B1(n_138), .B2(n_0_1), .ZN(n_0_47));
   NAND2_X1 i_0_28 (.A1(n_99), .A2(n_0_3), .ZN(n_0_48));
   AOI22_X1 i_0_29 (.A1(n_83), .A2(n_0_2), .B1(n_139), .B2(n_0_1), .ZN(n_0_49));
   OAI21_X1 i_0_30 (.A(n_0_52), .B1(n_0_156), .B2(A[3]), .ZN(n_0_51));
   NAND2_X1 i_0_31 (.A1(n_0_53), .A2(n_0_54), .ZN(n_0_52));
   INV_X1 i_0_32 (.A(n_0_155), .ZN(n_0_53));
   INV_X1 i_0_33 (.A(A[4]), .ZN(n_0_54));
   INV_X1 i_0_34 (.A(n_0_230), .ZN(n_135));
   INV_X1 i_0_35 (.A(n_0_231), .ZN(n_136));
   INV_X1 i_0_36 (.A(n_0_234), .ZN(n_137));
   OAI211_X1 i_0_37 (.A(n_0_56), .B(n_0_63), .C1(n_0_27), .C2(n_0_65), .ZN(n_138));
   NAND2_X1 i_0_38 (.A1(n_50), .A2(n_0_22), .ZN(n_0_56));
   NAND2_X1 i_0_39 (.A1(n_66), .A2(n_0_23), .ZN(n_0_63));
   OAI211_X1 i_0_40 (.A(n_0_66), .B(n_0_64), .C1(n_0_67), .C2(n_0_65), .ZN(n_139));
   NAND2_X1 i_0_41 (.A1(n_52), .A2(n_0_22), .ZN(n_0_64));
   INV_X1 i_0_42 (.A(n_0_21), .ZN(n_0_65));
   NAND2_X1 i_0_43 (.A1(n_68), .A2(n_0_23), .ZN(n_0_66));
   INV_X1 i_0_44 (.A(n_141), .ZN(n_0_67));
   NAND2_X1 i_0_45 (.A1(n_0_81), .A2(n_0_76), .ZN(n_140));
   NAND2_X1 i_0_46 (.A1(n_34), .A2(n_0_43), .ZN(n_0_76));
   AOI22_X1 i_0_47 (.A1(n_18), .A2(n_0_42), .B1(n_144), .B2(n_0_41), .ZN(n_0_81));
   NAND2_X1 i_0_48 (.A1(n_0_83), .A2(n_0_82), .ZN(n_141));
   NAND2_X1 i_0_49 (.A1(n_21), .A2(n_0_42), .ZN(n_0_82));
   AOI22_X1 i_0_50 (.A1(n_37), .A2(n_0_43), .B1(n_145), .B2(n_0_41), .ZN(n_0_83));
   OAI21_X1 i_0_51 (.A(n_0_88), .B1(n_0_104), .B2(n_0_84), .ZN(n_142));
   INV_X1 i_0_52 (.A(n_0_85), .ZN(n_0_84));
   NAND2_X1 i_0_53 (.A1(n_0_87), .A2(n_0_86), .ZN(n_0_85));
   NAND2_X1 i_0_54 (.A1(A[1]), .A2(n_147), .ZN(n_0_86));
   NAND2_X1 i_0_55 (.A1(n_0_92), .A2(n_1), .ZN(n_0_87));
   NAND3_X1 i_0_56 (.A1(n_0_96), .A2(n_0_104), .A3(n_146), .ZN(n_0_88));
   OAI21_X1 i_0_57 (.A(n_0_94), .B1(n_0_104), .B2(n_0_89), .ZN(n_143));
   INV_X1 i_0_58 (.A(n_0_90), .ZN(n_0_89));
   NAND2_X1 i_0_59 (.A1(n_0_91), .A2(n_0_93), .ZN(n_0_90));
   NAND2_X1 i_0_60 (.A1(n_0_92), .A2(n_2), .ZN(n_0_91));
   INV_X1 i_0_61 (.A(A[1]), .ZN(n_0_92));
   NAND2_X1 i_0_62 (.A1(A[1]), .A2(n_148), .ZN(n_0_93));
   NAND3_X1 i_0_63 (.A1(n_0_96), .A2(n_0_104), .A3(n_147), .ZN(n_0_94));
   NAND3_X1 i_0_64 (.A1(n_0_103), .A2(n_0_101), .A3(n_0_95), .ZN(n_144));
   NAND3_X1 i_0_65 (.A1(n_0_96), .A2(n_0_104), .A3(n_148), .ZN(n_0_95));
   INV_X1 i_0_66 (.A(n_0_153), .ZN(n_0_96));
   NAND2_X1 i_0_67 (.A1(n_0_68), .A2(n_255), .ZN(n_0_101));
   NAND2_X1 i_0_68 (.A1(A[1]), .A2(A[0]), .ZN(n_0_102));
   NAND2_X1 i_0_69 (.A1(n_3), .A2(n_0_70), .ZN(n_0_103));
   INV_X1 i_0_70 (.A(A[0]), .ZN(n_0_104));
   INV_X1 i_0_71 (.A(n_0_50), .ZN(n_145));
   AOI21_X1 i_0_72 (.A(n_0_136), .B1(B[1]), .B2(B[0]), .ZN(n_146));
   AOI21_X1 i_0_73 (.A(n_0_134), .B1(B[2]), .B2(n_0_135), .ZN(n_147));
   AOI21_X1 i_0_74 (.A(n_0_132), .B1(B[3]), .B2(n_0_133), .ZN(n_148));
   INV_X1 i_0_75 (.A(n_0_105), .ZN(n_0_75));
   OR2_X1 i_0_76 (.A1(n_0_391), .A2(B[15]), .ZN(n_0_105));
   INV_X1 i_0_77 (.A(n_239), .ZN(n_0_27));
   OAI21_X1 i_0_78 (.A(n_0_106), .B1(n_0_107), .B2(n_0_113), .ZN(product[15]));
   AOI22_X1 i_0_79 (.A1(n_426), .A2(n_0_79), .B1(n_152), .B2(n_0_77), .ZN(
      n_0_106));
   INV_X1 i_0_80 (.A(n_419), .ZN(n_0_107));
   OAI21_X1 i_0_81 (.A(n_0_108), .B1(n_0_109), .B2(n_0_113), .ZN(product[16]));
   AOI22_X1 i_0_82 (.A1(n_427), .A2(n_0_79), .B1(n_153), .B2(n_0_77), .ZN(
      n_0_108));
   INV_X1 i_0_83 (.A(n_420), .ZN(n_0_109));
   OAI21_X1 i_0_84 (.A(n_0_110), .B1(n_0_111), .B2(n_0_113), .ZN(product[17]));
   AOI22_X1 i_0_85 (.A1(n_428), .A2(n_0_79), .B1(n_154), .B2(n_0_77), .ZN(
      n_0_110));
   INV_X1 i_0_86 (.A(n_421), .ZN(n_0_111));
   OAI21_X1 i_0_87 (.A(n_0_112), .B1(n_0_114), .B2(n_0_113), .ZN(product[18]));
   AOI22_X1 i_0_88 (.A1(n_429), .A2(n_0_79), .B1(n_155), .B2(n_0_77), .ZN(
      n_0_112));
   NOR2_X1 i_0_89 (.A1(n_0_79), .A2(n_0_78), .ZN(n_0_77));
   NOR2_X1 i_0_90 (.A1(n_0_215), .A2(A[11]), .ZN(n_0_79));
   INV_X1 i_0_91 (.A(n_0_78), .ZN(n_0_113));
   NOR2_X1 i_0_92 (.A1(A[15]), .A2(n_0_196), .ZN(n_0_78));
   INV_X1 i_0_93 (.A(n_422), .ZN(n_0_114));
   NAND2_X1 i_0_94 (.A1(n_0_115), .A2(n_0_116), .ZN(n_149));
   AOI22_X1 i_0_95 (.A1(n_409), .A2(n_0_99), .B1(n_0_97), .B2(n_157), .ZN(
      n_0_115));
   NAND2_X1 i_0_96 (.A1(n_401), .A2(n_0_98), .ZN(n_0_116));
   OAI21_X1 i_0_97 (.A(n_0_121), .B1(n_0_122), .B2(n_0_141), .ZN(n_150));
   AOI22_X1 i_0_98 (.A1(n_402), .A2(n_0_98), .B1(n_0_97), .B2(n_158), .ZN(
      n_0_121));
   INV_X1 i_0_99 (.A(n_410), .ZN(n_0_122));
   OAI21_X1 i_0_100 (.A(n_0_123), .B1(n_0_124), .B2(n_0_141), .ZN(n_151));
   AOI22_X1 i_0_101 (.A1(n_403), .A2(n_0_98), .B1(n_0_97), .B2(n_159), .ZN(
      n_0_123));
   INV_X1 i_0_102 (.A(n_411), .ZN(n_0_124));
   OAI21_X1 i_0_103 (.A(n_0_125), .B1(n_0_126), .B2(n_0_141), .ZN(n_152));
   AOI22_X1 i_0_104 (.A1(n_404), .A2(n_0_98), .B1(n_0_97), .B2(n_160), .ZN(
      n_0_125));
   INV_X1 i_0_105 (.A(n_412), .ZN(n_0_126));
   OAI21_X1 i_0_106 (.A(n_0_127), .B1(n_0_128), .B2(n_0_141), .ZN(n_153));
   AOI22_X1 i_0_107 (.A1(n_405), .A2(n_0_98), .B1(n_0_97), .B2(n_161), .ZN(
      n_0_127));
   INV_X1 i_0_114 (.A(n_413), .ZN(n_0_128));
   OAI21_X1 i_0_115 (.A(n_0_129), .B1(n_0_130), .B2(n_0_141), .ZN(n_154));
   AOI22_X1 i_0_116 (.A1(n_406), .A2(n_0_98), .B1(n_0_97), .B2(n_162), .ZN(
      n_0_129));
   INV_X1 i_0_117 (.A(n_414), .ZN(n_0_130));
   OAI21_X1 i_0_118 (.A(n_0_131), .B1(n_0_142), .B2(n_0_141), .ZN(n_155));
   AOI22_X1 i_0_119 (.A1(n_407), .A2(n_0_98), .B1(n_0_97), .B2(n_163), .ZN(
      n_0_131));
   NOR2_X1 i_0_120 (.A1(n_0_195), .A2(A[11]), .ZN(n_0_98));
   INV_X1 i_0_121 (.A(n_0_10), .ZN(n_0_97));
   INV_X1 i_0_122 (.A(n_0_99), .ZN(n_0_141));
   NOR2_X1 i_0_123 (.A1(n_0_196), .A2(A[10]), .ZN(n_0_99));
   INV_X1 i_0_124 (.A(n_415), .ZN(n_0_142));
   OAI21_X1 i_0_125 (.A(n_0_143), .B1(n_0_144), .B2(n_0_166), .ZN(n_156));
   AOI22_X1 i_0_126 (.A1(n_383), .A2(n_0_118), .B1(n_165), .B2(n_0_117), 
      .ZN(n_0_143));
   INV_X1 i_0_127 (.A(n_392), .ZN(n_0_144));
   OAI21_X1 i_0_128 (.A(n_0_145), .B1(n_0_146), .B2(n_0_166), .ZN(n_157));
   AOI22_X1 i_0_129 (.A1(n_384), .A2(n_0_118), .B1(n_166), .B2(n_0_117), 
      .ZN(n_0_145));
   INV_X1 i_0_130 (.A(n_393), .ZN(n_0_146));
   OAI21_X1 i_0_131 (.A(n_0_147), .B1(n_0_148), .B2(n_0_166), .ZN(n_158));
   AOI22_X1 i_0_132 (.A1(n_385), .A2(n_0_118), .B1(n_167), .B2(n_0_117), 
      .ZN(n_0_147));
   INV_X1 i_0_133 (.A(n_394), .ZN(n_0_148));
   OAI21_X1 i_0_134 (.A(n_0_149), .B1(n_0_150), .B2(n_0_166), .ZN(n_159));
   AOI22_X1 i_0_135 (.A1(n_386), .A2(n_0_118), .B1(n_168), .B2(n_0_117), 
      .ZN(n_0_149));
   INV_X1 i_0_136 (.A(n_395), .ZN(n_0_150));
   OAI21_X1 i_0_137 (.A(n_0_151), .B1(n_0_152), .B2(n_0_166), .ZN(n_160));
   AOI22_X1 i_0_138 (.A1(n_387), .A2(n_0_118), .B1(n_169), .B2(n_0_117), 
      .ZN(n_0_151));
   INV_X1 i_0_139 (.A(n_396), .ZN(n_0_152));
   OAI21_X1 i_0_140 (.A(n_0_161), .B1(n_0_162), .B2(n_0_166), .ZN(n_161));
   AOI22_X1 i_0_141 (.A1(n_388), .A2(n_0_118), .B1(n_170), .B2(n_0_117), 
      .ZN(n_0_161));
   INV_X1 i_0_142 (.A(n_397), .ZN(n_0_162));
   OAI21_X1 i_0_143 (.A(n_0_163), .B1(n_0_164), .B2(n_0_166), .ZN(n_162));
   AOI22_X1 i_0_146 (.A1(n_389), .A2(n_0_118), .B1(n_171), .B2(n_0_117), 
      .ZN(n_0_163));
   INV_X1 i_0_147 (.A(n_398), .ZN(n_0_164));
   OAI21_X1 i_0_148 (.A(n_0_165), .B1(n_0_167), .B2(n_0_166), .ZN(n_163));
   AOI22_X1 i_0_149 (.A1(n_390), .A2(n_0_118), .B1(n_172), .B2(n_0_117), 
      .ZN(n_0_165));
   NOR2_X1 i_0_150 (.A1(n_0_119), .A2(n_0_118), .ZN(n_0_117));
   NOR2_X1 i_0_151 (.A1(A[10]), .A2(n_0_194), .ZN(n_0_118));
   INV_X1 i_0_152 (.A(n_0_119), .ZN(n_0_166));
   NOR2_X1 i_0_153 (.A1(n_0_195), .A2(A[9]), .ZN(n_0_119));
   INV_X1 i_0_154 (.A(n_399), .ZN(n_0_167));
   OAI21_X1 i_0_155 (.A(n_0_168), .B1(n_0_169), .B2(n_0_193), .ZN(n_164));
   AOI22_X1 i_0_156 (.A1(n_363), .A2(n_0_138), .B1(n_174), .B2(n_0_137), 
      .ZN(n_0_168));
   INV_X1 i_0_157 (.A(n_373), .ZN(n_0_169));
   NAND2_X1 i_0_158 (.A1(n_0_171), .A2(n_0_170), .ZN(n_165));
   AOI22_X1 i_0_159 (.A1(n_374), .A2(n_0_139), .B1(n_175), .B2(n_0_137), 
      .ZN(n_0_170));
   NAND2_X1 i_0_160 (.A1(n_364), .A2(n_0_138), .ZN(n_0_171));
   NAND2_X1 i_0_161 (.A1(n_0_181), .A2(n_0_172), .ZN(n_166));
   AOI22_X1 i_0_162 (.A1(n_375), .A2(n_0_139), .B1(n_176), .B2(n_0_137), 
      .ZN(n_0_172));
   NAND2_X1 i_0_163 (.A1(n_365), .A2(n_0_138), .ZN(n_0_181));
   OAI21_X1 i_0_164 (.A(n_0_182), .B1(n_0_183), .B2(n_0_193), .ZN(n_167));
   AOI22_X1 i_0_165 (.A1(n_366), .A2(n_0_138), .B1(n_177), .B2(n_0_137), 
      .ZN(n_0_182));
   INV_X1 i_0_166 (.A(n_376), .ZN(n_0_183));
   OAI21_X1 i_0_167 (.A(n_0_184), .B1(n_0_185), .B2(n_0_193), .ZN(n_168));
   AOI22_X1 i_0_168 (.A1(n_367), .A2(n_0_138), .B1(n_178), .B2(n_0_137), 
      .ZN(n_0_184));
   INV_X1 i_0_169 (.A(n_377), .ZN(n_0_185));
   OAI21_X1 i_0_170 (.A(n_0_186), .B1(n_0_187), .B2(n_0_193), .ZN(n_169));
   AOI22_X1 i_0_171 (.A1(n_368), .A2(n_0_138), .B1(n_179), .B2(n_0_137), 
      .ZN(n_0_186));
   INV_X1 i_0_172 (.A(n_378), .ZN(n_0_187));
   OAI21_X1 i_0_173 (.A(n_0_188), .B1(n_0_189), .B2(n_0_193), .ZN(n_170));
   AOI22_X1 i_0_174 (.A1(n_369), .A2(n_0_138), .B1(n_180), .B2(n_0_137), 
      .ZN(n_0_188));
   INV_X1 i_0_175 (.A(n_379), .ZN(n_0_189));
   OAI21_X1 i_0_176 (.A(n_0_190), .B1(n_0_191), .B2(n_0_193), .ZN(n_171));
   AOI22_X1 i_0_177 (.A1(n_370), .A2(n_0_138), .B1(n_181), .B2(n_0_137), 
      .ZN(n_0_190));
   INV_X1 i_0_178 (.A(n_380), .ZN(n_0_191));
   OAI21_X1 i_0_179 (.A(n_0_192), .B1(n_0_201), .B2(n_0_193), .ZN(n_172));
   AOI22_X1 i_0_182 (.A1(n_371), .A2(n_0_138), .B1(n_182), .B2(n_0_137), 
      .ZN(n_0_192));
   NOR2_X1 i_0_183 (.A1(n_0_139), .A2(n_0_138), .ZN(n_0_137));
   NOR2_X1 i_0_184 (.A1(n_0_176), .A2(A[9]), .ZN(n_0_138));
   INV_X1 i_0_185 (.A(n_0_139), .ZN(n_0_193));
   NOR2_X1 i_0_186 (.A1(n_0_194), .A2(A[8]), .ZN(n_0_139));
   INV_X1 i_0_187 (.A(n_381), .ZN(n_0_201));
   OAI21_X1 i_0_188 (.A(n_0_202), .B1(n_0_203), .B2(n_0_229), .ZN(n_173));
   AOI22_X1 i_0_189 (.A1(n_341), .A2(n_0_158), .B1(n_184), .B2(n_0_157), 
      .ZN(n_0_202));
   INV_X1 i_0_190 (.A(n_352), .ZN(n_0_203));
   OAI21_X1 i_0_191 (.A(n_0_204), .B1(n_0_205), .B2(n_0_209), .ZN(n_174));
   AOI22_X1 i_0_192 (.A1(n_353), .A2(n_0_159), .B1(n_185), .B2(n_0_157), 
      .ZN(n_0_204));
   INV_X1 i_0_193 (.A(n_342), .ZN(n_0_205));
   OAI21_X1 i_0_194 (.A(n_0_206), .B1(n_0_207), .B2(n_0_209), .ZN(n_175));
   AOI22_X1 i_0_195 (.A1(n_354), .A2(n_0_159), .B1(n_186), .B2(n_0_157), 
      .ZN(n_0_206));
   INV_X1 i_0_196 (.A(n_343), .ZN(n_0_207));
   OAI21_X1 i_0_197 (.A(n_0_208), .B1(n_0_210), .B2(n_0_209), .ZN(n_176));
   AOI22_X1 i_0_198 (.A1(n_355), .A2(n_0_159), .B1(n_187), .B2(n_0_157), 
      .ZN(n_0_208));
   INV_X1 i_0_199 (.A(n_0_158), .ZN(n_0_209));
   INV_X1 i_0_200 (.A(n_344), .ZN(n_0_210));
   OAI21_X1 i_0_201 (.A(n_0_211), .B1(n_0_212), .B2(n_0_229), .ZN(n_177));
   AOI22_X1 i_0_202 (.A1(n_345), .A2(n_0_158), .B1(n_188), .B2(n_0_157), 
      .ZN(n_0_211));
   INV_X1 i_0_203 (.A(n_356), .ZN(n_0_212));
   OAI21_X1 i_0_204 (.A(n_0_213), .B1(n_0_221), .B2(n_0_229), .ZN(n_178));
   AOI22_X1 i_0_205 (.A1(n_346), .A2(n_0_158), .B1(n_189), .B2(n_0_157), 
      .ZN(n_0_213));
   INV_X1 i_0_206 (.A(n_357), .ZN(n_0_221));
   OAI21_X1 i_0_207 (.A(n_0_222), .B1(n_0_223), .B2(n_0_229), .ZN(n_179));
   AOI22_X1 i_0_208 (.A1(n_347), .A2(n_0_158), .B1(n_190), .B2(n_0_157), 
      .ZN(n_0_222));
   INV_X1 i_0_209 (.A(n_358), .ZN(n_0_223));
   OAI21_X1 i_0_210 (.A(n_0_224), .B1(n_0_225), .B2(n_0_229), .ZN(n_180));
   AOI22_X1 i_0_211 (.A1(n_348), .A2(n_0_158), .B1(n_191), .B2(n_0_157), 
      .ZN(n_0_224));
   INV_X1 i_0_212 (.A(n_359), .ZN(n_0_225));
   OAI21_X1 i_0_213 (.A(n_0_226), .B1(n_0_227), .B2(n_0_229), .ZN(n_181));
   AOI22_X1 i_0_214 (.A1(n_349), .A2(n_0_158), .B1(n_192), .B2(n_0_157), 
      .ZN(n_0_226));
   INV_X1 i_0_215 (.A(n_360), .ZN(n_0_227));
   OAI21_X1 i_0_218 (.A(n_0_228), .B1(n_0_232), .B2(n_0_229), .ZN(n_182));
   AOI22_X1 i_0_219 (.A1(n_350), .A2(n_0_158), .B1(n_193), .B2(n_0_157), 
      .ZN(n_0_228));
   NOR2_X1 i_0_220 (.A1(n_0_159), .A2(n_0_158), .ZN(n_0_157));
   NOR2_X1 i_0_221 (.A1(A[8]), .A2(n_0_175), .ZN(n_0_158));
   INV_X1 i_0_222 (.A(n_0_159), .ZN(n_0_229));
   NOR2_X1 i_0_223 (.A1(n_0_176), .A2(A[7]), .ZN(n_0_159));
   INV_X1 i_0_224 (.A(n_361), .ZN(n_0_232));
   OAI21_X1 i_0_225 (.A(n_0_233), .B1(n_0_236), .B2(n_0_257), .ZN(n_183));
   AOI22_X1 i_0_226 (.A1(n_317), .A2(n_0_178), .B1(n_0_177), .B2(n_195), 
      .ZN(n_0_233));
   INV_X1 i_0_227 (.A(n_329), .ZN(n_0_236));
   OAI21_X1 i_0_228 (.A(n_0_237), .B1(n_0_238), .B2(n_0_246), .ZN(n_184));
   AOI22_X1 i_0_229 (.A1(n_330), .A2(n_0_179), .B1(n_0_177), .B2(n_196), 
      .ZN(n_0_237));
   INV_X1 i_0_230 (.A(n_318), .ZN(n_0_238));
   OAI21_X1 i_0_231 (.A(n_0_239), .B1(n_0_240), .B2(n_0_246), .ZN(n_185));
   AOI22_X1 i_0_232 (.A1(n_331), .A2(n_0_179), .B1(n_0_177), .B2(n_197), 
      .ZN(n_0_239));
   INV_X1 i_0_233 (.A(n_319), .ZN(n_0_240));
   OAI21_X1 i_0_234 (.A(n_0_241), .B1(n_0_242), .B2(n_0_246), .ZN(n_186));
   AOI22_X1 i_0_235 (.A1(n_332), .A2(n_0_179), .B1(n_0_177), .B2(n_198), 
      .ZN(n_0_241));
   INV_X1 i_0_236 (.A(n_320), .ZN(n_0_242));
   OAI21_X1 i_0_237 (.A(n_0_243), .B1(n_0_244), .B2(n_0_246), .ZN(n_187));
   AOI22_X1 i_0_238 (.A1(n_333), .A2(n_0_179), .B1(n_0_177), .B2(n_199), 
      .ZN(n_0_243));
   INV_X1 i_0_239 (.A(n_321), .ZN(n_0_244));
   OAI21_X1 i_0_240 (.A(n_0_245), .B1(n_0_247), .B2(n_0_246), .ZN(n_188));
   AOI22_X1 i_0_241 (.A1(n_334), .A2(n_0_179), .B1(n_0_177), .B2(n_200), 
      .ZN(n_0_245));
   INV_X1 i_0_242 (.A(n_0_178), .ZN(n_0_246));
   INV_X1 i_0_243 (.A(n_322), .ZN(n_0_247));
   OAI21_X1 i_0_244 (.A(n_0_248), .B1(n_0_249), .B2(n_0_257), .ZN(n_189));
   AOI22_X1 i_0_245 (.A1(n_323), .A2(n_0_178), .B1(n_0_177), .B2(n_201), 
      .ZN(n_0_248));
   INV_X1 i_0_246 (.A(n_335), .ZN(n_0_249));
   OAI21_X1 i_0_247 (.A(n_0_250), .B1(n_0_251), .B2(n_0_257), .ZN(n_190));
   AOI22_X1 i_0_248 (.A1(n_324), .A2(n_0_178), .B1(n_0_177), .B2(n_202), 
      .ZN(n_0_250));
   INV_X1 i_0_249 (.A(n_336), .ZN(n_0_251));
   OAI21_X1 i_0_250 (.A(n_0_252), .B1(n_0_253), .B2(n_0_257), .ZN(n_191));
   AOI22_X1 i_0_251 (.A1(n_325), .A2(n_0_178), .B1(n_0_177), .B2(n_203), 
      .ZN(n_0_252));
   INV_X1 i_0_254 (.A(n_337), .ZN(n_0_253));
   OAI21_X1 i_0_255 (.A(n_0_254), .B1(n_0_255), .B2(n_0_257), .ZN(n_192));
   AOI22_X1 i_0_256 (.A1(n_326), .A2(n_0_178), .B1(n_0_177), .B2(n_204), 
      .ZN(n_0_254));
   INV_X1 i_0_257 (.A(n_338), .ZN(n_0_255));
   OAI21_X1 i_0_258 (.A(n_0_256), .B1(n_0_258), .B2(n_0_257), .ZN(n_193));
   AOI22_X1 i_0_259 (.A1(n_327), .A2(n_0_178), .B1(n_0_177), .B2(n_205), 
      .ZN(n_0_256));
   NOR2_X1 i_0_260 (.A1(n_0_174), .A2(A[7]), .ZN(n_0_178));
   INV_X1 i_0_261 (.A(n_0_32), .ZN(n_0_177));
   INV_X1 i_0_262 (.A(n_0_179), .ZN(n_0_257));
   NOR2_X1 i_0_263 (.A1(n_0_175), .A2(A[6]), .ZN(n_0_179));
   INV_X1 i_0_264 (.A(n_339), .ZN(n_0_258));
   OAI21_X1 i_0_265 (.A(n_0_259), .B1(n_0_260), .B2(n_0_283), .ZN(n_194));
   AOI22_X1 i_0_266 (.A1(n_291), .A2(n_0_198), .B1(n_207), .B2(n_0_197), 
      .ZN(n_0_259));
   INV_X1 i_0_267 (.A(n_304), .ZN(n_0_260));
   OAI21_X1 i_0_268 (.A(n_0_261), .B1(n_0_262), .B2(n_0_272), .ZN(n_195));
   AOI22_X1 i_0_269 (.A1(n_305), .A2(n_0_199), .B1(n_208), .B2(n_0_197), 
      .ZN(n_0_261));
   INV_X1 i_0_270 (.A(n_292), .ZN(n_0_262));
   OAI21_X1 i_0_271 (.A(n_0_263), .B1(n_0_264), .B2(n_0_272), .ZN(n_196));
   AOI22_X1 i_0_272 (.A1(n_306), .A2(n_0_199), .B1(n_209), .B2(n_0_197), 
      .ZN(n_0_263));
   INV_X1 i_0_273 (.A(n_293), .ZN(n_0_264));
   OAI21_X1 i_0_274 (.A(n_0_265), .B1(n_0_266), .B2(n_0_272), .ZN(n_197));
   AOI22_X1 i_0_275 (.A1(n_307), .A2(n_0_199), .B1(n_210), .B2(n_0_197), 
      .ZN(n_0_265));
   INV_X1 i_0_276 (.A(n_294), .ZN(n_0_266));
   OAI21_X1 i_0_277 (.A(n_0_267), .B1(n_0_268), .B2(n_0_272), .ZN(n_198));
   AOI22_X1 i_0_278 (.A1(n_308), .A2(n_0_199), .B1(n_211), .B2(n_0_197), 
      .ZN(n_0_267));
   INV_X1 i_0_279 (.A(n_295), .ZN(n_0_268));
   OAI21_X1 i_0_280 (.A(n_0_269), .B1(n_0_270), .B2(n_0_272), .ZN(n_199));
   AOI22_X1 i_0_281 (.A1(n_309), .A2(n_0_199), .B1(n_212), .B2(n_0_197), 
      .ZN(n_0_269));
   INV_X1 i_0_282 (.A(n_296), .ZN(n_0_270));
   OAI21_X1 i_0_283 (.A(n_0_271), .B1(n_0_273), .B2(n_0_272), .ZN(n_200));
   AOI22_X1 i_0_284 (.A1(n_310), .A2(n_0_199), .B1(n_213), .B2(n_0_197), 
      .ZN(n_0_271));
   INV_X1 i_0_285 (.A(n_0_198), .ZN(n_0_272));
   INV_X1 i_0_286 (.A(n_297), .ZN(n_0_273));
   OAI21_X1 i_0_287 (.A(n_0_274), .B1(n_0_275), .B2(n_0_283), .ZN(n_201));
   AOI22_X1 i_0_290 (.A1(n_298), .A2(n_0_198), .B1(n_214), .B2(n_0_197), 
      .ZN(n_0_274));
   INV_X1 i_0_291 (.A(n_311), .ZN(n_0_275));
   OAI21_X1 i_0_292 (.A(n_0_276), .B1(n_0_277), .B2(n_0_283), .ZN(n_202));
   AOI22_X1 i_0_293 (.A1(n_299), .A2(n_0_198), .B1(n_215), .B2(n_0_197), 
      .ZN(n_0_276));
   INV_X1 i_0_294 (.A(n_312), .ZN(n_0_277));
   OAI21_X1 i_0_295 (.A(n_0_278), .B1(n_0_279), .B2(n_0_283), .ZN(n_203));
   AOI22_X1 i_0_296 (.A1(n_300), .A2(n_0_198), .B1(n_216), .B2(n_0_197), 
      .ZN(n_0_278));
   INV_X1 i_0_297 (.A(n_313), .ZN(n_0_279));
   OAI21_X1 i_0_298 (.A(n_0_280), .B1(n_0_281), .B2(n_0_283), .ZN(n_204));
   AOI22_X1 i_0_299 (.A1(n_301), .A2(n_0_198), .B1(n_217), .B2(n_0_197), 
      .ZN(n_0_280));
   INV_X1 i_0_300 (.A(n_314), .ZN(n_0_281));
   OAI21_X1 i_0_301 (.A(n_0_282), .B1(n_0_284), .B2(n_0_283), .ZN(n_205));
   AOI22_X1 i_0_302 (.A1(n_302), .A2(n_0_198), .B1(n_218), .B2(n_0_197), 
      .ZN(n_0_282));
   NOR2_X1 i_0_303 (.A1(n_0_199), .A2(n_0_198), .ZN(n_0_197));
   NOR2_X1 i_0_304 (.A1(A[6]), .A2(n_0_173), .ZN(n_0_198));
   INV_X1 i_0_305 (.A(n_0_199), .ZN(n_0_283));
   NOR2_X1 i_0_306 (.A1(n_0_174), .A2(A[5]), .ZN(n_0_199));
   INV_X1 i_0_307 (.A(n_315), .ZN(n_0_284));
   OAI21_X1 i_0_308 (.A(n_0_285), .B1(n_0_286), .B2(n_0_312), .ZN(n_206));
   AOI22_X1 i_0_309 (.A1(n_265), .A2(n_0_218), .B1(n_219), .B2(n_0_217), 
      .ZN(n_0_285));
   INV_X1 i_0_310 (.A(n_278), .ZN(n_0_286));
   OAI21_X1 i_0_311 (.A(n_0_287), .B1(n_0_288), .B2(n_0_311), .ZN(n_207));
   AOI22_X1 i_0_312 (.A1(n_279), .A2(n_0_219), .B1(n_220), .B2(n_0_217), 
      .ZN(n_0_287));
   INV_X1 i_0_313 (.A(n_266), .ZN(n_0_288));
   OAI21_X1 i_0_314 (.A(n_0_289), .B1(n_0_290), .B2(n_0_311), .ZN(n_208));
   AOI22_X1 i_0_315 (.A1(n_280), .A2(n_0_219), .B1(n_221), .B2(n_0_217), 
      .ZN(n_0_289));
   INV_X1 i_0_316 (.A(n_267), .ZN(n_0_290));
   OAI21_X1 i_0_317 (.A(n_0_291), .B1(n_0_292), .B2(n_0_311), .ZN(n_209));
   AOI22_X1 i_0_318 (.A1(n_281), .A2(n_0_219), .B1(n_222), .B2(n_0_217), 
      .ZN(n_0_291));
   INV_X1 i_0_319 (.A(n_268), .ZN(n_0_292));
   OAI21_X1 i_0_320 (.A(n_0_293), .B1(n_0_294), .B2(n_0_311), .ZN(n_210));
   AOI22_X1 i_0_321 (.A1(n_282), .A2(n_0_219), .B1(n_223), .B2(n_0_217), 
      .ZN(n_0_293));
   INV_X1 i_0_322 (.A(n_269), .ZN(n_0_294));
   OAI21_X1 i_0_323 (.A(n_0_295), .B1(n_0_296), .B2(n_0_311), .ZN(n_211));
   AOI22_X1 i_0_326 (.A1(n_283), .A2(n_0_219), .B1(n_224), .B2(n_0_217), 
      .ZN(n_0_295));
   INV_X1 i_0_327 (.A(n_270), .ZN(n_0_296));
   OAI21_X1 i_0_328 (.A(n_0_297), .B1(n_0_298), .B2(n_0_311), .ZN(n_212));
   AOI22_X1 i_0_329 (.A1(n_284), .A2(n_0_219), .B1(n_225), .B2(n_0_217), 
      .ZN(n_0_297));
   INV_X1 i_0_330 (.A(n_271), .ZN(n_0_298));
   OAI21_X1 i_0_331 (.A(n_0_299), .B1(n_0_300), .B2(n_0_311), .ZN(n_213));
   AOI22_X1 i_0_332 (.A1(n_285), .A2(n_0_219), .B1(n_226), .B2(n_0_217), 
      .ZN(n_0_299));
   INV_X1 i_0_333 (.A(n_272), .ZN(n_0_300));
   OAI21_X1 i_0_334 (.A(n_0_301), .B1(n_0_302), .B2(n_0_312), .ZN(n_214));
   AOI22_X1 i_0_335 (.A1(n_273), .A2(n_0_218), .B1(n_135), .B2(n_0_217), 
      .ZN(n_0_301));
   INV_X1 i_0_336 (.A(n_286), .ZN(n_0_302));
   OAI21_X1 i_0_337 (.A(n_0_303), .B1(n_0_304), .B2(n_0_312), .ZN(n_215));
   AOI22_X1 i_0_338 (.A1(n_274), .A2(n_0_218), .B1(n_136), .B2(n_0_217), 
      .ZN(n_0_303));
   INV_X1 i_0_339 (.A(n_287), .ZN(n_0_304));
   OAI21_X1 i_0_340 (.A(n_0_305), .B1(n_0_306), .B2(n_0_312), .ZN(n_216));
   AOI22_X1 i_0_341 (.A1(n_275), .A2(n_0_218), .B1(n_227), .B2(n_0_217), 
      .ZN(n_0_305));
   INV_X1 i_0_342 (.A(n_288), .ZN(n_0_306));
   OAI21_X1 i_0_343 (.A(n_0_307), .B1(n_0_308), .B2(n_0_312), .ZN(n_217));
   AOI22_X1 i_0_344 (.A1(n_276), .A2(n_0_218), .B1(n_228), .B2(n_0_217), 
      .ZN(n_0_307));
   INV_X1 i_0_345 (.A(n_289), .ZN(n_0_308));
   OAI21_X1 i_0_346 (.A(n_0_309), .B1(n_0_313), .B2(n_0_312), .ZN(n_218));
   AOI22_X1 i_0_347 (.A1(n_277), .A2(n_0_218), .B1(n_137), .B2(n_0_217), 
      .ZN(n_0_309));
   INV_X1 i_0_348 (.A(n_0_310), .ZN(n_0_217));
   NAND2_X1 i_0_349 (.A1(n_0_312), .A2(n_0_311), .ZN(n_0_310));
   INV_X1 i_0_350 (.A(n_0_218), .ZN(n_0_311));
   NOR2_X1 i_0_351 (.A1(n_0_156), .A2(A[5]), .ZN(n_0_218));
   INV_X1 i_0_352 (.A(n_0_219), .ZN(n_0_312));
   NOR2_X1 i_0_353 (.A1(n_0_173), .A2(A[4]), .ZN(n_0_219));
   INV_X1 i_0_354 (.A(n_290), .ZN(n_0_313));
   OAI211_X1 i_0_355 (.A(n_0_314), .B(n_0_315), .C1(n_0_51), .C2(n_0_316), 
      .ZN(n_219));
   NAND2_X1 i_0_356 (.A1(n_82), .A2(n_0_2), .ZN(n_0_314));
   NAND2_X1 i_0_357 (.A1(n_98), .A2(n_0_3), .ZN(n_0_315));
   INV_X1 i_0_358 (.A(n_229), .ZN(n_0_316));
   NAND2_X1 i_0_359 (.A1(n_0_48), .A2(n_0_49), .ZN(n_220));
   OAI21_X1 i_0_362 (.A(n_0_317), .B1(n_0_318), .B2(n_0_332), .ZN(n_221));
   AOI22_X1 i_0_363 (.A1(n_84), .A2(n_0_2), .B1(n_0_1), .B2(n_230), .ZN(n_0_317));
   INV_X1 i_0_364 (.A(n_100), .ZN(n_0_318));
   OAI21_X1 i_0_365 (.A(n_0_319), .B1(n_0_320), .B2(n_0_332), .ZN(n_222));
   AOI22_X1 i_0_366 (.A1(n_85), .A2(n_0_2), .B1(n_0_1), .B2(n_231), .ZN(n_0_319));
   INV_X1 i_0_367 (.A(n_101), .ZN(n_0_320));
   OAI21_X1 i_0_368 (.A(n_0_321), .B1(n_0_322), .B2(n_0_332), .ZN(n_223));
   AOI22_X1 i_0_369 (.A1(n_86), .A2(n_0_2), .B1(n_0_1), .B2(n_232), .ZN(n_0_321));
   INV_X1 i_0_370 (.A(n_102), .ZN(n_0_322));
   OAI21_X1 i_0_371 (.A(n_0_323), .B1(n_0_324), .B2(n_0_332), .ZN(n_224));
   AOI22_X1 i_0_372 (.A1(n_87), .A2(n_0_2), .B1(n_0_1), .B2(n_233), .ZN(n_0_323));
   INV_X1 i_0_373 (.A(n_103), .ZN(n_0_324));
   OAI21_X1 i_0_374 (.A(n_0_325), .B1(n_0_326), .B2(n_0_332), .ZN(n_225));
   AOI22_X1 i_0_375 (.A1(n_88), .A2(n_0_2), .B1(n_234), .B2(n_0_1), .ZN(n_0_325));
   INV_X1 i_0_376 (.A(n_104), .ZN(n_0_326));
   OAI21_X1 i_0_377 (.A(n_0_327), .B1(n_0_328), .B2(n_0_332), .ZN(n_226));
   AOI22_X1 i_0_378 (.A1(n_89), .A2(n_0_2), .B1(n_235), .B2(n_0_1), .ZN(n_0_327));
   INV_X1 i_0_379 (.A(n_105), .ZN(n_0_328));
   OAI21_X1 i_0_380 (.A(n_0_329), .B1(n_0_330), .B2(n_0_332), .ZN(n_227));
   AOI22_X1 i_0_381 (.A1(n_92), .A2(n_0_2), .B1(n_237), .B2(n_0_1), .ZN(n_0_329));
   INV_X1 i_0_382 (.A(n_108), .ZN(n_0_330));
   OAI21_X1 i_0_383 (.A(n_0_331), .B1(n_0_333), .B2(n_0_332), .ZN(n_228));
   AOI22_X1 i_0_384 (.A1(n_93), .A2(n_0_2), .B1(n_238), .B2(n_0_1), .ZN(n_0_331));
   INV_X1 i_0_385 (.A(n_0_52), .ZN(n_0_2));
   INV_X1 i_0_386 (.A(n_0_51), .ZN(n_0_1));
   INV_X1 i_0_387 (.A(n_0_3), .ZN(n_0_332));
   NOR2_X1 i_0_388 (.A1(n_0_156), .A2(A[3]), .ZN(n_0_3));
   INV_X1 i_0_390 (.A(n_109), .ZN(n_0_333));
   NAND2_X1 i_0_391 (.A1(n_0_334), .A2(n_0_335), .ZN(n_229));
   AOI22_X1 i_0_393 (.A1(n_51), .A2(n_0_22), .B1(n_240), .B2(n_0_21), .ZN(
      n_0_334));
   NAND2_X1 i_0_394 (.A1(n_67), .A2(n_0_23), .ZN(n_0_335));
   OAI21_X1 i_0_395 (.A(n_0_336), .B1(n_0_337), .B2(n_0_346), .ZN(n_230));
   AOI22_X1 i_0_398 (.A1(n_69), .A2(n_0_23), .B1(n_241), .B2(n_0_21), .ZN(
      n_0_336));
   INV_X1 i_0_399 (.A(n_53), .ZN(n_0_337));
   OAI21_X1 i_0_400 (.A(n_0_338), .B1(n_0_339), .B2(n_0_347), .ZN(n_231));
   AOI22_X1 i_0_401 (.A1(n_54), .A2(n_0_22), .B1(n_242), .B2(n_0_21), .ZN(
      n_0_338));
   INV_X1 i_0_402 (.A(n_70), .ZN(n_0_339));
   NAND2_X1 i_0_403 (.A1(n_0_340), .A2(n_0_341), .ZN(n_232));
   AOI22_X1 i_0_404 (.A1(n_55), .A2(n_0_22), .B1(n_243), .B2(n_0_21), .ZN(
      n_0_340));
   NAND2_X1 i_0_405 (.A1(n_71), .A2(n_0_23), .ZN(n_0_341));
   OAI21_X1 i_0_406 (.A(n_0_342), .B1(n_0_343), .B2(n_0_346), .ZN(n_233));
   AOI22_X1 i_0_407 (.A1(n_72), .A2(n_0_23), .B1(n_244), .B2(n_0_21), .ZN(
      n_0_342));
   INV_X1 i_0_408 (.A(n_56), .ZN(n_0_343));
   INV_X1 i_0_409 (.A(n_0_13), .ZN(n_234));
   INV_X1 i_0_410 (.A(n_0_14), .ZN(n_235));
   OAI21_X1 i_0_411 (.A(n_0_344), .B1(n_0_348), .B2(n_0_347), .ZN(n_236));
   AOI22_X1 i_0_412 (.A1(n_60), .A2(n_0_22), .B1(n_246), .B2(n_0_21), .ZN(
      n_0_344));
   INV_X1 i_0_413 (.A(n_0_345), .ZN(n_0_21));
   NAND2_X1 i_0_414 (.A1(n_0_347), .A2(n_0_346), .ZN(n_0_345));
   INV_X1 i_0_415 (.A(n_0_22), .ZN(n_0_346));
   NOR2_X1 i_0_416 (.A1(A[3]), .A2(n_0_154), .ZN(n_0_22));
   INV_X1 i_0_418 (.A(n_0_23), .ZN(n_0_347));
   NOR2_X1 i_0_420 (.A1(n_0_155), .A2(A[2]), .ZN(n_0_23));
   INV_X1 i_0_421 (.A(n_76), .ZN(n_0_348));
   INV_X1 i_0_422 (.A(n_0_17), .ZN(n_237));
   INV_X1 i_0_423 (.A(n_0_18), .ZN(n_238));
   OAI21_X1 i_0_424 (.A(n_0_349), .B1(n_0_350), .B2(n_0_363), .ZN(n_239));
   AOI22_X1 i_0_429 (.A1(n_35), .A2(n_0_43), .B1(n_247), .B2(n_0_41), .ZN(
      n_0_349));
   INV_X1 i_0_430 (.A(n_19), .ZN(n_0_350));
   OAI21_X1 i_0_431 (.A(n_0_351), .B1(n_0_352), .B2(n_0_360), .ZN(n_240));
   AOI22_X1 i_0_436 (.A1(n_20), .A2(n_0_42), .B1(n_248), .B2(n_0_41), .ZN(
      n_0_351));
   INV_X1 i_0_437 (.A(n_36), .ZN(n_0_352));
   OAI21_X1 i_0_438 (.A(n_0_353), .B1(n_0_354), .B2(n_0_360), .ZN(n_241));
   AOI22_X1 i_0_439 (.A1(n_22), .A2(n_0_42), .B1(n_249), .B2(n_0_41), .ZN(
      n_0_353));
   INV_X1 i_0_440 (.A(n_38), .ZN(n_0_354));
   OAI21_X1 i_0_441 (.A(n_0_355), .B1(n_0_356), .B2(n_0_360), .ZN(n_242));
   AOI22_X1 i_0_442 (.A1(n_23), .A2(n_0_42), .B1(n_250), .B2(n_0_41), .ZN(
      n_0_355));
   INV_X1 i_0_443 (.A(n_39), .ZN(n_0_356));
   OAI21_X1 i_0_444 (.A(n_0_357), .B1(n_0_358), .B2(n_0_360), .ZN(n_243));
   AOI22_X1 i_0_445 (.A1(n_24), .A2(n_0_42), .B1(n_251), .B2(n_0_41), .ZN(
      n_0_357));
   INV_X1 i_0_446 (.A(n_40), .ZN(n_0_358));
   OAI21_X1 i_0_447 (.A(n_0_359), .B1(n_0_361), .B2(n_0_360), .ZN(n_244));
   AOI22_X1 i_0_448 (.A1(n_25), .A2(n_0_42), .B1(n_252), .B2(n_0_41), .ZN(
      n_0_359));
   INV_X1 i_0_449 (.A(n_0_43), .ZN(n_0_360));
   INV_X1 i_0_450 (.A(n_41), .ZN(n_0_361));
   OAI21_X1 i_0_452 (.A(n_0_362), .B1(n_0_364), .B2(n_0_363), .ZN(n_245));
   AOI22_X1 i_0_456 (.A1(n_44), .A2(n_0_43), .B1(n_254), .B2(n_0_41), .ZN(
      n_0_362));
   NOR2_X1 i_0_457 (.A1(n_0_43), .A2(n_0_42), .ZN(n_0_41));
   NOR2_X1 i_0_458 (.A1(n_0_154), .A2(A[1]), .ZN(n_0_43));
   INV_X1 i_0_460 (.A(n_0_42), .ZN(n_0_363));
   NOR2_X1 i_0_465 (.A1(A[2]), .A2(n_0_153), .ZN(n_0_42));
   INV_X1 i_0_466 (.A(n_28), .ZN(n_0_364));
   INV_X1 i_0_467 (.A(n_0_37), .ZN(n_246));
   OAI211_X1 i_0_472 (.A(n_0_366), .B(n_0_365), .C1(n_0_378), .C2(n_0_375), 
      .ZN(n_247));
   NAND2_X1 i_0_473 (.A1(n_0_68), .A2(n_256), .ZN(n_0_365));
   NAND2_X1 i_0_474 (.A1(n_4), .A2(n_0_70), .ZN(n_0_366));
   OAI211_X1 i_0_475 (.A(n_0_368), .B(n_0_367), .C1(n_0_102), .C2(n_0_380), 
      .ZN(n_248));
   NAND2_X1 i_0_476 (.A1(n_0_59), .A2(n_256), .ZN(n_0_367));
   NAND2_X1 i_0_477 (.A1(n_5), .A2(n_0_70), .ZN(n_0_368));
   OAI221_X1 i_0_478 (.A(n_0_369), .B1(n_0_102), .B2(n_0_371), .C1(n_0_382), 
      .C2(n_0_375), .ZN(n_249));
   NAND2_X1 i_0_479 (.A1(n_7), .A2(n_0_70), .ZN(n_0_369));
   OAI221_X1 i_0_480 (.A(n_0_370), .B1(n_0_102), .B2(n_0_385), .C1(n_0_371), 
      .C2(n_0_375), .ZN(n_250));
   NAND2_X1 i_0_481 (.A1(n_8), .A2(n_0_70), .ZN(n_0_370));
   INV_X1 i_0_482 (.A(n_259), .ZN(n_0_371));
   OAI221_X1 i_0_483 (.A(n_0_372), .B1(n_0_102), .B2(n_0_387), .C1(n_0_385), 
      .C2(n_0_375), .ZN(n_251));
   NAND2_X1 i_0_484 (.A1(n_9), .A2(n_0_70), .ZN(n_0_372));
   OAI211_X1 i_0_485 (.A(n_0_374), .B(n_0_373), .C1(n_0_387), .C2(n_0_375), 
      .ZN(n_252));
   NAND2_X1 i_0_486 (.A1(n_0_68), .A2(n_262), .ZN(n_0_373));
   NAND2_X1 i_0_487 (.A1(n_10), .A2(n_0_70), .ZN(n_0_374));
   INV_X1 i_0_492 (.A(n_0_59), .ZN(n_0_375));
   NAND2_X1 i_0_493 (.A1(n_0_377), .A2(n_0_376), .ZN(n_253));
   AOI22_X1 i_0_494 (.A1(n_264), .A2(n_0_68), .B1(n_263), .B2(n_0_59), .ZN(
      n_0_376));
   NOR2_X1 i_0_501 (.A1(n_0_153), .A2(A[0]), .ZN(n_0_59));
   INV_X1 i_0_502 (.A(n_0_102), .ZN(n_0_68));
   NAND2_X1 i_0_503 (.A1(n_12), .A2(n_0_70), .ZN(n_0_377));
   NOR2_X1 i_0_506 (.A1(A[1]), .A2(n_0_104), .ZN(n_0_70));
   INV_X1 i_0_507 (.A(n_0_57), .ZN(n_254));
   INV_X1 i_0_508 (.A(n_0_378), .ZN(n_255));
   NAND2_X1 i_0_509 (.A1(n_0_403), .A2(n_0_379), .ZN(n_0_378));
   NAND2_X1 i_0_510 (.A1(n_0_404), .A2(B[4]), .ZN(n_0_379));
   XNOR2_X1 i_0_511 (.A(n_0_403), .B(n_0_410), .ZN(n_256));
   INV_X1 i_0_512 (.A(n_0_380), .ZN(n_257));
   NAND2_X1 i_0_513 (.A1(n_0_399), .A2(n_0_381), .ZN(n_0_380));
   NAND2_X1 i_0_514 (.A1(n_0_401), .A2(B[6]), .ZN(n_0_381));
   INV_X1 i_0_515 (.A(n_0_382), .ZN(n_258));
   NAND2_X1 i_0_516 (.A1(n_0_397), .A2(n_0_383), .ZN(n_0_382));
   NAND2_X1 i_0_518 (.A1(n_0_399), .A2(B[7]), .ZN(n_0_383));
   AND2_X1 i_0_519 (.A1(n_0_395), .A2(n_0_384), .ZN(n_259));
   NAND2_X1 i_0_520 (.A1(n_0_397), .A2(B[8]), .ZN(n_0_384));
   INV_X1 i_0_521 (.A(n_0_385), .ZN(n_260));
   NAND2_X1 i_0_522 (.A1(n_0_393), .A2(n_0_386), .ZN(n_0_385));
   NAND2_X1 i_0_523 (.A1(n_0_395), .A2(B[9]), .ZN(n_0_386));
   INV_X1 i_0_524 (.A(n_0_387), .ZN(n_261));
   NAND2_X1 i_0_525 (.A1(n_0_389), .A2(n_0_388), .ZN(n_0_387));
   NAND2_X1 i_0_528 (.A1(n_0_393), .A2(B[10]), .ZN(n_0_388));
   XNOR2_X1 i_0_529 (.A(n_0_389), .B(n_0_416), .ZN(n_262));
   NAND2_X1 i_0_530 (.A1(n_0_392), .A2(n_0_415), .ZN(n_0_389));
   INV_X1 i_0_534 (.A(n_0_390), .ZN(n_263));
   XNOR2_X1 i_0_535 (.A(n_0_391), .B(B[15]), .ZN(n_0_390));
   NAND3_X1 i_0_538 (.A1(n_0_392), .A2(n_0_416), .A3(n_0_415), .ZN(n_0_391));
   INV_X1 i_0_541 (.A(n_0_393), .ZN(n_0_392));
   NAND2_X1 i_0_542 (.A1(n_0_394), .A2(n_0_414), .ZN(n_0_393));
   INV_X1 i_0_543 (.A(n_0_395), .ZN(n_0_394));
   NAND2_X1 i_0_544 (.A1(n_0_396), .A2(n_0_413), .ZN(n_0_395));
   INV_X1 i_0_545 (.A(n_0_397), .ZN(n_0_396));
   NAND2_X1 i_0_546 (.A1(n_0_398), .A2(n_0_412), .ZN(n_0_397));
   INV_X1 i_0_547 (.A(n_0_399), .ZN(n_0_398));
   NAND2_X1 i_0_548 (.A1(n_0_400), .A2(n_0_411), .ZN(n_0_399));
   INV_X1 i_0_549 (.A(n_0_401), .ZN(n_0_400));
   NAND2_X1 i_0_550 (.A1(n_0_402), .A2(n_0_410), .ZN(n_0_401));
   INV_X1 i_0_551 (.A(n_0_403), .ZN(n_0_402));
   NAND2_X1 i_0_552 (.A1(n_0_132), .A2(n_0_409), .ZN(n_0_403));
   INV_X1 i_0_553 (.A(n_0_404), .ZN(n_0_132));
   NAND2_X1 i_0_560 (.A1(n_0_134), .A2(n_0_408), .ZN(n_0_404));
   INV_X1 i_0_561 (.A(n_0_133), .ZN(n_0_134));
   NAND2_X1 i_0_562 (.A1(n_0_136), .A2(n_0_407), .ZN(n_0_133));
   INV_X1 i_0_563 (.A(n_0_135), .ZN(n_0_136));
   NAND2_X1 i_0_564 (.A1(n_0_406), .A2(n_0_405), .ZN(n_0_135));
   INV_X1 i_0_565 (.A(B[0]), .ZN(n_0_405));
   INV_X1 i_0_566 (.A(B[1]), .ZN(n_0_406));
   INV_X1 i_0_567 (.A(B[2]), .ZN(n_0_407));
   INV_X1 i_0_568 (.A(B[3]), .ZN(n_0_408));
   INV_X1 i_0_569 (.A(B[4]), .ZN(n_0_409));
   INV_X1 i_0_570 (.A(B[5]), .ZN(n_0_410));
   INV_X1 i_0_571 (.A(B[6]), .ZN(n_0_411));
   INV_X1 i_0_572 (.A(B[7]), .ZN(n_0_412));
   INV_X1 i_0_573 (.A(B[8]), .ZN(n_0_413));
   INV_X1 i_0_574 (.A(B[9]), .ZN(n_0_414));
   INV_X1 i_0_575 (.A(B[10]), .ZN(n_0_415));
   INV_X1 i_0_576 (.A(B[11]), .ZN(n_0_416));
   AOI21_X1 i_0_577 (.A(n_0_73), .B1(B[15]), .B2(n_0_74), .ZN(n_264));
   FA_X1 i_1_0 (.A(B[1]), .B(n_219), .CI(n_1_166), .CO(n_1_2), .S(n_265));
   FA_X1 i_1_1 (.A(B[2]), .B(n_220), .CI(n_1_2), .CO(n_1_3), .S(n_266));
   FA_X1 i_1_2 (.A(B[3]), .B(n_221), .CI(n_1_3), .CO(n_1_4), .S(n_267));
   FA_X1 i_1_3 (.A(B[4]), .B(n_222), .CI(n_1_4), .CO(n_1_5), .S(n_268));
   FA_X1 i_1_4 (.A(B[5]), .B(n_223), .CI(n_1_5), .CO(n_1_6), .S(n_269));
   FA_X1 i_1_5 (.A(B[6]), .B(n_224), .CI(n_1_6), .CO(n_1_7), .S(n_270));
   FA_X1 i_1_6 (.A(B[7]), .B(n_225), .CI(n_1_7), .CO(n_1_8), .S(n_271));
   FA_X1 i_1_7 (.A(B[8]), .B(n_226), .CI(n_1_8), .CO(n_1_9), .S(n_272));
   FA_X1 i_1_8 (.A(B[9]), .B(n_135), .CI(n_1_9), .CO(n_1_10), .S(n_273));
   FA_X1 i_1_9 (.A(B[10]), .B(n_136), .CI(n_1_10), .CO(n_1_11), .S(n_274));
   FA_X1 i_1_10 (.A(B[11]), .B(n_227), .CI(n_1_11), .CO(n_1_12), .S(n_275));
   FA_X1 i_1_11 (.A(B[15]), .B(n_228), .CI(n_1_12), .CO(n_1_13), .S(n_276));
   FA_X1 i_1_12 (.A(B[15]), .B(n_137), .CI(n_1_13), .CO(n_1_14), .S(n_277));
   FA_X1 i_1_13 (.A(n_146), .B(n_219), .CI(n_1_166), .CO(n_1_0), .S(n_278));
   FA_X1 i_1_14 (.A(n_147), .B(n_220), .CI(n_1_0), .CO(n_1_1), .S(n_279));
   FA_X1 i_1_15 (.A(n_148), .B(n_221), .CI(n_1_1), .CO(n_1_15), .S(n_280));
   FA_X1 i_1_16 (.A(n_255), .B(n_222), .CI(n_1_15), .CO(n_1_16), .S(n_281));
   FA_X1 i_1_17 (.A(n_256), .B(n_223), .CI(n_1_16), .CO(n_1_17), .S(n_282));
   FA_X1 i_1_18 (.A(n_257), .B(n_224), .CI(n_1_17), .CO(n_1_18), .S(n_283));
   FA_X1 i_1_19 (.A(n_258), .B(n_225), .CI(n_1_18), .CO(n_1_19), .S(n_284));
   FA_X1 i_1_20 (.A(n_259), .B(n_226), .CI(n_1_19), .CO(n_1_20), .S(n_285));
   FA_X1 i_1_21 (.A(n_260), .B(n_135), .CI(n_1_20), .CO(n_1_21), .S(n_286));
   FA_X1 i_1_22 (.A(n_261), .B(n_136), .CI(n_1_21), .CO(n_1_22), .S(n_287));
   FA_X1 i_1_23 (.A(n_262), .B(n_227), .CI(n_1_22), .CO(n_1_23), .S(n_288));
   FA_X1 i_1_24 (.A(n_263), .B(n_228), .CI(n_1_23), .CO(n_1_24), .S(n_289));
   FA_X1 i_1_25 (.A(n_264), .B(n_137), .CI(n_1_24), .CO(n_1_25), .S(n_290));
   FA_X1 i_1_26 (.A(B[1]), .B(n_207), .CI(n_1_167), .CO(n_1_26), .S(n_291));
   FA_X1 i_1_27 (.A(B[2]), .B(n_208), .CI(n_1_26), .CO(n_1_27), .S(n_292));
   FA_X1 i_1_28 (.A(B[3]), .B(n_209), .CI(n_1_27), .CO(n_1_28), .S(n_293));
   FA_X1 i_1_29 (.A(B[4]), .B(n_210), .CI(n_1_28), .CO(n_1_29), .S(n_294));
   FA_X1 i_1_30 (.A(B[5]), .B(n_211), .CI(n_1_29), .CO(n_1_30), .S(n_295));
   FA_X1 i_1_31 (.A(B[6]), .B(n_212), .CI(n_1_30), .CO(n_1_31), .S(n_296));
   FA_X1 i_1_32 (.A(B[7]), .B(n_213), .CI(n_1_31), .CO(n_1_32), .S(n_297));
   FA_X1 i_1_33 (.A(B[8]), .B(n_214), .CI(n_1_32), .CO(n_1_33), .S(n_298));
   FA_X1 i_1_34 (.A(B[9]), .B(n_215), .CI(n_1_33), .CO(n_1_34), .S(n_299));
   FA_X1 i_1_35 (.A(B[10]), .B(n_216), .CI(n_1_34), .CO(n_1_35), .S(n_300));
   FA_X1 i_1_36 (.A(B[11]), .B(n_217), .CI(n_1_35), .CO(n_1_36), .S(n_301));
   FA_X1 i_1_37 (.A(B[15]), .B(n_218), .CI(n_1_36), .CO(n_1_37), .S(n_302));
   FA_X1 i_1_38 (.A(B[15]), .B(n_133), .CI(n_1_37), .CO(n_1_38), .S(n_303));
   FA_X1 i_1_39 (.A(n_146), .B(n_207), .CI(n_1_167), .CO(n_1_39), .S(n_304));
   FA_X1 i_1_40 (.A(n_147), .B(n_208), .CI(n_1_39), .CO(n_1_40), .S(n_305));
   FA_X1 i_1_41 (.A(n_148), .B(n_209), .CI(n_1_40), .CO(n_1_41), .S(n_306));
   FA_X1 i_1_42 (.A(n_255), .B(n_210), .CI(n_1_41), .CO(n_1_42), .S(n_307));
   FA_X1 i_1_43 (.A(n_256), .B(n_211), .CI(n_1_42), .CO(n_1_43), .S(n_308));
   FA_X1 i_1_44 (.A(n_257), .B(n_212), .CI(n_1_43), .CO(n_1_44), .S(n_309));
   FA_X1 i_1_45 (.A(n_258), .B(n_213), .CI(n_1_44), .CO(n_1_45), .S(n_310));
   FA_X1 i_1_46 (.A(n_259), .B(n_214), .CI(n_1_45), .CO(n_1_46), .S(n_311));
   FA_X1 i_1_47 (.A(n_260), .B(n_215), .CI(n_1_46), .CO(n_1_47), .S(n_312));
   FA_X1 i_1_48 (.A(n_261), .B(n_216), .CI(n_1_47), .CO(n_1_48), .S(n_313));
   FA_X1 i_1_49 (.A(n_262), .B(n_217), .CI(n_1_48), .CO(n_1_49), .S(n_314));
   FA_X1 i_1_50 (.A(n_263), .B(n_218), .CI(n_1_49), .CO(n_1_50), .S(n_315));
   FA_X1 i_1_51 (.A(n_264), .B(n_133), .CI(n_1_50), .CO(n_1_51), .S(n_316));
   FA_X1 i_1_52 (.A(B[1]), .B(n_195), .CI(n_1_168), .CO(n_1_52), .S(n_317));
   FA_X1 i_1_53 (.A(B[2]), .B(n_196), .CI(n_1_52), .CO(n_1_53), .S(n_318));
   FA_X1 i_1_54 (.A(B[3]), .B(n_197), .CI(n_1_53), .CO(n_1_54), .S(n_319));
   FA_X1 i_1_55 (.A(B[4]), .B(n_198), .CI(n_1_54), .CO(n_1_55), .S(n_320));
   FA_X1 i_1_56 (.A(B[5]), .B(n_199), .CI(n_1_55), .CO(n_1_56), .S(n_321));
   FA_X1 i_1_57 (.A(B[6]), .B(n_200), .CI(n_1_56), .CO(n_1_57), .S(n_322));
   FA_X1 i_1_58 (.A(B[7]), .B(n_201), .CI(n_1_57), .CO(n_1_58), .S(n_323));
   FA_X1 i_1_59 (.A(B[8]), .B(n_202), .CI(n_1_58), .CO(n_1_59), .S(n_324));
   FA_X1 i_1_60 (.A(B[9]), .B(n_203), .CI(n_1_59), .CO(n_1_60), .S(n_325));
   FA_X1 i_1_61 (.A(B[10]), .B(n_204), .CI(n_1_60), .CO(n_1_61), .S(n_326));
   FA_X1 i_1_62 (.A(B[11]), .B(n_205), .CI(n_1_61), .CO(n_1_62), .S(n_327));
   FA_X1 i_1_63 (.A(B[15]), .B(n_132), .CI(n_1_62), .CO(n_1_63), .S(n_328));
   FA_X1 i_1_64 (.A(n_146), .B(n_195), .CI(n_1_168), .CO(n_1_64), .S(n_329));
   FA_X1 i_1_65 (.A(n_147), .B(n_196), .CI(n_1_64), .CO(n_1_65), .S(n_330));
   FA_X1 i_1_66 (.A(n_148), .B(n_197), .CI(n_1_65), .CO(n_1_66), .S(n_331));
   FA_X1 i_1_67 (.A(n_255), .B(n_198), .CI(n_1_66), .CO(n_1_67), .S(n_332));
   FA_X1 i_1_68 (.A(n_256), .B(n_199), .CI(n_1_67), .CO(n_1_68), .S(n_333));
   FA_X1 i_1_69 (.A(n_257), .B(n_200), .CI(n_1_68), .CO(n_1_69), .S(n_334));
   FA_X1 i_1_70 (.A(n_258), .B(n_201), .CI(n_1_69), .CO(n_1_70), .S(n_335));
   FA_X1 i_1_71 (.A(n_259), .B(n_202), .CI(n_1_70), .CO(n_1_71), .S(n_336));
   FA_X1 i_1_72 (.A(n_260), .B(n_203), .CI(n_1_71), .CO(n_1_72), .S(n_337));
   FA_X1 i_1_73 (.A(n_261), .B(n_204), .CI(n_1_72), .CO(n_1_73), .S(n_338));
   FA_X1 i_1_74 (.A(n_262), .B(n_205), .CI(n_1_73), .CO(n_1_74), .S(n_339));
   FA_X1 i_1_75 (.A(n_263), .B(n_132), .CI(n_1_74), .CO(n_1_75), .S(n_340));
   FA_X1 i_1_76 (.A(B[1]), .B(n_184), .CI(n_1_169), .CO(n_1_76), .S(n_341));
   FA_X1 i_1_77 (.A(B[2]), .B(n_185), .CI(n_1_76), .CO(n_1_77), .S(n_342));
   FA_X1 i_1_78 (.A(B[3]), .B(n_186), .CI(n_1_77), .CO(n_1_78), .S(n_343));
   FA_X1 i_1_79 (.A(B[4]), .B(n_187), .CI(n_1_78), .CO(n_1_79), .S(n_344));
   FA_X1 i_1_80 (.A(B[5]), .B(n_188), .CI(n_1_79), .CO(n_1_80), .S(n_345));
   FA_X1 i_1_81 (.A(B[6]), .B(n_189), .CI(n_1_80), .CO(n_1_81), .S(n_346));
   FA_X1 i_1_82 (.A(B[7]), .B(n_190), .CI(n_1_81), .CO(n_1_82), .S(n_347));
   FA_X1 i_1_83 (.A(B[8]), .B(n_191), .CI(n_1_82), .CO(n_1_83), .S(n_348));
   FA_X1 i_1_84 (.A(B[9]), .B(n_192), .CI(n_1_83), .CO(n_1_84), .S(n_349));
   FA_X1 i_1_85 (.A(B[10]), .B(n_193), .CI(n_1_84), .CO(n_1_85), .S(n_350));
   FA_X1 i_1_86 (.A(B[11]), .B(n_131), .CI(n_1_85), .CO(n_1_86), .S(n_351));
   FA_X1 i_1_87 (.A(n_146), .B(n_184), .CI(n_1_169), .CO(n_1_87), .S(n_352));
   FA_X1 i_1_88 (.A(n_147), .B(n_185), .CI(n_1_87), .CO(n_1_88), .S(n_353));
   FA_X1 i_1_89 (.A(n_148), .B(n_186), .CI(n_1_88), .CO(n_1_89), .S(n_354));
   FA_X1 i_1_90 (.A(n_255), .B(n_187), .CI(n_1_89), .CO(n_1_90), .S(n_355));
   FA_X1 i_1_91 (.A(n_256), .B(n_188), .CI(n_1_90), .CO(n_1_91), .S(n_356));
   FA_X1 i_1_92 (.A(n_257), .B(n_189), .CI(n_1_91), .CO(n_1_92), .S(n_357));
   FA_X1 i_1_93 (.A(n_258), .B(n_190), .CI(n_1_92), .CO(n_1_93), .S(n_358));
   FA_X1 i_1_94 (.A(n_259), .B(n_191), .CI(n_1_93), .CO(n_1_94), .S(n_359));
   FA_X1 i_1_95 (.A(n_260), .B(n_192), .CI(n_1_94), .CO(n_1_95), .S(n_360));
   FA_X1 i_1_96 (.A(n_261), .B(n_193), .CI(n_1_95), .CO(n_1_96), .S(n_361));
   FA_X1 i_1_97 (.A(n_262), .B(n_131), .CI(n_1_96), .CO(n_1_97), .S(n_362));
   FA_X1 i_1_98 (.A(B[1]), .B(n_174), .CI(n_1_170), .CO(n_1_98), .S(n_363));
   FA_X1 i_1_99 (.A(B[2]), .B(n_175), .CI(n_1_98), .CO(n_1_99), .S(n_364));
   FA_X1 i_1_100 (.A(B[3]), .B(n_176), .CI(n_1_99), .CO(n_1_100), .S(n_365));
   FA_X1 i_1_101 (.A(B[4]), .B(n_177), .CI(n_1_100), .CO(n_1_101), .S(n_366));
   FA_X1 i_1_102 (.A(B[5]), .B(n_178), .CI(n_1_101), .CO(n_1_102), .S(n_367));
   FA_X1 i_1_103 (.A(B[6]), .B(n_179), .CI(n_1_102), .CO(n_1_103), .S(n_368));
   FA_X1 i_1_104 (.A(B[7]), .B(n_180), .CI(n_1_103), .CO(n_1_104), .S(n_369));
   FA_X1 i_1_105 (.A(B[8]), .B(n_181), .CI(n_1_104), .CO(n_1_105), .S(n_370));
   FA_X1 i_1_106 (.A(B[9]), .B(n_182), .CI(n_1_105), .CO(n_1_106), .S(n_371));
   FA_X1 i_1_107 (.A(B[10]), .B(n_130), .CI(n_1_106), .CO(n_1_107), .S(n_372));
   FA_X1 i_1_108 (.A(n_146), .B(n_174), .CI(n_1_170), .CO(n_1_108), .S(n_373));
   FA_X1 i_1_109 (.A(n_147), .B(n_175), .CI(n_1_108), .CO(n_1_109), .S(n_374));
   FA_X1 i_1_110 (.A(n_148), .B(n_176), .CI(n_1_109), .CO(n_1_110), .S(n_375));
   FA_X1 i_1_111 (.A(n_255), .B(n_177), .CI(n_1_110), .CO(n_1_111), .S(n_376));
   FA_X1 i_1_112 (.A(n_256), .B(n_178), .CI(n_1_111), .CO(n_1_112), .S(n_377));
   FA_X1 i_1_113 (.A(n_257), .B(n_179), .CI(n_1_112), .CO(n_1_113), .S(n_378));
   FA_X1 i_1_114 (.A(n_258), .B(n_180), .CI(n_1_113), .CO(n_1_114), .S(n_379));
   FA_X1 i_1_115 (.A(n_259), .B(n_181), .CI(n_1_114), .CO(n_1_115), .S(n_380));
   FA_X1 i_1_116 (.A(n_260), .B(n_182), .CI(n_1_115), .CO(n_1_116), .S(n_381));
   FA_X1 i_1_117 (.A(n_261), .B(n_130), .CI(n_1_116), .CO(n_1_117), .S(n_382));
   FA_X1 i_1_118 (.A(B[1]), .B(n_165), .CI(n_1_171), .CO(n_1_118), .S(n_383));
   FA_X1 i_1_119 (.A(B[2]), .B(n_166), .CI(n_1_118), .CO(n_1_119), .S(n_384));
   FA_X1 i_1_120 (.A(B[3]), .B(n_167), .CI(n_1_119), .CO(n_1_120), .S(n_385));
   FA_X1 i_1_121 (.A(B[4]), .B(n_168), .CI(n_1_120), .CO(n_1_121), .S(n_386));
   FA_X1 i_1_122 (.A(B[5]), .B(n_169), .CI(n_1_121), .CO(n_1_122), .S(n_387));
   FA_X1 i_1_123 (.A(B[6]), .B(n_170), .CI(n_1_122), .CO(n_1_123), .S(n_388));
   FA_X1 i_1_124 (.A(B[7]), .B(n_171), .CI(n_1_123), .CO(n_1_124), .S(n_389));
   FA_X1 i_1_125 (.A(B[8]), .B(n_172), .CI(n_1_124), .CO(n_1_125), .S(n_390));
   FA_X1 i_1_126 (.A(B[9]), .B(n_129), .CI(n_1_125), .CO(n_1_126), .S(n_391));
   FA_X1 i_1_127 (.A(n_146), .B(n_165), .CI(n_1_171), .CO(n_1_127), .S(n_392));
   FA_X1 i_1_128 (.A(n_147), .B(n_166), .CI(n_1_127), .CO(n_1_128), .S(n_393));
   FA_X1 i_1_129 (.A(n_148), .B(n_167), .CI(n_1_128), .CO(n_1_129), .S(n_394));
   FA_X1 i_1_130 (.A(n_255), .B(n_168), .CI(n_1_129), .CO(n_1_130), .S(n_395));
   FA_X1 i_1_131 (.A(n_256), .B(n_169), .CI(n_1_130), .CO(n_1_131), .S(n_396));
   FA_X1 i_1_132 (.A(n_257), .B(n_170), .CI(n_1_131), .CO(n_1_132), .S(n_397));
   FA_X1 i_1_133 (.A(n_258), .B(n_171), .CI(n_1_132), .CO(n_1_133), .S(n_398));
   FA_X1 i_1_134 (.A(n_259), .B(n_172), .CI(n_1_133), .CO(n_1_134), .S(n_399));
   FA_X1 i_1_135 (.A(n_260), .B(n_129), .CI(n_1_134), .CO(n_1_135), .S(n_400));
   FA_X1 i_1_136 (.A(B[1]), .B(n_157), .CI(n_1_172), .CO(n_1_136), .S(n_401));
   FA_X1 i_1_137 (.A(B[2]), .B(n_158), .CI(n_1_136), .CO(n_1_137), .S(n_402));
   FA_X1 i_1_138 (.A(B[3]), .B(n_159), .CI(n_1_137), .CO(n_1_138), .S(n_403));
   FA_X1 i_1_139 (.A(B[4]), .B(n_160), .CI(n_1_138), .CO(n_1_139), .S(n_404));
   FA_X1 i_1_140 (.A(B[5]), .B(n_161), .CI(n_1_139), .CO(n_1_140), .S(n_405));
   FA_X1 i_1_141 (.A(B[6]), .B(n_162), .CI(n_1_140), .CO(n_1_141), .S(n_406));
   FA_X1 i_1_142 (.A(B[7]), .B(n_163), .CI(n_1_141), .CO(n_1_142), .S(n_407));
   FA_X1 i_1_143 (.A(B[8]), .B(n_128), .CI(n_1_142), .CO(n_1_143), .S(n_408));
   FA_X1 i_1_144 (.A(n_146), .B(n_157), .CI(n_1_172), .CO(n_1_144), .S(n_409));
   FA_X1 i_1_145 (.A(n_147), .B(n_158), .CI(n_1_144), .CO(n_1_145), .S(n_410));
   FA_X1 i_1_146 (.A(n_148), .B(n_159), .CI(n_1_145), .CO(n_1_146), .S(n_411));
   FA_X1 i_1_147 (.A(n_255), .B(n_160), .CI(n_1_146), .CO(n_1_147), .S(n_412));
   FA_X1 i_1_148 (.A(n_256), .B(n_161), .CI(n_1_147), .CO(n_1_148), .S(n_413));
   FA_X1 i_1_149 (.A(n_257), .B(n_162), .CI(n_1_148), .CO(n_1_149), .S(n_414));
   FA_X1 i_1_150 (.A(n_258), .B(n_163), .CI(n_1_149), .CO(n_1_150), .S(n_415));
   FA_X1 i_1_151 (.A(n_259), .B(n_128), .CI(n_1_150), .CO(n_1_151), .S(n_416));
   FA_X1 i_1_152 (.A(B[1]), .B(n_150), .CI(n_1_173), .CO(n_1_152), .S(n_417));
   FA_X1 i_1_153 (.A(B[2]), .B(n_151), .CI(n_1_152), .CO(n_1_153), .S(n_418));
   FA_X1 i_1_154 (.A(B[3]), .B(n_152), .CI(n_1_153), .CO(n_1_154), .S(n_419));
   FA_X1 i_1_155 (.A(B[4]), .B(n_153), .CI(n_1_154), .CO(n_1_155), .S(n_420));
   FA_X1 i_1_156 (.A(B[5]), .B(n_154), .CI(n_1_155), .CO(n_1_156), .S(n_421));
   FA_X1 i_1_157 (.A(B[6]), .B(n_155), .CI(n_1_156), .CO(n_1_157), .S(n_422));
   FA_X1 i_1_158 (.A(B[7]), .B(n_127), .CI(n_1_157), .CO(n_1_158), .S(n_423));
   FA_X1 i_1_159 (.A(n_146), .B(n_150), .CI(n_1_173), .CO(n_1_159), .S(n_424));
   FA_X1 i_1_160 (.A(n_147), .B(n_151), .CI(n_1_159), .CO(n_1_160), .S(n_425));
   FA_X1 i_1_161 (.A(n_148), .B(n_152), .CI(n_1_160), .CO(n_1_161), .S(n_426));
   FA_X1 i_1_162 (.A(n_255), .B(n_153), .CI(n_1_161), .CO(n_1_162), .S(n_427));
   FA_X1 i_1_163 (.A(n_256), .B(n_154), .CI(n_1_162), .CO(n_1_163), .S(n_428));
   FA_X1 i_1_164 (.A(n_257), .B(n_155), .CI(n_1_163), .CO(n_1_164), .S(n_429));
   FA_X1 i_1_165 (.A(n_258), .B(n_127), .CI(n_1_164), .CO(n_1_165), .S(n_430));
   HA_X1 i_1_166 (.A(B[0]), .B(n_134), .CO(n_1_166), .S(n_431));
   HA_X1 i_1_167 (.A(B[0]), .B(n_206), .CO(n_1_167), .S(n_432));
   HA_X1 i_1_168 (.A(B[0]), .B(n_194), .CO(n_1_168), .S(n_433));
   HA_X1 i_1_169 (.A(B[0]), .B(n_183), .CO(n_1_169), .S(n_434));
   HA_X1 i_1_170 (.A(B[0]), .B(n_173), .CO(n_1_170), .S(n_435));
   HA_X1 i_1_171 (.A(B[0]), .B(n_164), .CO(n_1_171), .S(n_436));
   HA_X1 i_1_172 (.A(B[0]), .B(n_156), .CO(n_1_172), .S(n_437));
   HA_X1 i_1_173 (.A(B[0]), .B(n_149), .CO(n_1_173), .S(n_438));
   XNOR2_X1 i_1_174 (.A(n_112), .B(n_1_174), .ZN(n_439));
   XNOR2_X1 i_1_175 (.A(n_125), .B(n_1_25), .ZN(n_1_174));
   INV_X1 i_1_176 (.A(n_1_14), .ZN(n_1_175));
   XNOR2_X1 i_1_177 (.A(n_112), .B(B[15]), .ZN(n_1_176));
   INV_X1 i_1_178 (.A(n_1_176), .ZN(n_1_177));
   AOI22_X1 i_1_179 (.A1(n_1_175), .A2(n_1_176), .B1(n_1_14), .B2(n_1_177), 
      .ZN(n_440));
endmodule

module multiplier_16bit__0_1434(first_operand, second_operand, out, enable, 
      overflow);
   input [15:0]first_operand;
   input [15:0]second_operand;
   output [15:0]out;
   input enable;
   output overflow;

   wire [31:0]temp_result_wire;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_9;
   wire n_0_0_39;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_29;
   wire n_0_0_18;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_30;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_28;

   booth_16bit_multiplier__1 mult (.A({first_operand[12], uc_0, uc_1, uc_2, 
      first_operand[11], first_operand[10], first_operand[9], first_operand[8], 
      first_operand[7], first_operand[6], first_operand[5], first_operand[4], 
      first_operand[3], first_operand[2], first_operand[1], first_operand[0]}), 
      .B({second_operand[12], uc_3, uc_4, uc_5, second_operand[11], 
      second_operand[10], second_operand[9], second_operand[8], 
      second_operand[7], second_operand[6], second_operand[5], second_operand[4], 
      second_operand[3], second_operand[2], second_operand[1], second_operand[0]}), 
      .product({uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, 
      uc_16, uc_17, temp_result_wire[19], temp_result_wire[18], 
      temp_result_wire[17], temp_result_wire[16], temp_result_wire[15], 
      temp_result_wire[14], temp_result_wire[13], temp_result_wire[12], 
      temp_result_wire[11], temp_result_wire[10], temp_result_wire[9], 
      temp_result_wire[8], temp_result_wire[7], temp_result_wire[6], 
      temp_result_wire[5], temp_result_wire[4], temp_result_wire[3], 
      temp_result_wire[2], temp_result_wire[1], temp_result_wire[0]}));
   MUX2_X1 i_0_0_0 (.A(temp_result_wire[0]), .B(temp_result_wire[4]), .S(
      n_0_0_30), .Z(n_0_0_0));
   MUX2_X1 i_0_0_1 (.A(temp_result_wire[1]), .B(temp_result_wire[5]), .S(
      n_0_0_30), .Z(n_0_0_1));
   MUX2_X1 i_0_0_2 (.A(temp_result_wire[2]), .B(temp_result_wire[6]), .S(
      n_0_0_30), .Z(n_0_0_2));
   MUX2_X1 i_0_0_3 (.A(temp_result_wire[3]), .B(temp_result_wire[7]), .S(
      n_0_0_30), .Z(n_0_0_3));
   MUX2_X1 i_0_0_4 (.A(temp_result_wire[4]), .B(temp_result_wire[8]), .S(
      n_0_0_30), .Z(n_0_0_4));
   MUX2_X1 i_0_0_5 (.A(temp_result_wire[5]), .B(temp_result_wire[9]), .S(
      n_0_0_30), .Z(n_0_0_5));
   MUX2_X1 i_0_0_6 (.A(temp_result_wire[6]), .B(temp_result_wire[10]), .S(
      n_0_0_30), .Z(n_0_0_6));
   MUX2_X1 i_0_0_7 (.A(temp_result_wire[7]), .B(temp_result_wire[11]), .S(
      n_0_0_30), .Z(n_0_0_7));
   MUX2_X1 i_0_0_8 (.A(temp_result_wire[8]), .B(temp_result_wire[12]), .S(
      n_0_0_30), .Z(n_0_0_8));
   MUX2_X1 i_0_0_16 (.A(n_0_0_0), .B(n_0_0_2), .S(n_0_0_29), .Z(n_0_0_31));
   MUX2_X1 i_0_0_17 (.A(n_0_0_1), .B(n_0_0_3), .S(n_0_0_29), .Z(n_0_0_32));
   MUX2_X1 i_0_0_18 (.A(n_0_0_2), .B(n_0_0_4), .S(n_0_0_29), .Z(n_0_0_33));
   MUX2_X1 i_0_0_19 (.A(n_0_0_3), .B(n_0_0_5), .S(n_0_0_29), .Z(n_0_0_34));
   MUX2_X1 i_0_0_20 (.A(n_0_0_4), .B(n_0_0_6), .S(n_0_0_29), .Z(n_0_0_35));
   MUX2_X1 i_0_0_21 (.A(n_0_0_5), .B(n_0_0_7), .S(n_0_0_29), .Z(n_0_0_36));
   MUX2_X1 i_0_0_22 (.A(n_0_0_6), .B(n_0_0_8), .S(n_0_0_29), .Z(n_0_0_37));
   MUX2_X1 i_0_0_23 (.A(n_0_0_7), .B(n_0_0_9), .S(n_0_0_29), .Z(n_0_0_38));
   MUX2_X1 i_0_0_30 (.A(n_0_0_31), .B(n_0_0_32), .S(n_0_0_28), .Z(out[0]));
   MUX2_X1 i_0_0_31 (.A(n_0_0_32), .B(n_0_0_33), .S(n_0_0_28), .Z(out[1]));
   MUX2_X1 i_0_0_32 (.A(n_0_0_33), .B(n_0_0_34), .S(n_0_0_28), .Z(out[2]));
   MUX2_X1 i_0_0_33 (.A(n_0_0_34), .B(n_0_0_35), .S(n_0_0_28), .Z(out[3]));
   MUX2_X1 i_0_0_34 (.A(n_0_0_35), .B(n_0_0_36), .S(n_0_0_28), .Z(out[4]));
   MUX2_X1 i_0_0_35 (.A(n_0_0_36), .B(n_0_0_37), .S(n_0_0_28), .Z(out[5]));
   MUX2_X1 i_0_0_36 (.A(n_0_0_37), .B(n_0_0_38), .S(n_0_0_28), .Z(out[6]));
   MUX2_X1 i_0_0_37 (.A(n_0_0_38), .B(n_0_0_39), .S(n_0_0_28), .Z(out[7]));
   INV_X1 i_0_0_43 (.A(second_operand[13]), .ZN(n_0_0_19));
   INV_X1 i_0_0_44 (.A(second_operand[14]), .ZN(n_0_0_20));
   OAI211_X1 i_0_0_45 (.A(n_0_0_19), .B(first_operand[13]), .C1(n_0_0_20), 
      .C2(first_operand[14]), .ZN(n_0_0_21));
   INV_X1 i_0_0_46 (.A(first_operand[14]), .ZN(n_0_0_22));
   OAI21_X1 i_0_0_47 (.A(n_0_0_21), .B1(second_operand[14]), .B2(n_0_0_22), 
      .ZN(n_0_0_23));
   INV_X1 i_0_0_48 (.A(second_operand[15]), .ZN(n_0_0_24));
   OAI21_X1 i_0_0_49 (.A(n_0_0_23), .B1(first_operand[15]), .B2(n_0_0_24), 
      .ZN(n_0_0_25));
   INV_X1 i_0_0_50 (.A(first_operand[15]), .ZN(n_0_0_26));
   OAI21_X1 i_0_0_51 (.A(n_0_0_25), .B1(second_operand[15]), .B2(n_0_0_26), 
      .ZN(n_0_0_27));
   MUX2_X1 i_0_0_55 (.A(second_operand[13]), .B(first_operand[13]), .S(n_0_0_27), 
      .Z(out[13]));
   MUX2_X1 i_0_0_56 (.A(second_operand[14]), .B(first_operand[14]), .S(n_0_0_27), 
      .Z(out[14]));
   MUX2_X1 i_0_0_57 (.A(second_operand[15]), .B(first_operand[15]), .S(n_0_0_27), 
      .Z(out[15]));
   NOR2_X1 i_0_0_9 (.A1(n_0_0_12), .A2(n_0_0_13), .ZN(n_0_0_9));
   AOI21_X1 i_0_0_10 (.A(n_0_0_10), .B1(n_0_0_16), .B2(n_0_0_29), .ZN(n_0_0_39));
   NOR2_X1 i_0_0_11 (.A1(n_0_0_8), .A2(n_0_0_29), .ZN(n_0_0_10));
   AOI21_X1 i_0_0_12 (.A(n_0_0_11), .B1(n_0_0_14), .B2(n_0_0_28), .ZN(out[9]));
   AND2_X1 i_0_0_13 (.A1(n_0_0_58), .A2(n_0_0_52), .ZN(n_0_0_11));
   NOR2_X1 i_0_0_14 (.A1(temp_result_wire[13]), .A2(n_0_0_82), .ZN(n_0_0_12));
   NOR2_X1 i_0_0_15 (.A1(temp_result_wire[9]), .A2(n_0_0_30), .ZN(n_0_0_13));
   OAI21_X1 i_0_0_24 (.A(n_0_0_15), .B1(n_0_0_40), .B2(n_0_0_84), .ZN(n_0_0_14));
   NAND2_X1 i_0_0_25 (.A1(n_0_0_16), .A2(n_0_0_84), .ZN(n_0_0_15));
   OAI21_X1 i_0_0_26 (.A(n_0_0_17), .B1(temp_result_wire[14]), .B2(n_0_0_82), 
      .ZN(n_0_0_16));
   OR2_X1 i_0_0_27 (.A1(temp_result_wire[10]), .A2(n_0_0_30), .ZN(n_0_0_17));
   INV_X1 i_0_0_28 (.A(n_0_0_84), .ZN(n_0_0_29));
   NAND2_X1 i_0_0_29 (.A1(n_0_0_42), .A2(n_0_0_18), .ZN(out[12]));
   NAND2_X1 i_0_0_38 (.A1(n_0_0_55), .A2(n_0_0_52), .ZN(n_0_0_18));
   MUX2_X1 i_0_0_39 (.A(temp_result_wire[16]), .B(temp_result_wire[12]), 
      .S(n_0_0_82), .Z(n_0_0_40));
   NAND2_X1 i_0_0_40 (.A1(temp_result_wire[14]), .A2(n_0_0_82), .ZN(n_0_0_41));
   NAND2_X1 i_0_0_41 (.A1(n_0_0_43), .A2(n_0_0_28), .ZN(n_0_0_42));
   OAI21_X1 i_0_0_42 (.A(n_0_0_44), .B1(n_0_0_45), .B2(n_0_0_84), .ZN(n_0_0_43));
   NAND2_X1 i_0_0_52 (.A1(n_0_0_57), .A2(n_0_0_84), .ZN(n_0_0_44));
   AOI21_X1 i_0_0_53 (.A(n_0_0_46), .B1(temp_result_wire[19]), .B2(n_0_0_30), 
      .ZN(n_0_0_45));
   INV_X1 i_0_0_54 (.A(n_0_0_47), .ZN(n_0_0_46));
   NAND2_X1 i_0_0_58 (.A1(temp_result_wire[15]), .A2(n_0_0_82), .ZN(n_0_0_47));
   NAND2_X1 i_0_0_59 (.A1(n_0_0_27), .A2(n_0_0_49), .ZN(n_0_0_48));
   INV_X1 i_0_0_60 (.A(second_operand[15]), .ZN(n_0_0_49));
   NAND2_X1 i_0_0_61 (.A1(n_0_0_27), .A2(n_0_0_51), .ZN(n_0_0_50));
   INV_X1 i_0_0_62 (.A(second_operand[14]), .ZN(n_0_0_51));
   OAI21_X1 i_0_0_63 (.A(n_0_0_53), .B1(first_operand[13]), .B2(n_0_0_27), 
      .ZN(n_0_0_52));
   NAND2_X1 i_0_0_64 (.A1(n_0_0_27), .A2(n_0_0_54), .ZN(n_0_0_53));
   INV_X1 i_0_0_65 (.A(second_operand[13]), .ZN(n_0_0_54));
   OAI21_X1 i_0_0_66 (.A(n_0_0_68), .B1(n_0_0_56), .B2(n_0_0_84), .ZN(n_0_0_55));
   AOI21_X1 i_0_0_67 (.A(n_0_0_69), .B1(temp_result_wire[18]), .B2(n_0_0_30), 
      .ZN(n_0_0_56));
   OAI21_X1 i_0_0_68 (.A(n_0_0_72), .B1(n_0_0_73), .B2(n_0_0_82), .ZN(n_0_0_57));
   OAI21_X1 i_0_0_69 (.A(n_0_0_61), .B1(n_0_0_58), .B2(n_0_0_52), .ZN(out[8]));
   INV_X1 i_0_0_70 (.A(n_0_0_59), .ZN(n_0_0_58));
   OAI21_X1 i_0_0_71 (.A(n_0_0_60), .B1(n_0_0_75), .B2(n_0_0_84), .ZN(n_0_0_59));
   OR3_X1 i_0_0_72 (.A1(n_0_0_12), .A2(n_0_0_13), .A3(n_0_0_83), .ZN(n_0_0_60));
   NAND2_X1 i_0_0_73 (.A1(n_0_0_39), .A2(n_0_0_52), .ZN(n_0_0_61));
   INV_X1 i_0_0_74 (.A(n_0_0_62), .ZN(out[10]));
   OAI221_X1 i_0_0_75 (.A(n_0_0_65), .B1(temp_result_wire[17]), .B2(n_0_0_81), 
      .C1(n_0_0_52), .C2(n_0_0_63), .ZN(n_0_0_62));
   AOI21_X1 i_0_0_76 (.A(n_0_0_64), .B1(n_0_0_75), .B2(n_0_0_78), .ZN(n_0_0_63));
   NOR3_X1 i_0_0_77 (.A1(temp_result_wire[13]), .A2(n_0_0_84), .A3(n_0_0_30), 
      .ZN(n_0_0_64));
   NAND2_X1 i_0_0_78 (.A1(n_0_0_14), .A2(n_0_0_52), .ZN(n_0_0_65));
   OAI211_X1 i_0_0_79 (.A(n_0_0_79), .B(n_0_0_70), .C1(n_0_0_52), .C2(n_0_0_66), 
      .ZN(out[11]));
   AOI21_X1 i_0_0_80 (.A(n_0_0_67), .B1(n_0_0_69), .B2(n_0_0_83), .ZN(n_0_0_66));
   INV_X1 i_0_0_81 (.A(n_0_0_68), .ZN(n_0_0_67));
   NAND2_X1 i_0_0_82 (.A1(n_0_0_40), .A2(n_0_0_84), .ZN(n_0_0_68));
   INV_X1 i_0_0_83 (.A(n_0_0_41), .ZN(n_0_0_69));
   NAND2_X1 i_0_0_84 (.A1(n_0_0_71), .A2(n_0_0_74), .ZN(n_0_0_70));
   OAI211_X1 i_0_0_85 (.A(n_0_0_83), .B(n_0_0_72), .C1(n_0_0_73), .C2(n_0_0_82), 
      .ZN(n_0_0_71));
   NAND2_X1 i_0_0_86 (.A1(temp_result_wire[13]), .A2(n_0_0_82), .ZN(n_0_0_72));
   INV_X1 i_0_0_87 (.A(temp_result_wire[17]), .ZN(n_0_0_73));
   AOI21_X1 i_0_0_88 (.A(n_0_0_28), .B1(n_0_0_75), .B2(n_0_0_78), .ZN(n_0_0_74));
   AOI21_X1 i_0_0_89 (.A(n_0_0_76), .B1(temp_result_wire[15]), .B2(n_0_0_30), 
      .ZN(n_0_0_75));
   INV_X1 i_0_0_90 (.A(n_0_0_77), .ZN(n_0_0_76));
   NAND2_X1 i_0_0_91 (.A1(temp_result_wire[11]), .A2(n_0_0_82), .ZN(n_0_0_77));
   INV_X1 i_0_0_92 (.A(n_0_0_29), .ZN(n_0_0_78));
   NAND2_X1 i_0_0_93 (.A1(temp_result_wire[18]), .A2(n_0_0_80), .ZN(n_0_0_79));
   INV_X1 i_0_0_94 (.A(n_0_0_81), .ZN(n_0_0_80));
   NAND3_X1 i_0_0_95 (.A1(n_0_0_28), .A2(n_0_0_83), .A3(n_0_0_30), .ZN(n_0_0_81));
   INV_X1 i_0_0_96 (.A(n_0_0_82), .ZN(n_0_0_30));
   OAI21_X1 i_0_0_97 (.A(n_0_0_48), .B1(n_0_0_27), .B2(first_operand[15]), 
      .ZN(n_0_0_82));
   INV_X1 i_0_0_98 (.A(n_0_0_84), .ZN(n_0_0_83));
   OAI21_X1 i_0_0_99 (.A(n_0_0_50), .B1(n_0_0_27), .B2(first_operand[14]), 
      .ZN(n_0_0_84));
   INV_X1 i_0_0_100 (.A(n_0_0_52), .ZN(n_0_0_28));
endmodule

module booth_16bit_multiplier(A, B, product);
   input [15:0]A;
   input [15:0]B;
   output [31:0]product;

   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_80;
   wire n_0_100;
   wire n_0_120;
   wire n_0_140;
   wire n_0_160;
   wire n_0_180;
   wire n_0_200;
   wire n_0_214;
   wire n_0_216;
   wire n_0_220;
   wire n_0_230;
   wire n_0_231;
   wire n_0_234;
   wire n_0_235;
   wire n_0_0;
   wire n_0_4;
   wire n_0_5;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_24;
   wire n_0_25;
   wire n_0_34;
   wire n_0_35;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_44;
   wire n_0_50;
   wire n_0_55;
   wire n_0_57;
   wire n_0_58;
   wire n_0_69;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_215;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_16;
   wire n_0_26;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_36;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_56;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_76;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_75;
   wire n_0_105;
   wire n_0_27;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_77;
   wire n_0_79;
   wire n_0_113;
   wire n_0_78;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_98;
   wire n_0_97;
   wire n_0_141;
   wire n_0_99;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_117;
   wire n_0_118;
   wire n_0_166;
   wire n_0_119;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_137;
   wire n_0_138;
   wire n_0_193;
   wire n_0_139;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_157;
   wire n_0_158;
   wire n_0_229;
   wire n_0_159;
   wire n_0_232;
   wire n_0_233;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_178;
   wire n_0_177;
   wire n_0_257;
   wire n_0_179;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_197;
   wire n_0_198;
   wire n_0_283;
   wire n_0_199;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_217;
   wire n_0_310;
   wire n_0_311;
   wire n_0_218;
   wire n_0_312;
   wire n_0_219;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_2;
   wire n_0_1;
   wire n_0_332;
   wire n_0_3;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_21;
   wire n_0_345;
   wire n_0_346;
   wire n_0_22;
   wire n_0_347;
   wire n_0_23;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_41;
   wire n_0_43;
   wire n_0_363;
   wire n_0_42;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_59;
   wire n_0_68;
   wire n_0_377;
   wire n_0_70;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_132;
   wire n_0_404;
   wire n_0_134;
   wire n_0_133;
   wire n_0_136;
   wire n_0_135;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_0;
   wire n_1_1;
   wire n_1_15;
   wire n_1_16;
   wire n_1_17;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;
   wire n_1_28;
   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire n_1_60;
   wire n_1_61;
   wire n_1_62;
   wire n_1_63;
   wire n_1_64;
   wire n_1_65;
   wire n_1_66;
   wire n_1_67;
   wire n_1_68;
   wire n_1_69;
   wire n_1_70;
   wire n_1_71;
   wire n_1_72;
   wire n_1_73;
   wire n_1_74;
   wire n_1_75;
   wire n_1_76;
   wire n_1_77;
   wire n_1_78;
   wire n_1_79;
   wire n_1_80;
   wire n_1_81;
   wire n_1_82;
   wire n_1_83;
   wire n_1_84;
   wire n_1_85;
   wire n_1_86;
   wire n_1_87;
   wire n_1_88;
   wire n_1_89;
   wire n_1_90;
   wire n_1_91;
   wire n_1_92;
   wire n_1_93;
   wire n_1_94;
   wire n_1_95;
   wire n_1_96;
   wire n_1_97;
   wire n_1_98;
   wire n_1_99;
   wire n_1_100;
   wire n_1_101;
   wire n_1_102;
   wire n_1_103;
   wire n_1_104;
   wire n_1_105;
   wire n_1_106;
   wire n_1_107;
   wire n_1_108;
   wire n_1_109;
   wire n_1_110;
   wire n_1_111;
   wire n_1_112;
   wire n_1_113;
   wire n_1_114;
   wire n_1_115;
   wire n_1_116;
   wire n_1_117;
   wire n_1_118;
   wire n_1_119;
   wire n_1_120;
   wire n_1_121;
   wire n_1_122;
   wire n_1_123;
   wire n_1_124;
   wire n_1_125;
   wire n_1_126;
   wire n_1_127;
   wire n_1_128;
   wire n_1_129;
   wire n_1_130;
   wire n_1_131;
   wire n_1_132;
   wire n_1_133;
   wire n_1_134;
   wire n_1_135;
   wire n_1_136;
   wire n_1_137;
   wire n_1_138;
   wire n_1_139;
   wire n_1_140;
   wire n_1_141;
   wire n_1_142;
   wire n_1_143;
   wire n_1_144;
   wire n_1_145;
   wire n_1_146;
   wire n_1_147;
   wire n_1_148;
   wire n_1_149;
   wire n_1_150;
   wire n_1_151;
   wire n_1_152;
   wire n_1_153;
   wire n_1_154;
   wire n_1_155;
   wire n_1_156;
   wire n_1_157;
   wire n_1_158;
   wire n_1_159;
   wire n_1_160;
   wire n_1_161;
   wire n_1_162;
   wire n_1_163;
   wire n_1_164;
   wire n_1_165;
   wire n_1_166;
   wire n_1_167;
   wire n_1_168;
   wire n_1_169;
   wire n_1_170;
   wire n_1_171;
   wire n_1_172;
   wire n_1_173;
   wire n_1_174;
   wire n_1_175;
   wire n_1_176;
   wire n_1_177;

   datapath__0_1 i_2 (.B({B[15], uc_0, uc_1, uc_2, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({n_124, n_126, 
      n_125, n_264, n_263, n_262, n_261, n_260, n_259, n_258, n_257, n_256, 
      n_255, n_148, n_147, n_146}), .p_1({n_15, n_14, n_13, n_12, n_11, n_10, 
      n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0}));
   datapath__0_6 i_5 (.B({B[15], uc_3, uc_4, uc_5, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_6, n_123, n_122, 
      n_254, n_253, n_121, n_252, n_251, n_250, n_249, n_145, n_248, n_247, 
      n_144, n_143, n_142}), .p_1({n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
      n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16}));
   datapath__0_7 i_6 (.p_0({n_126, n_125, n_264, n_263, n_262, n_261, n_260, 
      n_259, n_258, n_257, n_256, n_255, n_148, n_147, n_146, B[0]}), .p_1({uc_7, 
      n_123, n_122, n_254, n_253, n_121, n_252, n_251, n_250, n_249, n_145, 
      n_248, n_247, n_144, n_143, n_142}), .p_2({n_47, n_46, n_45, n_44, n_43, 
      n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32}));
   datapath__0_12 i_9 (.B({B[15], uc_8, uc_9, uc_10, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_11, n_120, 
      n_119, n_246, n_245, n_118, n_117, n_244, n_243, n_242, n_241, n_141, 
      n_240, n_239, n_140, n_116}), .p_1({n_63, n_62, n_61, n_60, n_59, n_58, 
      n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48}));
   datapath__0_13 i_10 (.p_0({n_126, n_125, n_264, n_263, n_262, n_261, n_260, 
      n_259, n_258, n_257, n_256, n_255, n_148, n_147, n_146, B[0]}), .p_1({
      uc_12, n_120, n_119, n_246, n_245, n_118, n_117, n_244, n_243, n_242, 
      n_241, n_141, n_240, n_239, n_140, n_116}), .p_2({n_79, n_78, n_77, n_76, 
      n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64}));
   datapath__0_18 i_13 (.B({B[15], uc_13, uc_14, uc_15, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_16, n_115, 
      n_238, n_237, n_236, n_114, n_235, n_234, n_233, n_232, n_231, n_230, 
      n_139, n_229, n_138, n_113}), .p_1({n_95, n_94, n_93, n_92, n_91, n_90, 
      n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80}));
   datapath__0_19 i_14 (.p_0({n_126, n_125, n_264, n_263, n_262, n_261, n_260, 
      n_259, n_258, n_257, n_256, n_255, n_148, n_147, n_146, B[0]}), .p_1({
      uc_17, n_115, n_238, n_237, n_236, n_114, n_235, n_234, n_233, n_232, 
      n_231, n_230, n_139, n_229, n_138, n_113}), .p_2({n_111, n_110, n_109, 
      n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
      n_97, n_96}));
   INV_X1 i_0_108 (.A(n_0_60), .ZN(product[12]));
   AOI222_X1 i_0_109 (.A1(n_438), .A2(n_0_79), .B1(n_438), .B2(n_0_78), .C1(
      n_149), .C2(n_0_77), .ZN(n_0_60));
   INV_X1 i_0_110 (.A(n_0_61), .ZN(product[13]));
   AOI222_X1 i_0_111 (.A1(n_424), .A2(n_0_79), .B1(n_417), .B2(n_0_78), .C1(
      n_150), .C2(n_0_77), .ZN(n_0_61));
   INV_X1 i_0_112 (.A(n_0_62), .ZN(product[14]));
   AOI222_X1 i_0_113 (.A1(n_425), .A2(n_0_79), .B1(n_418), .B2(n_0_78), .C1(
      n_151), .C2(n_0_77), .ZN(n_0_62));
   INV_X1 i_0_144 (.A(n_0_80), .ZN(product[11]));
   AOI222_X1 i_0_145 (.A1(n_437), .A2(n_0_98), .B1(n_437), .B2(n_0_99), .C1(
      n_156), .C2(n_0_97), .ZN(n_0_80));
   INV_X1 i_0_180 (.A(n_0_100), .ZN(product[10]));
   AOI222_X1 i_0_181 (.A1(n_436), .A2(n_0_118), .B1(n_436), .B2(n_0_119), 
      .C1(n_164), .C2(n_0_117), .ZN(n_0_100));
   INV_X1 i_0_216 (.A(n_0_120), .ZN(product[9]));
   AOI222_X1 i_0_217 (.A1(n_435), .A2(n_0_138), .B1(n_435), .B2(n_0_139), 
      .C1(n_173), .C2(n_0_137), .ZN(n_0_120));
   INV_X1 i_0_252 (.A(n_0_140), .ZN(product[8]));
   AOI222_X1 i_0_253 (.A1(n_434), .A2(n_0_158), .B1(n_434), .B2(n_0_159), 
      .C1(n_183), .C2(n_0_157), .ZN(n_0_140));
   INV_X1 i_0_288 (.A(n_0_160), .ZN(product[7]));
   AOI222_X1 i_0_289 (.A1(n_433), .A2(n_0_178), .B1(n_433), .B2(n_0_179), 
      .C1(n_194), .C2(n_0_177), .ZN(n_0_160));
   INV_X1 i_0_324 (.A(n_0_180), .ZN(product[6]));
   AOI222_X1 i_0_325 (.A1(n_432), .A2(n_0_198), .B1(n_432), .B2(n_0_199), 
      .C1(n_206), .C2(n_0_197), .ZN(n_0_180));
   INV_X1 i_0_360 (.A(n_0_200), .ZN(product[5]));
   AOI222_X1 i_0_361 (.A1(n_431), .A2(n_0_218), .B1(n_431), .B2(n_0_219), 
      .C1(n_134), .C2(n_0_217), .ZN(n_0_200));
   AOI221_X1 i_0_389 (.A(n_0_216), .B1(n_440), .B2(n_0_218), .C1(n_439), 
      .C2(n_0_219), .ZN(n_0_214));
   AND2_X1 i_0_392 (.A1(n_112), .A2(n_0_217), .ZN(n_0_216));
   INV_X1 i_0_396 (.A(n_0_220), .ZN(product[4]));
   AOI222_X1 i_0_397 (.A1(n_80), .A2(n_0_2), .B1(n_96), .B2(n_0_3), .C1(n_113), 
      .C2(n_0_1), .ZN(n_0_220));
   AOI222_X1 i_0_417 (.A1(n_90), .A2(n_0_2), .B1(n_106), .B2(n_0_3), .C1(n_114), 
      .C2(n_0_1), .ZN(n_0_230));
   AOI222_X1 i_0_419 (.A1(n_107), .A2(n_0_3), .B1(n_91), .B2(n_0_2), .C1(n_236), 
      .C2(n_0_1), .ZN(n_0_231));
   AOI221_X1 i_0_425 (.A(n_0_0), .B1(n_94), .B2(n_0_2), .C1(n_110), .C2(n_0_3), 
      .ZN(n_0_234));
   INV_X1 i_0_426 (.A(n_0_235), .ZN(n_112));
   AOI221_X1 i_0_427 (.A(n_0_0), .B1(n_95), .B2(n_0_2), .C1(n_111), .C2(n_0_3), 
      .ZN(n_0_235));
   AND2_X1 i_0_428 (.A1(n_115), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_432 (.A(n_0_4), .ZN(product[3]));
   AOI222_X1 i_0_433 (.A1(n_48), .A2(n_0_22), .B1(n_64), .B2(n_0_23), .C1(n_116), 
      .C2(n_0_21), .ZN(n_0_4));
   INV_X1 i_0_434 (.A(n_0_5), .ZN(n_113));
   AOI222_X1 i_0_435 (.A1(n_49), .A2(n_0_22), .B1(n_65), .B2(n_0_23), .C1(n_140), 
      .C2(n_0_21), .ZN(n_0_5));
   AOI222_X1 i_0_451 (.A1(n_57), .A2(n_0_22), .B1(n_73), .B2(n_0_23), .C1(n_117), 
      .C2(n_0_21), .ZN(n_0_13));
   AOI222_X1 i_0_453 (.A1(n_58), .A2(n_0_22), .B1(n_74), .B2(n_0_23), .C1(n_118), 
      .C2(n_0_21), .ZN(n_0_14));
   INV_X1 i_0_454 (.A(n_0_15), .ZN(n_114));
   AOI222_X1 i_0_455 (.A1(n_59), .A2(n_0_22), .B1(n_75), .B2(n_0_23), .C1(n_245), 
      .C2(n_0_21), .ZN(n_0_15));
   AOI222_X1 i_0_459 (.A1(n_77), .A2(n_0_23), .B1(n_61), .B2(n_0_22), .C1(n_119), 
      .C2(n_0_21), .ZN(n_0_17));
   AOI221_X1 i_0_461 (.A(n_0_20), .B1(n_62), .B2(n_0_22), .C1(n_78), .C2(n_0_23), 
      .ZN(n_0_18));
   INV_X1 i_0_462 (.A(n_0_19), .ZN(n_115));
   AOI221_X1 i_0_463 (.A(n_0_20), .B1(n_63), .B2(n_0_22), .C1(n_79), .C2(n_0_23), 
      .ZN(n_0_19));
   AND2_X1 i_0_464 (.A1(n_120), .A2(n_0_21), .ZN(n_0_20));
   INV_X1 i_0_468 (.A(n_0_24), .ZN(product[2]));
   AOI222_X1 i_0_469 (.A1(n_16), .A2(n_0_42), .B1(n_32), .B2(n_0_43), .C1(n_142), 
      .C2(n_0_41), .ZN(n_0_24));
   INV_X1 i_0_470 (.A(n_0_25), .ZN(n_116));
   AOI222_X1 i_0_471 (.A1(n_17), .A2(n_0_42), .B1(n_33), .B2(n_0_43), .C1(n_143), 
      .C2(n_0_41), .ZN(n_0_25));
   INV_X1 i_0_488 (.A(n_0_34), .ZN(n_117));
   AOI222_X1 i_0_489 (.A1(n_26), .A2(n_0_42), .B1(n_42), .B2(n_0_43), .C1(n_121), 
      .C2(n_0_41), .ZN(n_0_34));
   INV_X1 i_0_490 (.A(n_0_35), .ZN(n_118));
   AOI222_X1 i_0_491 (.A1(n_27), .A2(n_0_42), .B1(n_43), .B2(n_0_43), .C1(n_253), 
      .C2(n_0_41), .ZN(n_0_35));
   AOI222_X1 i_0_495 (.A1(n_45), .A2(n_0_43), .B1(n_29), .B2(n_0_42), .C1(n_122), 
      .C2(n_0_41), .ZN(n_0_37));
   INV_X1 i_0_496 (.A(n_0_38), .ZN(n_119));
   AOI221_X1 i_0_497 (.A(n_0_40), .B1(n_30), .B2(n_0_42), .C1(n_46), .C2(n_0_43), 
      .ZN(n_0_38));
   INV_X1 i_0_498 (.A(n_0_39), .ZN(n_120));
   AOI221_X1 i_0_499 (.A(n_0_40), .B1(n_31), .B2(n_0_42), .C1(n_47), .C2(n_0_43), 
      .ZN(n_0_39));
   AND2_X1 i_0_500 (.A1(n_123), .A2(n_0_41), .ZN(n_0_40));
   INV_X1 i_0_504 (.A(n_0_44), .ZN(product[1]));
   AOI222_X1 i_0_505 (.A1(n_0), .A2(n_0_70), .B1(B[0]), .B2(n_0_59), .C1(n_146), 
      .C2(n_0_68), .ZN(n_0_44));
   AOI222_X1 i_0_517 (.A1(n_6), .A2(n_0_70), .B1(n_257), .B2(n_0_59), .C1(n_258), 
      .C2(n_0_68), .ZN(n_0_50));
   INV_X1 i_0_526 (.A(n_0_55), .ZN(n_121));
   AOI222_X1 i_0_527 (.A1(n_262), .A2(n_0_59), .B1(n_11), .B2(n_0_70), .C1(n_263), 
      .C2(n_0_68), .ZN(n_0_55));
   AOI222_X1 i_0_531 (.A1(n_13), .A2(n_0_70), .B1(n_264), .B2(n_0_59), .C1(n_125), 
      .C2(n_0_68), .ZN(n_0_57));
   INV_X1 i_0_532 (.A(n_0_58), .ZN(n_122));
   AOI222_X1 i_0_533 (.A1(n_125), .A2(n_0_59), .B1(n_14), .B2(n_0_70), .C1(n_126), 
      .C2(n_0_68), .ZN(n_0_58));
   INV_X1 i_0_536 (.A(n_0_69), .ZN(n_123));
   AOI22_X1 i_0_537 (.A1(n_15), .A2(n_0_70), .B1(A[1]), .B2(n_126), .ZN(n_0_69));
   AND2_X1 i_0_539 (.A1(B[0]), .A2(A[0]), .ZN(product[0]));
   AND2_X1 i_0_540 (.A1(A[0]), .A2(n_126), .ZN(n_124));
   AOI21_X1 i_0_554 (.A(n_0_71), .B1(B[15]), .B2(n_0_72), .ZN(n_125));
   XNOR2_X1 i_0_555 (.A(B[15]), .B(n_0_71), .ZN(n_126));
   NOR2_X1 i_0_556 (.A1(B[15]), .A2(n_0_72), .ZN(n_0_71));
   INV_X1 i_0_557 (.A(n_0_73), .ZN(n_0_72));
   NOR2_X1 i_0_558 (.A1(B[15]), .A2(n_0_74), .ZN(n_0_73));
   INV_X1 i_0_559 (.A(n_0_75), .ZN(n_0_74));
   INV_X1 i_0_584 (.A(A[1]), .ZN(n_0_153));
   INV_X1 i_0_585 (.A(A[2]), .ZN(n_0_154));
   INV_X1 i_0_586 (.A(A[3]), .ZN(n_0_155));
   INV_X1 i_0_587 (.A(A[4]), .ZN(n_0_156));
   INV_X1 i_0_588 (.A(A[5]), .ZN(n_0_173));
   INV_X1 i_0_589 (.A(A[6]), .ZN(n_0_174));
   INV_X1 i_0_590 (.A(A[7]), .ZN(n_0_175));
   INV_X1 i_0_591 (.A(A[8]), .ZN(n_0_176));
   INV_X1 i_0_592 (.A(A[9]), .ZN(n_0_194));
   INV_X1 i_0_593 (.A(A[10]), .ZN(n_0_195));
   INV_X1 i_0_594 (.A(A[11]), .ZN(n_0_196));
   INV_X1 i_0_595 (.A(A[15]), .ZN(n_0_215));
   NAND3_X1 i_0_0 (.A1(n_0_6), .A2(n_0_8), .A3(n_0_7), .ZN(product[19]));
   NAND2_X1 i_0_1 (.A1(n_430), .A2(n_0_79), .ZN(n_0_6));
   NAND2_X1 i_0_2 (.A1(n_127), .A2(n_0_77), .ZN(n_0_7));
   NAND2_X1 i_0_3 (.A1(n_423), .A2(n_0_78), .ZN(n_0_8));
   OAI21_X1 i_0_4 (.A(n_0_9), .B1(n_0_11), .B2(n_0_141), .ZN(n_127));
   AOI22_X1 i_0_5 (.A1(n_408), .A2(n_0_98), .B1(n_128), .B2(n_0_97), .ZN(n_0_9));
   OR2_X1 i_0_6 (.A1(n_0_99), .A2(n_0_98), .ZN(n_0_10));
   INV_X1 i_0_7 (.A(n_416), .ZN(n_0_11));
   OAI21_X1 i_0_8 (.A(n_0_12), .B1(n_0_16), .B2(n_0_166), .ZN(n_128));
   AOI22_X1 i_0_9 (.A1(n_391), .A2(n_0_118), .B1(n_129), .B2(n_0_117), .ZN(
      n_0_12));
   INV_X1 i_0_10 (.A(n_400), .ZN(n_0_16));
   OAI21_X1 i_0_11 (.A(n_0_26), .B1(n_0_28), .B2(n_0_193), .ZN(n_129));
   AOI22_X1 i_0_12 (.A1(n_372), .A2(n_0_138), .B1(n_130), .B2(n_0_137), .ZN(
      n_0_26));
   INV_X1 i_0_13 (.A(n_382), .ZN(n_0_28));
   OAI21_X1 i_0_14 (.A(n_0_29), .B1(n_0_30), .B2(n_0_229), .ZN(n_130));
   AOI22_X1 i_0_15 (.A1(n_351), .A2(n_0_158), .B1(n_131), .B2(n_0_157), .ZN(
      n_0_29));
   INV_X1 i_0_16 (.A(n_362), .ZN(n_0_30));
   OAI21_X1 i_0_17 (.A(n_0_31), .B1(n_0_33), .B2(n_0_257), .ZN(n_131));
   AOI22_X1 i_0_18 (.A1(n_328), .A2(n_0_178), .B1(n_132), .B2(n_0_177), .ZN(
      n_0_31));
   NAND2_X1 i_0_19 (.A1(n_0_257), .A2(n_0_246), .ZN(n_0_32));
   INV_X1 i_0_20 (.A(n_340), .ZN(n_0_33));
   OAI21_X1 i_0_21 (.A(n_0_36), .B1(n_0_45), .B2(n_0_283), .ZN(n_132));
   AOI22_X1 i_0_22 (.A1(n_303), .A2(n_0_198), .B1(n_133), .B2(n_0_197), .ZN(
      n_0_36));
   INV_X1 i_0_23 (.A(n_316), .ZN(n_0_45));
   INV_X1 i_0_24 (.A(n_0_214), .ZN(n_133));
   NAND2_X1 i_0_25 (.A1(n_0_47), .A2(n_0_46), .ZN(n_134));
   NAND2_X1 i_0_26 (.A1(n_97), .A2(n_0_3), .ZN(n_0_46));
   AOI22_X1 i_0_27 (.A1(n_81), .A2(n_0_2), .B1(n_138), .B2(n_0_1), .ZN(n_0_47));
   NAND2_X1 i_0_28 (.A1(n_99), .A2(n_0_3), .ZN(n_0_48));
   AOI22_X1 i_0_29 (.A1(n_83), .A2(n_0_2), .B1(n_139), .B2(n_0_1), .ZN(n_0_49));
   OAI21_X1 i_0_30 (.A(n_0_52), .B1(n_0_156), .B2(A[3]), .ZN(n_0_51));
   NAND2_X1 i_0_31 (.A1(n_0_53), .A2(n_0_54), .ZN(n_0_52));
   INV_X1 i_0_32 (.A(n_0_155), .ZN(n_0_53));
   INV_X1 i_0_33 (.A(A[4]), .ZN(n_0_54));
   INV_X1 i_0_34 (.A(n_0_230), .ZN(n_135));
   INV_X1 i_0_35 (.A(n_0_231), .ZN(n_136));
   INV_X1 i_0_36 (.A(n_0_234), .ZN(n_137));
   OAI211_X1 i_0_37 (.A(n_0_56), .B(n_0_63), .C1(n_0_27), .C2(n_0_65), .ZN(n_138));
   NAND2_X1 i_0_38 (.A1(n_50), .A2(n_0_22), .ZN(n_0_56));
   NAND2_X1 i_0_39 (.A1(n_66), .A2(n_0_23), .ZN(n_0_63));
   OAI211_X1 i_0_40 (.A(n_0_66), .B(n_0_64), .C1(n_0_67), .C2(n_0_65), .ZN(n_139));
   NAND2_X1 i_0_41 (.A1(n_52), .A2(n_0_22), .ZN(n_0_64));
   INV_X1 i_0_42 (.A(n_0_21), .ZN(n_0_65));
   NAND2_X1 i_0_43 (.A1(n_68), .A2(n_0_23), .ZN(n_0_66));
   INV_X1 i_0_44 (.A(n_141), .ZN(n_0_67));
   NAND2_X1 i_0_45 (.A1(n_0_81), .A2(n_0_76), .ZN(n_140));
   NAND2_X1 i_0_46 (.A1(n_34), .A2(n_0_43), .ZN(n_0_76));
   AOI22_X1 i_0_47 (.A1(n_18), .A2(n_0_42), .B1(n_144), .B2(n_0_41), .ZN(n_0_81));
   NAND2_X1 i_0_48 (.A1(n_0_83), .A2(n_0_82), .ZN(n_141));
   NAND2_X1 i_0_49 (.A1(n_21), .A2(n_0_42), .ZN(n_0_82));
   AOI22_X1 i_0_50 (.A1(n_37), .A2(n_0_43), .B1(n_145), .B2(n_0_41), .ZN(n_0_83));
   OAI21_X1 i_0_51 (.A(n_0_88), .B1(n_0_104), .B2(n_0_84), .ZN(n_142));
   INV_X1 i_0_52 (.A(n_0_85), .ZN(n_0_84));
   NAND2_X1 i_0_53 (.A1(n_0_87), .A2(n_0_86), .ZN(n_0_85));
   NAND2_X1 i_0_54 (.A1(A[1]), .A2(n_147), .ZN(n_0_86));
   NAND2_X1 i_0_55 (.A1(n_0_92), .A2(n_1), .ZN(n_0_87));
   NAND3_X1 i_0_56 (.A1(n_0_96), .A2(n_0_104), .A3(n_146), .ZN(n_0_88));
   OAI21_X1 i_0_57 (.A(n_0_94), .B1(n_0_104), .B2(n_0_89), .ZN(n_143));
   INV_X1 i_0_58 (.A(n_0_90), .ZN(n_0_89));
   NAND2_X1 i_0_59 (.A1(n_0_91), .A2(n_0_93), .ZN(n_0_90));
   NAND2_X1 i_0_60 (.A1(n_0_92), .A2(n_2), .ZN(n_0_91));
   INV_X1 i_0_61 (.A(A[1]), .ZN(n_0_92));
   NAND2_X1 i_0_62 (.A1(A[1]), .A2(n_148), .ZN(n_0_93));
   NAND3_X1 i_0_63 (.A1(n_0_96), .A2(n_0_104), .A3(n_147), .ZN(n_0_94));
   NAND3_X1 i_0_64 (.A1(n_0_103), .A2(n_0_101), .A3(n_0_95), .ZN(n_144));
   NAND3_X1 i_0_65 (.A1(n_0_96), .A2(n_0_104), .A3(n_148), .ZN(n_0_95));
   INV_X1 i_0_66 (.A(n_0_153), .ZN(n_0_96));
   NAND2_X1 i_0_67 (.A1(n_0_68), .A2(n_255), .ZN(n_0_101));
   NAND2_X1 i_0_68 (.A1(A[1]), .A2(A[0]), .ZN(n_0_102));
   NAND2_X1 i_0_69 (.A1(n_3), .A2(n_0_70), .ZN(n_0_103));
   INV_X1 i_0_70 (.A(A[0]), .ZN(n_0_104));
   INV_X1 i_0_71 (.A(n_0_50), .ZN(n_145));
   AOI21_X1 i_0_72 (.A(n_0_136), .B1(B[1]), .B2(B[0]), .ZN(n_146));
   AOI21_X1 i_0_73 (.A(n_0_134), .B1(B[2]), .B2(n_0_135), .ZN(n_147));
   AOI21_X1 i_0_74 (.A(n_0_132), .B1(B[3]), .B2(n_0_133), .ZN(n_148));
   INV_X1 i_0_75 (.A(n_0_105), .ZN(n_0_75));
   OR2_X1 i_0_76 (.A1(n_0_391), .A2(B[15]), .ZN(n_0_105));
   INV_X1 i_0_77 (.A(n_239), .ZN(n_0_27));
   OAI21_X1 i_0_78 (.A(n_0_106), .B1(n_0_107), .B2(n_0_113), .ZN(product[15]));
   AOI22_X1 i_0_79 (.A1(n_426), .A2(n_0_79), .B1(n_152), .B2(n_0_77), .ZN(
      n_0_106));
   INV_X1 i_0_80 (.A(n_419), .ZN(n_0_107));
   OAI21_X1 i_0_81 (.A(n_0_108), .B1(n_0_109), .B2(n_0_113), .ZN(product[16]));
   AOI22_X1 i_0_82 (.A1(n_427), .A2(n_0_79), .B1(n_153), .B2(n_0_77), .ZN(
      n_0_108));
   INV_X1 i_0_83 (.A(n_420), .ZN(n_0_109));
   OAI21_X1 i_0_84 (.A(n_0_110), .B1(n_0_111), .B2(n_0_113), .ZN(product[17]));
   AOI22_X1 i_0_85 (.A1(n_428), .A2(n_0_79), .B1(n_154), .B2(n_0_77), .ZN(
      n_0_110));
   INV_X1 i_0_86 (.A(n_421), .ZN(n_0_111));
   OAI21_X1 i_0_87 (.A(n_0_112), .B1(n_0_114), .B2(n_0_113), .ZN(product[18]));
   AOI22_X1 i_0_88 (.A1(n_429), .A2(n_0_79), .B1(n_155), .B2(n_0_77), .ZN(
      n_0_112));
   NOR2_X1 i_0_89 (.A1(n_0_79), .A2(n_0_78), .ZN(n_0_77));
   NOR2_X1 i_0_90 (.A1(n_0_215), .A2(A[11]), .ZN(n_0_79));
   INV_X1 i_0_91 (.A(n_0_78), .ZN(n_0_113));
   NOR2_X1 i_0_92 (.A1(A[15]), .A2(n_0_196), .ZN(n_0_78));
   INV_X1 i_0_93 (.A(n_422), .ZN(n_0_114));
   NAND2_X1 i_0_94 (.A1(n_0_115), .A2(n_0_116), .ZN(n_149));
   AOI22_X1 i_0_95 (.A1(n_409), .A2(n_0_99), .B1(n_0_97), .B2(n_157), .ZN(
      n_0_115));
   NAND2_X1 i_0_96 (.A1(n_401), .A2(n_0_98), .ZN(n_0_116));
   OAI21_X1 i_0_97 (.A(n_0_121), .B1(n_0_122), .B2(n_0_141), .ZN(n_150));
   AOI22_X1 i_0_98 (.A1(n_402), .A2(n_0_98), .B1(n_0_97), .B2(n_158), .ZN(
      n_0_121));
   INV_X1 i_0_99 (.A(n_410), .ZN(n_0_122));
   OAI21_X1 i_0_100 (.A(n_0_123), .B1(n_0_124), .B2(n_0_141), .ZN(n_151));
   AOI22_X1 i_0_101 (.A1(n_403), .A2(n_0_98), .B1(n_0_97), .B2(n_159), .ZN(
      n_0_123));
   INV_X1 i_0_102 (.A(n_411), .ZN(n_0_124));
   OAI21_X1 i_0_103 (.A(n_0_125), .B1(n_0_126), .B2(n_0_141), .ZN(n_152));
   AOI22_X1 i_0_104 (.A1(n_404), .A2(n_0_98), .B1(n_0_97), .B2(n_160), .ZN(
      n_0_125));
   INV_X1 i_0_105 (.A(n_412), .ZN(n_0_126));
   OAI21_X1 i_0_106 (.A(n_0_127), .B1(n_0_128), .B2(n_0_141), .ZN(n_153));
   AOI22_X1 i_0_107 (.A1(n_405), .A2(n_0_98), .B1(n_0_97), .B2(n_161), .ZN(
      n_0_127));
   INV_X1 i_0_114 (.A(n_413), .ZN(n_0_128));
   OAI21_X1 i_0_115 (.A(n_0_129), .B1(n_0_130), .B2(n_0_141), .ZN(n_154));
   AOI22_X1 i_0_116 (.A1(n_406), .A2(n_0_98), .B1(n_0_97), .B2(n_162), .ZN(
      n_0_129));
   INV_X1 i_0_117 (.A(n_414), .ZN(n_0_130));
   OAI21_X1 i_0_118 (.A(n_0_131), .B1(n_0_142), .B2(n_0_141), .ZN(n_155));
   AOI22_X1 i_0_119 (.A1(n_407), .A2(n_0_98), .B1(n_0_97), .B2(n_163), .ZN(
      n_0_131));
   NOR2_X1 i_0_120 (.A1(n_0_195), .A2(A[11]), .ZN(n_0_98));
   INV_X1 i_0_121 (.A(n_0_10), .ZN(n_0_97));
   INV_X1 i_0_122 (.A(n_0_99), .ZN(n_0_141));
   NOR2_X1 i_0_123 (.A1(n_0_196), .A2(A[10]), .ZN(n_0_99));
   INV_X1 i_0_124 (.A(n_415), .ZN(n_0_142));
   OAI21_X1 i_0_125 (.A(n_0_143), .B1(n_0_144), .B2(n_0_166), .ZN(n_156));
   AOI22_X1 i_0_126 (.A1(n_383), .A2(n_0_118), .B1(n_165), .B2(n_0_117), 
      .ZN(n_0_143));
   INV_X1 i_0_127 (.A(n_392), .ZN(n_0_144));
   OAI21_X1 i_0_128 (.A(n_0_145), .B1(n_0_146), .B2(n_0_166), .ZN(n_157));
   AOI22_X1 i_0_129 (.A1(n_384), .A2(n_0_118), .B1(n_166), .B2(n_0_117), 
      .ZN(n_0_145));
   INV_X1 i_0_130 (.A(n_393), .ZN(n_0_146));
   OAI21_X1 i_0_131 (.A(n_0_147), .B1(n_0_148), .B2(n_0_166), .ZN(n_158));
   AOI22_X1 i_0_132 (.A1(n_385), .A2(n_0_118), .B1(n_167), .B2(n_0_117), 
      .ZN(n_0_147));
   INV_X1 i_0_133 (.A(n_394), .ZN(n_0_148));
   OAI21_X1 i_0_134 (.A(n_0_149), .B1(n_0_150), .B2(n_0_166), .ZN(n_159));
   AOI22_X1 i_0_135 (.A1(n_386), .A2(n_0_118), .B1(n_168), .B2(n_0_117), 
      .ZN(n_0_149));
   INV_X1 i_0_136 (.A(n_395), .ZN(n_0_150));
   OAI21_X1 i_0_137 (.A(n_0_151), .B1(n_0_152), .B2(n_0_166), .ZN(n_160));
   AOI22_X1 i_0_138 (.A1(n_387), .A2(n_0_118), .B1(n_169), .B2(n_0_117), 
      .ZN(n_0_151));
   INV_X1 i_0_139 (.A(n_396), .ZN(n_0_152));
   OAI21_X1 i_0_140 (.A(n_0_161), .B1(n_0_162), .B2(n_0_166), .ZN(n_161));
   AOI22_X1 i_0_141 (.A1(n_388), .A2(n_0_118), .B1(n_170), .B2(n_0_117), 
      .ZN(n_0_161));
   INV_X1 i_0_142 (.A(n_397), .ZN(n_0_162));
   OAI21_X1 i_0_143 (.A(n_0_163), .B1(n_0_164), .B2(n_0_166), .ZN(n_162));
   AOI22_X1 i_0_146 (.A1(n_389), .A2(n_0_118), .B1(n_171), .B2(n_0_117), 
      .ZN(n_0_163));
   INV_X1 i_0_147 (.A(n_398), .ZN(n_0_164));
   OAI21_X1 i_0_148 (.A(n_0_165), .B1(n_0_167), .B2(n_0_166), .ZN(n_163));
   AOI22_X1 i_0_149 (.A1(n_390), .A2(n_0_118), .B1(n_172), .B2(n_0_117), 
      .ZN(n_0_165));
   NOR2_X1 i_0_150 (.A1(n_0_119), .A2(n_0_118), .ZN(n_0_117));
   NOR2_X1 i_0_151 (.A1(A[10]), .A2(n_0_194), .ZN(n_0_118));
   INV_X1 i_0_152 (.A(n_0_119), .ZN(n_0_166));
   NOR2_X1 i_0_153 (.A1(n_0_195), .A2(A[9]), .ZN(n_0_119));
   INV_X1 i_0_154 (.A(n_399), .ZN(n_0_167));
   OAI21_X1 i_0_155 (.A(n_0_168), .B1(n_0_169), .B2(n_0_193), .ZN(n_164));
   AOI22_X1 i_0_156 (.A1(n_363), .A2(n_0_138), .B1(n_174), .B2(n_0_137), 
      .ZN(n_0_168));
   INV_X1 i_0_157 (.A(n_373), .ZN(n_0_169));
   NAND2_X1 i_0_158 (.A1(n_0_171), .A2(n_0_170), .ZN(n_165));
   AOI22_X1 i_0_159 (.A1(n_374), .A2(n_0_139), .B1(n_175), .B2(n_0_137), 
      .ZN(n_0_170));
   NAND2_X1 i_0_160 (.A1(n_364), .A2(n_0_138), .ZN(n_0_171));
   NAND2_X1 i_0_161 (.A1(n_0_181), .A2(n_0_172), .ZN(n_166));
   AOI22_X1 i_0_162 (.A1(n_375), .A2(n_0_139), .B1(n_176), .B2(n_0_137), 
      .ZN(n_0_172));
   NAND2_X1 i_0_163 (.A1(n_365), .A2(n_0_138), .ZN(n_0_181));
   OAI21_X1 i_0_164 (.A(n_0_182), .B1(n_0_183), .B2(n_0_193), .ZN(n_167));
   AOI22_X1 i_0_165 (.A1(n_366), .A2(n_0_138), .B1(n_177), .B2(n_0_137), 
      .ZN(n_0_182));
   INV_X1 i_0_166 (.A(n_376), .ZN(n_0_183));
   OAI21_X1 i_0_167 (.A(n_0_184), .B1(n_0_185), .B2(n_0_193), .ZN(n_168));
   AOI22_X1 i_0_168 (.A1(n_367), .A2(n_0_138), .B1(n_178), .B2(n_0_137), 
      .ZN(n_0_184));
   INV_X1 i_0_169 (.A(n_377), .ZN(n_0_185));
   OAI21_X1 i_0_170 (.A(n_0_186), .B1(n_0_187), .B2(n_0_193), .ZN(n_169));
   AOI22_X1 i_0_171 (.A1(n_368), .A2(n_0_138), .B1(n_179), .B2(n_0_137), 
      .ZN(n_0_186));
   INV_X1 i_0_172 (.A(n_378), .ZN(n_0_187));
   OAI21_X1 i_0_173 (.A(n_0_188), .B1(n_0_189), .B2(n_0_193), .ZN(n_170));
   AOI22_X1 i_0_174 (.A1(n_369), .A2(n_0_138), .B1(n_180), .B2(n_0_137), 
      .ZN(n_0_188));
   INV_X1 i_0_175 (.A(n_379), .ZN(n_0_189));
   OAI21_X1 i_0_176 (.A(n_0_190), .B1(n_0_191), .B2(n_0_193), .ZN(n_171));
   AOI22_X1 i_0_177 (.A1(n_370), .A2(n_0_138), .B1(n_181), .B2(n_0_137), 
      .ZN(n_0_190));
   INV_X1 i_0_178 (.A(n_380), .ZN(n_0_191));
   OAI21_X1 i_0_179 (.A(n_0_192), .B1(n_0_201), .B2(n_0_193), .ZN(n_172));
   AOI22_X1 i_0_182 (.A1(n_371), .A2(n_0_138), .B1(n_182), .B2(n_0_137), 
      .ZN(n_0_192));
   NOR2_X1 i_0_183 (.A1(n_0_139), .A2(n_0_138), .ZN(n_0_137));
   NOR2_X1 i_0_184 (.A1(n_0_176), .A2(A[9]), .ZN(n_0_138));
   INV_X1 i_0_185 (.A(n_0_139), .ZN(n_0_193));
   NOR2_X1 i_0_186 (.A1(n_0_194), .A2(A[8]), .ZN(n_0_139));
   INV_X1 i_0_187 (.A(n_381), .ZN(n_0_201));
   OAI21_X1 i_0_188 (.A(n_0_202), .B1(n_0_203), .B2(n_0_229), .ZN(n_173));
   AOI22_X1 i_0_189 (.A1(n_341), .A2(n_0_158), .B1(n_184), .B2(n_0_157), 
      .ZN(n_0_202));
   INV_X1 i_0_190 (.A(n_352), .ZN(n_0_203));
   OAI21_X1 i_0_191 (.A(n_0_204), .B1(n_0_205), .B2(n_0_209), .ZN(n_174));
   AOI22_X1 i_0_192 (.A1(n_353), .A2(n_0_159), .B1(n_185), .B2(n_0_157), 
      .ZN(n_0_204));
   INV_X1 i_0_193 (.A(n_342), .ZN(n_0_205));
   OAI21_X1 i_0_194 (.A(n_0_206), .B1(n_0_207), .B2(n_0_209), .ZN(n_175));
   AOI22_X1 i_0_195 (.A1(n_354), .A2(n_0_159), .B1(n_186), .B2(n_0_157), 
      .ZN(n_0_206));
   INV_X1 i_0_196 (.A(n_343), .ZN(n_0_207));
   OAI21_X1 i_0_197 (.A(n_0_208), .B1(n_0_210), .B2(n_0_209), .ZN(n_176));
   AOI22_X1 i_0_198 (.A1(n_355), .A2(n_0_159), .B1(n_187), .B2(n_0_157), 
      .ZN(n_0_208));
   INV_X1 i_0_199 (.A(n_0_158), .ZN(n_0_209));
   INV_X1 i_0_200 (.A(n_344), .ZN(n_0_210));
   OAI21_X1 i_0_201 (.A(n_0_211), .B1(n_0_212), .B2(n_0_229), .ZN(n_177));
   AOI22_X1 i_0_202 (.A1(n_345), .A2(n_0_158), .B1(n_188), .B2(n_0_157), 
      .ZN(n_0_211));
   INV_X1 i_0_203 (.A(n_356), .ZN(n_0_212));
   OAI21_X1 i_0_204 (.A(n_0_213), .B1(n_0_221), .B2(n_0_229), .ZN(n_178));
   AOI22_X1 i_0_205 (.A1(n_346), .A2(n_0_158), .B1(n_189), .B2(n_0_157), 
      .ZN(n_0_213));
   INV_X1 i_0_206 (.A(n_357), .ZN(n_0_221));
   OAI21_X1 i_0_207 (.A(n_0_222), .B1(n_0_223), .B2(n_0_229), .ZN(n_179));
   AOI22_X1 i_0_208 (.A1(n_347), .A2(n_0_158), .B1(n_190), .B2(n_0_157), 
      .ZN(n_0_222));
   INV_X1 i_0_209 (.A(n_358), .ZN(n_0_223));
   OAI21_X1 i_0_210 (.A(n_0_224), .B1(n_0_225), .B2(n_0_229), .ZN(n_180));
   AOI22_X1 i_0_211 (.A1(n_348), .A2(n_0_158), .B1(n_191), .B2(n_0_157), 
      .ZN(n_0_224));
   INV_X1 i_0_212 (.A(n_359), .ZN(n_0_225));
   OAI21_X1 i_0_213 (.A(n_0_226), .B1(n_0_227), .B2(n_0_229), .ZN(n_181));
   AOI22_X1 i_0_214 (.A1(n_349), .A2(n_0_158), .B1(n_192), .B2(n_0_157), 
      .ZN(n_0_226));
   INV_X1 i_0_215 (.A(n_360), .ZN(n_0_227));
   OAI21_X1 i_0_218 (.A(n_0_228), .B1(n_0_232), .B2(n_0_229), .ZN(n_182));
   AOI22_X1 i_0_219 (.A1(n_350), .A2(n_0_158), .B1(n_193), .B2(n_0_157), 
      .ZN(n_0_228));
   NOR2_X1 i_0_220 (.A1(n_0_159), .A2(n_0_158), .ZN(n_0_157));
   NOR2_X1 i_0_221 (.A1(A[8]), .A2(n_0_175), .ZN(n_0_158));
   INV_X1 i_0_222 (.A(n_0_159), .ZN(n_0_229));
   NOR2_X1 i_0_223 (.A1(n_0_176), .A2(A[7]), .ZN(n_0_159));
   INV_X1 i_0_224 (.A(n_361), .ZN(n_0_232));
   OAI21_X1 i_0_225 (.A(n_0_233), .B1(n_0_236), .B2(n_0_257), .ZN(n_183));
   AOI22_X1 i_0_226 (.A1(n_317), .A2(n_0_178), .B1(n_0_177), .B2(n_195), 
      .ZN(n_0_233));
   INV_X1 i_0_227 (.A(n_329), .ZN(n_0_236));
   OAI21_X1 i_0_228 (.A(n_0_237), .B1(n_0_238), .B2(n_0_246), .ZN(n_184));
   AOI22_X1 i_0_229 (.A1(n_330), .A2(n_0_179), .B1(n_0_177), .B2(n_196), 
      .ZN(n_0_237));
   INV_X1 i_0_230 (.A(n_318), .ZN(n_0_238));
   OAI21_X1 i_0_231 (.A(n_0_239), .B1(n_0_240), .B2(n_0_246), .ZN(n_185));
   AOI22_X1 i_0_232 (.A1(n_331), .A2(n_0_179), .B1(n_0_177), .B2(n_197), 
      .ZN(n_0_239));
   INV_X1 i_0_233 (.A(n_319), .ZN(n_0_240));
   OAI21_X1 i_0_234 (.A(n_0_241), .B1(n_0_242), .B2(n_0_246), .ZN(n_186));
   AOI22_X1 i_0_235 (.A1(n_332), .A2(n_0_179), .B1(n_0_177), .B2(n_198), 
      .ZN(n_0_241));
   INV_X1 i_0_236 (.A(n_320), .ZN(n_0_242));
   OAI21_X1 i_0_237 (.A(n_0_243), .B1(n_0_244), .B2(n_0_246), .ZN(n_187));
   AOI22_X1 i_0_238 (.A1(n_333), .A2(n_0_179), .B1(n_0_177), .B2(n_199), 
      .ZN(n_0_243));
   INV_X1 i_0_239 (.A(n_321), .ZN(n_0_244));
   OAI21_X1 i_0_240 (.A(n_0_245), .B1(n_0_247), .B2(n_0_246), .ZN(n_188));
   AOI22_X1 i_0_241 (.A1(n_334), .A2(n_0_179), .B1(n_0_177), .B2(n_200), 
      .ZN(n_0_245));
   INV_X1 i_0_242 (.A(n_0_178), .ZN(n_0_246));
   INV_X1 i_0_243 (.A(n_322), .ZN(n_0_247));
   OAI21_X1 i_0_244 (.A(n_0_248), .B1(n_0_249), .B2(n_0_257), .ZN(n_189));
   AOI22_X1 i_0_245 (.A1(n_323), .A2(n_0_178), .B1(n_0_177), .B2(n_201), 
      .ZN(n_0_248));
   INV_X1 i_0_246 (.A(n_335), .ZN(n_0_249));
   OAI21_X1 i_0_247 (.A(n_0_250), .B1(n_0_251), .B2(n_0_257), .ZN(n_190));
   AOI22_X1 i_0_248 (.A1(n_324), .A2(n_0_178), .B1(n_0_177), .B2(n_202), 
      .ZN(n_0_250));
   INV_X1 i_0_249 (.A(n_336), .ZN(n_0_251));
   OAI21_X1 i_0_250 (.A(n_0_252), .B1(n_0_253), .B2(n_0_257), .ZN(n_191));
   AOI22_X1 i_0_251 (.A1(n_325), .A2(n_0_178), .B1(n_0_177), .B2(n_203), 
      .ZN(n_0_252));
   INV_X1 i_0_254 (.A(n_337), .ZN(n_0_253));
   OAI21_X1 i_0_255 (.A(n_0_254), .B1(n_0_255), .B2(n_0_257), .ZN(n_192));
   AOI22_X1 i_0_256 (.A1(n_326), .A2(n_0_178), .B1(n_0_177), .B2(n_204), 
      .ZN(n_0_254));
   INV_X1 i_0_257 (.A(n_338), .ZN(n_0_255));
   OAI21_X1 i_0_258 (.A(n_0_256), .B1(n_0_258), .B2(n_0_257), .ZN(n_193));
   AOI22_X1 i_0_259 (.A1(n_327), .A2(n_0_178), .B1(n_0_177), .B2(n_205), 
      .ZN(n_0_256));
   NOR2_X1 i_0_260 (.A1(n_0_174), .A2(A[7]), .ZN(n_0_178));
   INV_X1 i_0_261 (.A(n_0_32), .ZN(n_0_177));
   INV_X1 i_0_262 (.A(n_0_179), .ZN(n_0_257));
   NOR2_X1 i_0_263 (.A1(n_0_175), .A2(A[6]), .ZN(n_0_179));
   INV_X1 i_0_264 (.A(n_339), .ZN(n_0_258));
   OAI21_X1 i_0_265 (.A(n_0_259), .B1(n_0_260), .B2(n_0_283), .ZN(n_194));
   AOI22_X1 i_0_266 (.A1(n_291), .A2(n_0_198), .B1(n_207), .B2(n_0_197), 
      .ZN(n_0_259));
   INV_X1 i_0_267 (.A(n_304), .ZN(n_0_260));
   OAI21_X1 i_0_268 (.A(n_0_261), .B1(n_0_262), .B2(n_0_272), .ZN(n_195));
   AOI22_X1 i_0_269 (.A1(n_305), .A2(n_0_199), .B1(n_208), .B2(n_0_197), 
      .ZN(n_0_261));
   INV_X1 i_0_270 (.A(n_292), .ZN(n_0_262));
   OAI21_X1 i_0_271 (.A(n_0_263), .B1(n_0_264), .B2(n_0_272), .ZN(n_196));
   AOI22_X1 i_0_272 (.A1(n_306), .A2(n_0_199), .B1(n_209), .B2(n_0_197), 
      .ZN(n_0_263));
   INV_X1 i_0_273 (.A(n_293), .ZN(n_0_264));
   OAI21_X1 i_0_274 (.A(n_0_265), .B1(n_0_266), .B2(n_0_272), .ZN(n_197));
   AOI22_X1 i_0_275 (.A1(n_307), .A2(n_0_199), .B1(n_210), .B2(n_0_197), 
      .ZN(n_0_265));
   INV_X1 i_0_276 (.A(n_294), .ZN(n_0_266));
   OAI21_X1 i_0_277 (.A(n_0_267), .B1(n_0_268), .B2(n_0_272), .ZN(n_198));
   AOI22_X1 i_0_278 (.A1(n_308), .A2(n_0_199), .B1(n_211), .B2(n_0_197), 
      .ZN(n_0_267));
   INV_X1 i_0_279 (.A(n_295), .ZN(n_0_268));
   OAI21_X1 i_0_280 (.A(n_0_269), .B1(n_0_270), .B2(n_0_272), .ZN(n_199));
   AOI22_X1 i_0_281 (.A1(n_309), .A2(n_0_199), .B1(n_212), .B2(n_0_197), 
      .ZN(n_0_269));
   INV_X1 i_0_282 (.A(n_296), .ZN(n_0_270));
   OAI21_X1 i_0_283 (.A(n_0_271), .B1(n_0_273), .B2(n_0_272), .ZN(n_200));
   AOI22_X1 i_0_284 (.A1(n_310), .A2(n_0_199), .B1(n_213), .B2(n_0_197), 
      .ZN(n_0_271));
   INV_X1 i_0_285 (.A(n_0_198), .ZN(n_0_272));
   INV_X1 i_0_286 (.A(n_297), .ZN(n_0_273));
   OAI21_X1 i_0_287 (.A(n_0_274), .B1(n_0_275), .B2(n_0_283), .ZN(n_201));
   AOI22_X1 i_0_290 (.A1(n_298), .A2(n_0_198), .B1(n_214), .B2(n_0_197), 
      .ZN(n_0_274));
   INV_X1 i_0_291 (.A(n_311), .ZN(n_0_275));
   OAI21_X1 i_0_292 (.A(n_0_276), .B1(n_0_277), .B2(n_0_283), .ZN(n_202));
   AOI22_X1 i_0_293 (.A1(n_299), .A2(n_0_198), .B1(n_215), .B2(n_0_197), 
      .ZN(n_0_276));
   INV_X1 i_0_294 (.A(n_312), .ZN(n_0_277));
   OAI21_X1 i_0_295 (.A(n_0_278), .B1(n_0_279), .B2(n_0_283), .ZN(n_203));
   AOI22_X1 i_0_296 (.A1(n_300), .A2(n_0_198), .B1(n_216), .B2(n_0_197), 
      .ZN(n_0_278));
   INV_X1 i_0_297 (.A(n_313), .ZN(n_0_279));
   OAI21_X1 i_0_298 (.A(n_0_280), .B1(n_0_281), .B2(n_0_283), .ZN(n_204));
   AOI22_X1 i_0_299 (.A1(n_301), .A2(n_0_198), .B1(n_217), .B2(n_0_197), 
      .ZN(n_0_280));
   INV_X1 i_0_300 (.A(n_314), .ZN(n_0_281));
   OAI21_X1 i_0_301 (.A(n_0_282), .B1(n_0_284), .B2(n_0_283), .ZN(n_205));
   AOI22_X1 i_0_302 (.A1(n_302), .A2(n_0_198), .B1(n_218), .B2(n_0_197), 
      .ZN(n_0_282));
   NOR2_X1 i_0_303 (.A1(n_0_199), .A2(n_0_198), .ZN(n_0_197));
   NOR2_X1 i_0_304 (.A1(A[6]), .A2(n_0_173), .ZN(n_0_198));
   INV_X1 i_0_305 (.A(n_0_199), .ZN(n_0_283));
   NOR2_X1 i_0_306 (.A1(n_0_174), .A2(A[5]), .ZN(n_0_199));
   INV_X1 i_0_307 (.A(n_315), .ZN(n_0_284));
   OAI21_X1 i_0_308 (.A(n_0_285), .B1(n_0_286), .B2(n_0_312), .ZN(n_206));
   AOI22_X1 i_0_309 (.A1(n_265), .A2(n_0_218), .B1(n_219), .B2(n_0_217), 
      .ZN(n_0_285));
   INV_X1 i_0_310 (.A(n_278), .ZN(n_0_286));
   OAI21_X1 i_0_311 (.A(n_0_287), .B1(n_0_288), .B2(n_0_311), .ZN(n_207));
   AOI22_X1 i_0_312 (.A1(n_279), .A2(n_0_219), .B1(n_220), .B2(n_0_217), 
      .ZN(n_0_287));
   INV_X1 i_0_313 (.A(n_266), .ZN(n_0_288));
   OAI21_X1 i_0_314 (.A(n_0_289), .B1(n_0_290), .B2(n_0_311), .ZN(n_208));
   AOI22_X1 i_0_315 (.A1(n_280), .A2(n_0_219), .B1(n_221), .B2(n_0_217), 
      .ZN(n_0_289));
   INV_X1 i_0_316 (.A(n_267), .ZN(n_0_290));
   OAI21_X1 i_0_317 (.A(n_0_291), .B1(n_0_292), .B2(n_0_311), .ZN(n_209));
   AOI22_X1 i_0_318 (.A1(n_281), .A2(n_0_219), .B1(n_222), .B2(n_0_217), 
      .ZN(n_0_291));
   INV_X1 i_0_319 (.A(n_268), .ZN(n_0_292));
   OAI21_X1 i_0_320 (.A(n_0_293), .B1(n_0_294), .B2(n_0_311), .ZN(n_210));
   AOI22_X1 i_0_321 (.A1(n_282), .A2(n_0_219), .B1(n_223), .B2(n_0_217), 
      .ZN(n_0_293));
   INV_X1 i_0_322 (.A(n_269), .ZN(n_0_294));
   OAI21_X1 i_0_323 (.A(n_0_295), .B1(n_0_296), .B2(n_0_311), .ZN(n_211));
   AOI22_X1 i_0_326 (.A1(n_283), .A2(n_0_219), .B1(n_224), .B2(n_0_217), 
      .ZN(n_0_295));
   INV_X1 i_0_327 (.A(n_270), .ZN(n_0_296));
   OAI21_X1 i_0_328 (.A(n_0_297), .B1(n_0_298), .B2(n_0_311), .ZN(n_212));
   AOI22_X1 i_0_329 (.A1(n_284), .A2(n_0_219), .B1(n_225), .B2(n_0_217), 
      .ZN(n_0_297));
   INV_X1 i_0_330 (.A(n_271), .ZN(n_0_298));
   OAI21_X1 i_0_331 (.A(n_0_299), .B1(n_0_300), .B2(n_0_311), .ZN(n_213));
   AOI22_X1 i_0_332 (.A1(n_285), .A2(n_0_219), .B1(n_226), .B2(n_0_217), 
      .ZN(n_0_299));
   INV_X1 i_0_333 (.A(n_272), .ZN(n_0_300));
   OAI21_X1 i_0_334 (.A(n_0_301), .B1(n_0_302), .B2(n_0_312), .ZN(n_214));
   AOI22_X1 i_0_335 (.A1(n_273), .A2(n_0_218), .B1(n_135), .B2(n_0_217), 
      .ZN(n_0_301));
   INV_X1 i_0_336 (.A(n_286), .ZN(n_0_302));
   OAI21_X1 i_0_337 (.A(n_0_303), .B1(n_0_304), .B2(n_0_312), .ZN(n_215));
   AOI22_X1 i_0_338 (.A1(n_274), .A2(n_0_218), .B1(n_136), .B2(n_0_217), 
      .ZN(n_0_303));
   INV_X1 i_0_339 (.A(n_287), .ZN(n_0_304));
   OAI21_X1 i_0_340 (.A(n_0_305), .B1(n_0_306), .B2(n_0_312), .ZN(n_216));
   AOI22_X1 i_0_341 (.A1(n_275), .A2(n_0_218), .B1(n_227), .B2(n_0_217), 
      .ZN(n_0_305));
   INV_X1 i_0_342 (.A(n_288), .ZN(n_0_306));
   OAI21_X1 i_0_343 (.A(n_0_307), .B1(n_0_308), .B2(n_0_312), .ZN(n_217));
   AOI22_X1 i_0_344 (.A1(n_276), .A2(n_0_218), .B1(n_228), .B2(n_0_217), 
      .ZN(n_0_307));
   INV_X1 i_0_345 (.A(n_289), .ZN(n_0_308));
   OAI21_X1 i_0_346 (.A(n_0_309), .B1(n_0_313), .B2(n_0_312), .ZN(n_218));
   AOI22_X1 i_0_347 (.A1(n_277), .A2(n_0_218), .B1(n_137), .B2(n_0_217), 
      .ZN(n_0_309));
   INV_X1 i_0_348 (.A(n_0_310), .ZN(n_0_217));
   NAND2_X1 i_0_349 (.A1(n_0_312), .A2(n_0_311), .ZN(n_0_310));
   INV_X1 i_0_350 (.A(n_0_218), .ZN(n_0_311));
   NOR2_X1 i_0_351 (.A1(n_0_156), .A2(A[5]), .ZN(n_0_218));
   INV_X1 i_0_352 (.A(n_0_219), .ZN(n_0_312));
   NOR2_X1 i_0_353 (.A1(n_0_173), .A2(A[4]), .ZN(n_0_219));
   INV_X1 i_0_354 (.A(n_290), .ZN(n_0_313));
   OAI211_X1 i_0_355 (.A(n_0_314), .B(n_0_315), .C1(n_0_51), .C2(n_0_316), 
      .ZN(n_219));
   NAND2_X1 i_0_356 (.A1(n_82), .A2(n_0_2), .ZN(n_0_314));
   NAND2_X1 i_0_357 (.A1(n_98), .A2(n_0_3), .ZN(n_0_315));
   INV_X1 i_0_358 (.A(n_229), .ZN(n_0_316));
   NAND2_X1 i_0_359 (.A1(n_0_48), .A2(n_0_49), .ZN(n_220));
   OAI21_X1 i_0_362 (.A(n_0_317), .B1(n_0_318), .B2(n_0_332), .ZN(n_221));
   AOI22_X1 i_0_363 (.A1(n_84), .A2(n_0_2), .B1(n_0_1), .B2(n_230), .ZN(n_0_317));
   INV_X1 i_0_364 (.A(n_100), .ZN(n_0_318));
   OAI21_X1 i_0_365 (.A(n_0_319), .B1(n_0_320), .B2(n_0_332), .ZN(n_222));
   AOI22_X1 i_0_366 (.A1(n_85), .A2(n_0_2), .B1(n_0_1), .B2(n_231), .ZN(n_0_319));
   INV_X1 i_0_367 (.A(n_101), .ZN(n_0_320));
   OAI21_X1 i_0_368 (.A(n_0_321), .B1(n_0_322), .B2(n_0_332), .ZN(n_223));
   AOI22_X1 i_0_369 (.A1(n_86), .A2(n_0_2), .B1(n_0_1), .B2(n_232), .ZN(n_0_321));
   INV_X1 i_0_370 (.A(n_102), .ZN(n_0_322));
   OAI21_X1 i_0_371 (.A(n_0_323), .B1(n_0_324), .B2(n_0_332), .ZN(n_224));
   AOI22_X1 i_0_372 (.A1(n_87), .A2(n_0_2), .B1(n_0_1), .B2(n_233), .ZN(n_0_323));
   INV_X1 i_0_373 (.A(n_103), .ZN(n_0_324));
   OAI21_X1 i_0_374 (.A(n_0_325), .B1(n_0_326), .B2(n_0_332), .ZN(n_225));
   AOI22_X1 i_0_375 (.A1(n_88), .A2(n_0_2), .B1(n_234), .B2(n_0_1), .ZN(n_0_325));
   INV_X1 i_0_376 (.A(n_104), .ZN(n_0_326));
   OAI21_X1 i_0_377 (.A(n_0_327), .B1(n_0_328), .B2(n_0_332), .ZN(n_226));
   AOI22_X1 i_0_378 (.A1(n_89), .A2(n_0_2), .B1(n_235), .B2(n_0_1), .ZN(n_0_327));
   INV_X1 i_0_379 (.A(n_105), .ZN(n_0_328));
   OAI21_X1 i_0_380 (.A(n_0_329), .B1(n_0_330), .B2(n_0_332), .ZN(n_227));
   AOI22_X1 i_0_381 (.A1(n_92), .A2(n_0_2), .B1(n_237), .B2(n_0_1), .ZN(n_0_329));
   INV_X1 i_0_382 (.A(n_108), .ZN(n_0_330));
   OAI21_X1 i_0_383 (.A(n_0_331), .B1(n_0_333), .B2(n_0_332), .ZN(n_228));
   AOI22_X1 i_0_384 (.A1(n_93), .A2(n_0_2), .B1(n_238), .B2(n_0_1), .ZN(n_0_331));
   INV_X1 i_0_385 (.A(n_0_52), .ZN(n_0_2));
   INV_X1 i_0_386 (.A(n_0_51), .ZN(n_0_1));
   INV_X1 i_0_387 (.A(n_0_3), .ZN(n_0_332));
   NOR2_X1 i_0_388 (.A1(n_0_156), .A2(A[3]), .ZN(n_0_3));
   INV_X1 i_0_390 (.A(n_109), .ZN(n_0_333));
   NAND2_X1 i_0_391 (.A1(n_0_334), .A2(n_0_335), .ZN(n_229));
   AOI22_X1 i_0_393 (.A1(n_51), .A2(n_0_22), .B1(n_240), .B2(n_0_21), .ZN(
      n_0_334));
   NAND2_X1 i_0_394 (.A1(n_67), .A2(n_0_23), .ZN(n_0_335));
   OAI21_X1 i_0_395 (.A(n_0_336), .B1(n_0_337), .B2(n_0_346), .ZN(n_230));
   AOI22_X1 i_0_398 (.A1(n_69), .A2(n_0_23), .B1(n_241), .B2(n_0_21), .ZN(
      n_0_336));
   INV_X1 i_0_399 (.A(n_53), .ZN(n_0_337));
   OAI21_X1 i_0_400 (.A(n_0_338), .B1(n_0_339), .B2(n_0_347), .ZN(n_231));
   AOI22_X1 i_0_401 (.A1(n_54), .A2(n_0_22), .B1(n_242), .B2(n_0_21), .ZN(
      n_0_338));
   INV_X1 i_0_402 (.A(n_70), .ZN(n_0_339));
   NAND2_X1 i_0_403 (.A1(n_0_340), .A2(n_0_341), .ZN(n_232));
   AOI22_X1 i_0_404 (.A1(n_55), .A2(n_0_22), .B1(n_243), .B2(n_0_21), .ZN(
      n_0_340));
   NAND2_X1 i_0_405 (.A1(n_71), .A2(n_0_23), .ZN(n_0_341));
   OAI21_X1 i_0_406 (.A(n_0_342), .B1(n_0_343), .B2(n_0_346), .ZN(n_233));
   AOI22_X1 i_0_407 (.A1(n_72), .A2(n_0_23), .B1(n_244), .B2(n_0_21), .ZN(
      n_0_342));
   INV_X1 i_0_408 (.A(n_56), .ZN(n_0_343));
   INV_X1 i_0_409 (.A(n_0_13), .ZN(n_234));
   INV_X1 i_0_410 (.A(n_0_14), .ZN(n_235));
   OAI21_X1 i_0_411 (.A(n_0_344), .B1(n_0_348), .B2(n_0_347), .ZN(n_236));
   AOI22_X1 i_0_412 (.A1(n_60), .A2(n_0_22), .B1(n_246), .B2(n_0_21), .ZN(
      n_0_344));
   INV_X1 i_0_413 (.A(n_0_345), .ZN(n_0_21));
   NAND2_X1 i_0_414 (.A1(n_0_347), .A2(n_0_346), .ZN(n_0_345));
   INV_X1 i_0_415 (.A(n_0_22), .ZN(n_0_346));
   NOR2_X1 i_0_416 (.A1(A[3]), .A2(n_0_154), .ZN(n_0_22));
   INV_X1 i_0_418 (.A(n_0_23), .ZN(n_0_347));
   NOR2_X1 i_0_420 (.A1(n_0_155), .A2(A[2]), .ZN(n_0_23));
   INV_X1 i_0_421 (.A(n_76), .ZN(n_0_348));
   INV_X1 i_0_422 (.A(n_0_17), .ZN(n_237));
   INV_X1 i_0_423 (.A(n_0_18), .ZN(n_238));
   OAI21_X1 i_0_424 (.A(n_0_349), .B1(n_0_350), .B2(n_0_363), .ZN(n_239));
   AOI22_X1 i_0_429 (.A1(n_35), .A2(n_0_43), .B1(n_247), .B2(n_0_41), .ZN(
      n_0_349));
   INV_X1 i_0_430 (.A(n_19), .ZN(n_0_350));
   OAI21_X1 i_0_431 (.A(n_0_351), .B1(n_0_352), .B2(n_0_360), .ZN(n_240));
   AOI22_X1 i_0_436 (.A1(n_20), .A2(n_0_42), .B1(n_248), .B2(n_0_41), .ZN(
      n_0_351));
   INV_X1 i_0_437 (.A(n_36), .ZN(n_0_352));
   OAI21_X1 i_0_438 (.A(n_0_353), .B1(n_0_354), .B2(n_0_360), .ZN(n_241));
   AOI22_X1 i_0_439 (.A1(n_22), .A2(n_0_42), .B1(n_249), .B2(n_0_41), .ZN(
      n_0_353));
   INV_X1 i_0_440 (.A(n_38), .ZN(n_0_354));
   OAI21_X1 i_0_441 (.A(n_0_355), .B1(n_0_356), .B2(n_0_360), .ZN(n_242));
   AOI22_X1 i_0_442 (.A1(n_23), .A2(n_0_42), .B1(n_250), .B2(n_0_41), .ZN(
      n_0_355));
   INV_X1 i_0_443 (.A(n_39), .ZN(n_0_356));
   OAI21_X1 i_0_444 (.A(n_0_357), .B1(n_0_358), .B2(n_0_360), .ZN(n_243));
   AOI22_X1 i_0_445 (.A1(n_24), .A2(n_0_42), .B1(n_251), .B2(n_0_41), .ZN(
      n_0_357));
   INV_X1 i_0_446 (.A(n_40), .ZN(n_0_358));
   OAI21_X1 i_0_447 (.A(n_0_359), .B1(n_0_361), .B2(n_0_360), .ZN(n_244));
   AOI22_X1 i_0_448 (.A1(n_25), .A2(n_0_42), .B1(n_252), .B2(n_0_41), .ZN(
      n_0_359));
   INV_X1 i_0_449 (.A(n_0_43), .ZN(n_0_360));
   INV_X1 i_0_450 (.A(n_41), .ZN(n_0_361));
   OAI21_X1 i_0_452 (.A(n_0_362), .B1(n_0_364), .B2(n_0_363), .ZN(n_245));
   AOI22_X1 i_0_456 (.A1(n_44), .A2(n_0_43), .B1(n_254), .B2(n_0_41), .ZN(
      n_0_362));
   NOR2_X1 i_0_457 (.A1(n_0_43), .A2(n_0_42), .ZN(n_0_41));
   NOR2_X1 i_0_458 (.A1(n_0_154), .A2(A[1]), .ZN(n_0_43));
   INV_X1 i_0_460 (.A(n_0_42), .ZN(n_0_363));
   NOR2_X1 i_0_465 (.A1(A[2]), .A2(n_0_153), .ZN(n_0_42));
   INV_X1 i_0_466 (.A(n_28), .ZN(n_0_364));
   INV_X1 i_0_467 (.A(n_0_37), .ZN(n_246));
   OAI211_X1 i_0_472 (.A(n_0_366), .B(n_0_365), .C1(n_0_378), .C2(n_0_375), 
      .ZN(n_247));
   NAND2_X1 i_0_473 (.A1(n_0_68), .A2(n_256), .ZN(n_0_365));
   NAND2_X1 i_0_474 (.A1(n_4), .A2(n_0_70), .ZN(n_0_366));
   OAI211_X1 i_0_475 (.A(n_0_368), .B(n_0_367), .C1(n_0_102), .C2(n_0_380), 
      .ZN(n_248));
   NAND2_X1 i_0_476 (.A1(n_0_59), .A2(n_256), .ZN(n_0_367));
   NAND2_X1 i_0_477 (.A1(n_5), .A2(n_0_70), .ZN(n_0_368));
   OAI221_X1 i_0_478 (.A(n_0_369), .B1(n_0_102), .B2(n_0_371), .C1(n_0_382), 
      .C2(n_0_375), .ZN(n_249));
   NAND2_X1 i_0_479 (.A1(n_7), .A2(n_0_70), .ZN(n_0_369));
   OAI221_X1 i_0_480 (.A(n_0_370), .B1(n_0_102), .B2(n_0_385), .C1(n_0_371), 
      .C2(n_0_375), .ZN(n_250));
   NAND2_X1 i_0_481 (.A1(n_8), .A2(n_0_70), .ZN(n_0_370));
   INV_X1 i_0_482 (.A(n_259), .ZN(n_0_371));
   OAI221_X1 i_0_483 (.A(n_0_372), .B1(n_0_102), .B2(n_0_387), .C1(n_0_385), 
      .C2(n_0_375), .ZN(n_251));
   NAND2_X1 i_0_484 (.A1(n_9), .A2(n_0_70), .ZN(n_0_372));
   OAI211_X1 i_0_485 (.A(n_0_374), .B(n_0_373), .C1(n_0_387), .C2(n_0_375), 
      .ZN(n_252));
   NAND2_X1 i_0_486 (.A1(n_0_68), .A2(n_262), .ZN(n_0_373));
   NAND2_X1 i_0_487 (.A1(n_10), .A2(n_0_70), .ZN(n_0_374));
   INV_X1 i_0_492 (.A(n_0_59), .ZN(n_0_375));
   NAND2_X1 i_0_493 (.A1(n_0_377), .A2(n_0_376), .ZN(n_253));
   AOI22_X1 i_0_494 (.A1(n_264), .A2(n_0_68), .B1(n_263), .B2(n_0_59), .ZN(
      n_0_376));
   NOR2_X1 i_0_501 (.A1(n_0_153), .A2(A[0]), .ZN(n_0_59));
   INV_X1 i_0_502 (.A(n_0_102), .ZN(n_0_68));
   NAND2_X1 i_0_503 (.A1(n_12), .A2(n_0_70), .ZN(n_0_377));
   NOR2_X1 i_0_506 (.A1(A[1]), .A2(n_0_104), .ZN(n_0_70));
   INV_X1 i_0_507 (.A(n_0_57), .ZN(n_254));
   INV_X1 i_0_508 (.A(n_0_378), .ZN(n_255));
   NAND2_X1 i_0_509 (.A1(n_0_403), .A2(n_0_379), .ZN(n_0_378));
   NAND2_X1 i_0_510 (.A1(n_0_404), .A2(B[4]), .ZN(n_0_379));
   XNOR2_X1 i_0_511 (.A(n_0_403), .B(n_0_410), .ZN(n_256));
   INV_X1 i_0_512 (.A(n_0_380), .ZN(n_257));
   NAND2_X1 i_0_513 (.A1(n_0_399), .A2(n_0_381), .ZN(n_0_380));
   NAND2_X1 i_0_514 (.A1(n_0_401), .A2(B[6]), .ZN(n_0_381));
   INV_X1 i_0_515 (.A(n_0_382), .ZN(n_258));
   NAND2_X1 i_0_516 (.A1(n_0_397), .A2(n_0_383), .ZN(n_0_382));
   NAND2_X1 i_0_518 (.A1(n_0_399), .A2(B[7]), .ZN(n_0_383));
   AND2_X1 i_0_519 (.A1(n_0_395), .A2(n_0_384), .ZN(n_259));
   NAND2_X1 i_0_520 (.A1(n_0_397), .A2(B[8]), .ZN(n_0_384));
   INV_X1 i_0_521 (.A(n_0_385), .ZN(n_260));
   NAND2_X1 i_0_522 (.A1(n_0_393), .A2(n_0_386), .ZN(n_0_385));
   NAND2_X1 i_0_523 (.A1(n_0_395), .A2(B[9]), .ZN(n_0_386));
   INV_X1 i_0_524 (.A(n_0_387), .ZN(n_261));
   NAND2_X1 i_0_525 (.A1(n_0_389), .A2(n_0_388), .ZN(n_0_387));
   NAND2_X1 i_0_528 (.A1(n_0_393), .A2(B[10]), .ZN(n_0_388));
   XNOR2_X1 i_0_529 (.A(n_0_389), .B(n_0_416), .ZN(n_262));
   NAND2_X1 i_0_530 (.A1(n_0_392), .A2(n_0_415), .ZN(n_0_389));
   INV_X1 i_0_534 (.A(n_0_390), .ZN(n_263));
   XNOR2_X1 i_0_535 (.A(n_0_391), .B(B[15]), .ZN(n_0_390));
   NAND3_X1 i_0_538 (.A1(n_0_392), .A2(n_0_416), .A3(n_0_415), .ZN(n_0_391));
   INV_X1 i_0_541 (.A(n_0_393), .ZN(n_0_392));
   NAND2_X1 i_0_542 (.A1(n_0_394), .A2(n_0_414), .ZN(n_0_393));
   INV_X1 i_0_543 (.A(n_0_395), .ZN(n_0_394));
   NAND2_X1 i_0_544 (.A1(n_0_396), .A2(n_0_413), .ZN(n_0_395));
   INV_X1 i_0_545 (.A(n_0_397), .ZN(n_0_396));
   NAND2_X1 i_0_546 (.A1(n_0_398), .A2(n_0_412), .ZN(n_0_397));
   INV_X1 i_0_547 (.A(n_0_399), .ZN(n_0_398));
   NAND2_X1 i_0_548 (.A1(n_0_400), .A2(n_0_411), .ZN(n_0_399));
   INV_X1 i_0_549 (.A(n_0_401), .ZN(n_0_400));
   NAND2_X1 i_0_550 (.A1(n_0_402), .A2(n_0_410), .ZN(n_0_401));
   INV_X1 i_0_551 (.A(n_0_403), .ZN(n_0_402));
   NAND2_X1 i_0_552 (.A1(n_0_132), .A2(n_0_409), .ZN(n_0_403));
   INV_X1 i_0_553 (.A(n_0_404), .ZN(n_0_132));
   NAND2_X1 i_0_560 (.A1(n_0_134), .A2(n_0_408), .ZN(n_0_404));
   INV_X1 i_0_561 (.A(n_0_133), .ZN(n_0_134));
   NAND2_X1 i_0_562 (.A1(n_0_136), .A2(n_0_407), .ZN(n_0_133));
   INV_X1 i_0_563 (.A(n_0_135), .ZN(n_0_136));
   NAND2_X1 i_0_564 (.A1(n_0_406), .A2(n_0_405), .ZN(n_0_135));
   INV_X1 i_0_565 (.A(B[0]), .ZN(n_0_405));
   INV_X1 i_0_566 (.A(B[1]), .ZN(n_0_406));
   INV_X1 i_0_567 (.A(B[2]), .ZN(n_0_407));
   INV_X1 i_0_568 (.A(B[3]), .ZN(n_0_408));
   INV_X1 i_0_569 (.A(B[4]), .ZN(n_0_409));
   INV_X1 i_0_570 (.A(B[5]), .ZN(n_0_410));
   INV_X1 i_0_571 (.A(B[6]), .ZN(n_0_411));
   INV_X1 i_0_572 (.A(B[7]), .ZN(n_0_412));
   INV_X1 i_0_573 (.A(B[8]), .ZN(n_0_413));
   INV_X1 i_0_574 (.A(B[9]), .ZN(n_0_414));
   INV_X1 i_0_575 (.A(B[10]), .ZN(n_0_415));
   INV_X1 i_0_576 (.A(B[11]), .ZN(n_0_416));
   AOI21_X1 i_0_577 (.A(n_0_73), .B1(B[15]), .B2(n_0_74), .ZN(n_264));
   FA_X1 i_1_0 (.A(B[1]), .B(n_219), .CI(n_1_166), .CO(n_1_2), .S(n_265));
   FA_X1 i_1_1 (.A(B[2]), .B(n_220), .CI(n_1_2), .CO(n_1_3), .S(n_266));
   FA_X1 i_1_2 (.A(B[3]), .B(n_221), .CI(n_1_3), .CO(n_1_4), .S(n_267));
   FA_X1 i_1_3 (.A(B[4]), .B(n_222), .CI(n_1_4), .CO(n_1_5), .S(n_268));
   FA_X1 i_1_4 (.A(B[5]), .B(n_223), .CI(n_1_5), .CO(n_1_6), .S(n_269));
   FA_X1 i_1_5 (.A(B[6]), .B(n_224), .CI(n_1_6), .CO(n_1_7), .S(n_270));
   FA_X1 i_1_6 (.A(B[7]), .B(n_225), .CI(n_1_7), .CO(n_1_8), .S(n_271));
   FA_X1 i_1_7 (.A(B[8]), .B(n_226), .CI(n_1_8), .CO(n_1_9), .S(n_272));
   FA_X1 i_1_8 (.A(B[9]), .B(n_135), .CI(n_1_9), .CO(n_1_10), .S(n_273));
   FA_X1 i_1_9 (.A(B[10]), .B(n_136), .CI(n_1_10), .CO(n_1_11), .S(n_274));
   FA_X1 i_1_10 (.A(B[11]), .B(n_227), .CI(n_1_11), .CO(n_1_12), .S(n_275));
   FA_X1 i_1_11 (.A(B[15]), .B(n_228), .CI(n_1_12), .CO(n_1_13), .S(n_276));
   FA_X1 i_1_12 (.A(B[15]), .B(n_137), .CI(n_1_13), .CO(n_1_14), .S(n_277));
   FA_X1 i_1_13 (.A(n_146), .B(n_219), .CI(n_1_166), .CO(n_1_0), .S(n_278));
   FA_X1 i_1_14 (.A(n_147), .B(n_220), .CI(n_1_0), .CO(n_1_1), .S(n_279));
   FA_X1 i_1_15 (.A(n_148), .B(n_221), .CI(n_1_1), .CO(n_1_15), .S(n_280));
   FA_X1 i_1_16 (.A(n_255), .B(n_222), .CI(n_1_15), .CO(n_1_16), .S(n_281));
   FA_X1 i_1_17 (.A(n_256), .B(n_223), .CI(n_1_16), .CO(n_1_17), .S(n_282));
   FA_X1 i_1_18 (.A(n_257), .B(n_224), .CI(n_1_17), .CO(n_1_18), .S(n_283));
   FA_X1 i_1_19 (.A(n_258), .B(n_225), .CI(n_1_18), .CO(n_1_19), .S(n_284));
   FA_X1 i_1_20 (.A(n_259), .B(n_226), .CI(n_1_19), .CO(n_1_20), .S(n_285));
   FA_X1 i_1_21 (.A(n_260), .B(n_135), .CI(n_1_20), .CO(n_1_21), .S(n_286));
   FA_X1 i_1_22 (.A(n_261), .B(n_136), .CI(n_1_21), .CO(n_1_22), .S(n_287));
   FA_X1 i_1_23 (.A(n_262), .B(n_227), .CI(n_1_22), .CO(n_1_23), .S(n_288));
   FA_X1 i_1_24 (.A(n_263), .B(n_228), .CI(n_1_23), .CO(n_1_24), .S(n_289));
   FA_X1 i_1_25 (.A(n_264), .B(n_137), .CI(n_1_24), .CO(n_1_25), .S(n_290));
   FA_X1 i_1_26 (.A(B[1]), .B(n_207), .CI(n_1_167), .CO(n_1_26), .S(n_291));
   FA_X1 i_1_27 (.A(B[2]), .B(n_208), .CI(n_1_26), .CO(n_1_27), .S(n_292));
   FA_X1 i_1_28 (.A(B[3]), .B(n_209), .CI(n_1_27), .CO(n_1_28), .S(n_293));
   FA_X1 i_1_29 (.A(B[4]), .B(n_210), .CI(n_1_28), .CO(n_1_29), .S(n_294));
   FA_X1 i_1_30 (.A(B[5]), .B(n_211), .CI(n_1_29), .CO(n_1_30), .S(n_295));
   FA_X1 i_1_31 (.A(B[6]), .B(n_212), .CI(n_1_30), .CO(n_1_31), .S(n_296));
   FA_X1 i_1_32 (.A(B[7]), .B(n_213), .CI(n_1_31), .CO(n_1_32), .S(n_297));
   FA_X1 i_1_33 (.A(B[8]), .B(n_214), .CI(n_1_32), .CO(n_1_33), .S(n_298));
   FA_X1 i_1_34 (.A(B[9]), .B(n_215), .CI(n_1_33), .CO(n_1_34), .S(n_299));
   FA_X1 i_1_35 (.A(B[10]), .B(n_216), .CI(n_1_34), .CO(n_1_35), .S(n_300));
   FA_X1 i_1_36 (.A(B[11]), .B(n_217), .CI(n_1_35), .CO(n_1_36), .S(n_301));
   FA_X1 i_1_37 (.A(B[15]), .B(n_218), .CI(n_1_36), .CO(n_1_37), .S(n_302));
   FA_X1 i_1_38 (.A(B[15]), .B(n_133), .CI(n_1_37), .CO(n_1_38), .S(n_303));
   FA_X1 i_1_39 (.A(n_146), .B(n_207), .CI(n_1_167), .CO(n_1_39), .S(n_304));
   FA_X1 i_1_40 (.A(n_147), .B(n_208), .CI(n_1_39), .CO(n_1_40), .S(n_305));
   FA_X1 i_1_41 (.A(n_148), .B(n_209), .CI(n_1_40), .CO(n_1_41), .S(n_306));
   FA_X1 i_1_42 (.A(n_255), .B(n_210), .CI(n_1_41), .CO(n_1_42), .S(n_307));
   FA_X1 i_1_43 (.A(n_256), .B(n_211), .CI(n_1_42), .CO(n_1_43), .S(n_308));
   FA_X1 i_1_44 (.A(n_257), .B(n_212), .CI(n_1_43), .CO(n_1_44), .S(n_309));
   FA_X1 i_1_45 (.A(n_258), .B(n_213), .CI(n_1_44), .CO(n_1_45), .S(n_310));
   FA_X1 i_1_46 (.A(n_259), .B(n_214), .CI(n_1_45), .CO(n_1_46), .S(n_311));
   FA_X1 i_1_47 (.A(n_260), .B(n_215), .CI(n_1_46), .CO(n_1_47), .S(n_312));
   FA_X1 i_1_48 (.A(n_261), .B(n_216), .CI(n_1_47), .CO(n_1_48), .S(n_313));
   FA_X1 i_1_49 (.A(n_262), .B(n_217), .CI(n_1_48), .CO(n_1_49), .S(n_314));
   FA_X1 i_1_50 (.A(n_263), .B(n_218), .CI(n_1_49), .CO(n_1_50), .S(n_315));
   FA_X1 i_1_51 (.A(n_264), .B(n_133), .CI(n_1_50), .CO(n_1_51), .S(n_316));
   FA_X1 i_1_52 (.A(B[1]), .B(n_195), .CI(n_1_168), .CO(n_1_52), .S(n_317));
   FA_X1 i_1_53 (.A(B[2]), .B(n_196), .CI(n_1_52), .CO(n_1_53), .S(n_318));
   FA_X1 i_1_54 (.A(B[3]), .B(n_197), .CI(n_1_53), .CO(n_1_54), .S(n_319));
   FA_X1 i_1_55 (.A(B[4]), .B(n_198), .CI(n_1_54), .CO(n_1_55), .S(n_320));
   FA_X1 i_1_56 (.A(B[5]), .B(n_199), .CI(n_1_55), .CO(n_1_56), .S(n_321));
   FA_X1 i_1_57 (.A(B[6]), .B(n_200), .CI(n_1_56), .CO(n_1_57), .S(n_322));
   FA_X1 i_1_58 (.A(B[7]), .B(n_201), .CI(n_1_57), .CO(n_1_58), .S(n_323));
   FA_X1 i_1_59 (.A(B[8]), .B(n_202), .CI(n_1_58), .CO(n_1_59), .S(n_324));
   FA_X1 i_1_60 (.A(B[9]), .B(n_203), .CI(n_1_59), .CO(n_1_60), .S(n_325));
   FA_X1 i_1_61 (.A(B[10]), .B(n_204), .CI(n_1_60), .CO(n_1_61), .S(n_326));
   FA_X1 i_1_62 (.A(B[11]), .B(n_205), .CI(n_1_61), .CO(n_1_62), .S(n_327));
   FA_X1 i_1_63 (.A(B[15]), .B(n_132), .CI(n_1_62), .CO(n_1_63), .S(n_328));
   FA_X1 i_1_64 (.A(n_146), .B(n_195), .CI(n_1_168), .CO(n_1_64), .S(n_329));
   FA_X1 i_1_65 (.A(n_147), .B(n_196), .CI(n_1_64), .CO(n_1_65), .S(n_330));
   FA_X1 i_1_66 (.A(n_148), .B(n_197), .CI(n_1_65), .CO(n_1_66), .S(n_331));
   FA_X1 i_1_67 (.A(n_255), .B(n_198), .CI(n_1_66), .CO(n_1_67), .S(n_332));
   FA_X1 i_1_68 (.A(n_256), .B(n_199), .CI(n_1_67), .CO(n_1_68), .S(n_333));
   FA_X1 i_1_69 (.A(n_257), .B(n_200), .CI(n_1_68), .CO(n_1_69), .S(n_334));
   FA_X1 i_1_70 (.A(n_258), .B(n_201), .CI(n_1_69), .CO(n_1_70), .S(n_335));
   FA_X1 i_1_71 (.A(n_259), .B(n_202), .CI(n_1_70), .CO(n_1_71), .S(n_336));
   FA_X1 i_1_72 (.A(n_260), .B(n_203), .CI(n_1_71), .CO(n_1_72), .S(n_337));
   FA_X1 i_1_73 (.A(n_261), .B(n_204), .CI(n_1_72), .CO(n_1_73), .S(n_338));
   FA_X1 i_1_74 (.A(n_262), .B(n_205), .CI(n_1_73), .CO(n_1_74), .S(n_339));
   FA_X1 i_1_75 (.A(n_263), .B(n_132), .CI(n_1_74), .CO(n_1_75), .S(n_340));
   FA_X1 i_1_76 (.A(B[1]), .B(n_184), .CI(n_1_169), .CO(n_1_76), .S(n_341));
   FA_X1 i_1_77 (.A(B[2]), .B(n_185), .CI(n_1_76), .CO(n_1_77), .S(n_342));
   FA_X1 i_1_78 (.A(B[3]), .B(n_186), .CI(n_1_77), .CO(n_1_78), .S(n_343));
   FA_X1 i_1_79 (.A(B[4]), .B(n_187), .CI(n_1_78), .CO(n_1_79), .S(n_344));
   FA_X1 i_1_80 (.A(B[5]), .B(n_188), .CI(n_1_79), .CO(n_1_80), .S(n_345));
   FA_X1 i_1_81 (.A(B[6]), .B(n_189), .CI(n_1_80), .CO(n_1_81), .S(n_346));
   FA_X1 i_1_82 (.A(B[7]), .B(n_190), .CI(n_1_81), .CO(n_1_82), .S(n_347));
   FA_X1 i_1_83 (.A(B[8]), .B(n_191), .CI(n_1_82), .CO(n_1_83), .S(n_348));
   FA_X1 i_1_84 (.A(B[9]), .B(n_192), .CI(n_1_83), .CO(n_1_84), .S(n_349));
   FA_X1 i_1_85 (.A(B[10]), .B(n_193), .CI(n_1_84), .CO(n_1_85), .S(n_350));
   FA_X1 i_1_86 (.A(B[11]), .B(n_131), .CI(n_1_85), .CO(n_1_86), .S(n_351));
   FA_X1 i_1_87 (.A(n_146), .B(n_184), .CI(n_1_169), .CO(n_1_87), .S(n_352));
   FA_X1 i_1_88 (.A(n_147), .B(n_185), .CI(n_1_87), .CO(n_1_88), .S(n_353));
   FA_X1 i_1_89 (.A(n_148), .B(n_186), .CI(n_1_88), .CO(n_1_89), .S(n_354));
   FA_X1 i_1_90 (.A(n_255), .B(n_187), .CI(n_1_89), .CO(n_1_90), .S(n_355));
   FA_X1 i_1_91 (.A(n_256), .B(n_188), .CI(n_1_90), .CO(n_1_91), .S(n_356));
   FA_X1 i_1_92 (.A(n_257), .B(n_189), .CI(n_1_91), .CO(n_1_92), .S(n_357));
   FA_X1 i_1_93 (.A(n_258), .B(n_190), .CI(n_1_92), .CO(n_1_93), .S(n_358));
   FA_X1 i_1_94 (.A(n_259), .B(n_191), .CI(n_1_93), .CO(n_1_94), .S(n_359));
   FA_X1 i_1_95 (.A(n_260), .B(n_192), .CI(n_1_94), .CO(n_1_95), .S(n_360));
   FA_X1 i_1_96 (.A(n_261), .B(n_193), .CI(n_1_95), .CO(n_1_96), .S(n_361));
   FA_X1 i_1_97 (.A(n_262), .B(n_131), .CI(n_1_96), .CO(n_1_97), .S(n_362));
   FA_X1 i_1_98 (.A(B[1]), .B(n_174), .CI(n_1_170), .CO(n_1_98), .S(n_363));
   FA_X1 i_1_99 (.A(B[2]), .B(n_175), .CI(n_1_98), .CO(n_1_99), .S(n_364));
   FA_X1 i_1_100 (.A(B[3]), .B(n_176), .CI(n_1_99), .CO(n_1_100), .S(n_365));
   FA_X1 i_1_101 (.A(B[4]), .B(n_177), .CI(n_1_100), .CO(n_1_101), .S(n_366));
   FA_X1 i_1_102 (.A(B[5]), .B(n_178), .CI(n_1_101), .CO(n_1_102), .S(n_367));
   FA_X1 i_1_103 (.A(B[6]), .B(n_179), .CI(n_1_102), .CO(n_1_103), .S(n_368));
   FA_X1 i_1_104 (.A(B[7]), .B(n_180), .CI(n_1_103), .CO(n_1_104), .S(n_369));
   FA_X1 i_1_105 (.A(B[8]), .B(n_181), .CI(n_1_104), .CO(n_1_105), .S(n_370));
   FA_X1 i_1_106 (.A(B[9]), .B(n_182), .CI(n_1_105), .CO(n_1_106), .S(n_371));
   FA_X1 i_1_107 (.A(B[10]), .B(n_130), .CI(n_1_106), .CO(n_1_107), .S(n_372));
   FA_X1 i_1_108 (.A(n_146), .B(n_174), .CI(n_1_170), .CO(n_1_108), .S(n_373));
   FA_X1 i_1_109 (.A(n_147), .B(n_175), .CI(n_1_108), .CO(n_1_109), .S(n_374));
   FA_X1 i_1_110 (.A(n_148), .B(n_176), .CI(n_1_109), .CO(n_1_110), .S(n_375));
   FA_X1 i_1_111 (.A(n_255), .B(n_177), .CI(n_1_110), .CO(n_1_111), .S(n_376));
   FA_X1 i_1_112 (.A(n_256), .B(n_178), .CI(n_1_111), .CO(n_1_112), .S(n_377));
   FA_X1 i_1_113 (.A(n_257), .B(n_179), .CI(n_1_112), .CO(n_1_113), .S(n_378));
   FA_X1 i_1_114 (.A(n_258), .B(n_180), .CI(n_1_113), .CO(n_1_114), .S(n_379));
   FA_X1 i_1_115 (.A(n_259), .B(n_181), .CI(n_1_114), .CO(n_1_115), .S(n_380));
   FA_X1 i_1_116 (.A(n_260), .B(n_182), .CI(n_1_115), .CO(n_1_116), .S(n_381));
   FA_X1 i_1_117 (.A(n_261), .B(n_130), .CI(n_1_116), .CO(n_1_117), .S(n_382));
   FA_X1 i_1_118 (.A(B[1]), .B(n_165), .CI(n_1_171), .CO(n_1_118), .S(n_383));
   FA_X1 i_1_119 (.A(B[2]), .B(n_166), .CI(n_1_118), .CO(n_1_119), .S(n_384));
   FA_X1 i_1_120 (.A(B[3]), .B(n_167), .CI(n_1_119), .CO(n_1_120), .S(n_385));
   FA_X1 i_1_121 (.A(B[4]), .B(n_168), .CI(n_1_120), .CO(n_1_121), .S(n_386));
   FA_X1 i_1_122 (.A(B[5]), .B(n_169), .CI(n_1_121), .CO(n_1_122), .S(n_387));
   FA_X1 i_1_123 (.A(B[6]), .B(n_170), .CI(n_1_122), .CO(n_1_123), .S(n_388));
   FA_X1 i_1_124 (.A(B[7]), .B(n_171), .CI(n_1_123), .CO(n_1_124), .S(n_389));
   FA_X1 i_1_125 (.A(B[8]), .B(n_172), .CI(n_1_124), .CO(n_1_125), .S(n_390));
   FA_X1 i_1_126 (.A(B[9]), .B(n_129), .CI(n_1_125), .CO(n_1_126), .S(n_391));
   FA_X1 i_1_127 (.A(n_146), .B(n_165), .CI(n_1_171), .CO(n_1_127), .S(n_392));
   FA_X1 i_1_128 (.A(n_147), .B(n_166), .CI(n_1_127), .CO(n_1_128), .S(n_393));
   FA_X1 i_1_129 (.A(n_148), .B(n_167), .CI(n_1_128), .CO(n_1_129), .S(n_394));
   FA_X1 i_1_130 (.A(n_255), .B(n_168), .CI(n_1_129), .CO(n_1_130), .S(n_395));
   FA_X1 i_1_131 (.A(n_256), .B(n_169), .CI(n_1_130), .CO(n_1_131), .S(n_396));
   FA_X1 i_1_132 (.A(n_257), .B(n_170), .CI(n_1_131), .CO(n_1_132), .S(n_397));
   FA_X1 i_1_133 (.A(n_258), .B(n_171), .CI(n_1_132), .CO(n_1_133), .S(n_398));
   FA_X1 i_1_134 (.A(n_259), .B(n_172), .CI(n_1_133), .CO(n_1_134), .S(n_399));
   FA_X1 i_1_135 (.A(n_260), .B(n_129), .CI(n_1_134), .CO(n_1_135), .S(n_400));
   FA_X1 i_1_136 (.A(B[1]), .B(n_157), .CI(n_1_172), .CO(n_1_136), .S(n_401));
   FA_X1 i_1_137 (.A(B[2]), .B(n_158), .CI(n_1_136), .CO(n_1_137), .S(n_402));
   FA_X1 i_1_138 (.A(B[3]), .B(n_159), .CI(n_1_137), .CO(n_1_138), .S(n_403));
   FA_X1 i_1_139 (.A(B[4]), .B(n_160), .CI(n_1_138), .CO(n_1_139), .S(n_404));
   FA_X1 i_1_140 (.A(B[5]), .B(n_161), .CI(n_1_139), .CO(n_1_140), .S(n_405));
   FA_X1 i_1_141 (.A(B[6]), .B(n_162), .CI(n_1_140), .CO(n_1_141), .S(n_406));
   FA_X1 i_1_142 (.A(B[7]), .B(n_163), .CI(n_1_141), .CO(n_1_142), .S(n_407));
   FA_X1 i_1_143 (.A(B[8]), .B(n_128), .CI(n_1_142), .CO(n_1_143), .S(n_408));
   FA_X1 i_1_144 (.A(n_146), .B(n_157), .CI(n_1_172), .CO(n_1_144), .S(n_409));
   FA_X1 i_1_145 (.A(n_147), .B(n_158), .CI(n_1_144), .CO(n_1_145), .S(n_410));
   FA_X1 i_1_146 (.A(n_148), .B(n_159), .CI(n_1_145), .CO(n_1_146), .S(n_411));
   FA_X1 i_1_147 (.A(n_255), .B(n_160), .CI(n_1_146), .CO(n_1_147), .S(n_412));
   FA_X1 i_1_148 (.A(n_256), .B(n_161), .CI(n_1_147), .CO(n_1_148), .S(n_413));
   FA_X1 i_1_149 (.A(n_257), .B(n_162), .CI(n_1_148), .CO(n_1_149), .S(n_414));
   FA_X1 i_1_150 (.A(n_258), .B(n_163), .CI(n_1_149), .CO(n_1_150), .S(n_415));
   FA_X1 i_1_151 (.A(n_259), .B(n_128), .CI(n_1_150), .CO(n_1_151), .S(n_416));
   FA_X1 i_1_152 (.A(B[1]), .B(n_150), .CI(n_1_173), .CO(n_1_152), .S(n_417));
   FA_X1 i_1_153 (.A(B[2]), .B(n_151), .CI(n_1_152), .CO(n_1_153), .S(n_418));
   FA_X1 i_1_154 (.A(B[3]), .B(n_152), .CI(n_1_153), .CO(n_1_154), .S(n_419));
   FA_X1 i_1_155 (.A(B[4]), .B(n_153), .CI(n_1_154), .CO(n_1_155), .S(n_420));
   FA_X1 i_1_156 (.A(B[5]), .B(n_154), .CI(n_1_155), .CO(n_1_156), .S(n_421));
   FA_X1 i_1_157 (.A(B[6]), .B(n_155), .CI(n_1_156), .CO(n_1_157), .S(n_422));
   FA_X1 i_1_158 (.A(B[7]), .B(n_127), .CI(n_1_157), .CO(n_1_158), .S(n_423));
   FA_X1 i_1_159 (.A(n_146), .B(n_150), .CI(n_1_173), .CO(n_1_159), .S(n_424));
   FA_X1 i_1_160 (.A(n_147), .B(n_151), .CI(n_1_159), .CO(n_1_160), .S(n_425));
   FA_X1 i_1_161 (.A(n_148), .B(n_152), .CI(n_1_160), .CO(n_1_161), .S(n_426));
   FA_X1 i_1_162 (.A(n_255), .B(n_153), .CI(n_1_161), .CO(n_1_162), .S(n_427));
   FA_X1 i_1_163 (.A(n_256), .B(n_154), .CI(n_1_162), .CO(n_1_163), .S(n_428));
   FA_X1 i_1_164 (.A(n_257), .B(n_155), .CI(n_1_163), .CO(n_1_164), .S(n_429));
   FA_X1 i_1_165 (.A(n_258), .B(n_127), .CI(n_1_164), .CO(n_1_165), .S(n_430));
   HA_X1 i_1_166 (.A(B[0]), .B(n_134), .CO(n_1_166), .S(n_431));
   HA_X1 i_1_167 (.A(B[0]), .B(n_206), .CO(n_1_167), .S(n_432));
   HA_X1 i_1_168 (.A(B[0]), .B(n_194), .CO(n_1_168), .S(n_433));
   HA_X1 i_1_169 (.A(B[0]), .B(n_183), .CO(n_1_169), .S(n_434));
   HA_X1 i_1_170 (.A(B[0]), .B(n_173), .CO(n_1_170), .S(n_435));
   HA_X1 i_1_171 (.A(B[0]), .B(n_164), .CO(n_1_171), .S(n_436));
   HA_X1 i_1_172 (.A(B[0]), .B(n_156), .CO(n_1_172), .S(n_437));
   HA_X1 i_1_173 (.A(B[0]), .B(n_149), .CO(n_1_173), .S(n_438));
   XNOR2_X1 i_1_174 (.A(n_112), .B(n_1_174), .ZN(n_439));
   XNOR2_X1 i_1_175 (.A(n_125), .B(n_1_25), .ZN(n_1_174));
   INV_X1 i_1_176 (.A(n_1_14), .ZN(n_1_175));
   XNOR2_X1 i_1_177 (.A(n_112), .B(B[15]), .ZN(n_1_176));
   INV_X1 i_1_178 (.A(n_1_176), .ZN(n_1_177));
   AOI22_X1 i_1_179 (.A1(n_1_175), .A2(n_1_176), .B1(n_1_14), .B2(n_1_177), 
      .ZN(n_440));
endmodule

module multiplier_16bit(first_operand, second_operand, out, enable, overflow);
   input [15:0]first_operand;
   input [15:0]second_operand;
   output [15:0]out;
   input enable;
   output overflow;

   wire [31:0]temp_result_wire;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_9;
   wire n_0_0_39;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_29;
   wire n_0_0_18;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_30;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_28;

   booth_16bit_multiplier mult (.A({first_operand[12], uc_0, uc_1, uc_2, 
      first_operand[11], first_operand[10], first_operand[9], first_operand[8], 
      first_operand[7], first_operand[6], first_operand[5], first_operand[4], 
      first_operand[3], first_operand[2], first_operand[1], first_operand[0]}), 
      .B({second_operand[12], uc_3, uc_4, uc_5, second_operand[11], 
      second_operand[10], second_operand[9], second_operand[8], 
      second_operand[7], second_operand[6], second_operand[5], second_operand[4], 
      second_operand[3], second_operand[2], second_operand[1], second_operand[0]}), 
      .product({uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, 
      uc_16, uc_17, temp_result_wire[19], temp_result_wire[18], 
      temp_result_wire[17], temp_result_wire[16], temp_result_wire[15], 
      temp_result_wire[14], temp_result_wire[13], temp_result_wire[12], 
      temp_result_wire[11], temp_result_wire[10], temp_result_wire[9], 
      temp_result_wire[8], temp_result_wire[7], temp_result_wire[6], 
      temp_result_wire[5], temp_result_wire[4], temp_result_wire[3], 
      temp_result_wire[2], temp_result_wire[1], temp_result_wire[0]}));
   MUX2_X1 i_0_0_0 (.A(temp_result_wire[0]), .B(temp_result_wire[4]), .S(
      n_0_0_30), .Z(n_0_0_0));
   MUX2_X1 i_0_0_1 (.A(temp_result_wire[1]), .B(temp_result_wire[5]), .S(
      n_0_0_30), .Z(n_0_0_1));
   MUX2_X1 i_0_0_2 (.A(temp_result_wire[2]), .B(temp_result_wire[6]), .S(
      n_0_0_30), .Z(n_0_0_2));
   MUX2_X1 i_0_0_3 (.A(temp_result_wire[3]), .B(temp_result_wire[7]), .S(
      n_0_0_30), .Z(n_0_0_3));
   MUX2_X1 i_0_0_4 (.A(temp_result_wire[4]), .B(temp_result_wire[8]), .S(
      n_0_0_30), .Z(n_0_0_4));
   MUX2_X1 i_0_0_5 (.A(temp_result_wire[5]), .B(temp_result_wire[9]), .S(
      n_0_0_30), .Z(n_0_0_5));
   MUX2_X1 i_0_0_6 (.A(temp_result_wire[6]), .B(temp_result_wire[10]), .S(
      n_0_0_30), .Z(n_0_0_6));
   MUX2_X1 i_0_0_7 (.A(temp_result_wire[7]), .B(temp_result_wire[11]), .S(
      n_0_0_30), .Z(n_0_0_7));
   MUX2_X1 i_0_0_8 (.A(temp_result_wire[8]), .B(temp_result_wire[12]), .S(
      n_0_0_30), .Z(n_0_0_8));
   MUX2_X1 i_0_0_16 (.A(n_0_0_0), .B(n_0_0_2), .S(n_0_0_29), .Z(n_0_0_31));
   MUX2_X1 i_0_0_17 (.A(n_0_0_1), .B(n_0_0_3), .S(n_0_0_29), .Z(n_0_0_32));
   MUX2_X1 i_0_0_18 (.A(n_0_0_2), .B(n_0_0_4), .S(n_0_0_29), .Z(n_0_0_33));
   MUX2_X1 i_0_0_19 (.A(n_0_0_3), .B(n_0_0_5), .S(n_0_0_29), .Z(n_0_0_34));
   MUX2_X1 i_0_0_20 (.A(n_0_0_4), .B(n_0_0_6), .S(n_0_0_29), .Z(n_0_0_35));
   MUX2_X1 i_0_0_21 (.A(n_0_0_5), .B(n_0_0_7), .S(n_0_0_29), .Z(n_0_0_36));
   MUX2_X1 i_0_0_22 (.A(n_0_0_6), .B(n_0_0_8), .S(n_0_0_29), .Z(n_0_0_37));
   MUX2_X1 i_0_0_23 (.A(n_0_0_7), .B(n_0_0_9), .S(n_0_0_29), .Z(n_0_0_38));
   MUX2_X1 i_0_0_30 (.A(n_0_0_31), .B(n_0_0_32), .S(n_0_0_28), .Z(out[0]));
   MUX2_X1 i_0_0_31 (.A(n_0_0_32), .B(n_0_0_33), .S(n_0_0_28), .Z(out[1]));
   MUX2_X1 i_0_0_32 (.A(n_0_0_33), .B(n_0_0_34), .S(n_0_0_28), .Z(out[2]));
   MUX2_X1 i_0_0_33 (.A(n_0_0_34), .B(n_0_0_35), .S(n_0_0_28), .Z(out[3]));
   MUX2_X1 i_0_0_34 (.A(n_0_0_35), .B(n_0_0_36), .S(n_0_0_28), .Z(out[4]));
   MUX2_X1 i_0_0_35 (.A(n_0_0_36), .B(n_0_0_37), .S(n_0_0_28), .Z(out[5]));
   MUX2_X1 i_0_0_36 (.A(n_0_0_37), .B(n_0_0_38), .S(n_0_0_28), .Z(out[6]));
   MUX2_X1 i_0_0_37 (.A(n_0_0_38), .B(n_0_0_39), .S(n_0_0_28), .Z(out[7]));
   INV_X1 i_0_0_43 (.A(second_operand[13]), .ZN(n_0_0_19));
   INV_X1 i_0_0_44 (.A(second_operand[14]), .ZN(n_0_0_20));
   OAI211_X1 i_0_0_45 (.A(n_0_0_19), .B(first_operand[13]), .C1(n_0_0_20), 
      .C2(first_operand[14]), .ZN(n_0_0_21));
   INV_X1 i_0_0_46 (.A(first_operand[14]), .ZN(n_0_0_22));
   OAI21_X1 i_0_0_47 (.A(n_0_0_21), .B1(second_operand[14]), .B2(n_0_0_22), 
      .ZN(n_0_0_23));
   INV_X1 i_0_0_48 (.A(second_operand[15]), .ZN(n_0_0_24));
   OAI21_X1 i_0_0_49 (.A(n_0_0_23), .B1(first_operand[15]), .B2(n_0_0_24), 
      .ZN(n_0_0_25));
   INV_X1 i_0_0_50 (.A(first_operand[15]), .ZN(n_0_0_26));
   OAI21_X1 i_0_0_51 (.A(n_0_0_25), .B1(second_operand[15]), .B2(n_0_0_26), 
      .ZN(n_0_0_27));
   MUX2_X1 i_0_0_55 (.A(second_operand[13]), .B(first_operand[13]), .S(n_0_0_27), 
      .Z(out[13]));
   MUX2_X1 i_0_0_56 (.A(second_operand[14]), .B(first_operand[14]), .S(n_0_0_27), 
      .Z(out[14]));
   MUX2_X1 i_0_0_57 (.A(second_operand[15]), .B(first_operand[15]), .S(n_0_0_27), 
      .Z(out[15]));
   NOR2_X1 i_0_0_9 (.A1(n_0_0_12), .A2(n_0_0_13), .ZN(n_0_0_9));
   AOI21_X1 i_0_0_10 (.A(n_0_0_10), .B1(n_0_0_16), .B2(n_0_0_29), .ZN(n_0_0_39));
   NOR2_X1 i_0_0_11 (.A1(n_0_0_8), .A2(n_0_0_29), .ZN(n_0_0_10));
   AOI21_X1 i_0_0_12 (.A(n_0_0_11), .B1(n_0_0_14), .B2(n_0_0_28), .ZN(out[9]));
   AND2_X1 i_0_0_13 (.A1(n_0_0_58), .A2(n_0_0_52), .ZN(n_0_0_11));
   NOR2_X1 i_0_0_14 (.A1(temp_result_wire[13]), .A2(n_0_0_82), .ZN(n_0_0_12));
   NOR2_X1 i_0_0_15 (.A1(temp_result_wire[9]), .A2(n_0_0_30), .ZN(n_0_0_13));
   OAI21_X1 i_0_0_24 (.A(n_0_0_15), .B1(n_0_0_40), .B2(n_0_0_84), .ZN(n_0_0_14));
   NAND2_X1 i_0_0_25 (.A1(n_0_0_16), .A2(n_0_0_84), .ZN(n_0_0_15));
   OAI21_X1 i_0_0_26 (.A(n_0_0_17), .B1(temp_result_wire[14]), .B2(n_0_0_82), 
      .ZN(n_0_0_16));
   OR2_X1 i_0_0_27 (.A1(temp_result_wire[10]), .A2(n_0_0_30), .ZN(n_0_0_17));
   INV_X1 i_0_0_28 (.A(n_0_0_84), .ZN(n_0_0_29));
   NAND2_X1 i_0_0_29 (.A1(n_0_0_42), .A2(n_0_0_18), .ZN(out[12]));
   NAND2_X1 i_0_0_38 (.A1(n_0_0_55), .A2(n_0_0_52), .ZN(n_0_0_18));
   MUX2_X1 i_0_0_39 (.A(temp_result_wire[16]), .B(temp_result_wire[12]), 
      .S(n_0_0_82), .Z(n_0_0_40));
   NAND2_X1 i_0_0_40 (.A1(temp_result_wire[14]), .A2(n_0_0_82), .ZN(n_0_0_41));
   NAND2_X1 i_0_0_41 (.A1(n_0_0_43), .A2(n_0_0_28), .ZN(n_0_0_42));
   OAI21_X1 i_0_0_42 (.A(n_0_0_44), .B1(n_0_0_45), .B2(n_0_0_84), .ZN(n_0_0_43));
   NAND2_X1 i_0_0_52 (.A1(n_0_0_57), .A2(n_0_0_84), .ZN(n_0_0_44));
   AOI21_X1 i_0_0_53 (.A(n_0_0_46), .B1(temp_result_wire[19]), .B2(n_0_0_30), 
      .ZN(n_0_0_45));
   INV_X1 i_0_0_54 (.A(n_0_0_47), .ZN(n_0_0_46));
   NAND2_X1 i_0_0_58 (.A1(temp_result_wire[15]), .A2(n_0_0_82), .ZN(n_0_0_47));
   NAND2_X1 i_0_0_59 (.A1(n_0_0_27), .A2(n_0_0_49), .ZN(n_0_0_48));
   INV_X1 i_0_0_60 (.A(second_operand[15]), .ZN(n_0_0_49));
   NAND2_X1 i_0_0_61 (.A1(n_0_0_27), .A2(n_0_0_51), .ZN(n_0_0_50));
   INV_X1 i_0_0_62 (.A(second_operand[14]), .ZN(n_0_0_51));
   OAI21_X1 i_0_0_63 (.A(n_0_0_53), .B1(first_operand[13]), .B2(n_0_0_27), 
      .ZN(n_0_0_52));
   NAND2_X1 i_0_0_64 (.A1(n_0_0_27), .A2(n_0_0_54), .ZN(n_0_0_53));
   INV_X1 i_0_0_65 (.A(second_operand[13]), .ZN(n_0_0_54));
   OAI21_X1 i_0_0_66 (.A(n_0_0_68), .B1(n_0_0_56), .B2(n_0_0_84), .ZN(n_0_0_55));
   AOI21_X1 i_0_0_67 (.A(n_0_0_69), .B1(temp_result_wire[18]), .B2(n_0_0_30), 
      .ZN(n_0_0_56));
   OAI21_X1 i_0_0_68 (.A(n_0_0_72), .B1(n_0_0_73), .B2(n_0_0_82), .ZN(n_0_0_57));
   OAI21_X1 i_0_0_69 (.A(n_0_0_61), .B1(n_0_0_58), .B2(n_0_0_52), .ZN(out[8]));
   INV_X1 i_0_0_70 (.A(n_0_0_59), .ZN(n_0_0_58));
   OAI21_X1 i_0_0_71 (.A(n_0_0_60), .B1(n_0_0_75), .B2(n_0_0_84), .ZN(n_0_0_59));
   OR3_X1 i_0_0_72 (.A1(n_0_0_12), .A2(n_0_0_13), .A3(n_0_0_83), .ZN(n_0_0_60));
   NAND2_X1 i_0_0_73 (.A1(n_0_0_39), .A2(n_0_0_52), .ZN(n_0_0_61));
   INV_X1 i_0_0_74 (.A(n_0_0_62), .ZN(out[10]));
   OAI221_X1 i_0_0_75 (.A(n_0_0_65), .B1(temp_result_wire[17]), .B2(n_0_0_81), 
      .C1(n_0_0_52), .C2(n_0_0_63), .ZN(n_0_0_62));
   AOI21_X1 i_0_0_76 (.A(n_0_0_64), .B1(n_0_0_75), .B2(n_0_0_78), .ZN(n_0_0_63));
   NOR3_X1 i_0_0_77 (.A1(temp_result_wire[13]), .A2(n_0_0_84), .A3(n_0_0_30), 
      .ZN(n_0_0_64));
   NAND2_X1 i_0_0_78 (.A1(n_0_0_14), .A2(n_0_0_52), .ZN(n_0_0_65));
   OAI211_X1 i_0_0_79 (.A(n_0_0_79), .B(n_0_0_70), .C1(n_0_0_52), .C2(n_0_0_66), 
      .ZN(out[11]));
   AOI21_X1 i_0_0_80 (.A(n_0_0_67), .B1(n_0_0_69), .B2(n_0_0_83), .ZN(n_0_0_66));
   INV_X1 i_0_0_81 (.A(n_0_0_68), .ZN(n_0_0_67));
   NAND2_X1 i_0_0_82 (.A1(n_0_0_40), .A2(n_0_0_84), .ZN(n_0_0_68));
   INV_X1 i_0_0_83 (.A(n_0_0_41), .ZN(n_0_0_69));
   NAND2_X1 i_0_0_84 (.A1(n_0_0_71), .A2(n_0_0_74), .ZN(n_0_0_70));
   OAI211_X1 i_0_0_85 (.A(n_0_0_83), .B(n_0_0_72), .C1(n_0_0_73), .C2(n_0_0_82), 
      .ZN(n_0_0_71));
   NAND2_X1 i_0_0_86 (.A1(temp_result_wire[13]), .A2(n_0_0_82), .ZN(n_0_0_72));
   INV_X1 i_0_0_87 (.A(temp_result_wire[17]), .ZN(n_0_0_73));
   AOI21_X1 i_0_0_88 (.A(n_0_0_28), .B1(n_0_0_75), .B2(n_0_0_78), .ZN(n_0_0_74));
   AOI21_X1 i_0_0_89 (.A(n_0_0_76), .B1(temp_result_wire[15]), .B2(n_0_0_30), 
      .ZN(n_0_0_75));
   INV_X1 i_0_0_90 (.A(n_0_0_77), .ZN(n_0_0_76));
   NAND2_X1 i_0_0_91 (.A1(temp_result_wire[11]), .A2(n_0_0_82), .ZN(n_0_0_77));
   INV_X1 i_0_0_92 (.A(n_0_0_29), .ZN(n_0_0_78));
   NAND2_X1 i_0_0_93 (.A1(temp_result_wire[18]), .A2(n_0_0_80), .ZN(n_0_0_79));
   INV_X1 i_0_0_94 (.A(n_0_0_81), .ZN(n_0_0_80));
   NAND3_X1 i_0_0_95 (.A1(n_0_0_28), .A2(n_0_0_83), .A3(n_0_0_30), .ZN(n_0_0_81));
   INV_X1 i_0_0_96 (.A(n_0_0_82), .ZN(n_0_0_30));
   OAI21_X1 i_0_0_97 (.A(n_0_0_48), .B1(n_0_0_27), .B2(first_operand[15]), 
      .ZN(n_0_0_82));
   INV_X1 i_0_0_98 (.A(n_0_0_84), .ZN(n_0_0_83));
   OAI21_X1 i_0_0_99 (.A(n_0_0_50), .B1(n_0_0_27), .B2(first_operand[14]), 
      .ZN(n_0_0_84));
   INV_X1 i_0_0_100 (.A(n_0_0_52), .ZN(n_0_0_28));
endmodule

module carry_lookahead_adder_4bit__3_97(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_0;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_6;

   AOI21_X1 i_0_0 (.A(n_0_11), .B1(n_0_10), .B2(n_0_2), .ZN(cout));
   XNOR2_X1 i_0_4 (.A(n_0_5), .B(n_0_1), .ZN(sum[2]));
   XNOR2_X1 i_0_5 (.A(in1[2]), .B(in0[2]), .ZN(n_0_1));
   XNOR2_X1 i_0_6 (.A(n_0_9), .B(n_0_2), .ZN(sum[3]));
   OAI21_X1 i_0_7 (.A(n_0_3), .B1(in0[2]), .B2(in1[2]), .ZN(n_0_2));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_9 (.A(n_0_5), .B1(in0[2]), .B2(in1[2]), .ZN(n_0_4));
   OAI21_X1 i_0_10 (.A(n_0_7), .B1(n_0_8), .B2(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_12 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_7));
   NOR2_X1 i_0_13 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(in1[3]), .B(in0[3]), .Z(n_0_9));
   NAND2_X1 i_0_15 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_10));
   NOR2_X1 i_0_16 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_11));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(sum[0]));
   XNOR2_X1 i_0_2 (.A(in0[0]), .B(in1[0]), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(n_0_12), .A2(n_0_16), .ZN(sum[1]));
   NAND3_X1 i_0_11 (.A1(n_0_14), .A2(n_0_13), .A3(n_0_15), .ZN(n_0_12));
   NAND2_X1 i_0_17 (.A1(n_0_19), .A2(in1[1]), .ZN(n_0_13));
   NAND2_X1 i_0_18 (.A1(n_0_20), .A2(in0[1]), .ZN(n_0_14));
   INV_X1 i_0_19 (.A(n_0_6), .ZN(n_0_15));
   NAND3_X1 i_0_20 (.A1(n_0_18), .A2(n_0_6), .A3(n_0_17), .ZN(n_0_16));
   NAND2_X1 i_0_21 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_17));
   NAND2_X1 i_0_22 (.A1(n_0_20), .A2(n_0_19), .ZN(n_0_18));
   INV_X1 i_0_23 (.A(in0[1]), .ZN(n_0_19));
   INV_X1 i_0_24 (.A(in1[1]), .ZN(n_0_20));
   NAND2_X1 i_0_25 (.A1(in0[0]), .A2(in1[0]), .ZN(n_0_6));
endmodule

module carry_lookahead_adder_4bit__3_88(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;

   AOI21_X1 i_0_0 (.A(n_0_13), .B1(n_0_1), .B2(n_0_12), .ZN(cout));
   XNOR2_X1 i_0_1 (.A(cin), .B(n_0_7), .ZN(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_6), .B(n_0_0), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(in1[1]), .B(in0[1]), .ZN(n_0_0));
   XOR2_X1 i_0_4 (.A(n_0_9), .B(n_0_3), .Z(sum[2]));
   XNOR2_X1 i_0_5 (.A(n_0_10), .B(n_0_1), .ZN(sum[3]));
   AOI21_X1 i_0_6 (.A(n_0_2), .B1(in0[2]), .B2(in1[2]), .ZN(n_0_1));
   NOR2_X1 i_0_7 (.A1(n_0_9), .A2(n_0_3), .ZN(n_0_2));
   OAI21_X1 i_0_8 (.A(n_0_4), .B1(in0[1]), .B2(in1[1]), .ZN(n_0_3));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(n_0_4));
   AOI21_X1 i_0_10 (.A(n_0_6), .B1(in0[1]), .B2(in1[1]), .ZN(n_0_5));
   OAI21_X1 i_0_11 (.A(n_0_8), .B1(n_0_7), .B2(n_0_14), .ZN(n_0_6));
   XNOR2_X1 i_0_12 (.A(in1[0]), .B(in0[0]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_8));
   XNOR2_X1 i_0_14 (.A(in1[2]), .B(in0[2]), .ZN(n_0_9));
   NOR2_X1 i_0_15 (.A1(n_0_13), .A2(n_0_11), .ZN(n_0_10));
   INV_X1 i_0_16 (.A(n_0_12), .ZN(n_0_11));
   NAND2_X1 i_0_17 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_12));
   NOR2_X1 i_0_18 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_13));
   INV_X1 i_0_19 (.A(cin), .ZN(n_0_14));
endmodule

module carry_lookahead_adder_4bit__3_79(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;

   AOI21_X1 i_0_0 (.A(n_0_13), .B1(n_0_1), .B2(n_0_12), .ZN(cout));
   XNOR2_X1 i_0_1 (.A(cin), .B(n_0_7), .ZN(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_6), .B(n_0_0), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(in1[1]), .B(in0[1]), .ZN(n_0_0));
   XOR2_X1 i_0_4 (.A(n_0_9), .B(n_0_3), .Z(sum[2]));
   XNOR2_X1 i_0_5 (.A(n_0_10), .B(n_0_1), .ZN(sum[3]));
   AOI21_X1 i_0_6 (.A(n_0_2), .B1(in0[2]), .B2(in1[2]), .ZN(n_0_1));
   NOR2_X1 i_0_7 (.A1(n_0_9), .A2(n_0_3), .ZN(n_0_2));
   OAI21_X1 i_0_8 (.A(n_0_4), .B1(in0[1]), .B2(in1[1]), .ZN(n_0_3));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(n_0_4));
   AOI21_X1 i_0_10 (.A(n_0_6), .B1(in0[1]), .B2(in1[1]), .ZN(n_0_5));
   OAI21_X1 i_0_11 (.A(n_0_8), .B1(n_0_7), .B2(n_0_14), .ZN(n_0_6));
   XNOR2_X1 i_0_12 (.A(in1[0]), .B(in0[0]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_8));
   XNOR2_X1 i_0_14 (.A(in1[2]), .B(in0[2]), .ZN(n_0_9));
   NOR2_X1 i_0_15 (.A1(n_0_13), .A2(n_0_11), .ZN(n_0_10));
   INV_X1 i_0_16 (.A(n_0_12), .ZN(n_0_11));
   NAND2_X1 i_0_17 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_12));
   NOR2_X1 i_0_18 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_13));
   INV_X1 i_0_19 (.A(cin), .ZN(n_0_14));
endmodule

module carry_lookahead_adder_4bit__3_70(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire [3:0]p;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .Z(p[0]));
   XOR2_X1 i_0_1 (.A(p[0]), .B(cin), .Z(sum[0]));
endmodule

module carry_lookahead_adder_20bit__3_98(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [19:0]in0;
   input [19:0]in1;
   input cin;
   output [19:0]sum;
   output cout;
   output v;

   wire c1;
   wire c2;
   wire c3;

   carry_lookahead_adder_4bit__3_97 cla0 (.in0({in0[3], in0[2], in0[1], in0[0]}), 
      .in1({in1[3], in1[2], in1[1], in1[0]}), .cin(), .sum({sum[3], sum[2], 
      sum[1], sum[0]}), .cout(c1), .v());
   carry_lookahead_adder_4bit__3_88 cla1 (.in0({in0[7], in0[6], in0[5], in0[4]}), 
      .in1({in1[7], in1[6], in1[5], in1[4]}), .cin(c1), .sum({sum[7], sum[6], 
      sum[5], sum[4]}), .cout(c2), .v());
   carry_lookahead_adder_4bit__3_79 cla2 (.in0({in0[11], in0[10], in0[9], in0[8]}), 
      .in1({in1[11], in1[10], in1[9], in1[8]}), .cin(c2), .sum({sum[11], sum[10], 
      sum[9], sum[8]}), .cout(c3), .v());
   carry_lookahead_adder_4bit__3_70 cla3 (.in0({uc_0, uc_1, uc_2, in0[12]}), 
      .in1({uc_3, uc_4, uc_5, in1[12]}), .cin(c3), .sum({uc_6, uc_7, uc_8, 
      sum[12]}), .cout(), .v());
endmodule

module add_sub_cla__3_99(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   wire n_0_28;
   wire n_0_29;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire [19:0]tempIn11;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire [19:0]tempIn22;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_83;
   wire n_0_81;
   wire n_0_1;
   wire n_0_80;
   wire n_0_2;
   wire n_0_25;
   wire n_0_4;
   wire n_0_23;
   wire n_0_6;
   wire n_0_8;
   wire n_0_31;
   wire n_0_30;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_16;
   wire n_0_22;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_21;
   wire n_0_20;
   wire n_0_24;
   wire n_0_26;
   wire n_0_27;
   wire n_0_82;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_78;
   wire n_0_134;
   wire n_0_79;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_0;
   wire n_0_141;
   wire n_0_14;
   wire n_0_15;
   wire n_0_142;
   wire n_0_143;
   wire n_0_7;
   wire n_0_144;
   wire n_0_145;
   wire n_0_5;
   wire n_0_146;
   wire n_0_3;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;

   carry_lookahead_adder_20bit__3_98 cs0 (.sub(), .in0({uc_0, uc_1, uc_2, uc_3, 
      uc_4, uc_5, uc_6, tempIn11[12], tempIn11[11], tempIn11[10], tempIn11[9], 
      tempIn11[8], tempIn11[7], tempIn11[6], tempIn11[5], tempIn11[4], 
      tempIn11[3], tempIn11[2], tempIn11[1], tempIn11[0]}), .in1({uc_7, uc_8, 
      uc_9, uc_10, uc_11, uc_12, uc_13, tempIn22[12], tempIn22[11], tempIn22[10], 
      tempIn22[9], tempIn22[8], tempIn22[7], tempIn22[6], tempIn22[5], 
      tempIn22[4], tempIn22[3], tempIn22[2], tempIn22[1], tempIn22[0]}), .cin(), 
      .sum({uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, out[12], out[11], 
      out[10], out[9], out[8], out[7], out[6], out[5], out[4], out[3], out[2], 
      out[1], out[0]}), .cout(), .v());
   AOI22_X1 i_0_16 (.A1(n_0_0), .A2(n_0_15), .B1(n_0_14), .B2(n_0_5), .ZN(
      out[13]));
   AOI22_X1 i_0_17 (.A1(n_0_7), .A2(n_0_15), .B1(n_0_14), .B2(n_0_3), .ZN(
      out[14]));
   OR2_X1 i_0_18 (.A1(in1[15]), .A2(in2[15]), .ZN(out[15]));
   NAND2_X1 i_0_33 (.A1(n_0_25), .A2(in1[1]), .ZN(n_0_28));
   INV_X1 i_0_34 (.A(n_0_28), .ZN(n_0_29));
   INV_X1 i_0_37 (.A(n_0_25), .ZN(n_0_32));
   AOI22_X1 i_0_38 (.A1(n_0_25), .A2(in1[2]), .B1(n_0_32), .B2(in1[0]), .ZN(
      n_0_33));
   INV_X1 i_0_39 (.A(n_0_33), .ZN(n_0_34));
   OAI221_X1 i_0_40 (.A(n_0_23), .B1(n_0_29), .B2(n_0_31), .C1(n_0_34), .C2(
      n_0_30), .ZN(n_0_35));
   INV_X1 i_0_41 (.A(in1[2]), .ZN(n_0_36));
   OAI22_X1 i_0_42 (.A1(n_0_35), .A2(n_0_21), .B1(n_0_36), .B2(n_0_20), .ZN(
      tempIn11[2]));
   AOI22_X1 i_0_43 (.A1(n_0_25), .A2(in1[3]), .B1(n_0_32), .B2(in1[1]), .ZN(
      n_0_37));
   OAI33_X1 i_0_44 (.A1(n_0_37), .A2(n_0_30), .A3(n_0_22), .B1(n_0_33), .B2(
      n_0_31), .B3(n_0_22), .ZN(n_0_38));
   AOI22_X1 i_0_45 (.A1(n_0_38), .A2(n_0_20), .B1(in1[3]), .B2(n_0_21), .ZN(
      n_0_39));
   INV_X1 i_0_46 (.A(n_0_39), .ZN(tempIn11[3]));
   OAI21_X1 i_0_47 (.A(n_0_30), .B1(n_0_37), .B2(n_0_22), .ZN(n_0_40));
   AOI22_X1 i_0_48 (.A1(n_0_25), .A2(in1[4]), .B1(n_0_32), .B2(in1[2]), .ZN(
      n_0_41));
   NAND2_X1 i_0_49 (.A1(n_0_25), .A2(in1[0]), .ZN(n_0_42));
   AOI22_X1 i_0_50 (.A1(n_0_41), .A2(n_0_23), .B1(n_0_42), .B2(n_0_22), .ZN(
      n_0_43));
   OAI21_X1 i_0_51 (.A(n_0_40), .B1(n_0_43), .B2(n_0_30), .ZN(n_0_44));
   INV_X1 i_0_52 (.A(in1[4]), .ZN(n_0_45));
   AOI22_X1 i_0_53 (.A1(n_0_44), .A2(n_0_20), .B1(n_0_21), .B2(n_0_45), .ZN(
      tempIn11[4]));
   OAI22_X1 i_0_54 (.A1(n_0_25), .A2(in1[3]), .B1(n_0_32), .B2(in1[5]), .ZN(
      n_0_46));
   AOI22_X1 i_0_55 (.A1(n_0_46), .A2(n_0_23), .B1(n_0_28), .B2(n_0_22), .ZN(
      n_0_47));
   OAI221_X1 i_0_56 (.A(n_0_20), .B1(n_0_47), .B2(n_0_30), .C1(n_0_43), .C2(
      n_0_31), .ZN(n_0_48));
   INV_X1 i_0_57 (.A(in1[5]), .ZN(n_0_49));
   OAI21_X1 i_0_58 (.A(n_0_48), .B1(n_0_49), .B2(n_0_20), .ZN(tempIn11[5]));
   AOI22_X1 i_0_59 (.A1(n_0_25), .A2(in1[6]), .B1(n_0_32), .B2(in1[4]), .ZN(
      n_0_50));
   AOI22_X1 i_0_60 (.A1(n_0_50), .A2(n_0_23), .B1(n_0_33), .B2(n_0_22), .ZN(
      n_0_51));
   AOI221_X1 i_0_61 (.A(n_0_21), .B1(n_0_47), .B2(n_0_30), .C1(n_0_51), .C2(
      n_0_31), .ZN(n_0_52));
   INV_X1 i_0_62 (.A(in1[6]), .ZN(n_0_53));
   AOI21_X1 i_0_63 (.A(n_0_52), .B1(n_0_53), .B2(n_0_21), .ZN(tempIn11[6]));
   AOI22_X1 i_0_64 (.A1(n_0_25), .A2(in1[7]), .B1(n_0_32), .B2(in1[5]), .ZN(
      n_0_54));
   OAI22_X1 i_0_65 (.A1(n_0_37), .A2(n_0_23), .B1(n_0_54), .B2(n_0_22), .ZN(
      n_0_55));
   AOI221_X1 i_0_66 (.A(n_0_21), .B1(n_0_55), .B2(n_0_31), .C1(n_0_51), .C2(
      n_0_30), .ZN(n_0_56));
   INV_X1 i_0_67 (.A(in1[7]), .ZN(n_0_57));
   AOI21_X1 i_0_68 (.A(n_0_56), .B1(n_0_57), .B2(n_0_21), .ZN(tempIn11[7]));
   OAI22_X1 i_0_69 (.A1(n_0_32), .A2(in1[8]), .B1(n_0_25), .B2(in1[6]), .ZN(
      n_0_58));
   OAI22_X1 i_0_70 (.A1(n_0_41), .A2(n_0_23), .B1(n_0_58), .B2(n_0_22), .ZN(
      n_0_59));
   OAI221_X1 i_0_71 (.A(n_0_20), .B1(n_0_59), .B2(n_0_30), .C1(n_0_55), .C2(
      n_0_31), .ZN(n_0_60));
   INV_X1 i_0_72 (.A(in1[8]), .ZN(n_0_61));
   OAI21_X1 i_0_73 (.A(n_0_60), .B1(n_0_61), .B2(n_0_20), .ZN(tempIn11[8]));
   AOI221_X1 i_0_74 (.A(n_0_22), .B1(n_0_25), .B2(in1[9]), .C1(in1[7]), .C2(
      n_0_32), .ZN(n_0_62));
   AOI21_X1 i_0_75 (.A(n_0_62), .B1(n_0_46), .B2(n_0_22), .ZN(n_0_63));
   OAI221_X1 i_0_76 (.A(n_0_20), .B1(n_0_31), .B2(n_0_59), .C1(n_0_63), .C2(
      n_0_30), .ZN(n_0_64));
   INV_X1 i_0_77 (.A(in1[9]), .ZN(n_0_65));
   OAI21_X1 i_0_78 (.A(n_0_64), .B1(n_0_65), .B2(n_0_20), .ZN(tempIn11[9]));
   OAI22_X1 i_0_79 (.A1(n_0_25), .A2(in1[8]), .B1(n_0_32), .B2(in1[10]), 
      .ZN(n_0_66));
   OAI22_X1 i_0_80 (.A1(n_0_50), .A2(n_0_23), .B1(n_0_66), .B2(n_0_22), .ZN(
      n_0_67));
   OAI221_X1 i_0_81 (.A(n_0_20), .B1(n_0_67), .B2(n_0_30), .C1(n_0_63), .C2(
      n_0_31), .ZN(n_0_68));
   INV_X1 i_0_82 (.A(in1[10]), .ZN(n_0_69));
   OAI21_X1 i_0_83 (.A(n_0_68), .B1(n_0_69), .B2(n_0_20), .ZN(tempIn11[10]));
   AOI22_X1 i_0_84 (.A1(n_0_25), .A2(in1[11]), .B1(n_0_32), .B2(in1[9]), 
      .ZN(n_0_70));
   OAI22_X1 i_0_85 (.A1(n_0_54), .A2(n_0_23), .B1(n_0_70), .B2(n_0_22), .ZN(
      n_0_71));
   OAI221_X1 i_0_86 (.A(n_0_20), .B1(n_0_67), .B2(n_0_31), .C1(n_0_71), .C2(
      n_0_30), .ZN(n_0_72));
   INV_X1 i_0_87 (.A(in1[11]), .ZN(n_0_73));
   OAI21_X1 i_0_88 (.A(n_0_72), .B1(n_0_73), .B2(n_0_20), .ZN(tempIn11[11]));
   AOI221_X1 i_0_89 (.A(n_0_22), .B1(n_0_32), .B2(in1[10]), .C1(in1[12]), 
      .C2(n_0_25), .ZN(n_0_74));
   AOI211_X1 i_0_90 (.A(n_0_30), .B(n_0_74), .C1(n_0_58), .C2(n_0_22), .ZN(
      n_0_75));
   AOI211_X1 i_0_91 (.A(n_0_21), .B(n_0_75), .C1(n_0_30), .C2(n_0_71), .ZN(
      n_0_76));
   INV_X1 i_0_92 (.A(in1[12]), .ZN(n_0_77));
   AOI21_X1 i_0_93 (.A(n_0_76), .B1(n_0_77), .B2(n_0_21), .ZN(tempIn11[12]));
   INV_X1 i_0_102 (.A(n_0_80), .ZN(n_0_84));
   AOI22_X1 i_0_103 (.A1(n_0_80), .A2(in2[0]), .B1(n_0_84), .B2(in2[2]), 
      .ZN(n_0_85));
   NOR2_X1 i_0_104 (.A1(n_0_85), .A2(n_0_79), .ZN(n_0_86));
   AOI221_X1 i_0_105 (.A(n_0_14), .B1(in2[1]), .B2(n_0_81), .C1(n_0_86), 
      .C2(n_0_31), .ZN(n_0_87));
   INV_X1 i_0_106 (.A(in2[2]), .ZN(n_0_88));
   AOI21_X1 i_0_107 (.A(n_0_87), .B1(n_0_88), .B2(n_0_14), .ZN(tempIn22[2]));
   AOI22_X1 i_0_108 (.A1(n_0_84), .A2(in2[3]), .B1(n_0_80), .B2(in2[1]), 
      .ZN(n_0_89));
   NOR2_X1 i_0_109 (.A1(n_0_89), .A2(n_0_79), .ZN(n_0_90));
   AOI221_X1 i_0_110 (.A(n_0_14), .B1(n_0_86), .B2(n_0_30), .C1(n_0_31), 
      .C2(n_0_90), .ZN(n_0_91));
   INV_X1 i_0_111 (.A(in2[3]), .ZN(n_0_92));
   AOI21_X1 i_0_112 (.A(n_0_91), .B1(n_0_92), .B2(n_0_14), .ZN(tempIn22[3]));
   AOI22_X1 i_0_113 (.A1(n_0_84), .A2(in2[4]), .B1(n_0_80), .B2(in2[2]), 
      .ZN(n_0_93));
   NAND2_X1 i_0_114 (.A1(n_0_79), .A2(n_0_84), .ZN(n_0_94));
   OAI22_X1 i_0_115 (.A1(n_0_93), .A2(n_0_79), .B1(n_0_94), .B2(n_0_78), 
      .ZN(n_0_95));
   OAI221_X1 i_0_116 (.A(n_0_15), .B1(n_0_90), .B2(n_0_31), .C1(n_0_95), 
      .C2(n_0_30), .ZN(n_0_96));
   INV_X1 i_0_117 (.A(in2[4]), .ZN(n_0_97));
   OAI21_X1 i_0_118 (.A(n_0_96), .B1(n_0_97), .B2(n_0_15), .ZN(tempIn22[4]));
   AOI22_X1 i_0_119 (.A1(n_0_84), .A2(in2[5]), .B1(n_0_80), .B2(in2[3]), 
      .ZN(n_0_98));
   OAI22_X1 i_0_120 (.A1(n_0_98), .A2(n_0_79), .B1(n_0_94), .B2(n_0_83), 
      .ZN(n_0_99));
   OAI221_X1 i_0_121 (.A(n_0_15), .B1(n_0_95), .B2(n_0_31), .C1(n_0_30), 
      .C2(n_0_99), .ZN(n_0_100));
   INV_X1 i_0_122 (.A(in2[5]), .ZN(n_0_101));
   OAI21_X1 i_0_123 (.A(n_0_100), .B1(n_0_101), .B2(n_0_15), .ZN(tempIn22[5]));
   INV_X1 i_0_124 (.A(n_0_79), .ZN(n_0_102));
   AOI22_X1 i_0_125 (.A1(n_0_80), .A2(in2[4]), .B1(n_0_84), .B2(in2[6]), 
      .ZN(n_0_103));
   OAI22_X1 i_0_126 (.A1(n_0_85), .A2(n_0_102), .B1(n_0_103), .B2(n_0_79), 
      .ZN(n_0_104));
   AOI221_X1 i_0_127 (.A(n_0_14), .B1(n_0_99), .B2(n_0_30), .C1(n_0_104), 
      .C2(n_0_31), .ZN(n_0_105));
   INV_X1 i_0_128 (.A(in2[6]), .ZN(n_0_106));
   AOI21_X1 i_0_129 (.A(n_0_105), .B1(n_0_106), .B2(n_0_14), .ZN(tempIn22[6]));
   AOI22_X1 i_0_130 (.A1(n_0_84), .A2(in2[7]), .B1(n_0_80), .B2(in2[5]), 
      .ZN(n_0_107));
   AOI22_X1 i_0_131 (.A1(n_0_107), .A2(n_0_102), .B1(n_0_89), .B2(n_0_79), 
      .ZN(n_0_108));
   AOI221_X1 i_0_132 (.A(n_0_14), .B1(n_0_104), .B2(n_0_30), .C1(n_0_31), 
      .C2(n_0_108), .ZN(n_0_109));
   INV_X1 i_0_133 (.A(in2[7]), .ZN(n_0_110));
   AOI21_X1 i_0_134 (.A(n_0_109), .B1(n_0_110), .B2(n_0_14), .ZN(tempIn22[7]));
   AOI22_X1 i_0_135 (.A1(n_0_84), .A2(in2[8]), .B1(n_0_80), .B2(in2[6]), 
      .ZN(n_0_111));
   OAI22_X1 i_0_136 (.A1(n_0_93), .A2(n_0_102), .B1(n_0_111), .B2(n_0_79), 
      .ZN(n_0_112));
   AOI221_X1 i_0_137 (.A(n_0_14), .B1(n_0_112), .B2(n_0_31), .C1(n_0_30), 
      .C2(n_0_108), .ZN(n_0_113));
   INV_X1 i_0_138 (.A(in2[8]), .ZN(n_0_114));
   AOI21_X1 i_0_139 (.A(n_0_113), .B1(n_0_114), .B2(n_0_14), .ZN(tempIn22[8]));
   OAI221_X1 i_0_140 (.A(n_0_102), .B1(n_0_80), .B2(in2[9]), .C1(in2[7]), 
      .C2(n_0_84), .ZN(n_0_115));
   OAI21_X1 i_0_141 (.A(n_0_115), .B1(n_0_102), .B2(n_0_98), .ZN(n_0_116));
   OAI221_X1 i_0_142 (.A(n_0_15), .B1(n_0_31), .B2(n_0_112), .C1(n_0_116), 
      .C2(n_0_30), .ZN(n_0_117));
   INV_X1 i_0_143 (.A(in2[9]), .ZN(n_0_118));
   OAI21_X1 i_0_144 (.A(n_0_117), .B1(n_0_118), .B2(n_0_15), .ZN(tempIn22[9]));
   OAI221_X1 i_0_145 (.A(n_0_102), .B1(n_0_84), .B2(in2[8]), .C1(in2[10]), 
      .C2(n_0_80), .ZN(n_0_119));
   OAI21_X1 i_0_146 (.A(n_0_119), .B1(n_0_102), .B2(n_0_103), .ZN(n_0_120));
   OAI221_X1 i_0_147 (.A(n_0_15), .B1(n_0_116), .B2(n_0_31), .C1(n_0_30), 
      .C2(n_0_120), .ZN(n_0_121));
   INV_X1 i_0_148 (.A(in2[10]), .ZN(n_0_122));
   OAI21_X1 i_0_149 (.A(n_0_121), .B1(n_0_122), .B2(n_0_15), .ZN(tempIn22[10]));
   OAI22_X1 i_0_150 (.A1(n_0_84), .A2(in2[9]), .B1(n_0_80), .B2(in2[11]), 
      .ZN(n_0_123));
   OAI22_X1 i_0_151 (.A1(n_0_107), .A2(n_0_102), .B1(n_0_123), .B2(n_0_79), 
      .ZN(n_0_124));
   OAI221_X1 i_0_152 (.A(n_0_15), .B1(n_0_30), .B2(n_0_124), .C1(n_0_120), 
      .C2(n_0_31), .ZN(n_0_125));
   INV_X1 i_0_153 (.A(in2[11]), .ZN(n_0_126));
   OAI21_X1 i_0_154 (.A(n_0_125), .B1(n_0_126), .B2(n_0_15), .ZN(tempIn22[11]));
   NOR2_X1 i_0_155 (.A1(n_0_15), .A2(in2[12]), .ZN(n_0_127));
   NOR2_X1 i_0_156 (.A1(n_0_84), .A2(in2[10]), .ZN(n_0_128));
   AOI22_X1 i_0_157 (.A1(n_0_111), .A2(n_0_79), .B1(n_0_128), .B2(n_0_102), 
      .ZN(n_0_129));
   OAI22_X1 i_0_158 (.A1(n_0_124), .A2(n_0_31), .B1(n_0_129), .B2(n_0_30), 
      .ZN(n_0_130));
   AOI21_X1 i_0_159 (.A(n_0_127), .B1(n_0_130), .B2(n_0_15), .ZN(tempIn22[12]));
   INV_X1 i_0_0 (.A(in2[1]), .ZN(n_0_83));
   INV_X1 i_0_1 (.A(n_0_1), .ZN(n_0_81));
   NAND2_X1 i_0_2 (.A1(n_0_134), .A2(n_0_8), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(n_0_80));
   NAND2_X1 i_0_4 (.A1(n_0_132), .A2(n_0_6), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(n_0_4), .ZN(n_0_25));
   NAND2_X1 i_0_6 (.A1(n_0_13), .A2(n_0_82), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(n_0_22), .ZN(n_0_23));
   NAND3_X1 i_0_8 (.A1(n_0_146), .A2(n_0_143), .A3(n_0_140), .ZN(n_0_6));
   NAND2_X1 i_0_9 (.A1(n_0_132), .A2(n_0_82), .ZN(n_0_8));
   INV_X1 i_0_10 (.A(n_0_30), .ZN(n_0_31));
   NAND2_X1 i_0_11 (.A1(n_0_145), .A2(n_0_140), .ZN(n_0_30));
   INV_X1 i_0_12 (.A(n_0_9), .ZN(tempIn11[0]));
   NAND2_X1 i_0_13 (.A1(n_0_21), .A2(in1[0]), .ZN(n_0_9));
   NAND2_X1 i_0_14 (.A1(n_0_10), .A2(n_0_19), .ZN(tempIn11[1]));
   NAND3_X1 i_0_15 (.A1(n_0_16), .A2(n_0_20), .A3(n_0_11), .ZN(n_0_10));
   INV_X1 i_0_19 (.A(n_0_12), .ZN(n_0_11));
   NAND3_X1 i_0_20 (.A1(n_0_13), .A2(in1[0]), .A3(n_0_82), .ZN(n_0_12));
   NAND2_X1 i_0_21 (.A1(n_0_133), .A2(n_0_145), .ZN(n_0_13));
   INV_X1 i_0_22 (.A(n_0_22), .ZN(n_0_16));
   NAND2_X1 i_0_23 (.A1(n_0_142), .A2(n_0_17), .ZN(n_0_22));
   NAND3_X1 i_0_24 (.A1(n_0_18), .A2(n_0_148), .A3(n_0_146), .ZN(n_0_17));
   NAND2_X1 i_0_25 (.A1(n_0_131), .A2(n_0_143), .ZN(n_0_18));
   NAND2_X1 i_0_26 (.A1(n_0_21), .A2(in1[1]), .ZN(n_0_19));
   INV_X1 i_0_27 (.A(n_0_20), .ZN(n_0_21));
   NAND2_X1 i_0_28 (.A1(n_0_138), .A2(n_0_149), .ZN(n_0_20));
   INV_X1 i_0_29 (.A(n_0_24), .ZN(tempIn22[0]));
   NAND2_X1 i_0_30 (.A1(n_0_14), .A2(in2[0]), .ZN(n_0_24));
   NAND2_X1 i_0_31 (.A1(n_0_26), .A2(n_0_141), .ZN(tempIn22[1]));
   NAND3_X1 i_0_32 (.A1(n_0_134), .A2(n_0_27), .A3(n_0_15), .ZN(n_0_26));
   AOI21_X1 i_0_35 (.A(n_0_78), .B1(n_0_132), .B2(n_0_82), .ZN(n_0_27));
   NAND3_X1 i_0_36 (.A1(n_0_131), .A2(n_0_146), .A3(n_0_143), .ZN(n_0_82));
   INV_X1 i_0_94 (.A(n_0_145), .ZN(n_0_131));
   NAND2_X1 i_0_95 (.A1(n_0_133), .A2(n_0_137), .ZN(n_0_132));
   NAND2_X1 i_0_96 (.A1(n_0_146), .A2(n_0_143), .ZN(n_0_133));
   INV_X1 i_0_97 (.A(in2[0]), .ZN(n_0_78));
   INV_X1 i_0_98 (.A(n_0_79), .ZN(n_0_134));
   NAND2_X1 i_0_99 (.A1(n_0_138), .A2(n_0_135), .ZN(n_0_79));
   NAND3_X1 i_0_100 (.A1(n_0_136), .A2(n_0_148), .A3(n_0_143), .ZN(n_0_135));
   NAND2_X1 i_0_101 (.A1(n_0_137), .A2(n_0_146), .ZN(n_0_136));
   INV_X1 i_0_160 (.A(n_0_140), .ZN(n_0_137));
   NAND3_X1 i_0_161 (.A1(n_0_147), .A2(n_0_146), .A3(n_0_139), .ZN(n_0_138));
   NAND2_X1 i_0_162 (.A1(n_0_143), .A2(n_0_140), .ZN(n_0_139));
   NAND2_X1 i_0_163 (.A1(n_0_0), .A2(in2[13]), .ZN(n_0_140));
   INV_X1 i_0_164 (.A(in1[13]), .ZN(n_0_0));
   NAND2_X1 i_0_165 (.A1(n_0_14), .A2(in2[1]), .ZN(n_0_141));
   INV_X1 i_0_166 (.A(n_0_15), .ZN(n_0_14));
   NAND2_X1 i_0_167 (.A1(n_0_142), .A2(n_0_151), .ZN(n_0_15));
   NAND3_X1 i_0_168 (.A1(n_0_147), .A2(n_0_144), .A3(n_0_143), .ZN(n_0_142));
   NAND2_X1 i_0_169 (.A1(n_0_7), .A2(in2[14]), .ZN(n_0_143));
   INV_X1 i_0_170 (.A(in1[14]), .ZN(n_0_7));
   NAND2_X1 i_0_171 (.A1(n_0_146), .A2(n_0_145), .ZN(n_0_144));
   NAND2_X1 i_0_172 (.A1(n_0_5), .A2(in1[13]), .ZN(n_0_145));
   INV_X1 i_0_173 (.A(in2[13]), .ZN(n_0_5));
   NAND2_X1 i_0_174 (.A1(n_0_3), .A2(in1[14]), .ZN(n_0_146));
   INV_X1 i_0_175 (.A(in2[14]), .ZN(n_0_3));
   INV_X1 i_0_176 (.A(n_0_148), .ZN(n_0_147));
   NAND2_X1 i_0_177 (.A1(n_0_151), .A2(n_0_149), .ZN(n_0_148));
   NAND2_X1 i_0_178 (.A1(n_0_150), .A2(in2[15]), .ZN(n_0_149));
   INV_X1 i_0_179 (.A(in1[15]), .ZN(n_0_150));
   NAND2_X1 i_0_180 (.A1(n_0_152), .A2(in1[15]), .ZN(n_0_151));
   INV_X1 i_0_181 (.A(in2[15]), .ZN(n_0_152));
endmodule

module carry_lookahead_adder_4bit__3_161(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   AOI21_X1 i_0_0 (.A(n_0_11), .B1(n_0_10), .B2(n_0_2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1[0]), .B(in0[0]), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_6), .B(n_0_0), .ZN(sum[1]));
   XOR2_X1 i_0_3 (.A(in1[1]), .B(in0[1]), .Z(n_0_0));
   XNOR2_X1 i_0_4 (.A(n_0_5), .B(n_0_1), .ZN(sum[2]));
   XNOR2_X1 i_0_5 (.A(in1[2]), .B(in0[2]), .ZN(n_0_1));
   XNOR2_X1 i_0_6 (.A(n_0_9), .B(n_0_2), .ZN(sum[3]));
   OAI21_X1 i_0_7 (.A(n_0_3), .B1(in0[2]), .B2(in1[2]), .ZN(n_0_2));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_9 (.A(n_0_5), .B1(in0[2]), .B2(in1[2]), .ZN(n_0_4));
   OAI21_X1 i_0_10 (.A(n_0_7), .B1(n_0_8), .B2(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_11 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_7));
   NOR2_X1 i_0_13 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(in1[3]), .B(in0[3]), .Z(n_0_9));
   NAND2_X1 i_0_15 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_10));
   NOR2_X1 i_0_16 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_11));
endmodule

module carry_lookahead_adder_4bit__3_152(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   AOI21_X1 i_0_0 (.A(n_0_13), .B1(n_0_1), .B2(n_0_12), .ZN(cout));
   XNOR2_X1 i_0_1 (.A(cin), .B(n_0_6), .ZN(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_5), .B(n_0_0), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(in1[1]), .B(in0[1]), .ZN(n_0_0));
   XOR2_X1 i_0_4 (.A(n_0_9), .B(n_0_3), .Z(sum[2]));
   XNOR2_X1 i_0_5 (.A(n_0_10), .B(n_0_1), .ZN(sum[3]));
   AOI21_X1 i_0_6 (.A(n_0_2), .B1(in0[2]), .B2(in1[2]), .ZN(n_0_1));
   NOR2_X1 i_0_7 (.A1(n_0_9), .A2(n_0_3), .ZN(n_0_2));
   XNOR2_X1 i_0_14 (.A(in1[2]), .B(in0[2]), .ZN(n_0_9));
   NOR2_X1 i_0_15 (.A1(n_0_13), .A2(n_0_11), .ZN(n_0_10));
   INV_X1 i_0_16 (.A(n_0_12), .ZN(n_0_11));
   NAND2_X1 i_0_17 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_12));
   NOR2_X1 i_0_18 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_13));
   OAI22_X1 i_0_8 (.A1(in1[1]), .A2(in0[1]), .B1(n_0_5), .B2(n_0_4), .ZN(n_0_3));
   AND2_X1 i_0_9 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_4));
   OAI21_X1 i_0_10 (.A(n_0_7), .B1(n_0_8), .B2(n_0_6), .ZN(n_0_5));
   OAI21_X1 i_0_11 (.A(n_0_7), .B1(in1[0]), .B2(in0[0]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_7));
   INV_X1 i_0_13 (.A(cin), .ZN(n_0_8));
endmodule

module carry_lookahead_adder_4bit__3_143(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;

   AOI21_X1 i_0_0 (.A(n_0_13), .B1(n_0_1), .B2(n_0_12), .ZN(cout));
   XNOR2_X1 i_0_1 (.A(cin), .B(n_0_7), .ZN(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_6), .B(n_0_0), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(in1[1]), .B(in0[1]), .ZN(n_0_0));
   XOR2_X1 i_0_4 (.A(n_0_9), .B(n_0_3), .Z(sum[2]));
   XNOR2_X1 i_0_5 (.A(n_0_11), .B(n_0_1), .ZN(sum[3]));
   AOI21_X1 i_0_6 (.A(n_0_2), .B1(in0[2]), .B2(in1[2]), .ZN(n_0_1));
   NOR2_X1 i_0_7 (.A1(n_0_9), .A2(n_0_3), .ZN(n_0_2));
   OAI21_X1 i_0_8 (.A(n_0_4), .B1(in0[1]), .B2(in1[1]), .ZN(n_0_3));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(n_0_4));
   AOI21_X1 i_0_10 (.A(n_0_6), .B1(in0[1]), .B2(in1[1]), .ZN(n_0_5));
   OAI21_X1 i_0_11 (.A(n_0_8), .B1(n_0_7), .B2(n_0_10), .ZN(n_0_6));
   XNOR2_X1 i_0_12 (.A(in1[0]), .B(in0[0]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_8));
   XNOR2_X1 i_0_14 (.A(in1[2]), .B(in0[2]), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(cin), .ZN(n_0_10));
   AOI21_X1 i_0_15 (.A(n_0_13), .B1(in1[3]), .B2(in0[3]), .ZN(n_0_11));
   NAND2_X1 i_0_16 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_12));
   NOR2_X1 i_0_17 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_13));
endmodule

module carry_lookahead_adder_4bit__3_134(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire [3:0]p;

   XOR2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .Z(p[0]));
   XOR2_X1 i_0_1 (.A(p[0]), .B(cin), .Z(sum[0]));
endmodule

module carry_lookahead_adder_20bit__3_162(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [19:0]in0;
   input [19:0]in1;
   input cin;
   output [19:0]sum;
   output cout;
   output v;

   wire c1;
   wire c2;
   wire c3;

   carry_lookahead_adder_4bit__3_161 cla0 (.in0({in0[3], in0[2], in0[1], in0[0]}), 
      .in1({in1[3], in1[2], in1[1], in1[0]}), .cin(), .sum({sum[3], sum[2], 
      sum[1], sum[0]}), .cout(c1), .v());
   carry_lookahead_adder_4bit__3_152 cla1 (.in0({in0[7], in0[6], in0[5], in0[4]}), 
      .in1({in1[7], in1[6], in1[5], in1[4]}), .cin(c1), .sum({sum[7], sum[6], 
      sum[5], sum[4]}), .cout(c2), .v());
   carry_lookahead_adder_4bit__3_143 cla2 (.in0({in0[11], in0[10], in0[9], 
      in0[8]}), .in1({in1[11], in1[10], in1[9], in1[8]}), .cin(c2), .sum({
      sum[11], sum[10], sum[9], sum[8]}), .cout(c3), .v());
   carry_lookahead_adder_4bit__3_134 cla3 (.in0({uc_0, uc_1, uc_2, in0[12]}), 
      .in1({uc_3, uc_4, uc_5, in1[12]}), .cin(c3), .sum({uc_6, uc_7, uc_8, 
      sum[12]}), .cout(), .v());
endmodule

module add_sub_cla__3_163(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   wire [19:0]tempIn11;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_72;
   wire n_0_73;
   wire n_0_78;
   wire [19:0]tempIn22;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_58;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_71;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;

   carry_lookahead_adder_20bit__3_162 cs0 (.sub(), .in0({uc_0, uc_1, uc_2, uc_3, 
      uc_4, uc_5, uc_6, tempIn11[12], tempIn11[11], tempIn11[10], tempIn11[9], 
      tempIn11[8], tempIn11[7], tempIn11[6], tempIn11[5], tempIn11[4], 
      tempIn11[3], tempIn11[2], tempIn11[1], tempIn11[0]}), .in1({uc_7, uc_8, 
      uc_9, uc_10, uc_11, uc_12, uc_13, tempIn22[12], tempIn22[11], tempIn22[10], 
      tempIn22[9], tempIn22[8], tempIn22[7], tempIn22[6], tempIn22[5], 
      tempIn22[4], tempIn22[3], tempIn22[2], tempIn22[1], tempIn22[0]}), .cin(), 
      .sum({uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, out[12], out[11], 
      out[10], out[9], out[8], out[7], out[6], out[5], out[4], out[3], out[2], 
      out[1], out[0]}), .cout(), .v());
   AOI22_X1 i_0_17 (.A1(n_0_15), .A2(n_0_2), .B1(n_0_3), .B2(n_0_13), .ZN(
      out[14]));
   OR2_X1 i_0_18 (.A1(in1[15]), .A2(in2[15]), .ZN(out[15]));
   AND2_X1 i_0_0 (.A1(n_0_35), .A2(in1[0]), .ZN(tempIn11[0]));
   AOI22_X1 i_0_1 (.A1(n_0_19), .A2(in1[3]), .B1(n_0_18), .B2(in1[1]), .ZN(
      n_0_37));
   OAI33_X1 i_0_2 (.A1(n_0_37), .A2(n_0_33), .A3(n_0_25), .B1(n_0_31), .B2(
      n_0_32), .B3(n_0_25), .ZN(n_0_38));
   AOI22_X1 i_0_3 (.A1(n_0_38), .A2(n_0_21), .B1(in1[3]), .B2(n_0_35), .ZN(
      n_0_39));
   INV_X1 i_0_4 (.A(n_0_39), .ZN(tempIn11[3]));
   OAI21_X1 i_0_5 (.A(n_0_33), .B1(n_0_37), .B2(n_0_25), .ZN(n_0_40));
   AOI22_X1 i_0_6 (.A1(n_0_19), .A2(in1[4]), .B1(n_0_18), .B2(in1[2]), .ZN(
      n_0_41));
   NAND2_X1 i_0_7 (.A1(n_0_19), .A2(in1[0]), .ZN(n_0_42));
   AOI22_X1 i_0_8 (.A1(n_0_41), .A2(n_0_26), .B1(n_0_42), .B2(n_0_25), .ZN(
      n_0_43));
   OAI21_X1 i_0_9 (.A(n_0_40), .B1(n_0_43), .B2(n_0_33), .ZN(n_0_44));
   INV_X1 i_0_10 (.A(in1[4]), .ZN(n_0_45));
   AOI22_X1 i_0_11 (.A1(n_0_44), .A2(n_0_21), .B1(n_0_35), .B2(n_0_45), .ZN(
      tempIn11[4]));
   OAI22_X1 i_0_12 (.A1(n_0_19), .A2(in1[3]), .B1(n_0_18), .B2(in1[5]), .ZN(
      n_0_46));
   AOI22_X1 i_0_13 (.A1(n_0_46), .A2(n_0_26), .B1(n_0_34), .B2(n_0_25), .ZN(
      n_0_47));
   OAI221_X1 i_0_14 (.A(n_0_21), .B1(n_0_47), .B2(n_0_33), .C1(n_0_43), .C2(
      n_0_32), .ZN(n_0_48));
   INV_X1 i_0_15 (.A(in1[5]), .ZN(n_0_49));
   OAI21_X1 i_0_16 (.A(n_0_48), .B1(n_0_49), .B2(n_0_21), .ZN(tempIn11[5]));
   AOI22_X1 i_0_59 (.A1(n_0_19), .A2(in1[6]), .B1(n_0_18), .B2(in1[4]), .ZN(
      n_0_50));
   AOI22_X1 i_0_60 (.A1(n_0_50), .A2(n_0_26), .B1(n_0_31), .B2(n_0_25), .ZN(
      n_0_51));
   AOI221_X1 i_0_61 (.A(n_0_35), .B1(n_0_47), .B2(n_0_33), .C1(n_0_51), .C2(
      n_0_32), .ZN(n_0_52));
   INV_X1 i_0_62 (.A(in1[6]), .ZN(n_0_53));
   AOI21_X1 i_0_63 (.A(n_0_52), .B1(n_0_53), .B2(n_0_35), .ZN(tempIn11[6]));
   AOI22_X1 i_0_64 (.A1(n_0_19), .A2(in1[7]), .B1(n_0_18), .B2(in1[5]), .ZN(
      n_0_54));
   OAI22_X1 i_0_65 (.A1(n_0_37), .A2(n_0_26), .B1(n_0_54), .B2(n_0_25), .ZN(
      n_0_55));
   AOI221_X1 i_0_66 (.A(n_0_35), .B1(n_0_55), .B2(n_0_32), .C1(n_0_51), .C2(
      n_0_33), .ZN(n_0_56));
   INV_X1 i_0_67 (.A(in1[7]), .ZN(n_0_57));
   AOI21_X1 i_0_68 (.A(n_0_56), .B1(n_0_57), .B2(n_0_35), .ZN(tempIn11[7]));
   OAI22_X1 i_0_70 (.A1(n_0_41), .A2(n_0_26), .B1(n_0_58), .B2(n_0_25), .ZN(
      n_0_59));
   OAI221_X1 i_0_71 (.A(n_0_21), .B1(n_0_59), .B2(n_0_33), .C1(n_0_55), .C2(
      n_0_32), .ZN(n_0_60));
   INV_X1 i_0_72 (.A(in1[8]), .ZN(n_0_61));
   OAI21_X1 i_0_73 (.A(n_0_60), .B1(n_0_61), .B2(n_0_21), .ZN(tempIn11[8]));
   AOI221_X1 i_0_74 (.A(n_0_25), .B1(n_0_19), .B2(in1[9]), .C1(in1[7]), .C2(
      n_0_18), .ZN(n_0_62));
   AOI21_X1 i_0_75 (.A(n_0_62), .B1(n_0_46), .B2(n_0_25), .ZN(n_0_63));
   OAI221_X1 i_0_76 (.A(n_0_21), .B1(n_0_32), .B2(n_0_59), .C1(n_0_63), .C2(
      n_0_33), .ZN(n_0_64));
   INV_X1 i_0_77 (.A(in1[9]), .ZN(n_0_65));
   OAI21_X1 i_0_78 (.A(n_0_64), .B1(n_0_65), .B2(n_0_21), .ZN(tempIn11[9]));
   OAI22_X1 i_0_79 (.A1(n_0_19), .A2(in1[8]), .B1(n_0_18), .B2(in1[10]), 
      .ZN(n_0_66));
   OAI22_X1 i_0_80 (.A1(n_0_50), .A2(n_0_26), .B1(n_0_66), .B2(n_0_25), .ZN(
      n_0_67));
   OAI221_X1 i_0_81 (.A(n_0_21), .B1(n_0_67), .B2(n_0_33), .C1(n_0_63), .C2(
      n_0_32), .ZN(n_0_68));
   INV_X1 i_0_82 (.A(in1[10]), .ZN(n_0_69));
   OAI21_X1 i_0_83 (.A(n_0_68), .B1(n_0_69), .B2(n_0_21), .ZN(tempIn11[10]));
   AOI22_X1 i_0_84 (.A1(n_0_19), .A2(in1[11]), .B1(n_0_18), .B2(in1[9]), 
      .ZN(n_0_70));
   OAI221_X1 i_0_86 (.A(n_0_21), .B1(n_0_67), .B2(n_0_32), .C1(n_0_71), .C2(
      n_0_33), .ZN(n_0_72));
   INV_X1 i_0_87 (.A(in1[11]), .ZN(n_0_73));
   OAI21_X1 i_0_88 (.A(n_0_72), .B1(n_0_73), .B2(n_0_21), .ZN(tempIn11[11]));
   INV_X1 i_0_19 (.A(in2[0]), .ZN(n_0_78));
   NOR2_X1 i_0_20 (.A1(n_0_2), .A2(n_0_78), .ZN(tempIn22[0]));
   OAI21_X1 i_0_21 (.A(n_0_22), .B1(n_0_4), .B2(n_0_23), .ZN(n_0_79));
   XNOR2_X1 i_0_22 (.A(n_0_20), .B(n_0_24), .ZN(n_0_80));
   NOR3_X1 i_0_23 (.A1(n_0_79), .A2(n_0_80), .A3(n_0_32), .ZN(n_0_81));
   NAND3_X1 i_0_25 (.A1(n_0_81), .A2(in2[0]), .A3(n_0_2), .ZN(n_0_82));
   INV_X1 i_0_27 (.A(in2[1]), .ZN(n_0_83));
   OAI21_X1 i_0_28 (.A(n_0_82), .B1(n_0_83), .B2(n_0_2), .ZN(tempIn22[1]));
   INV_X1 i_0_30 (.A(n_0_80), .ZN(n_0_84));
   AOI22_X1 i_0_31 (.A1(n_0_80), .A2(in2[0]), .B1(n_0_84), .B2(in2[2]), .ZN(
      n_0_85));
   NOR2_X1 i_0_32 (.A1(n_0_85), .A2(n_0_79), .ZN(n_0_86));
   AOI221_X1 i_0_33 (.A(n_0_3), .B1(in2[1]), .B2(n_0_81), .C1(n_0_86), .C2(
      n_0_32), .ZN(n_0_87));
   INV_X1 i_0_34 (.A(in2[2]), .ZN(n_0_88));
   AOI21_X1 i_0_36 (.A(n_0_87), .B1(n_0_88), .B2(n_0_3), .ZN(tempIn22[2]));
   AOI22_X1 i_0_38 (.A1(n_0_84), .A2(in2[3]), .B1(n_0_80), .B2(in2[1]), .ZN(
      n_0_89));
   NOR2_X1 i_0_39 (.A1(n_0_89), .A2(n_0_79), .ZN(n_0_90));
   AOI221_X1 i_0_40 (.A(n_0_3), .B1(n_0_86), .B2(n_0_33), .C1(n_0_32), .C2(
      n_0_90), .ZN(n_0_91));
   INV_X1 i_0_41 (.A(in2[3]), .ZN(n_0_92));
   AOI21_X1 i_0_42 (.A(n_0_91), .B1(n_0_92), .B2(n_0_3), .ZN(tempIn22[3]));
   AOI22_X1 i_0_43 (.A1(n_0_84), .A2(in2[4]), .B1(n_0_80), .B2(in2[2]), .ZN(
      n_0_93));
   NAND2_X1 i_0_44 (.A1(n_0_79), .A2(n_0_84), .ZN(n_0_94));
   OAI22_X1 i_0_45 (.A1(n_0_93), .A2(n_0_79), .B1(n_0_94), .B2(n_0_78), .ZN(
      n_0_95));
   OAI221_X1 i_0_46 (.A(n_0_2), .B1(n_0_90), .B2(n_0_32), .C1(n_0_95), .C2(
      n_0_33), .ZN(n_0_96));
   INV_X1 i_0_47 (.A(in2[4]), .ZN(n_0_97));
   OAI21_X1 i_0_48 (.A(n_0_96), .B1(n_0_97), .B2(n_0_2), .ZN(tempIn22[4]));
   AOI22_X1 i_0_119 (.A1(n_0_84), .A2(in2[5]), .B1(n_0_80), .B2(in2[3]), 
      .ZN(n_0_98));
   OAI22_X1 i_0_120 (.A1(n_0_98), .A2(n_0_79), .B1(n_0_94), .B2(n_0_83), 
      .ZN(n_0_99));
   OAI221_X1 i_0_121 (.A(n_0_2), .B1(n_0_95), .B2(n_0_32), .C1(n_0_33), .C2(
      n_0_99), .ZN(n_0_100));
   INV_X1 i_0_122 (.A(in2[5]), .ZN(n_0_101));
   OAI21_X1 i_0_123 (.A(n_0_100), .B1(n_0_101), .B2(n_0_2), .ZN(tempIn22[5]));
   INV_X1 i_0_49 (.A(n_0_79), .ZN(n_0_102));
   AOI22_X1 i_0_125 (.A1(n_0_80), .A2(in2[4]), .B1(n_0_84), .B2(in2[6]), 
      .ZN(n_0_103));
   OAI22_X1 i_0_126 (.A1(n_0_85), .A2(n_0_102), .B1(n_0_103), .B2(n_0_79), 
      .ZN(n_0_104));
   AOI221_X1 i_0_127 (.A(n_0_3), .B1(n_0_99), .B2(n_0_33), .C1(n_0_104), 
      .C2(n_0_32), .ZN(n_0_105));
   INV_X1 i_0_128 (.A(in2[6]), .ZN(n_0_106));
   AOI21_X1 i_0_129 (.A(n_0_105), .B1(n_0_106), .B2(n_0_3), .ZN(tempIn22[6]));
   AOI22_X1 i_0_50 (.A1(n_0_84), .A2(in2[7]), .B1(n_0_80), .B2(in2[5]), .ZN(
      n_0_107));
   AOI22_X1 i_0_131 (.A1(n_0_107), .A2(n_0_102), .B1(n_0_89), .B2(n_0_79), 
      .ZN(n_0_108));
   AOI221_X1 i_0_132 (.A(n_0_3), .B1(n_0_104), .B2(n_0_33), .C1(n_0_32), 
      .C2(n_0_108), .ZN(n_0_109));
   INV_X1 i_0_133 (.A(in2[7]), .ZN(n_0_110));
   AOI21_X1 i_0_134 (.A(n_0_109), .B1(n_0_110), .B2(n_0_3), .ZN(tempIn22[7]));
   AOI22_X1 i_0_135 (.A1(n_0_84), .A2(in2[8]), .B1(n_0_80), .B2(in2[6]), 
      .ZN(n_0_111));
   OAI22_X1 i_0_136 (.A1(n_0_93), .A2(n_0_102), .B1(n_0_111), .B2(n_0_79), 
      .ZN(n_0_112));
   AOI221_X1 i_0_137 (.A(n_0_3), .B1(n_0_112), .B2(n_0_32), .C1(n_0_33), 
      .C2(n_0_108), .ZN(n_0_113));
   INV_X1 i_0_138 (.A(in2[8]), .ZN(n_0_114));
   AOI21_X1 i_0_139 (.A(n_0_113), .B1(n_0_114), .B2(n_0_3), .ZN(tempIn22[8]));
   OAI221_X1 i_0_140 (.A(n_0_102), .B1(n_0_80), .B2(in2[9]), .C1(in2[7]), 
      .C2(n_0_84), .ZN(n_0_115));
   OAI21_X1 i_0_141 (.A(n_0_115), .B1(n_0_102), .B2(n_0_98), .ZN(n_0_116));
   OAI221_X1 i_0_142 (.A(n_0_2), .B1(n_0_32), .B2(n_0_112), .C1(n_0_116), 
      .C2(n_0_33), .ZN(n_0_117));
   INV_X1 i_0_143 (.A(in2[9]), .ZN(n_0_118));
   OAI21_X1 i_0_144 (.A(n_0_117), .B1(n_0_118), .B2(n_0_2), .ZN(tempIn22[9]));
   OAI221_X1 i_0_145 (.A(n_0_102), .B1(n_0_84), .B2(in2[8]), .C1(in2[10]), 
      .C2(n_0_80), .ZN(n_0_119));
   OAI21_X1 i_0_146 (.A(n_0_119), .B1(n_0_102), .B2(n_0_103), .ZN(n_0_120));
   OAI221_X1 i_0_147 (.A(n_0_2), .B1(n_0_116), .B2(n_0_32), .C1(n_0_33), 
      .C2(n_0_120), .ZN(n_0_121));
   INV_X1 i_0_148 (.A(in2[10]), .ZN(n_0_122));
   OAI21_X1 i_0_149 (.A(n_0_121), .B1(n_0_122), .B2(n_0_2), .ZN(tempIn22[10]));
   OAI22_X1 i_0_51 (.A1(n_0_84), .A2(in2[9]), .B1(n_0_80), .B2(in2[11]), 
      .ZN(n_0_123));
   OAI22_X1 i_0_52 (.A1(n_0_107), .A2(n_0_102), .B1(n_0_123), .B2(n_0_79), 
      .ZN(n_0_124));
   OAI221_X1 i_0_152 (.A(n_0_2), .B1(n_0_33), .B2(n_0_124), .C1(n_0_120), 
      .C2(n_0_32), .ZN(n_0_125));
   INV_X1 i_0_153 (.A(in2[11]), .ZN(n_0_126));
   OAI21_X1 i_0_154 (.A(n_0_125), .B1(n_0_126), .B2(n_0_2), .ZN(tempIn22[11]));
   NOR2_X1 i_0_155 (.A1(n_0_2), .A2(in2[12]), .ZN(n_0_127));
   NOR2_X1 i_0_156 (.A1(n_0_84), .A2(in2[10]), .ZN(n_0_128));
   AOI22_X1 i_0_157 (.A1(n_0_111), .A2(n_0_79), .B1(n_0_128), .B2(n_0_102), 
      .ZN(n_0_129));
   OAI22_X1 i_0_158 (.A1(n_0_124), .A2(n_0_32), .B1(n_0_129), .B2(n_0_33), 
      .ZN(n_0_130));
   AOI21_X1 i_0_159 (.A(n_0_127), .B1(n_0_130), .B2(n_0_2), .ZN(tempIn22[12]));
   INV_X1 i_0_24 (.A(n_0_133), .ZN(n_0_58));
   INV_X1 i_0_26 (.A(n_0_74), .ZN(tempIn11[12]));
   NAND2_X1 i_0_29 (.A1(n_0_76), .A2(n_0_75), .ZN(n_0_74));
   OR2_X1 i_0_35 (.A1(in1[12]), .A2(n_0_21), .ZN(n_0_75));
   OAI21_X1 i_0_37 (.A(n_0_77), .B1(n_0_136), .B2(n_0_132), .ZN(n_0_76));
   AOI21_X1 i_0_69 (.A(n_0_35), .B1(n_0_71), .B2(n_0_33), .ZN(n_0_77));
   OAI21_X1 i_0_85 (.A(n_0_131), .B1(n_0_70), .B2(n_0_25), .ZN(n_0_71));
   OR2_X1 i_0_89 (.A1(n_0_54), .A2(n_0_26), .ZN(n_0_131));
   OAI211_X1 i_0_93 (.A(n_0_10), .B(n_0_24), .C1(n_0_133), .C2(n_0_26), .ZN(
      n_0_132));
   AOI21_X1 i_0_160 (.A(n_0_134), .B1(n_0_135), .B2(n_0_18), .ZN(n_0_133));
   NOR2_X1 i_0_161 (.A1(in1[8]), .A2(n_0_18), .ZN(n_0_134));
   INV_X1 i_0_162 (.A(in1[6]), .ZN(n_0_135));
   AOI21_X1 i_0_53 (.A(n_0_0), .B1(in1[12]), .B2(n_0_19), .ZN(n_0_136));
   OAI21_X1 i_0_54 (.A(n_0_26), .B1(n_0_1), .B2(n_0_19), .ZN(n_0_0));
   INV_X1 i_0_55 (.A(in1[10]), .ZN(n_0_1));
   OAI22_X1 i_0_56 (.A1(n_0_14), .A2(n_0_3), .B1(n_0_12), .B2(n_0_2), .ZN(
      out[13]));
   INV_X1 i_0_57 (.A(n_0_3), .ZN(n_0_2));
   OAI21_X1 i_0_58 (.A(n_0_6), .B1(n_0_7), .B2(n_0_5), .ZN(n_0_3));
   AOI21_X1 i_0_90 (.A(n_0_5), .B1(n_0_16), .B2(in2[15]), .ZN(n_0_4));
   NOR2_X1 i_0_91 (.A1(n_0_16), .A2(in2[15]), .ZN(n_0_5));
   NAND2_X1 i_0_92 (.A1(n_0_16), .A2(in2[15]), .ZN(n_0_6));
   OAI21_X1 i_0_94 (.A(n_0_11), .B1(n_0_10), .B2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_95 (.A(n_0_9), .ZN(n_0_8));
   NOR2_X1 i_0_96 (.A1(in1[14]), .A2(n_0_13), .ZN(n_0_9));
   NAND2_X1 i_0_97 (.A1(in1[13]), .A2(n_0_12), .ZN(n_0_10));
   NAND2_X1 i_0_98 (.A1(in1[14]), .A2(n_0_13), .ZN(n_0_11));
   INV_X1 i_0_99 (.A(in2[13]), .ZN(n_0_12));
   INV_X1 i_0_100 (.A(in2[14]), .ZN(n_0_13));
   INV_X1 i_0_101 (.A(in1[13]), .ZN(n_0_14));
   INV_X1 i_0_102 (.A(in1[14]), .ZN(n_0_15));
   INV_X1 i_0_103 (.A(in1[15]), .ZN(n_0_16));
   OAI22_X1 i_0_104 (.A1(n_0_18), .A2(n_0_17), .B1(n_0_27), .B2(n_0_21), 
      .ZN(tempIn11[1]));
   NAND3_X1 i_0_105 (.A1(in1[0]), .A2(n_0_26), .A3(n_0_21), .ZN(n_0_17));
   INV_X1 i_0_106 (.A(n_0_19), .ZN(n_0_18));
   XOR2_X1 i_0_107 (.A(n_0_10), .B(n_0_20), .Z(n_0_19));
   NAND2_X1 i_0_108 (.A1(n_0_11), .A2(n_0_8), .ZN(n_0_20));
   NAND2_X1 i_0_109 (.A1(n_0_6), .A2(n_0_22), .ZN(n_0_21));
   NAND2_X1 i_0_110 (.A1(n_0_4), .A2(n_0_23), .ZN(n_0_22));
   OAI21_X1 i_0_111 (.A(n_0_8), .B1(n_0_28), .B2(n_0_24), .ZN(n_0_23));
   NAND2_X1 i_0_112 (.A1(n_0_14), .A2(in2[13]), .ZN(n_0_24));
   INV_X1 i_0_113 (.A(n_0_26), .ZN(n_0_25));
   XOR2_X1 i_0_114 (.A(n_0_4), .B(n_0_7), .Z(n_0_26));
   INV_X1 i_0_115 (.A(in1[1]), .ZN(n_0_27));
   INV_X1 i_0_116 (.A(n_0_11), .ZN(n_0_28));
   INV_X1 i_0_117 (.A(n_0_29), .ZN(tempIn11[2]));
   AOI22_X1 i_0_118 (.A1(in1[2]), .A2(n_0_35), .B1(n_0_21), .B2(n_0_30), 
      .ZN(n_0_29));
   AOI221_X1 i_0_124 (.A(n_0_36), .B1(n_0_32), .B2(n_0_31), .C1(n_0_34), 
      .C2(n_0_33), .ZN(n_0_30));
   AOI22_X1 i_0_130 (.A1(in1[0]), .A2(n_0_18), .B1(n_0_19), .B2(in1[2]), 
      .ZN(n_0_31));
   INV_X1 i_0_150 (.A(n_0_33), .ZN(n_0_32));
   NAND2_X1 i_0_151 (.A1(n_0_24), .A2(n_0_10), .ZN(n_0_33));
   NAND2_X1 i_0_163 (.A1(n_0_19), .A2(in1[1]), .ZN(n_0_34));
   INV_X1 i_0_164 (.A(n_0_21), .ZN(n_0_35));
   INV_X1 i_0_165 (.A(n_0_26), .ZN(n_0_36));
endmodule

module carry_lookahead_adder_4bit__3_8(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   AOI21_X1 i_0_0 (.A(n_0_11), .B1(n_0_10), .B2(n_0_2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(in1[0]), .B(in0[0]), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_6), .B(n_0_0), .ZN(sum[1]));
   XOR2_X1 i_0_3 (.A(in1[1]), .B(in0[1]), .Z(n_0_0));
   XNOR2_X1 i_0_4 (.A(n_0_5), .B(n_0_1), .ZN(sum[2]));
   XNOR2_X1 i_0_5 (.A(in1[2]), .B(in0[2]), .ZN(n_0_1));
   XNOR2_X1 i_0_6 (.A(n_0_9), .B(n_0_2), .ZN(sum[3]));
   OAI21_X1 i_0_7 (.A(n_0_3), .B1(in0[2]), .B2(in1[2]), .ZN(n_0_2));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_9 (.A(n_0_5), .B1(in0[2]), .B2(in1[2]), .ZN(n_0_4));
   OAI21_X1 i_0_10 (.A(n_0_7), .B1(n_0_8), .B2(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_11 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_7));
   NOR2_X1 i_0_13 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(in1[3]), .B(in0[3]), .Z(n_0_9));
   NAND2_X1 i_0_15 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_10));
   NOR2_X1 i_0_16 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_11));
endmodule

module carry_lookahead_adder_4bit__3_17(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_2;
   wire n_0_9;
   wire n_0_15;
   wire n_0_1;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;

   XNOR2_X1 i_0_0 (.A(cin), .B(n_0_10), .ZN(sum[0]));
   XNOR2_X1 i_0_1 (.A(n_0_8), .B(n_0_0), .ZN(sum[1]));
   XNOR2_X1 i_0_2 (.A(in1[1]), .B(in0[1]), .ZN(n_0_0));
   XOR2_X1 i_0_4 (.A(n_0_9), .B(n_0_6), .Z(sum[2]));
   XNOR2_X1 i_0_5 (.A(n_0_13), .B(n_0_3), .ZN(sum[3]));
   NOR2_X1 i_0_7 (.A1(n_0_9), .A2(n_0_6), .ZN(n_0_2));
   XNOR2_X1 i_0_14 (.A(in1[2]), .B(in0[2]), .ZN(n_0_9));
   NOR2_X1 i_0_6 (.A1(n_0_15), .A2(n_0_14), .ZN(cout));
   AOI21_X1 i_0_17 (.A(n_0_1), .B1(in1[3]), .B2(in0[3]), .ZN(n_0_15));
   INV_X1 i_0_18 (.A(n_0_3), .ZN(n_0_1));
   AND2_X1 i_0_20 (.A1(n_0_5), .A2(n_0_4), .ZN(n_0_3));
   NAND2_X1 i_0_21 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_4));
   INV_X1 i_0_22 (.A(n_0_2), .ZN(n_0_5));
   OAI22_X1 i_0_3 (.A1(in1[1]), .A2(in0[1]), .B1(n_0_8), .B2(n_0_7), .ZN(n_0_6));
   AND2_X1 i_0_8 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_7));
   OAI21_X1 i_0_9 (.A(n_0_11), .B1(n_0_12), .B2(n_0_10), .ZN(n_0_8));
   OAI21_X1 i_0_10 (.A(n_0_11), .B1(in1[0]), .B2(in0[0]), .ZN(n_0_10));
   NAND2_X1 i_0_11 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_11));
   INV_X1 i_0_12 (.A(cin), .ZN(n_0_12));
   AOI21_X1 i_0_13 (.A(n_0_14), .B1(in1[3]), .B2(in0[3]), .ZN(n_0_13));
   NOR2_X1 i_0_15 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_14));
endmodule

module carry_lookahead_adder_4bit__3_26(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_2;
   wire n_0_4;
   wire n_0_5;
   wire n_0_8;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_3;
   wire n_0_18;
   wire n_0_19;
   wire n_0_9;
   wire n_0_6;
   wire n_0_7;
   wire n_0_1;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_20;

   XNOR2_X1 i_0_0 (.A(cin), .B(n_0_7), .ZN(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_6), .B(n_0_0), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(in1[1]), .B(in0[1]), .ZN(n_0_0));
   XOR2_X1 i_0_4 (.A(n_0_9), .B(n_0_3), .Z(sum[2]));
   XNOR2_X1 i_0_5 (.A(n_0_12), .B(n_0_11), .ZN(sum[3]));
   NAND2_X1 i_0_1 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_2), .ZN(n_0_4));
   OR2_X1 i_0_7 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_5));
   AOI21_X1 i_0_8 (.A(n_0_4), .B1(cin), .B2(n_0_5), .ZN(n_0_8));
   NOR2_X1 i_0_9 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_14));
   INV_X1 i_0_10 (.A(in1[1]), .ZN(n_0_15));
   INV_X1 i_0_11 (.A(in0[1]), .ZN(n_0_16));
   OAI22_X1 i_0_12 (.A1(n_0_8), .A2(n_0_14), .B1(n_0_15), .B2(n_0_16), .ZN(
      n_0_17));
   INV_X1 i_0_13 (.A(n_0_17), .ZN(n_0_3));
   OR2_X1 i_0_14 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_18));
   NAND2_X1 i_0_17 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_19));
   NAND2_X1 i_0_18 (.A1(n_0_18), .A2(n_0_19), .ZN(n_0_9));
   INV_X1 i_0_19 (.A(n_0_8), .ZN(n_0_6));
   NAND2_X1 i_0_15 (.A1(n_0_5), .A2(n_0_2), .ZN(n_0_7));
   INV_X1 i_0_22 (.A(n_0_19), .ZN(n_0_1));
   AOI21_X1 i_0_23 (.A(n_0_1), .B1(n_0_17), .B2(n_0_18), .ZN(n_0_10));
   AOI21_X1 i_0_25 (.A(n_0_20), .B1(n_0_13), .B2(n_0_10), .ZN(cout));
   BUF_X1 i_0_27 (.A(n_0_10), .Z(n_0_11));
   AOI21_X1 i_0_16 (.A(n_0_20), .B1(in1[3]), .B2(in0[3]), .ZN(n_0_12));
   NAND2_X1 i_0_20 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_13));
   NOR2_X1 i_0_21 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_20));
endmodule

module carry_lookahead_adder_4bit__3_35(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(cin), .B(n_0_0), .Z(sum[0]));
   XOR2_X1 i_0_1 (.A(in1[0]), .B(in0[0]), .Z(n_0_0));
endmodule

module carry_lookahead_adder_20bit__0_1292(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [19:0]in0;
   input [19:0]in1;
   input cin;
   output [19:0]sum;
   output cout;
   output v;

   wire c1;
   wire c2;
   wire c3;

   carry_lookahead_adder_4bit__3_8 cla0 (.in0({in0[3], in0[2], in0[1], in0[0]}), 
      .in1({in1[3], in1[2], in1[1], in1[0]}), .cin(), .sum({sum[3], sum[2], 
      sum[1], sum[0]}), .cout(c1), .v());
   carry_lookahead_adder_4bit__3_17 cla1 (.in0({in0[7], in0[6], in0[5], in0[4]}), 
      .in1({in1[7], in1[6], in1[5], in1[4]}), .cin(c1), .sum({sum[7], sum[6], 
      sum[5], sum[4]}), .cout(c2), .v());
   carry_lookahead_adder_4bit__3_26 cla2 (.in0({in0[11], in0[10], in0[9], in0[8]}), 
      .in1({in1[11], in1[10], in1[9], in1[8]}), .cin(c2), .sum({sum[11], sum[10], 
      sum[9], sum[8]}), .cout(c3), .v());
   carry_lookahead_adder_4bit__3_35 cla3 (.in0({uc_0, uc_1, uc_2, in0[12]}), 
      .in1({uc_3, uc_4, uc_5, in1[12]}), .cin(c3), .sum({uc_6, uc_7, uc_8, 
      sum[12]}), .cout(), .v());
endmodule

module add_sub_cla__0_1293(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   wire n_0_0;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire [19:0]tempIn11;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire [19:0]tempIn22;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_109;
   wire n_0_110;
   wire n_0_128;
   wire n_0_108;
   wire n_0_107;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_93;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_129;
   wire n_0_98;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_103;
   wire n_0_141;
   wire n_0_142;
   wire n_0_102;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_31;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_80;
   wire n_0_84;
   wire n_0_160;
   wire n_0_79;
   wire n_0_30;
   wire n_0_1;
   wire n_0_15;
   wire n_0_14;
   wire n_0_2;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;

   carry_lookahead_adder_20bit__0_1292 cs0 (.sub(), .in0({uc_0, uc_1, uc_2, uc_3, 
      uc_4, uc_5, uc_6, tempIn11[12], tempIn11[11], tempIn11[10], tempIn11[9], 
      tempIn11[8], tempIn11[7], tempIn11[6], tempIn11[5], tempIn11[4], 
      tempIn11[3], tempIn11[2], tempIn11[1], tempIn11[0]}), .in1({uc_7, uc_8, 
      uc_9, uc_10, uc_11, uc_12, uc_13, tempIn22[12], tempIn22[11], tempIn22[10], 
      tempIn22[9], tempIn22[8], tempIn22[7], tempIn22[6], tempIn22[5], 
      tempIn22[4], tempIn22[3], tempIn22[2], tempIn22[1], tempIn22[0]}), .cin(), 
      .sum({uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, out[12], out[11], 
      out[10], out[9], out[8], out[7], out[6], out[5], out[4], out[3], out[2], 
      out[1], out[0]}), .cout(), .v());
   INV_X1 i_0_0 (.A(in1[13]), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(in2[14]), .ZN(n_0_3));
   NAND2_X1 i_0_2 (.A1(n_0_3), .A2(in1[14]), .ZN(n_0_4));
   INV_X1 i_0_3 (.A(in2[13]), .ZN(n_0_5));
   NAND2_X1 i_0_4 (.A1(n_0_5), .A2(in1[13]), .ZN(n_0_6));
   INV_X1 i_0_5 (.A(in1[14]), .ZN(n_0_7));
   NAND2_X1 i_0_6 (.A1(n_0_7), .A2(in2[14]), .ZN(n_0_8));
   INV_X1 i_0_7 (.A(n_0_8), .ZN(n_0_9));
   OAI21_X1 i_0_8 (.A(n_0_4), .B1(n_0_6), .B2(n_0_9), .ZN(n_0_10));
   AOI22_X1 i_0_9 (.A1(n_0_0), .A2(n_0_15), .B1(n_0_14), .B2(n_0_5), .ZN(out[13]));
   AOI22_X1 i_0_10 (.A1(n_0_7), .A2(n_0_15), .B1(n_0_14), .B2(n_0_3), .ZN(
      out[14]));
   OR2_X1 i_0_18 (.A1(in1[15]), .A2(in2[15]), .ZN(out[15]));
   NAND2_X1 i_0_11 (.A1(n_0_0), .A2(in2[13]), .ZN(n_0_16));
   INV_X1 i_0_12 (.A(n_0_4), .ZN(n_0_17));
   OAI21_X1 i_0_13 (.A(n_0_8), .B1(n_0_16), .B2(n_0_17), .ZN(n_0_18));
   NAND2_X1 i_0_16 (.A1(n_0_18), .A2(n_0_2), .ZN(n_0_19));
   NAND2_X1 i_0_17 (.A1(n_0_19), .A2(n_0_11), .ZN(n_0_20));
   INV_X1 i_0_19 (.A(n_0_20), .ZN(n_0_21));
   AND2_X1 i_0_20 (.A1(n_0_21), .A2(in1[0]), .ZN(tempIn11[0]));
   XNOR2_X1 i_0_21 (.A(n_0_10), .B(n_0_2), .ZN(n_0_22));
   INV_X1 i_0_22 (.A(n_0_22), .ZN(n_0_23));
   NAND2_X1 i_0_23 (.A1(n_0_4), .A2(n_0_8), .ZN(n_0_24));
   XOR2_X1 i_0_24 (.A(n_0_24), .B(n_0_6), .Z(n_0_25));
   NAND4_X1 i_0_25 (.A1(n_0_23), .A2(in1[0]), .A3(n_0_20), .A4(n_0_25), .ZN(
      n_0_26));
   INV_X1 i_0_26 (.A(in1[1]), .ZN(n_0_27));
   OAI21_X1 i_0_27 (.A(n_0_26), .B1(n_0_27), .B2(n_0_20), .ZN(tempIn11[1]));
   NAND2_X1 i_0_28 (.A1(n_0_25), .A2(in1[1]), .ZN(n_0_28));
   INV_X1 i_0_29 (.A(n_0_28), .ZN(n_0_29));
   INV_X1 i_0_30 (.A(n_0_25), .ZN(n_0_32));
   AOI22_X1 i_0_31 (.A1(n_0_25), .A2(in1[2]), .B1(n_0_32), .B2(in1[0]), .ZN(
      n_0_33));
   INV_X1 i_0_32 (.A(n_0_33), .ZN(n_0_34));
   OAI221_X1 i_0_33 (.A(n_0_23), .B1(n_0_29), .B2(n_0_31), .C1(n_0_34), .C2(
      n_0_30), .ZN(n_0_35));
   INV_X1 i_0_34 (.A(in1[2]), .ZN(n_0_36));
   OAI22_X1 i_0_35 (.A1(n_0_35), .A2(n_0_21), .B1(n_0_36), .B2(n_0_20), .ZN(
      tempIn11[2]));
   AOI22_X1 i_0_37 (.A1(n_0_25), .A2(in1[3]), .B1(n_0_32), .B2(in1[1]), .ZN(
      n_0_37));
   OAI33_X1 i_0_38 (.A1(n_0_37), .A2(n_0_30), .A3(n_0_22), .B1(n_0_33), .B2(
      n_0_31), .B3(n_0_22), .ZN(n_0_38));
   AOI22_X1 i_0_39 (.A1(n_0_38), .A2(n_0_20), .B1(in1[3]), .B2(n_0_21), .ZN(
      n_0_39));
   INV_X1 i_0_40 (.A(n_0_39), .ZN(tempIn11[3]));
   OAI21_X1 i_0_41 (.A(n_0_30), .B1(n_0_37), .B2(n_0_22), .ZN(n_0_40));
   AOI22_X1 i_0_42 (.A1(n_0_25), .A2(in1[4]), .B1(n_0_32), .B2(in1[2]), .ZN(
      n_0_41));
   NAND2_X1 i_0_43 (.A1(n_0_25), .A2(in1[0]), .ZN(n_0_42));
   AOI22_X1 i_0_44 (.A1(n_0_41), .A2(n_0_23), .B1(n_0_42), .B2(n_0_22), .ZN(
      n_0_43));
   OAI21_X1 i_0_45 (.A(n_0_40), .B1(n_0_43), .B2(n_0_30), .ZN(n_0_44));
   INV_X1 i_0_46 (.A(in1[4]), .ZN(n_0_45));
   AOI22_X1 i_0_47 (.A1(n_0_44), .A2(n_0_20), .B1(n_0_21), .B2(n_0_45), .ZN(
      tempIn11[4]));
   OAI22_X1 i_0_48 (.A1(n_0_25), .A2(in1[3]), .B1(n_0_32), .B2(in1[5]), .ZN(
      n_0_46));
   AOI22_X1 i_0_49 (.A1(n_0_46), .A2(n_0_23), .B1(n_0_28), .B2(n_0_22), .ZN(
      n_0_47));
   OAI221_X1 i_0_50 (.A(n_0_20), .B1(n_0_47), .B2(n_0_30), .C1(n_0_43), .C2(
      n_0_31), .ZN(n_0_48));
   INV_X1 i_0_51 (.A(in1[5]), .ZN(n_0_49));
   OAI21_X1 i_0_52 (.A(n_0_48), .B1(n_0_49), .B2(n_0_20), .ZN(tempIn11[5]));
   AOI22_X1 i_0_53 (.A1(n_0_25), .A2(in1[6]), .B1(n_0_32), .B2(in1[4]), .ZN(
      n_0_50));
   AOI22_X1 i_0_54 (.A1(n_0_50), .A2(n_0_23), .B1(n_0_33), .B2(n_0_22), .ZN(
      n_0_51));
   AOI221_X1 i_0_55 (.A(n_0_21), .B1(n_0_47), .B2(n_0_30), .C1(n_0_51), .C2(
      n_0_31), .ZN(n_0_52));
   INV_X1 i_0_56 (.A(in1[6]), .ZN(n_0_53));
   AOI21_X1 i_0_57 (.A(n_0_52), .B1(n_0_53), .B2(n_0_21), .ZN(tempIn11[6]));
   AOI22_X1 i_0_58 (.A1(n_0_25), .A2(in1[7]), .B1(n_0_32), .B2(in1[5]), .ZN(
      n_0_54));
   OAI22_X1 i_0_59 (.A1(n_0_37), .A2(n_0_23), .B1(n_0_54), .B2(n_0_22), .ZN(
      n_0_55));
   AOI221_X1 i_0_60 (.A(n_0_21), .B1(n_0_55), .B2(n_0_31), .C1(n_0_51), .C2(
      n_0_30), .ZN(n_0_56));
   INV_X1 i_0_61 (.A(in1[7]), .ZN(n_0_57));
   AOI21_X1 i_0_62 (.A(n_0_56), .B1(n_0_57), .B2(n_0_21), .ZN(tempIn11[7]));
   OAI22_X1 i_0_63 (.A1(n_0_32), .A2(in1[8]), .B1(n_0_25), .B2(in1[6]), .ZN(
      n_0_58));
   OAI22_X1 i_0_64 (.A1(n_0_41), .A2(n_0_23), .B1(n_0_58), .B2(n_0_22), .ZN(
      n_0_59));
   OAI221_X1 i_0_65 (.A(n_0_20), .B1(n_0_59), .B2(n_0_30), .C1(n_0_55), .C2(
      n_0_31), .ZN(n_0_60));
   INV_X1 i_0_66 (.A(in1[8]), .ZN(n_0_61));
   OAI21_X1 i_0_67 (.A(n_0_60), .B1(n_0_61), .B2(n_0_20), .ZN(tempIn11[8]));
   AOI221_X1 i_0_68 (.A(n_0_22), .B1(n_0_25), .B2(in1[9]), .C1(in1[7]), .C2(
      n_0_32), .ZN(n_0_62));
   AOI21_X1 i_0_69 (.A(n_0_62), .B1(n_0_46), .B2(n_0_22), .ZN(n_0_63));
   OAI221_X1 i_0_70 (.A(n_0_20), .B1(n_0_31), .B2(n_0_59), .C1(n_0_63), .C2(
      n_0_30), .ZN(n_0_64));
   INV_X1 i_0_71 (.A(in1[9]), .ZN(n_0_65));
   OAI21_X1 i_0_72 (.A(n_0_64), .B1(n_0_65), .B2(n_0_20), .ZN(tempIn11[9]));
   OAI22_X1 i_0_73 (.A1(n_0_25), .A2(in1[8]), .B1(n_0_32), .B2(in1[10]), 
      .ZN(n_0_66));
   OAI22_X1 i_0_74 (.A1(n_0_50), .A2(n_0_23), .B1(n_0_66), .B2(n_0_22), .ZN(
      n_0_67));
   OAI221_X1 i_0_75 (.A(n_0_20), .B1(n_0_67), .B2(n_0_30), .C1(n_0_63), .C2(
      n_0_31), .ZN(n_0_68));
   INV_X1 i_0_76 (.A(in1[10]), .ZN(n_0_69));
   OAI21_X1 i_0_77 (.A(n_0_68), .B1(n_0_69), .B2(n_0_20), .ZN(tempIn11[10]));
   AOI22_X1 i_0_78 (.A1(n_0_25), .A2(in1[11]), .B1(n_0_32), .B2(in1[9]), 
      .ZN(n_0_70));
   OAI22_X1 i_0_79 (.A1(n_0_54), .A2(n_0_23), .B1(n_0_70), .B2(n_0_22), .ZN(
      n_0_71));
   OAI221_X1 i_0_80 (.A(n_0_20), .B1(n_0_67), .B2(n_0_31), .C1(n_0_71), .C2(
      n_0_30), .ZN(n_0_72));
   INV_X1 i_0_81 (.A(in1[11]), .ZN(n_0_73));
   OAI21_X1 i_0_82 (.A(n_0_72), .B1(n_0_73), .B2(n_0_20), .ZN(tempIn11[11]));
   AOI221_X1 i_0_83 (.A(n_0_22), .B1(n_0_32), .B2(in1[10]), .C1(in1[12]), 
      .C2(n_0_25), .ZN(n_0_74));
   AOI211_X1 i_0_84 (.A(n_0_30), .B(n_0_74), .C1(n_0_58), .C2(n_0_22), .ZN(
      n_0_75));
   AOI211_X1 i_0_85 (.A(n_0_21), .B(n_0_75), .C1(n_0_30), .C2(n_0_71), .ZN(
      n_0_76));
   INV_X1 i_0_86 (.A(in1[12]), .ZN(n_0_77));
   AOI21_X1 i_0_87 (.A(n_0_76), .B1(n_0_77), .B2(n_0_21), .ZN(tempIn11[12]));
   INV_X1 i_0_94 (.A(in2[0]), .ZN(n_0_78));
   NOR2_X1 i_0_95 (.A1(n_0_15), .A2(n_0_78), .ZN(tempIn22[0]));
   NOR3_X1 i_0_98 (.A1(n_0_79), .A2(n_0_80), .A3(n_0_31), .ZN(n_0_81));
   NAND3_X1 i_0_99 (.A1(n_0_81), .A2(in2[0]), .A3(n_0_15), .ZN(n_0_82));
   INV_X1 i_0_100 (.A(in2[1]), .ZN(n_0_83));
   OAI21_X1 i_0_101 (.A(n_0_82), .B1(n_0_83), .B2(n_0_15), .ZN(tempIn22[1]));
   AOI22_X1 i_0_103 (.A1(n_0_80), .A2(in2[0]), .B1(n_0_84), .B2(in2[2]), 
      .ZN(n_0_85));
   NOR2_X1 i_0_104 (.A1(n_0_85), .A2(n_0_79), .ZN(n_0_86));
   AOI221_X1 i_0_105 (.A(n_0_14), .B1(in2[1]), .B2(n_0_81), .C1(n_0_86), 
      .C2(n_0_31), .ZN(n_0_87));
   INV_X1 i_0_106 (.A(in2[2]), .ZN(n_0_88));
   AOI21_X1 i_0_107 (.A(n_0_87), .B1(n_0_88), .B2(n_0_14), .ZN(tempIn22[2]));
   AOI22_X1 i_0_88 (.A1(n_0_84), .A2(in2[3]), .B1(n_0_80), .B2(in2[1]), .ZN(
      n_0_89));
   NOR2_X1 i_0_109 (.A1(n_0_89), .A2(n_0_79), .ZN(n_0_90));
   AOI221_X1 i_0_110 (.A(n_0_14), .B1(n_0_86), .B2(n_0_30), .C1(n_0_31), 
      .C2(n_0_90), .ZN(n_0_91));
   INV_X1 i_0_111 (.A(in2[3]), .ZN(n_0_92));
   AOI21_X1 i_0_112 (.A(n_0_91), .B1(n_0_92), .B2(n_0_14), .ZN(tempIn22[3]));
   NAND2_X1 i_0_114 (.A1(n_0_79), .A2(n_0_84), .ZN(n_0_94));
   OAI22_X1 i_0_115 (.A1(n_0_93), .A2(n_0_79), .B1(n_0_94), .B2(n_0_78), 
      .ZN(n_0_95));
   OAI221_X1 i_0_116 (.A(n_0_15), .B1(n_0_90), .B2(n_0_31), .C1(n_0_95), 
      .C2(n_0_30), .ZN(n_0_96));
   INV_X1 i_0_117 (.A(in2[4]), .ZN(n_0_97));
   OAI21_X1 i_0_118 (.A(n_0_96), .B1(n_0_97), .B2(n_0_15), .ZN(tempIn22[4]));
   OAI22_X1 i_0_120 (.A1(n_0_98), .A2(n_0_79), .B1(n_0_94), .B2(n_0_83), 
      .ZN(n_0_99));
   OAI221_X1 i_0_121 (.A(n_0_15), .B1(n_0_95), .B2(n_0_31), .C1(n_0_30), 
      .C2(n_0_99), .ZN(n_0_100));
   INV_X1 i_0_122 (.A(in2[5]), .ZN(n_0_101));
   OAI21_X1 i_0_123 (.A(n_0_100), .B1(n_0_101), .B2(n_0_15), .ZN(tempIn22[5]));
   OAI22_X1 i_0_126 (.A1(n_0_85), .A2(n_0_102), .B1(n_0_103), .B2(n_0_79), 
      .ZN(n_0_104));
   AOI221_X1 i_0_127 (.A(n_0_14), .B1(n_0_99), .B2(n_0_30), .C1(n_0_104), 
      .C2(n_0_31), .ZN(n_0_105));
   INV_X1 i_0_128 (.A(in2[6]), .ZN(n_0_106));
   AOI21_X1 i_0_129 (.A(n_0_105), .B1(n_0_106), .B2(n_0_14), .ZN(tempIn22[6]));
   AOI221_X1 i_0_132 (.A(n_0_14), .B1(n_0_104), .B2(n_0_30), .C1(n_0_31), 
      .C2(n_0_108), .ZN(n_0_109));
   INV_X1 i_0_133 (.A(in2[7]), .ZN(n_0_110));
   AOI21_X1 i_0_134 (.A(n_0_109), .B1(n_0_110), .B2(n_0_14), .ZN(tempIn22[7]));
   NOR2_X1 i_0_89 (.A1(n_0_84), .A2(in2[10]), .ZN(n_0_128));
   INV_X1 i_0_14 (.A(n_0_113), .ZN(n_0_108));
   AOI21_X1 i_0_15 (.A(n_0_107), .B1(n_0_111), .B2(n_0_15), .ZN(tempIn22[8]));
   NOR2_X1 i_0_90 (.A1(in2[8]), .A2(n_0_15), .ZN(n_0_107));
   OAI21_X1 i_0_36 (.A(n_0_112), .B1(n_0_119), .B2(n_0_30), .ZN(n_0_111));
   NAND2_X1 i_0_96 (.A1(n_0_113), .A2(n_0_30), .ZN(n_0_112));
   OAI21_X1 i_0_91 (.A(n_0_114), .B1(n_0_156), .B2(n_0_79), .ZN(n_0_113));
   NAND2_X1 i_0_92 (.A1(n_0_89), .A2(n_0_79), .ZN(n_0_114));
   OAI21_X1 i_0_93 (.A(n_0_115), .B1(n_0_116), .B2(n_0_14), .ZN(tempIn22[9]));
   NAND2_X1 i_0_97 (.A1(in2[9]), .A2(n_0_14), .ZN(n_0_115));
   AOI21_X1 i_0_102 (.A(n_0_117), .B1(n_0_127), .B2(n_0_31), .ZN(n_0_116));
   INV_X1 i_0_108 (.A(n_0_118), .ZN(n_0_117));
   NAND2_X1 i_0_113 (.A1(n_0_119), .A2(n_0_30), .ZN(n_0_118));
   OAI21_X1 i_0_119 (.A(n_0_120), .B1(n_0_150), .B2(n_0_79), .ZN(n_0_119));
   OR2_X1 i_0_124 (.A1(n_0_93), .A2(n_0_102), .ZN(n_0_120));
   AOI21_X1 i_0_125 (.A(n_0_121), .B1(in2[4]), .B2(n_0_84), .ZN(n_0_93));
   INV_X1 i_0_130 (.A(n_0_122), .ZN(n_0_121));
   NAND2_X1 i_0_131 (.A1(in2[2]), .A2(n_0_80), .ZN(n_0_122));
   OAI21_X1 i_0_139 (.A(n_0_123), .B1(n_0_124), .B2(n_0_14), .ZN(tempIn22[10]));
   NAND2_X1 i_0_140 (.A1(in2[10]), .A2(n_0_14), .ZN(n_0_123));
   AOI21_X1 i_0_141 (.A(n_0_125), .B1(n_0_139), .B2(n_0_31), .ZN(n_0_124));
   INV_X1 i_0_142 (.A(n_0_126), .ZN(n_0_125));
   NAND2_X1 i_0_143 (.A1(n_0_127), .A2(n_0_30), .ZN(n_0_126));
   OAI21_X1 i_0_135 (.A(n_0_129), .B1(n_0_132), .B2(n_0_79), .ZN(n_0_127));
   OR2_X1 i_0_136 (.A1(n_0_98), .A2(n_0_102), .ZN(n_0_129));
   AOI21_X1 i_0_137 (.A(n_0_130), .B1(in2[5]), .B2(n_0_84), .ZN(n_0_98));
   INV_X1 i_0_138 (.A(n_0_131), .ZN(n_0_130));
   NAND2_X1 i_0_144 (.A1(in2[3]), .A2(n_0_80), .ZN(n_0_131));
   AOI21_X1 i_0_145 (.A(n_0_133), .B1(in2[9]), .B2(n_0_84), .ZN(n_0_132));
   INV_X1 i_0_146 (.A(n_0_134), .ZN(n_0_133));
   NAND2_X1 i_0_147 (.A1(in2[7]), .A2(n_0_80), .ZN(n_0_134));
   OAI21_X1 i_0_152 (.A(n_0_135), .B1(n_0_136), .B2(n_0_14), .ZN(tempIn22[11]));
   NAND2_X1 i_0_153 (.A1(in2[11]), .A2(n_0_14), .ZN(n_0_135));
   AOI21_X1 i_0_154 (.A(n_0_137), .B1(n_0_154), .B2(n_0_31), .ZN(n_0_136));
   INV_X1 i_0_155 (.A(n_0_138), .ZN(n_0_137));
   NAND2_X1 i_0_157 (.A1(n_0_139), .A2(n_0_30), .ZN(n_0_138));
   OAI21_X1 i_0_158 (.A(n_0_140), .B1(n_0_143), .B2(n_0_79), .ZN(n_0_139));
   OR2_X1 i_0_159 (.A1(n_0_103), .A2(n_0_102), .ZN(n_0_140));
   AOI21_X1 i_0_160 (.A(n_0_141), .B1(in2[6]), .B2(n_0_84), .ZN(n_0_103));
   INV_X1 i_0_161 (.A(n_0_142), .ZN(n_0_141));
   NAND2_X1 i_0_162 (.A1(in2[4]), .A2(n_0_80), .ZN(n_0_142));
   INV_X1 i_0_148 (.A(n_0_79), .ZN(n_0_102));
   AOI21_X1 i_0_164 (.A(n_0_144), .B1(in2[10]), .B2(n_0_84), .ZN(n_0_143));
   INV_X1 i_0_165 (.A(n_0_145), .ZN(n_0_144));
   NAND2_X1 i_0_166 (.A1(in2[8]), .A2(n_0_80), .ZN(n_0_145));
   INV_X1 i_0_149 (.A(n_0_30), .ZN(n_0_31));
   NOR2_X1 i_0_168 (.A1(n_0_146), .A2(n_0_1), .ZN(tempIn22[12]));
   AOI21_X1 i_0_169 (.A(n_0_147), .B1(n_0_154), .B2(n_0_30), .ZN(n_0_146));
   NAND2_X1 i_0_170 (.A1(n_0_148), .A2(n_0_15), .ZN(n_0_147));
   OAI21_X1 i_0_150 (.A(n_0_149), .B1(n_0_153), .B2(n_0_79), .ZN(n_0_148));
   AOI21_X1 i_0_151 (.A(n_0_30), .B1(n_0_150), .B2(n_0_79), .ZN(n_0_149));
   AOI21_X1 i_0_156 (.A(n_0_151), .B1(in2[8]), .B2(n_0_84), .ZN(n_0_150));
   INV_X1 i_0_163 (.A(n_0_152), .ZN(n_0_151));
   NAND2_X1 i_0_167 (.A1(in2[6]), .A2(n_0_80), .ZN(n_0_152));
   INV_X1 i_0_171 (.A(n_0_128), .ZN(n_0_153));
   OAI21_X1 i_0_177 (.A(n_0_155), .B1(n_0_157), .B2(n_0_79), .ZN(n_0_154));
   NAND2_X1 i_0_178 (.A1(n_0_156), .A2(n_0_79), .ZN(n_0_155));
   MUX2_X1 i_0_172 (.A(in2[7]), .B(in2[5]), .S(n_0_80), .Z(n_0_156));
   AOI21_X1 i_0_180 (.A(n_0_158), .B1(in2[11]), .B2(n_0_84), .ZN(n_0_157));
   INV_X1 i_0_181 (.A(n_0_159), .ZN(n_0_158));
   NAND2_X1 i_0_182 (.A1(in2[9]), .A2(n_0_80), .ZN(n_0_159));
   INV_X1 i_0_173 (.A(n_0_84), .ZN(n_0_80));
   XNOR2_X1 i_0_174 (.A(n_0_24), .B(n_0_160), .ZN(n_0_84));
   INV_X1 i_0_175 (.A(n_0_16), .ZN(n_0_160));
   OAI21_X1 i_0_176 (.A(n_0_19), .B1(n_0_2), .B2(n_0_18), .ZN(n_0_79));
   NAND2_X1 i_0_179 (.A1(n_0_6), .A2(n_0_16), .ZN(n_0_30));
   NOR2_X1 i_0_188 (.A1(in2[12]), .A2(n_0_15), .ZN(n_0_1));
   INV_X1 i_0_183 (.A(n_0_14), .ZN(n_0_15));
   AOI21_X1 i_0_184 (.A(n_0_12), .B1(n_0_10), .B2(n_0_2), .ZN(n_0_14));
   AOI21_X1 i_0_185 (.A(n_0_12), .B1(n_0_13), .B2(in2[15]), .ZN(n_0_2));
   NAND2_X1 i_0_186 (.A1(n_0_13), .A2(in2[15]), .ZN(n_0_11));
   NOR2_X1 i_0_187 (.A1(n_0_13), .A2(in2[15]), .ZN(n_0_12));
   INV_X1 i_0_189 (.A(in1[15]), .ZN(n_0_13));
endmodule

module Euler(INT, CLK, RST, DONE, Interpolate_DONE, Interpolate_Enable, 
      RAM_DATA_RD1, RAM_DATA_RD2, RAM_ADD_RD1, RAM_ADD_RD2, RAM_ADD_WR, 
      RAM_DATA_WR, RAM_ENABLE_WR);
   input INT;
   input CLK;
   input RST;
   output DONE;
   input Interpolate_DONE;
   output Interpolate_Enable;
   input [63:0]RAM_DATA_RD1;
   input [63:0]RAM_DATA_RD2;
   output [12:0]RAM_ADD_RD1;
   output [12:0]RAM_ADD_RD2;
   output [12:0]RAM_ADD_WR;
   output [63:0]RAM_DATA_WR;
   output RAM_ENABLE_WR;

   wire [15:0]NEW_MATRIX_CNT;
   wire [15:0]NEW_VECTOR_CNT;
   wire [15:0]NEW_MATRIX_ADD;
   wire [15:0]NEW_VECTOR2_ADD;
   wire [15:0]NEW_VECTOR_ADD;
   wire [15:0]NEW_RESULT_ADD;
   wire [15:0]h_VECTOR_RESULT;
   wire [15:0]Multiplication_Result;
   wire [15:0]Addition_Result;
   wire [15:0]FINAL_RESULT;
   wire [15:0]Element_Result;
   wire [15:0]RESULT_ADD;
   wire [15:0]VECTOR_ADD;
   wire [15:0]VECTOR2_ADD;
   wire [15:0]MATRIX_ADD;
   wire [15:0]VECTOR_CNT;
   wire [15:0]MATRIX_CNT;
   wire Back;
   wire [2:0]next;
   wire [1:0]counter;
   wire Matrix_Multiplication1_Enable;
   wire Matrix_Multiplication2_Enable;
   wire Final_Calc_Enable;
   wire [63:0]n_val;
   wire [63:0]m_val;
   wire n_0_0;
   wire n_0_0_0;
   wire n_0_1;
   wire n_0_0_1;
   wire n_0_2;
   wire n_0_0_2;
   wire n_0_3;
   wire n_0_0_3;
   wire n_0_4;
   wire n_0_0_4;
   wire n_0_5;
   wire n_0_0_5;
   wire n_0_6;
   wire n_0_0_6;
   wire n_0_7;
   wire n_0_0_7;
   wire n_0_8;
   wire n_0_0_8;
   wire n_0_9;
   wire n_0_0_9;
   wire n_0_10;
   wire n_0_0_10;
   wire n_0_11;
   wire n_0_0_11;
   wire n_0_12;
   wire n_0_0_12;
   wire n_0_13;
   wire n_0_0_13;
   wire n_0_14;
   wire n_0_0_14;
   wire n_0_15;
   wire n_0_0_15;
   wire n_0_16;
   wire n_0_0_16;
   wire n_0_17;
   wire n_0_0_17;
   wire n_0_18;
   wire n_0_0_18;
   wire n_0_19;
   wire n_0_0_19;
   wire n_0_20;
   wire n_0_0_20;
   wire n_0_21;
   wire n_0_0_21;
   wire n_0_22;
   wire n_0_0_22;
   wire n_0_23;
   wire n_0_0_23;
   wire n_0_24;
   wire n_0_0_24;
   wire n_0_25;
   wire n_0_0_25;
   wire n_0_26;
   wire n_0_0_26;
   wire n_0_27;
   wire n_0_0_27;
   wire n_0_28;
   wire n_0_0_28;
   wire n_0_29;
   wire n_0_0_29;
   wire n_0_30;
   wire n_0_0_30;
   wire n_0_31;
   wire n_0_0_31;
   wire n_0_32;
   wire n_0_0_32;
   wire n_0_33;
   wire n_0_0_33;
   wire n_0_34;
   wire n_0_0_34;
   wire n_0_35;
   wire n_0_0_35;
   wire n_0_36;
   wire n_0_0_36;
   wire n_0_37;
   wire n_0_0_37;
   wire n_0_38;
   wire n_0_0_38;
   wire n_0_39;
   wire n_0_0_39;
   wire n_0_40;
   wire n_0_0_40;
   wire n_0_41;
   wire n_0_0_41;
   wire n_0_42;
   wire n_0_0_42;
   wire n_0_43;
   wire n_0_0_43;
   wire n_0_44;
   wire n_0_0_44;
   wire n_0_45;
   wire n_0_0_45;
   wire n_0_46;
   wire n_0_0_46;
   wire n_0_47;
   wire n_0_0_47;
   wire n_0_48;
   wire n_0_0_48;
   wire n_0_49;
   wire n_0_0_49;
   wire n_0_50;
   wire n_0_0_50;
   wire n_0_51;
   wire n_0_0_51;
   wire n_0_52;
   wire n_0_0_52;
   wire n_0_53;
   wire n_0_0_53;
   wire n_0_54;
   wire n_0_0_54;
   wire n_0_55;
   wire n_0_0_55;
   wire n_0_56;
   wire n_0_0_56;
   wire n_0_57;
   wire n_0_0_57;
   wire n_0_58;
   wire n_0_0_58;
   wire n_0_59;
   wire n_0_0_59;
   wire n_0_60;
   wire n_0_0_60;
   wire n_0_61;
   wire n_0_0_61;
   wire n_0_62;
   wire n_0_0_62;
   wire n_0_63;
   wire n_0_0_63;
   wire n_0_64;
   wire n_0_0_64;
   wire n_0_65;
   wire n_0_0_65;
   wire n_0_66;
   wire n_0_0_66;
   wire n_0_67;
   wire n_0_0_67;
   wire n_0_68;
   wire n_0_0_68;
   wire n_0_69;
   wire n_0_0_69;
   wire n_0_70;
   wire n_0_0_70;
   wire n_0_71;
   wire n_0_0_71;
   wire n_0_72;
   wire n_0_0_72;
   wire n_0_73;
   wire n_0_0_73;
   wire n_0_74;
   wire n_0_0_74;
   wire n_0_75;
   wire n_0_0_75;
   wire n_0_76;
   wire n_0_0_76;
   wire n_0_77;
   wire n_0_0_77;
   wire n_0_78;
   wire n_0_0_78;
   wire n_0_79;
   wire n_0_0_79;
   wire n_0_80;
   wire n_0_0_80;
   wire n_0_81;
   wire n_0_0_81;
   wire n_0_82;
   wire n_0_0_82;
   wire n_0_83;
   wire n_0_0_83;
   wire n_0_84;
   wire n_0_0_84;
   wire n_0_85;
   wire n_0_0_85;
   wire n_0_86;
   wire n_0_0_86;
   wire n_0_87;
   wire n_0_0_87;
   wire n_0_88;
   wire n_0_0_88;
   wire n_0_89;
   wire n_0_0_89;
   wire n_0_90;
   wire n_0_0_90;
   wire n_0_91;
   wire n_0_0_91;
   wire n_0_92;
   wire n_0_0_92;
   wire n_0_93;
   wire n_0_0_93;
   wire n_0_94;
   wire n_0_0_94;
   wire n_0_95;
   wire n_0_0_95;
   wire n_0_96;
   wire n_0_0_96;
   wire n_0_97;
   wire n_0_0_97;
   wire n_0_98;
   wire n_0_0_98;
   wire n_0_99;
   wire n_0_0_99;
   wire n_0_100;
   wire n_0_0_100;
   wire n_0_101;
   wire n_0_0_101;
   wire n_0_102;
   wire n_0_0_102;
   wire n_0_103;
   wire n_0_0_103;
   wire n_0_104;
   wire n_0_0_104;
   wire n_0_105;
   wire n_0_0_105;
   wire n_0_106;
   wire n_0_0_106;
   wire n_0_107;
   wire n_0_0_107;
   wire n_0_108;
   wire n_0_0_108;
   wire n_0_109;
   wire n_0_0_109;
   wire n_0_110;
   wire n_0_0_110;
   wire n_0_111;
   wire n_0_0_111;
   wire n_0_112;
   wire n_0_0_112;
   wire n_0_113;
   wire n_0_0_113;
   wire n_0_114;
   wire n_0_0_114;
   wire n_0_115;
   wire n_0_0_115;
   wire n_0_116;
   wire n_0_0_116;
   wire n_0_117;
   wire n_0_0_117;
   wire n_0_118;
   wire n_0_0_118;
   wire n_0_119;
   wire n_0_0_119;
   wire n_0_120;
   wire n_0_0_120;
   wire n_0_121;
   wire n_0_0_121;
   wire n_0_122;
   wire n_0_0_122;
   wire n_0_123;
   wire n_0_0_123;
   wire n_0_124;
   wire n_0_0_124;
   wire n_0_125;
   wire n_0_0_125;
   wire n_0_126;
   wire n_0_0_126;
   wire n_0_127;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_129;
   wire n_0_0_131;
   wire n_0_130;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_131;
   wire n_0_0_134;
   wire n_0_132;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_133;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_134;
   wire n_0_135;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_199;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_137;
   wire n_0_0_267;
   wire n_0_138;
   wire n_0_0_268;
   wire n_0_139;
   wire n_0_0_269;
   wire n_0_140;
   wire n_0_0_270;
   wire n_0_141;
   wire n_0_0_271;
   wire n_0_142;
   wire n_0_0_272;
   wire n_0_143;
   wire n_0_0_273;
   wire n_0_144;
   wire n_0_0_274;
   wire n_0_145;
   wire n_0_0_275;
   wire n_0_146;
   wire n_0_0_276;
   wire n_0_147;
   wire n_0_0_277;
   wire n_0_148;
   wire n_0_0_278;
   wire n_0_149;
   wire n_0_0_279;
   wire n_0_150;
   wire n_0_0_280;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_154;
   wire n_0_0_286;
   wire n_0_155;
   wire n_0_0_287;
   wire n_0_156;
   wire n_0_0_288;
   wire n_0_157;
   wire n_0_0_289;
   wire n_0_158;
   wire n_0_0_290;
   wire n_0_159;
   wire n_0_0_291;
   wire n_0_160;
   wire n_0_0_292;
   wire n_0_161;
   wire n_0_0_293;
   wire n_0_162;
   wire n_0_0_294;
   wire n_0_163;
   wire n_0_0_295;
   wire n_0_164;
   wire n_0_0_296;
   wire n_0_165;
   wire n_0_0_297;
   wire n_0_166;
   wire n_0_0_298;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_170;
   wire n_0_0_304;
   wire n_0_171;
   wire n_0_0_305;
   wire n_0_172;
   wire n_0_0_306;
   wire n_0_173;
   wire n_0_0_307;
   wire n_0_174;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_175;
   wire n_0_0_310;
   wire n_0_176;
   wire n_0_0_311;
   wire n_0_177;
   wire n_0_0_312;
   wire n_0_178;
   wire n_0_0_313;
   wire n_0_179;
   wire n_0_0_314;
   wire n_0_180;
   wire n_0_0_315;
   wire n_0_181;
   wire n_0_0_316;
   wire n_0_182;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_186;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_187;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_188;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_189;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_190;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_191;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_192;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_193;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_194;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_195;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_196;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_197;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_198;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_199;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_200;
   wire n_0_0_365;
   wire n_0_201;
   wire n_0_0_366;
   wire n_0_202;
   wire n_0_0_367;
   wire n_0_203;
   wire n_0_0_368;
   wire n_0_204;
   wire n_0_0_369;
   wire n_0_0_370;
   wire n_0_205;
   wire n_0_0_371;
   wire n_0_206;
   wire n_0_0_372;
   wire n_0_207;
   wire n_0_0_373;
   wire n_0_208;
   wire n_0_0_374;
   wire n_0_209;
   wire n_0_0_375;
   wire n_0_210;
   wire n_0_0_376;
   wire n_0_211;
   wire n_0_0_377;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_0_383;
   wire n_0_212;
   wire n_0_0_384;
   wire n_0_213;
   wire n_0_0_385;
   wire n_0_214;
   wire n_0_0_386;
   wire n_0_215;
   wire n_0_0_387;
   wire n_0_216;
   wire n_0_0_388;
   wire n_0_217;
   wire n_0_0_389;
   wire n_0_218;
   wire n_0_0_390;
   wire n_0_219;
   wire n_0_0_391;
   wire n_0_220;
   wire n_0_0_392;
   wire n_0_221;
   wire n_0_0_393;
   wire n_0_222;
   wire n_0_0_394;
   wire n_0_223;
   wire n_0_0_395;
   wire n_0_224;
   wire n_0_0_396;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_0_402;
   wire n_0_228;
   wire n_0_0_403;
   wire n_0_229;
   wire n_0_0_404;
   wire n_0_230;
   wire n_0_0_405;
   wire n_0_231;
   wire n_0_0_406;
   wire n_0_232;
   wire n_0_0_407;
   wire n_0_233;
   wire n_0_0_408;
   wire n_0_234;
   wire n_0_0_409;
   wire n_0_235;
   wire n_0_0_410;
   wire n_0_236;
   wire n_0_0_411;
   wire n_0_237;
   wire n_0_0_412;
   wire n_0_238;
   wire n_0_0_413;
   wire n_0_239;
   wire n_0_0_414;
   wire n_0_240;
   wire n_0_0_415;
   wire n_0_0_416;
   wire n_0_0_417;
   wire n_0_0_418;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_421;
   wire n_0_0_422;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_0_425;
   wire n_0_0_426;
   wire n_0_0_427;
   wire n_0_0_428;
   wire n_0_0_429;
   wire n_0_241;
   wire n_0_0_430;
   wire n_0_242;
   wire n_0_0_431;
   wire n_0_243;
   wire n_0_0_432;
   wire n_0_244;
   wire n_0_0_433;
   wire n_0_245;
   wire n_0_0_434;
   wire n_0_246;
   wire n_0_0_435;
   wire n_0_247;
   wire n_0_0_436;
   wire n_0_248;
   wire n_0_0_437;
   wire n_0_249;
   wire n_0_0_438;
   wire n_0_250;
   wire n_0_0_439;
   wire n_0_251;
   wire n_0_0_440;
   wire n_0_254;
   wire n_0_0_443;
   wire n_0_255;
   wire n_0_0_444;
   wire n_0_256;
   wire n_0_0_445;
   wire n_0_0_448;
   wire n_0_0_449;
   wire n_0_0_451;
   wire n_0_0_452;
   wire n_0_0_453;
   wire n_0_0_454;
   wire n_0_0_455;
   wire n_0_0_457;
   wire n_0_257;
   wire n_0_0_458;
   wire n_0_258;
   wire n_0_0_459;
   wire n_0_259;
   wire n_0_0_460;
   wire n_0_260;
   wire n_0_0_461;
   wire n_0_261;
   wire n_0_0_462;
   wire n_0_262;
   wire n_0_0_463;
   wire n_0_263;
   wire n_0_0_464;
   wire n_0_264;
   wire n_0_0_465;
   wire n_0_265;
   wire n_0_0_466;
   wire n_0_266;
   wire n_0_0_467;
   wire n_0_267;
   wire n_0_0_468;
   wire n_0_268;
   wire n_0_0_469;
   wire n_0_269;
   wire n_0_0_470;
   wire n_0_270;
   wire n_0_0_471;
   wire n_0_271;
   wire n_0_0_472;
   wire n_0_272;
   wire n_0_0_473;
   wire n_0_0_474;
   wire n_0_0_475;
   wire n_0_0_476;
   wire n_0_273;
   wire n_0_0_477;
   wire n_0_274;
   wire n_0_0_478;
   wire n_0_275;
   wire n_0_0_479;
   wire n_0_276;
   wire n_0_0_480;
   wire n_0_277;
   wire n_0_0_481;
   wire n_0_278;
   wire n_0_0_482;
   wire n_0_279;
   wire n_0_0_483;
   wire n_0_280;
   wire n_0_0_484;
   wire n_0_281;
   wire n_0_0_485;
   wire n_0_282;
   wire n_0_0_486;
   wire n_0_283;
   wire n_0_0_487;
   wire n_0_286;
   wire n_0_0_490;
   wire n_0_287;
   wire n_0_0_491;
   wire n_0_288;
   wire n_0_0_492;
   wire n_0_0_493;
   wire n_0_289;
   wire n_0_290;
   wire n_0_0_495;
   wire n_0_0_496;
   wire n_0_0_497;
   wire n_0_0_498;
   wire n_0_0_499;
   wire n_0_291;
   wire n_0_0_500;
   wire n_0_292;
   wire n_0_0_501;
   wire n_0_293;
   wire n_0_0_502;
   wire n_0_294;
   wire n_0_0_503;
   wire n_0_295;
   wire n_0_0_504;
   wire n_0_296;
   wire n_0_0_505;
   wire n_0_297;
   wire n_0_0_506;
   wire n_0_298;
   wire n_0_0_507;
   wire n_0_299;
   wire n_0_0_508;
   wire n_0_300;
   wire n_0_0_509;
   wire n_0_301;
   wire n_0_0_510;
   wire n_0_302;
   wire n_0_0_511;
   wire n_0_303;
   wire n_0_0_512;
   wire n_0_0_516;
   wire n_0_0_517;
   wire n_0_0_518;
   wire n_0_0_519;
   wire n_0_0_520;
   wire n_0_0_521;
   wire n_0_0_522;
   wire n_0_0_523;
   wire n_0_0_524;
   wire n_0_0_525;
   wire n_0_0_526;
   wire n_0_151;
   wire n_0_0_527;
   wire n_0_152;
   wire n_0_0_528;
   wire n_0_153;
   wire n_0_0_529;
   wire n_0_167;
   wire n_0_0_530;
   wire n_0_168;
   wire n_0_0_531;
   wire n_0_169;
   wire n_0_0_532;
   wire n_0_183;
   wire n_0_0_533;
   wire n_0_184;
   wire n_0_0_534;
   wire n_0_185;
   wire n_0_0_535;
   wire n_0_225;
   wire n_0_0_536;
   wire n_0_226;
   wire n_0_0_537;
   wire n_0_227;
   wire n_0_0_538;
   wire n_0_304;
   wire n_0_0_539;
   wire n_0_0_543;
   wire n_0_0_544;
   wire n_0_0_546;
   wire n_0_0_547;
   wire n_0_0_548;
   wire n_0_0_549;
   wire n_0_0_550;
   wire n_0_0_551;
   wire n_0_0_553;
   wire n_0_0_554;
   wire n_0_0_555;
   wire n_0_0_556;
   wire n_0_0_557;
   wire n_0_0_558;
   wire n_0_0_559;
   wire n_0_0_560;
   wire n_0_0_561;
   wire n_0_0_562;
   wire n_0_0_563;
   wire n_0_305;
   wire n_0_0_564;
   wire n_0_0_565;
   wire n_0_0_566;
   wire n_0_0_567;
   wire n_0_0_568;
   wire n_0_0_569;
   wire n_0_0_570;
   wire n_0_0_571;
   wire n_0_0_572;
   wire n_0_0_573;
   wire n_0_0_574;
   wire n_0_0_575;
   wire n_0_0_576;
   wire n_0_0_577;
   wire n_0_0_578;
   wire n_0_0_579;
   wire n_0_0_580;
   wire n_0_0_581;
   wire n_0_0_582;
   wire n_0_0_583;
   wire n_0_0_584;
   wire n_0_0_585;
   wire n_0_0_586;
   wire n_0_0_587;
   wire n_0_0_588;
   wire n_0_0_589;
   wire n_0_0_590;
   wire n_0_0_591;
   wire n_0_0_592;
   wire n_0_0_593;
   wire n_0_0_594;
   wire n_0_0_595;
   wire n_0_0_598;
   wire n_0_0_599;
   wire n_0_0_600;
   wire n_0_0_601;
   wire n_0_0_602;
   wire n_0_0_603;
   wire n_0_0_605;
   wire n_0_0_606;
   wire n_0_0_607;
   wire n_0_0_608;
   wire n_0_0_609;
   wire n_0_0_610;
   wire n_0_0_611;
   wire n_0_0_612;
   wire n_0_0_613;
   wire n_0_0_614;
   wire n_0_0_615;
   wire n_0_0_616;
   wire n_0_0_617;
   wire n_0_0_618;
   wire n_0_0_619;
   wire n_0_0_620;
   wire n_0_0_621;
   wire n_0_0_622;
   wire n_0_0_624;
   wire n_0_0_625;
   wire n_0_0_626;
   wire n_0_0_627;
   wire n_0_0_628;
   wire n_0_0_630;
   wire n_0_0_631;
   wire n_0_0_632;
   wire n_0_0_633;
   wire n_0_0_634;
   wire n_0_0_636;
   wire n_0_0_637;
   wire n_0_0_638;
   wire n_0_0_142;
   wire n_0_0_146;
   wire n_0_0_149;
   wire n_0_0_157;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_216;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_239;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_255;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_136;
   wire n_0_0_301;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_397;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_456;
   wire n_0_0_513;
   wire n_0_0_635;
   wire n_0_0_623;
   wire n_0_0_596;
   wire n_0_0_604;
   wire n_0_0_514;
   wire n_0_0_515;
   wire n_0_0_540;
   wire n_0_0_541;
   wire n_0_0_542;
   wire n_0_0_597;
   wire n_0_0_629;
   wire n_0_0_321;
   wire n_0_252;
   wire n_0_0_441;
   wire n_0_0_442;
   wire n_0_253;
   wire n_0_0_488;
   wire n_0_0_447;
   wire n_0_0_446;
   wire n_0_0_489;
   wire n_0_0_450;
   wire n_0_284;
   wire n_0_0_639;
   wire n_0_0_640;
   wire n_0_0_641;
   wire n_0_285;
   wire n_0_0_642;
   wire n_0_0_552;
   wire n_0_0_643;
   wire n_0_0_644;
   wire n_0_0_545;
   wire n_0_0_645;
   wire n_0_0_494;
   wire [15:0]NEW_Element_Result;

   assign RAM_DATA_WR[63] = 1'b0;
   assign RAM_DATA_WR[62] = 1'b0;
   assign RAM_DATA_WR[61] = 1'b0;
   assign RAM_DATA_WR[60] = 1'b0;
   assign RAM_DATA_WR[59] = 1'b0;
   assign RAM_DATA_WR[58] = 1'b0;
   assign RAM_DATA_WR[57] = 1'b0;
   assign RAM_DATA_WR[56] = 1'b0;
   assign RAM_DATA_WR[55] = 1'b0;
   assign RAM_DATA_WR[54] = 1'b0;
   assign RAM_DATA_WR[53] = 1'b0;
   assign RAM_DATA_WR[52] = 1'b0;
   assign RAM_DATA_WR[51] = 1'b0;
   assign RAM_DATA_WR[50] = 1'b0;
   assign RAM_DATA_WR[49] = 1'b0;
   assign RAM_DATA_WR[48] = 1'b0;
   assign RAM_DATA_WR[47] = 1'b0;
   assign RAM_DATA_WR[46] = 1'b0;
   assign RAM_DATA_WR[45] = 1'b0;
   assign RAM_DATA_WR[44] = 1'b0;
   assign RAM_DATA_WR[43] = 1'b0;
   assign RAM_DATA_WR[42] = 1'b0;
   assign RAM_DATA_WR[41] = 1'b0;
   assign RAM_DATA_WR[40] = 1'b0;
   assign RAM_DATA_WR[39] = 1'b0;
   assign RAM_DATA_WR[38] = 1'b0;
   assign RAM_DATA_WR[37] = 1'b0;
   assign RAM_DATA_WR[36] = 1'b0;
   assign RAM_DATA_WR[35] = 1'b0;
   assign RAM_DATA_WR[34] = 1'b0;
   assign RAM_DATA_WR[33] = 1'b0;
   assign RAM_DATA_WR[32] = 1'b0;
   assign RAM_DATA_WR[31] = 1'b0;
   assign RAM_DATA_WR[30] = 1'b0;
   assign RAM_DATA_WR[29] = 1'b0;
   assign RAM_DATA_WR[28] = 1'b0;
   assign RAM_DATA_WR[27] = 1'b0;
   assign RAM_DATA_WR[26] = 1'b0;
   assign RAM_DATA_WR[25] = 1'b0;
   assign RAM_DATA_WR[24] = 1'b0;
   assign RAM_DATA_WR[23] = 1'b0;
   assign RAM_DATA_WR[22] = 1'b0;
   assign RAM_DATA_WR[21] = 1'b0;
   assign RAM_DATA_WR[20] = 1'b0;
   assign RAM_DATA_WR[19] = 1'b0;
   assign RAM_DATA_WR[18] = 1'b0;
   assign RAM_DATA_WR[17] = 1'b0;
   assign RAM_DATA_WR[16] = 1'b0;

   add_sub_cla__0_1377__GU MATRIX_CNT_adder (.sub(), .in1({uc_0, uc_1, uc_2, 
      MATRIX_CNT[12], MATRIX_CNT[11], MATRIX_CNT[10], MATRIX_CNT[9], 
      MATRIX_CNT[8], MATRIX_CNT[7], MATRIX_CNT[6], MATRIX_CNT[5], MATRIX_CNT[4], 
      MATRIX_CNT[3], MATRIX_CNT[2], MATRIX_CNT[1], MATRIX_CNT[0]}), .in2(), 
      .cin(), .out({uc_3, uc_4, uc_5, NEW_MATRIX_CNT[12], NEW_MATRIX_CNT[11], 
      NEW_MATRIX_CNT[10], NEW_MATRIX_CNT[9], NEW_MATRIX_CNT[8], 
      NEW_MATRIX_CNT[7], NEW_MATRIX_CNT[6], NEW_MATRIX_CNT[5], NEW_MATRIX_CNT[4], 
      NEW_MATRIX_CNT[3], NEW_MATRIX_CNT[2], NEW_MATRIX_CNT[1], NEW_MATRIX_CNT[0]}), 
      .cout(), .invalid());
   add_sub_cla__0_1321__GU VECTOR_CNT_adder (.sub(), .in1({uc_6, uc_7, uc_8, 
      VECTOR_CNT[12], VECTOR_CNT[11], VECTOR_CNT[10], VECTOR_CNT[9], 
      VECTOR_CNT[8], VECTOR_CNT[7], VECTOR_CNT[6], VECTOR_CNT[5], VECTOR_CNT[4], 
      VECTOR_CNT[3], VECTOR_CNT[2], VECTOR_CNT[1], VECTOR_CNT[0]}), .in2(), 
      .cin(), .out({uc_9, uc_10, uc_11, NEW_VECTOR_CNT[12], NEW_VECTOR_CNT[11], 
      NEW_VECTOR_CNT[10], NEW_VECTOR_CNT[9], NEW_VECTOR_CNT[8], 
      NEW_VECTOR_CNT[7], NEW_VECTOR_CNT[6], NEW_VECTOR_CNT[5], NEW_VECTOR_CNT[4], 
      NEW_VECTOR_CNT[3], NEW_VECTOR_CNT[2], NEW_VECTOR_CNT[1], NEW_VECTOR_CNT[0]}), 
      .cout(), .invalid());
   add_sub_cla__GU MATRIX_ADD_adder (.sub(), .in1({uc_12, uc_13, uc_14, 
      MATRIX_ADD[12], MATRIX_ADD[11], MATRIX_ADD[10], MATRIX_ADD[9], 
      MATRIX_ADD[8], MATRIX_ADD[7], MATRIX_ADD[6], MATRIX_ADD[5], MATRIX_ADD[4], 
      MATRIX_ADD[3], MATRIX_ADD[2], MATRIX_ADD[1], MATRIX_ADD[0]}), .in2(), 
      .cin(), .out({uc_15, uc_16, uc_17, NEW_MATRIX_ADD[12], NEW_MATRIX_ADD[11], 
      NEW_MATRIX_ADD[10], NEW_MATRIX_ADD[9], NEW_MATRIX_ADD[8], 
      NEW_MATRIX_ADD[7], NEW_MATRIX_ADD[6], NEW_MATRIX_ADD[5], NEW_MATRIX_ADD[4], 
      NEW_MATRIX_ADD[3], NEW_MATRIX_ADD[2], NEW_MATRIX_ADD[1], NEW_MATRIX_ADD[0]}), 
      .cout(), .invalid());
   add_sub_cla__0_1433__GU VECTOR2_ADD_adder (.sub(), .in1({uc_18, uc_19, uc_20, 
      VECTOR2_ADD[12], VECTOR2_ADD[11], VECTOR2_ADD[10], VECTOR2_ADD[9], 
      VECTOR2_ADD[8], VECTOR2_ADD[7], VECTOR2_ADD[6], VECTOR2_ADD[5], 
      VECTOR2_ADD[4], VECTOR2_ADD[3], VECTOR2_ADD[2], VECTOR2_ADD[1], 
      VECTOR2_ADD[0]}), .in2(), .cin(), .out({uc_21, uc_22, uc_23, 
      NEW_VECTOR2_ADD[12], NEW_VECTOR2_ADD[11], NEW_VECTOR2_ADD[10], 
      NEW_VECTOR2_ADD[9], NEW_VECTOR2_ADD[8], NEW_VECTOR2_ADD[7], 
      NEW_VECTOR2_ADD[6], NEW_VECTOR2_ADD[5], NEW_VECTOR2_ADD[4], 
      NEW_VECTOR2_ADD[3], NEW_VECTOR2_ADD[2], NEW_VECTOR2_ADD[1], 
      NEW_VECTOR2_ADD[0]}), .cout(), .invalid());
   add_sub_cla__0_1405__GU VECTOR_ADD_adder (.sub(), .in1({uc_24, uc_25, uc_26, 
      VECTOR_ADD[12], VECTOR_ADD[11], VECTOR_ADD[10], VECTOR_ADD[9], 
      VECTOR_ADD[8], VECTOR_ADD[7], VECTOR_ADD[6], VECTOR_ADD[5], VECTOR_ADD[4], 
      VECTOR_ADD[3], VECTOR_ADD[2], VECTOR_ADD[1], VECTOR_ADD[0]}), .in2(), 
      .cin(), .out({uc_27, uc_28, uc_29, NEW_VECTOR_ADD[12], NEW_VECTOR_ADD[11], 
      NEW_VECTOR_ADD[10], NEW_VECTOR_ADD[9], NEW_VECTOR_ADD[8], 
      NEW_VECTOR_ADD[7], NEW_VECTOR_ADD[6], NEW_VECTOR_ADD[5], NEW_VECTOR_ADD[4], 
      NEW_VECTOR_ADD[3], NEW_VECTOR_ADD[2], NEW_VECTOR_ADD[1], NEW_VECTOR_ADD[0]}), 
      .cout(), .invalid());
   add_sub_cla__0_1349__GU RESULT_ADD_adder (.sub(), .in1({uc_30, uc_31, uc_32, 
      RESULT_ADD[12], RESULT_ADD[11], RESULT_ADD[10], RESULT_ADD[9], 
      RESULT_ADD[8], RESULT_ADD[7], RESULT_ADD[6], RESULT_ADD[5], RESULT_ADD[4], 
      RESULT_ADD[3], RESULT_ADD[2], RESULT_ADD[1], RESULT_ADD[0]}), .in2(), 
      .cin(), .out({uc_33, uc_34, uc_35, NEW_RESULT_ADD[12], NEW_RESULT_ADD[11], 
      NEW_RESULT_ADD[10], NEW_RESULT_ADD[9], NEW_RESULT_ADD[8], 
      NEW_RESULT_ADD[7], NEW_RESULT_ADD[6], NEW_RESULT_ADD[5], NEW_RESULT_ADD[4], 
      NEW_RESULT_ADD[3], NEW_RESULT_ADD[2], NEW_RESULT_ADD[1], NEW_RESULT_ADD[0]}), 
      .cout(), .invalid());
   multiplier_16bit__0_1434 h_MUL (.first_operand(Addition_Result), 
      .second_operand({n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, 
      n_11, n_12, n_13, n_14, n_15}), .out(h_VECTOR_RESULT), .enable(), 
      .overflow());
   multiplier_16bit MUL (.first_operand({RAM_DATA_RD1[15], RAM_DATA_RD1[14], 
      RAM_DATA_RD1[13], RAM_DATA_RD1[12], RAM_DATA_RD1[11], RAM_DATA_RD1[10], 
      RAM_DATA_RD1[9], RAM_DATA_RD1[8], RAM_DATA_RD1[7], RAM_DATA_RD1[6], 
      RAM_DATA_RD1[5], RAM_DATA_RD1[4], RAM_DATA_RD1[3], RAM_DATA_RD1[2], 
      RAM_DATA_RD1[1], RAM_DATA_RD1[0]}), .second_operand({RAM_DATA_RD2[15], 
      RAM_DATA_RD2[14], RAM_DATA_RD2[13], RAM_DATA_RD2[12], RAM_DATA_RD2[11], 
      RAM_DATA_RD2[10], RAM_DATA_RD2[9], RAM_DATA_RD2[8], RAM_DATA_RD2[7], 
      RAM_DATA_RD2[6], RAM_DATA_RD2[5], RAM_DATA_RD2[4], RAM_DATA_RD2[3], 
      RAM_DATA_RD2[2], RAM_DATA_RD2[1], RAM_DATA_RD2[0]}), .out(
      Multiplication_Result), .enable(), .overflow());
   add_sub_cla__3_99 VEC1_VEC2_adder (.sub(), .in1({RAM_DATA_RD1[15], 
      RAM_DATA_RD1[14], RAM_DATA_RD1[13], RAM_DATA_RD1[12], RAM_DATA_RD1[11], 
      RAM_DATA_RD1[10], RAM_DATA_RD1[9], RAM_DATA_RD1[8], RAM_DATA_RD1[7], 
      RAM_DATA_RD1[6], RAM_DATA_RD1[5], RAM_DATA_RD1[4], RAM_DATA_RD1[3], 
      RAM_DATA_RD1[2], RAM_DATA_RD1[1], RAM_DATA_RD1[0]}), .in2({
      RAM_DATA_RD2[15], RAM_DATA_RD2[14], RAM_DATA_RD2[13], RAM_DATA_RD2[12], 
      RAM_DATA_RD2[11], RAM_DATA_RD2[10], RAM_DATA_RD2[9], RAM_DATA_RD2[8], 
      RAM_DATA_RD2[7], RAM_DATA_RD2[6], RAM_DATA_RD2[5], RAM_DATA_RD2[4], 
      RAM_DATA_RD2[3], RAM_DATA_RD2[2], RAM_DATA_RD2[1], RAM_DATA_RD2[0]}), 
      .cin(), .out(Addition_Result), .cout(), .invalid());
   add_sub_cla__3_163 FINAL_RESULT_adder (.sub(), .in1(h_VECTOR_RESULT), 
      .in2(Element_Result), .cin(), .out(FINAL_RESULT), .cout(), .invalid());
   DFF_X1 RAM_ENABLE_WR_reg (.D(n_0_305), .CK(n_0_136), .Q(RAM_ENABLE_WR), .QN());
   DFF_X1 \RAM_DATA_WR_reg[15]  (.D(n_0_288), .CK(n_0_136), .Q(RAM_DATA_WR[15]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[14]  (.D(n_0_287), .CK(n_0_136), .Q(RAM_DATA_WR[14]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[13]  (.D(n_0_286), .CK(n_0_136), .Q(RAM_DATA_WR[13]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[12]  (.D(n_0_285), .CK(n_0_136), .Q(RAM_DATA_WR[12]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[11]  (.D(n_0_284), .CK(n_0_136), .Q(RAM_DATA_WR[11]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[10]  (.D(n_0_283), .CK(n_0_136), .Q(RAM_DATA_WR[10]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[9]  (.D(n_0_282), .CK(n_0_136), .Q(RAM_DATA_WR[9]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[8]  (.D(n_0_281), .CK(n_0_136), .Q(RAM_DATA_WR[8]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[7]  (.D(n_0_280), .CK(n_0_136), .Q(RAM_DATA_WR[7]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[6]  (.D(n_0_279), .CK(n_0_136), .Q(RAM_DATA_WR[6]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[5]  (.D(n_0_278), .CK(n_0_136), .Q(RAM_DATA_WR[5]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[4]  (.D(n_0_277), .CK(n_0_136), .Q(RAM_DATA_WR[4]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[3]  (.D(n_0_276), .CK(n_0_136), .Q(RAM_DATA_WR[3]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[2]  (.D(n_0_275), .CK(n_0_136), .Q(RAM_DATA_WR[2]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[1]  (.D(n_0_274), .CK(n_0_136), .Q(RAM_DATA_WR[1]), 
      .QN());
   DFF_X1 \RAM_DATA_WR_reg[0]  (.D(n_0_273), .CK(n_0_136), .Q(RAM_DATA_WR[0]), 
      .QN());
   DFF_X1 \h_val_reg[15]  (.D(n_0_272), .CK(n_0_136), .Q(n_0), .QN());
   DFF_X1 \h_val_reg[14]  (.D(n_0_271), .CK(n_0_136), .Q(n_1), .QN());
   DFF_X1 \h_val_reg[13]  (.D(n_0_270), .CK(n_0_136), .Q(n_2), .QN());
   DFF_X1 \h_val_reg[12]  (.D(n_0_269), .CK(n_0_136), .Q(n_3), .QN());
   DFF_X1 \h_val_reg[11]  (.D(n_0_268), .CK(n_0_136), .Q(n_4), .QN());
   DFF_X1 \h_val_reg[10]  (.D(n_0_267), .CK(n_0_136), .Q(n_5), .QN());
   DFF_X1 \h_val_reg[9]  (.D(n_0_266), .CK(n_0_136), .Q(n_6), .QN());
   DFF_X1 \h_val_reg[8]  (.D(n_0_265), .CK(n_0_136), .Q(n_7), .QN());
   DFF_X1 \h_val_reg[7]  (.D(n_0_264), .CK(n_0_136), .Q(n_8), .QN());
   DFF_X1 \h_val_reg[6]  (.D(n_0_263), .CK(n_0_136), .Q(n_9), .QN());
   DFF_X1 \h_val_reg[5]  (.D(n_0_262), .CK(n_0_136), .Q(n_10), .QN());
   DFF_X1 \h_val_reg[4]  (.D(n_0_261), .CK(n_0_136), .Q(n_11), .QN());
   DFF_X1 \h_val_reg[3]  (.D(n_0_260), .CK(n_0_136), .Q(n_12), .QN());
   DFF_X1 \h_val_reg[2]  (.D(n_0_259), .CK(n_0_136), .Q(n_13), .QN());
   DFF_X1 \h_val_reg[1]  (.D(n_0_258), .CK(n_0_136), .Q(n_14), .QN());
   DFF_X1 \h_val_reg[0]  (.D(n_0_257), .CK(n_0_136), .Q(n_15), .QN());
   DFF_X1 \Element_Result_reg[15]  (.D(n_0_256), .CK(n_0_136), .Q(
      Element_Result[15]), .QN());
   DFF_X1 \Element_Result_reg[14]  (.D(n_0_255), .CK(n_0_136), .Q(
      Element_Result[14]), .QN());
   DFF_X1 \Element_Result_reg[13]  (.D(n_0_254), .CK(n_0_136), .Q(
      Element_Result[13]), .QN());
   DFF_X1 \Element_Result_reg[12]  (.D(n_0_253), .CK(n_0_136), .Q(
      Element_Result[12]), .QN());
   DFF_X1 \Element_Result_reg[11]  (.D(n_0_252), .CK(n_0_136), .Q(
      Element_Result[11]), .QN());
   DFF_X1 \Element_Result_reg[10]  (.D(n_0_251), .CK(n_0_136), .Q(
      Element_Result[10]), .QN());
   DFF_X1 \Element_Result_reg[9]  (.D(n_0_250), .CK(n_0_136), .Q(
      Element_Result[9]), .QN());
   DFF_X1 \Element_Result_reg[8]  (.D(n_0_249), .CK(n_0_136), .Q(
      Element_Result[8]), .QN());
   DFF_X1 \Element_Result_reg[7]  (.D(n_0_248), .CK(n_0_136), .Q(
      Element_Result[7]), .QN());
   DFF_X1 \Element_Result_reg[6]  (.D(n_0_247), .CK(n_0_136), .Q(
      Element_Result[6]), .QN());
   DFF_X1 \Element_Result_reg[5]  (.D(n_0_246), .CK(n_0_136), .Q(
      Element_Result[5]), .QN());
   DFF_X1 \Element_Result_reg[4]  (.D(n_0_245), .CK(n_0_136), .Q(
      Element_Result[4]), .QN());
   DFF_X1 \Element_Result_reg[3]  (.D(n_0_244), .CK(n_0_136), .Q(
      Element_Result[3]), .QN());
   DFF_X1 \Element_Result_reg[2]  (.D(n_0_243), .CK(n_0_136), .Q(
      Element_Result[2]), .QN());
   DFF_X1 \Element_Result_reg[1]  (.D(n_0_242), .CK(n_0_136), .Q(
      Element_Result[1]), .QN());
   DFF_X1 \Element_Result_reg[0]  (.D(n_0_241), .CK(n_0_136), .Q(
      Element_Result[0]), .QN());
   DFF_X1 \RAM_ADD_WR_reg[12]  (.D(n_0_240), .CK(n_0_136), .Q(RAM_ADD_WR[12]), 
      .QN());
   DFF_X1 \RAM_ADD_WR_reg[11]  (.D(n_0_239), .CK(n_0_136), .Q(RAM_ADD_WR[11]), 
      .QN());
   DFF_X1 \RAM_ADD_WR_reg[10]  (.D(n_0_238), .CK(n_0_136), .Q(RAM_ADD_WR[10]), 
      .QN());
   DFF_X1 \RAM_ADD_WR_reg[9]  (.D(n_0_237), .CK(n_0_136), .Q(RAM_ADD_WR[9]), 
      .QN());
   DFF_X1 \RAM_ADD_WR_reg[8]  (.D(n_0_236), .CK(n_0_136), .Q(RAM_ADD_WR[8]), 
      .QN());
   DFF_X1 \RAM_ADD_WR_reg[7]  (.D(n_0_235), .CK(n_0_136), .Q(RAM_ADD_WR[7]), 
      .QN());
   DFF_X1 \RAM_ADD_WR_reg[6]  (.D(n_0_234), .CK(n_0_136), .Q(RAM_ADD_WR[6]), 
      .QN());
   DFF_X1 \RAM_ADD_WR_reg[5]  (.D(n_0_233), .CK(n_0_136), .Q(RAM_ADD_WR[5]), 
      .QN());
   DFF_X1 \RAM_ADD_WR_reg[4]  (.D(n_0_232), .CK(n_0_136), .Q(RAM_ADD_WR[4]), 
      .QN());
   DFF_X1 \RAM_ADD_WR_reg[3]  (.D(n_0_231), .CK(n_0_136), .Q(RAM_ADD_WR[3]), 
      .QN());
   DFF_X1 \RAM_ADD_WR_reg[2]  (.D(n_0_230), .CK(n_0_136), .Q(RAM_ADD_WR[2]), 
      .QN());
   DFF_X1 \RAM_ADD_WR_reg[1]  (.D(n_0_229), .CK(n_0_136), .Q(RAM_ADD_WR[1]), 
      .QN());
   DFF_X1 \RAM_ADD_WR_reg[0]  (.D(n_0_228), .CK(n_0_136), .Q(RAM_ADD_WR[0]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[12]  (.D(n_0_224), .CK(n_0_136), .Q(RESULT_ADD[12]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[11]  (.D(n_0_223), .CK(n_0_136), .Q(RESULT_ADD[11]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[10]  (.D(n_0_222), .CK(n_0_136), .Q(RESULT_ADD[10]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[9]  (.D(n_0_221), .CK(n_0_136), .Q(RESULT_ADD[9]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[8]  (.D(n_0_220), .CK(n_0_136), .Q(RESULT_ADD[8]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[7]  (.D(n_0_219), .CK(n_0_136), .Q(RESULT_ADD[7]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[6]  (.D(n_0_218), .CK(n_0_136), .Q(RESULT_ADD[6]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[5]  (.D(n_0_217), .CK(n_0_136), .Q(RESULT_ADD[5]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[4]  (.D(n_0_216), .CK(n_0_136), .Q(RESULT_ADD[4]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[3]  (.D(n_0_215), .CK(n_0_136), .Q(RESULT_ADD[3]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[2]  (.D(n_0_214), .CK(n_0_136), .Q(RESULT_ADD[2]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[1]  (.D(n_0_213), .CK(n_0_136), .Q(RESULT_ADD[1]), 
      .QN());
   DFF_X1 \RESULT_ADD_reg[0]  (.D(n_0_212), .CK(n_0_136), .Q(RESULT_ADD[0]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[12]  (.D(n_0_211), .CK(n_0_136), .Q(RAM_ADD_RD2[12]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[11]  (.D(n_0_210), .CK(n_0_136), .Q(RAM_ADD_RD2[11]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[10]  (.D(n_0_209), .CK(n_0_136), .Q(RAM_ADD_RD2[10]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[9]  (.D(n_0_208), .CK(n_0_136), .Q(RAM_ADD_RD2[9]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[8]  (.D(n_0_207), .CK(n_0_136), .Q(RAM_ADD_RD2[8]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[7]  (.D(n_0_206), .CK(n_0_136), .Q(RAM_ADD_RD2[7]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[6]  (.D(n_0_205), .CK(n_0_136), .Q(RAM_ADD_RD2[6]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[5]  (.D(n_0_204), .CK(n_0_136), .Q(RAM_ADD_RD2[5]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[4]  (.D(n_0_203), .CK(n_0_136), .Q(RAM_ADD_RD2[4]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[3]  (.D(n_0_202), .CK(n_0_136), .Q(RAM_ADD_RD2[3]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[2]  (.D(n_0_201), .CK(n_0_136), .Q(RAM_ADD_RD2[2]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[1]  (.D(n_0_200), .CK(n_0_136), .Q(RAM_ADD_RD2[1]), 
      .QN());
   DFF_X1 \RAM_ADD_RD2_reg[0]  (.D(n_0_199), .CK(n_0_136), .Q(RAM_ADD_RD2[0]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[12]  (.D(n_0_198), .CK(n_0_136), .Q(RAM_ADD_RD1[12]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[11]  (.D(n_0_197), .CK(n_0_136), .Q(RAM_ADD_RD1[11]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[10]  (.D(n_0_196), .CK(n_0_136), .Q(RAM_ADD_RD1[10]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[9]  (.D(n_0_195), .CK(n_0_136), .Q(RAM_ADD_RD1[9]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[8]  (.D(n_0_194), .CK(n_0_136), .Q(RAM_ADD_RD1[8]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[7]  (.D(n_0_193), .CK(n_0_136), .Q(RAM_ADD_RD1[7]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[6]  (.D(n_0_192), .CK(n_0_136), .Q(RAM_ADD_RD1[6]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[5]  (.D(n_0_191), .CK(n_0_136), .Q(RAM_ADD_RD1[5]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[4]  (.D(n_0_190), .CK(n_0_136), .Q(RAM_ADD_RD1[4]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[3]  (.D(n_0_189), .CK(n_0_136), .Q(RAM_ADD_RD1[3]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[2]  (.D(n_0_188), .CK(n_0_136), .Q(RAM_ADD_RD1[2]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[1]  (.D(n_0_187), .CK(n_0_136), .Q(RAM_ADD_RD1[1]), 
      .QN());
   DFF_X1 \RAM_ADD_RD1_reg[0]  (.D(n_0_186), .CK(n_0_136), .Q(RAM_ADD_RD1[0]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[12]  (.D(n_0_182), .CK(n_0_136), .Q(VECTOR_ADD[12]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[11]  (.D(n_0_181), .CK(n_0_136), .Q(VECTOR_ADD[11]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[10]  (.D(n_0_180), .CK(n_0_136), .Q(VECTOR_ADD[10]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[9]  (.D(n_0_179), .CK(n_0_136), .Q(VECTOR_ADD[9]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[8]  (.D(n_0_178), .CK(n_0_136), .Q(VECTOR_ADD[8]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[7]  (.D(n_0_177), .CK(n_0_136), .Q(VECTOR_ADD[7]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[6]  (.D(n_0_176), .CK(n_0_136), .Q(VECTOR_ADD[6]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[5]  (.D(n_0_175), .CK(n_0_136), .Q(VECTOR_ADD[5]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[4]  (.D(n_0_174), .CK(n_0_136), .Q(VECTOR_ADD[4]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[3]  (.D(n_0_173), .CK(n_0_136), .Q(VECTOR_ADD[3]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[2]  (.D(n_0_172), .CK(n_0_136), .Q(VECTOR_ADD[2]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[1]  (.D(n_0_171), .CK(n_0_136), .Q(VECTOR_ADD[1]), 
      .QN());
   DFF_X1 \VECTOR_ADD_reg[0]  (.D(n_0_170), .CK(n_0_136), .Q(VECTOR_ADD[0]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[12]  (.D(n_0_166), .CK(n_0_136), .Q(VECTOR2_ADD[12]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[11]  (.D(n_0_165), .CK(n_0_136), .Q(VECTOR2_ADD[11]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[10]  (.D(n_0_164), .CK(n_0_136), .Q(VECTOR2_ADD[10]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[9]  (.D(n_0_163), .CK(n_0_136), .Q(VECTOR2_ADD[9]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[8]  (.D(n_0_162), .CK(n_0_136), .Q(VECTOR2_ADD[8]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[7]  (.D(n_0_161), .CK(n_0_136), .Q(VECTOR2_ADD[7]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[6]  (.D(n_0_160), .CK(n_0_136), .Q(VECTOR2_ADD[6]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[5]  (.D(n_0_159), .CK(n_0_136), .Q(VECTOR2_ADD[5]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[4]  (.D(n_0_158), .CK(n_0_136), .Q(VECTOR2_ADD[4]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[3]  (.D(n_0_157), .CK(n_0_136), .Q(VECTOR2_ADD[3]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[2]  (.D(n_0_156), .CK(n_0_136), .Q(VECTOR2_ADD[2]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[1]  (.D(n_0_155), .CK(n_0_136), .Q(VECTOR2_ADD[1]), 
      .QN());
   DFF_X1 \VECTOR2_ADD_reg[0]  (.D(n_0_154), .CK(n_0_136), .Q(VECTOR2_ADD[0]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[12]  (.D(n_0_150), .CK(n_0_136), .Q(MATRIX_ADD[12]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[11]  (.D(n_0_149), .CK(n_0_136), .Q(MATRIX_ADD[11]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[10]  (.D(n_0_148), .CK(n_0_136), .Q(MATRIX_ADD[10]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[9]  (.D(n_0_147), .CK(n_0_136), .Q(MATRIX_ADD[9]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[8]  (.D(n_0_146), .CK(n_0_136), .Q(MATRIX_ADD[8]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[7]  (.D(n_0_145), .CK(n_0_136), .Q(MATRIX_ADD[7]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[6]  (.D(n_0_144), .CK(n_0_136), .Q(MATRIX_ADD[6]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[5]  (.D(n_0_143), .CK(n_0_136), .Q(MATRIX_ADD[5]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[4]  (.D(n_0_142), .CK(n_0_136), .Q(MATRIX_ADD[4]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[3]  (.D(n_0_141), .CK(n_0_136), .Q(MATRIX_ADD[3]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[2]  (.D(n_0_140), .CK(n_0_136), .Q(MATRIX_ADD[2]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[1]  (.D(n_0_139), .CK(n_0_136), .Q(MATRIX_ADD[1]), 
      .QN());
   DFF_X1 \MATRIX_ADD_reg[0]  (.D(n_0_138), .CK(n_0_136), .Q(MATRIX_ADD[0]), 
      .QN());
   DFF_X1 Interpolate_Enable_reg (.D(n_0_137), .CK(n_0_136), .Q(
      Interpolate_Enable), .QN());
   DFF_X1 DONE_reg (.D(n_0_289), .CK(n_0_136), .Q(DONE), .QN());
   DFF_X1 \VECTOR_CNT_reg[12]  (.D(n_0_304), .CK(n_0_136), .Q(VECTOR_CNT[12]), 
      .QN());
   DFF_X1 \VECTOR_CNT_reg[11]  (.D(n_0_227), .CK(n_0_136), .Q(VECTOR_CNT[11]), 
      .QN());
   DFF_X1 \VECTOR_CNT_reg[10]  (.D(n_0_226), .CK(n_0_136), .Q(VECTOR_CNT[10]), 
      .QN());
   DFF_X1 \VECTOR_CNT_reg[9]  (.D(n_0_225), .CK(n_0_136), .Q(VECTOR_CNT[9]), 
      .QN());
   DFF_X1 \VECTOR_CNT_reg[8]  (.D(n_0_185), .CK(n_0_136), .Q(VECTOR_CNT[8]), 
      .QN());
   DFF_X1 \VECTOR_CNT_reg[7]  (.D(n_0_184), .CK(n_0_136), .Q(VECTOR_CNT[7]), 
      .QN());
   DFF_X1 \VECTOR_CNT_reg[6]  (.D(n_0_183), .CK(n_0_136), .Q(VECTOR_CNT[6]), 
      .QN());
   DFF_X1 \VECTOR_CNT_reg[5]  (.D(n_0_169), .CK(n_0_136), .Q(VECTOR_CNT[5]), 
      .QN());
   DFF_X1 \VECTOR_CNT_reg[4]  (.D(n_0_168), .CK(n_0_136), .Q(VECTOR_CNT[4]), 
      .QN());
   DFF_X1 \VECTOR_CNT_reg[3]  (.D(n_0_167), .CK(n_0_136), .Q(VECTOR_CNT[3]), 
      .QN());
   DFF_X1 \VECTOR_CNT_reg[2]  (.D(n_0_153), .CK(n_0_136), .Q(VECTOR_CNT[2]), 
      .QN());
   DFF_X1 \VECTOR_CNT_reg[1]  (.D(n_0_152), .CK(n_0_136), .Q(VECTOR_CNT[1]), 
      .QN());
   DFF_X1 \VECTOR_CNT_reg[0]  (.D(n_0_151), .CK(n_0_136), .Q(VECTOR_CNT[0]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[12]  (.D(n_0_303), .CK(n_0_136), .Q(MATRIX_CNT[12]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[11]  (.D(n_0_302), .CK(n_0_136), .Q(MATRIX_CNT[11]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[10]  (.D(n_0_301), .CK(n_0_136), .Q(MATRIX_CNT[10]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[9]  (.D(n_0_300), .CK(n_0_136), .Q(MATRIX_CNT[9]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[8]  (.D(n_0_299), .CK(n_0_136), .Q(MATRIX_CNT[8]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[7]  (.D(n_0_298), .CK(n_0_136), .Q(MATRIX_CNT[7]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[6]  (.D(n_0_297), .CK(n_0_136), .Q(MATRIX_CNT[6]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[5]  (.D(n_0_296), .CK(n_0_136), .Q(MATRIX_CNT[5]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[4]  (.D(n_0_295), .CK(n_0_136), .Q(MATRIX_CNT[4]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[3]  (.D(n_0_294), .CK(n_0_136), .Q(MATRIX_CNT[3]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[2]  (.D(n_0_293), .CK(n_0_136), .Q(MATRIX_CNT[2]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[1]  (.D(n_0_292), .CK(n_0_136), .Q(MATRIX_CNT[1]), 
      .QN());
   DFF_X1 \MATRIX_CNT_reg[0]  (.D(n_0_291), .CK(n_0_136), .Q(MATRIX_CNT[0]), 
      .QN());
   DFF_X1 Back_reg (.D(n_0_290), .CK(n_0_136), .Q(Back), .QN());
   DFF_X1 \next_reg[2]  (.D(n_0_135), .CK(n_0_136), .Q(next[2]), .QN());
   DFF_X1 \next_reg[1]  (.D(n_0_134), .CK(n_0_136), .Q(next[1]), .QN());
   DFF_X1 \next_reg[0]  (.D(n_0_133), .CK(n_0_136), .Q(next[0]), .QN());
   DFF_X1 \counter_reg[1]  (.D(n_0_132), .CK(n_0_136), .Q(counter[1]), .QN());
   DFF_X1 \counter_reg[0]  (.D(n_0_131), .CK(n_0_136), .Q(counter[0]), .QN());
   DFF_X1 Matrix_Multiplication1_Enable_reg (.D(n_0_130), .CK(n_0_136), .Q(
      Matrix_Multiplication1_Enable), .QN());
   DFF_X1 Matrix_Multiplication2_Enable_reg (.D(n_0_129), .CK(n_0_136), .Q(
      Matrix_Multiplication2_Enable), .QN());
   DFF_X1 Final_Calc_Enable_reg (.D(n_0_128), .CK(n_0_136), .Q(Final_Calc_Enable), 
      .QN());
   DFF_X1 \n_val_reg[63]  (.D(n_0_127), .CK(n_0_136), .Q(n_val[63]), .QN());
   DFF_X1 \n_val_reg[62]  (.D(n_0_126), .CK(n_0_136), .Q(n_val[62]), .QN());
   DFF_X1 \n_val_reg[61]  (.D(n_0_125), .CK(n_0_136), .Q(n_val[61]), .QN());
   DFF_X1 \n_val_reg[60]  (.D(n_0_124), .CK(n_0_136), .Q(n_val[60]), .QN());
   DFF_X1 \n_val_reg[59]  (.D(n_0_123), .CK(n_0_136), .Q(n_val[59]), .QN());
   DFF_X1 \n_val_reg[58]  (.D(n_0_122), .CK(n_0_136), .Q(n_val[58]), .QN());
   DFF_X1 \n_val_reg[57]  (.D(n_0_121), .CK(n_0_136), .Q(n_val[57]), .QN());
   DFF_X1 \n_val_reg[56]  (.D(n_0_120), .CK(n_0_136), .Q(n_val[56]), .QN());
   DFF_X1 \n_val_reg[55]  (.D(n_0_119), .CK(n_0_136), .Q(n_val[55]), .QN());
   DFF_X1 \n_val_reg[54]  (.D(n_0_118), .CK(n_0_136), .Q(n_val[54]), .QN());
   DFF_X1 \n_val_reg[53]  (.D(n_0_117), .CK(n_0_136), .Q(n_val[53]), .QN());
   DFF_X1 \n_val_reg[52]  (.D(n_0_116), .CK(n_0_136), .Q(n_val[52]), .QN());
   DFF_X1 \n_val_reg[51]  (.D(n_0_115), .CK(n_0_136), .Q(n_val[51]), .QN());
   DFF_X1 \n_val_reg[50]  (.D(n_0_114), .CK(n_0_136), .Q(n_val[50]), .QN());
   DFF_X1 \n_val_reg[49]  (.D(n_0_113), .CK(n_0_136), .Q(n_val[49]), .QN());
   DFF_X1 \n_val_reg[48]  (.D(n_0_112), .CK(n_0_136), .Q(n_val[48]), .QN());
   DFF_X1 \n_val_reg[47]  (.D(n_0_111), .CK(n_0_136), .Q(n_val[47]), .QN());
   DFF_X1 \n_val_reg[46]  (.D(n_0_110), .CK(n_0_136), .Q(n_val[46]), .QN());
   DFF_X1 \n_val_reg[45]  (.D(n_0_109), .CK(n_0_136), .Q(n_val[45]), .QN());
   DFF_X1 \n_val_reg[44]  (.D(n_0_108), .CK(n_0_136), .Q(n_val[44]), .QN());
   DFF_X1 \n_val_reg[43]  (.D(n_0_107), .CK(n_0_136), .Q(n_val[43]), .QN());
   DFF_X1 \n_val_reg[42]  (.D(n_0_106), .CK(n_0_136), .Q(n_val[42]), .QN());
   DFF_X1 \n_val_reg[41]  (.D(n_0_105), .CK(n_0_136), .Q(n_val[41]), .QN());
   DFF_X1 \n_val_reg[40]  (.D(n_0_104), .CK(n_0_136), .Q(n_val[40]), .QN());
   DFF_X1 \n_val_reg[39]  (.D(n_0_103), .CK(n_0_136), .Q(n_val[39]), .QN());
   DFF_X1 \n_val_reg[38]  (.D(n_0_102), .CK(n_0_136), .Q(n_val[38]), .QN());
   DFF_X1 \n_val_reg[37]  (.D(n_0_101), .CK(n_0_136), .Q(n_val[37]), .QN());
   DFF_X1 \n_val_reg[36]  (.D(n_0_100), .CK(n_0_136), .Q(n_val[36]), .QN());
   DFF_X1 \n_val_reg[35]  (.D(n_0_99), .CK(n_0_136), .Q(n_val[35]), .QN());
   DFF_X1 \n_val_reg[34]  (.D(n_0_98), .CK(n_0_136), .Q(n_val[34]), .QN());
   DFF_X1 \n_val_reg[33]  (.D(n_0_97), .CK(n_0_136), .Q(n_val[33]), .QN());
   DFF_X1 \n_val_reg[32]  (.D(n_0_96), .CK(n_0_136), .Q(n_val[32]), .QN());
   DFF_X1 \n_val_reg[31]  (.D(n_0_95), .CK(n_0_136), .Q(n_val[31]), .QN());
   DFF_X1 \n_val_reg[30]  (.D(n_0_94), .CK(n_0_136), .Q(n_val[30]), .QN());
   DFF_X1 \n_val_reg[29]  (.D(n_0_93), .CK(n_0_136), .Q(n_val[29]), .QN());
   DFF_X1 \n_val_reg[28]  (.D(n_0_92), .CK(n_0_136), .Q(n_val[28]), .QN());
   DFF_X1 \n_val_reg[27]  (.D(n_0_91), .CK(n_0_136), .Q(n_val[27]), .QN());
   DFF_X1 \n_val_reg[26]  (.D(n_0_90), .CK(n_0_136), .Q(n_val[26]), .QN());
   DFF_X1 \n_val_reg[25]  (.D(n_0_89), .CK(n_0_136), .Q(n_val[25]), .QN());
   DFF_X1 \n_val_reg[24]  (.D(n_0_88), .CK(n_0_136), .Q(n_val[24]), .QN());
   DFF_X1 \n_val_reg[23]  (.D(n_0_87), .CK(n_0_136), .Q(n_val[23]), .QN());
   DFF_X1 \n_val_reg[22]  (.D(n_0_86), .CK(n_0_136), .Q(n_val[22]), .QN());
   DFF_X1 \n_val_reg[21]  (.D(n_0_85), .CK(n_0_136), .Q(n_val[21]), .QN());
   DFF_X1 \n_val_reg[20]  (.D(n_0_84), .CK(n_0_136), .Q(n_val[20]), .QN());
   DFF_X1 \n_val_reg[19]  (.D(n_0_83), .CK(n_0_136), .Q(n_val[19]), .QN());
   DFF_X1 \n_val_reg[18]  (.D(n_0_82), .CK(n_0_136), .Q(n_val[18]), .QN());
   DFF_X1 \n_val_reg[17]  (.D(n_0_81), .CK(n_0_136), .Q(n_val[17]), .QN());
   DFF_X1 \n_val_reg[16]  (.D(n_0_80), .CK(n_0_136), .Q(n_val[16]), .QN());
   DFF_X1 \n_val_reg[15]  (.D(n_0_79), .CK(n_0_136), .Q(n_val[15]), .QN());
   DFF_X1 \n_val_reg[14]  (.D(n_0_78), .CK(n_0_136), .Q(n_val[14]), .QN());
   DFF_X1 \n_val_reg[13]  (.D(n_0_77), .CK(n_0_136), .Q(n_val[13]), .QN());
   DFF_X1 \n_val_reg[12]  (.D(n_0_76), .CK(n_0_136), .Q(n_val[12]), .QN());
   DFF_X1 \n_val_reg[11]  (.D(n_0_75), .CK(n_0_136), .Q(n_val[11]), .QN());
   DFF_X1 \n_val_reg[10]  (.D(n_0_74), .CK(n_0_136), .Q(n_val[10]), .QN());
   DFF_X1 \n_val_reg[9]  (.D(n_0_73), .CK(n_0_136), .Q(n_val[9]), .QN());
   DFF_X1 \n_val_reg[8]  (.D(n_0_72), .CK(n_0_136), .Q(n_val[8]), .QN());
   DFF_X1 \n_val_reg[7]  (.D(n_0_71), .CK(n_0_136), .Q(n_val[7]), .QN());
   DFF_X1 \n_val_reg[6]  (.D(n_0_70), .CK(n_0_136), .Q(n_val[6]), .QN());
   DFF_X1 \n_val_reg[5]  (.D(n_0_69), .CK(n_0_136), .Q(n_val[5]), .QN());
   DFF_X1 \n_val_reg[4]  (.D(n_0_68), .CK(n_0_136), .Q(n_val[4]), .QN());
   DFF_X1 \n_val_reg[3]  (.D(n_0_67), .CK(n_0_136), .Q(n_val[3]), .QN());
   DFF_X1 \n_val_reg[2]  (.D(n_0_66), .CK(n_0_136), .Q(n_val[2]), .QN());
   DFF_X1 \n_val_reg[1]  (.D(n_0_65), .CK(n_0_136), .Q(n_val[1]), .QN());
   DFF_X1 \n_val_reg[0]  (.D(n_0_64), .CK(n_0_136), .Q(n_val[0]), .QN());
   DFF_X1 \m_val_reg[63]  (.D(n_0_63), .CK(n_0_136), .Q(m_val[63]), .QN());
   DFF_X1 \m_val_reg[62]  (.D(n_0_62), .CK(n_0_136), .Q(m_val[62]), .QN());
   DFF_X1 \m_val_reg[61]  (.D(n_0_61), .CK(n_0_136), .Q(m_val[61]), .QN());
   DFF_X1 \m_val_reg[60]  (.D(n_0_60), .CK(n_0_136), .Q(m_val[60]), .QN());
   DFF_X1 \m_val_reg[59]  (.D(n_0_59), .CK(n_0_136), .Q(m_val[59]), .QN());
   DFF_X1 \m_val_reg[58]  (.D(n_0_58), .CK(n_0_136), .Q(m_val[58]), .QN());
   DFF_X1 \m_val_reg[57]  (.D(n_0_57), .CK(n_0_136), .Q(m_val[57]), .QN());
   DFF_X1 \m_val_reg[56]  (.D(n_0_56), .CK(n_0_136), .Q(m_val[56]), .QN());
   DFF_X1 \m_val_reg[55]  (.D(n_0_55), .CK(n_0_136), .Q(m_val[55]), .QN());
   DFF_X1 \m_val_reg[54]  (.D(n_0_54), .CK(n_0_136), .Q(m_val[54]), .QN());
   DFF_X1 \m_val_reg[53]  (.D(n_0_53), .CK(n_0_136), .Q(m_val[53]), .QN());
   DFF_X1 \m_val_reg[52]  (.D(n_0_52), .CK(n_0_136), .Q(m_val[52]), .QN());
   DFF_X1 \m_val_reg[51]  (.D(n_0_51), .CK(n_0_136), .Q(m_val[51]), .QN());
   DFF_X1 \m_val_reg[50]  (.D(n_0_50), .CK(n_0_136), .Q(m_val[50]), .QN());
   DFF_X1 \m_val_reg[49]  (.D(n_0_49), .CK(n_0_136), .Q(m_val[49]), .QN());
   DFF_X1 \m_val_reg[48]  (.D(n_0_48), .CK(n_0_136), .Q(m_val[48]), .QN());
   DFF_X1 \m_val_reg[47]  (.D(n_0_47), .CK(n_0_136), .Q(m_val[47]), .QN());
   DFF_X1 \m_val_reg[46]  (.D(n_0_46), .CK(n_0_136), .Q(m_val[46]), .QN());
   DFF_X1 \m_val_reg[45]  (.D(n_0_45), .CK(n_0_136), .Q(m_val[45]), .QN());
   DFF_X1 \m_val_reg[44]  (.D(n_0_44), .CK(n_0_136), .Q(m_val[44]), .QN());
   DFF_X1 \m_val_reg[43]  (.D(n_0_43), .CK(n_0_136), .Q(m_val[43]), .QN());
   DFF_X1 \m_val_reg[42]  (.D(n_0_42), .CK(n_0_136), .Q(m_val[42]), .QN());
   DFF_X1 \m_val_reg[41]  (.D(n_0_41), .CK(n_0_136), .Q(m_val[41]), .QN());
   DFF_X1 \m_val_reg[40]  (.D(n_0_40), .CK(n_0_136), .Q(m_val[40]), .QN());
   DFF_X1 \m_val_reg[39]  (.D(n_0_39), .CK(n_0_136), .Q(m_val[39]), .QN());
   DFF_X1 \m_val_reg[38]  (.D(n_0_38), .CK(n_0_136), .Q(m_val[38]), .QN());
   DFF_X1 \m_val_reg[37]  (.D(n_0_37), .CK(n_0_136), .Q(m_val[37]), .QN());
   DFF_X1 \m_val_reg[36]  (.D(n_0_36), .CK(n_0_136), .Q(m_val[36]), .QN());
   DFF_X1 \m_val_reg[35]  (.D(n_0_35), .CK(n_0_136), .Q(m_val[35]), .QN());
   DFF_X1 \m_val_reg[34]  (.D(n_0_34), .CK(n_0_136), .Q(m_val[34]), .QN());
   DFF_X1 \m_val_reg[33]  (.D(n_0_33), .CK(n_0_136), .Q(m_val[33]), .QN());
   DFF_X1 \m_val_reg[32]  (.D(n_0_32), .CK(n_0_136), .Q(m_val[32]), .QN());
   DFF_X1 \m_val_reg[31]  (.D(n_0_31), .CK(n_0_136), .Q(m_val[31]), .QN());
   DFF_X1 \m_val_reg[30]  (.D(n_0_30), .CK(n_0_136), .Q(m_val[30]), .QN());
   DFF_X1 \m_val_reg[29]  (.D(n_0_29), .CK(n_0_136), .Q(m_val[29]), .QN());
   DFF_X1 \m_val_reg[28]  (.D(n_0_28), .CK(n_0_136), .Q(m_val[28]), .QN());
   DFF_X1 \m_val_reg[27]  (.D(n_0_27), .CK(n_0_136), .Q(m_val[27]), .QN());
   DFF_X1 \m_val_reg[26]  (.D(n_0_26), .CK(n_0_136), .Q(m_val[26]), .QN());
   DFF_X1 \m_val_reg[25]  (.D(n_0_25), .CK(n_0_136), .Q(m_val[25]), .QN());
   DFF_X1 \m_val_reg[24]  (.D(n_0_24), .CK(n_0_136), .Q(m_val[24]), .QN());
   DFF_X1 \m_val_reg[23]  (.D(n_0_23), .CK(n_0_136), .Q(m_val[23]), .QN());
   DFF_X1 \m_val_reg[22]  (.D(n_0_22), .CK(n_0_136), .Q(m_val[22]), .QN());
   DFF_X1 \m_val_reg[21]  (.D(n_0_21), .CK(n_0_136), .Q(m_val[21]), .QN());
   DFF_X1 \m_val_reg[20]  (.D(n_0_20), .CK(n_0_136), .Q(m_val[20]), .QN());
   DFF_X1 \m_val_reg[19]  (.D(n_0_19), .CK(n_0_136), .Q(m_val[19]), .QN());
   DFF_X1 \m_val_reg[18]  (.D(n_0_18), .CK(n_0_136), .Q(m_val[18]), .QN());
   DFF_X1 \m_val_reg[17]  (.D(n_0_17), .CK(n_0_136), .Q(m_val[17]), .QN());
   DFF_X1 \m_val_reg[16]  (.D(n_0_16), .CK(n_0_136), .Q(m_val[16]), .QN());
   DFF_X1 \m_val_reg[15]  (.D(n_0_15), .CK(n_0_136), .Q(m_val[15]), .QN());
   DFF_X1 \m_val_reg[14]  (.D(n_0_14), .CK(n_0_136), .Q(m_val[14]), .QN());
   DFF_X1 \m_val_reg[13]  (.D(n_0_13), .CK(n_0_136), .Q(m_val[13]), .QN());
   DFF_X1 \m_val_reg[12]  (.D(n_0_12), .CK(n_0_136), .Q(m_val[12]), .QN());
   DFF_X1 \m_val_reg[11]  (.D(n_0_11), .CK(n_0_136), .Q(m_val[11]), .QN());
   DFF_X1 \m_val_reg[10]  (.D(n_0_10), .CK(n_0_136), .Q(m_val[10]), .QN());
   DFF_X1 \m_val_reg[9]  (.D(n_0_9), .CK(n_0_136), .Q(m_val[9]), .QN());
   DFF_X1 \m_val_reg[8]  (.D(n_0_8), .CK(n_0_136), .Q(m_val[8]), .QN());
   DFF_X1 \m_val_reg[7]  (.D(n_0_7), .CK(n_0_136), .Q(m_val[7]), .QN());
   DFF_X1 \m_val_reg[6]  (.D(n_0_6), .CK(n_0_136), .Q(m_val[6]), .QN());
   DFF_X1 \m_val_reg[5]  (.D(n_0_5), .CK(n_0_136), .Q(m_val[5]), .QN());
   DFF_X1 \m_val_reg[4]  (.D(n_0_4), .CK(n_0_136), .Q(m_val[4]), .QN());
   DFF_X1 \m_val_reg[3]  (.D(n_0_3), .CK(n_0_136), .Q(m_val[3]), .QN());
   DFF_X1 \m_val_reg[2]  (.D(n_0_2), .CK(n_0_136), .Q(m_val[2]), .QN());
   DFF_X1 \m_val_reg[1]  (.D(n_0_1), .CK(n_0_136), .Q(m_val[1]), .QN());
   DFF_X1 \m_val_reg[0]  (.D(n_0_0), .CK(n_0_136), .Q(m_val[0]), .QN());
   INV_X1 i_0_0_0 (.A(n_0_0_0), .ZN(n_0_0));
   AOI22_X1 i_0_0_1 (.A1(RAM_DATA_RD2[0]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[0]), .ZN(n_0_0_0));
   INV_X1 i_0_0_2 (.A(n_0_0_1), .ZN(n_0_1));
   AOI22_X1 i_0_0_3 (.A1(RAM_DATA_RD2[1]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[1]), .ZN(n_0_0_1));
   INV_X1 i_0_0_4 (.A(n_0_0_2), .ZN(n_0_2));
   AOI22_X1 i_0_0_5 (.A1(RAM_DATA_RD2[2]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[2]), .ZN(n_0_0_2));
   INV_X1 i_0_0_6 (.A(n_0_0_3), .ZN(n_0_3));
   AOI22_X1 i_0_0_7 (.A1(RAM_DATA_RD2[3]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[3]), .ZN(n_0_0_3));
   INV_X1 i_0_0_8 (.A(n_0_0_4), .ZN(n_0_4));
   AOI22_X1 i_0_0_9 (.A1(RAM_DATA_RD2[4]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[4]), .ZN(n_0_0_4));
   INV_X1 i_0_0_10 (.A(n_0_0_5), .ZN(n_0_5));
   AOI22_X1 i_0_0_11 (.A1(RAM_DATA_RD2[5]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[5]), .ZN(n_0_0_5));
   INV_X1 i_0_0_12 (.A(n_0_0_6), .ZN(n_0_6));
   AOI22_X1 i_0_0_13 (.A1(RAM_DATA_RD2[6]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[6]), .ZN(n_0_0_6));
   INV_X1 i_0_0_14 (.A(n_0_0_7), .ZN(n_0_7));
   AOI22_X1 i_0_0_15 (.A1(RAM_DATA_RD2[7]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[7]), .ZN(n_0_0_7));
   INV_X1 i_0_0_16 (.A(n_0_0_8), .ZN(n_0_8));
   AOI22_X1 i_0_0_17 (.A1(RAM_DATA_RD2[8]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[8]), .ZN(n_0_0_8));
   INV_X1 i_0_0_18 (.A(n_0_0_9), .ZN(n_0_9));
   AOI22_X1 i_0_0_19 (.A1(RAM_DATA_RD2[9]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[9]), .ZN(n_0_0_9));
   INV_X1 i_0_0_20 (.A(n_0_0_10), .ZN(n_0_10));
   AOI22_X1 i_0_0_21 (.A1(RAM_DATA_RD2[10]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[10]), .ZN(n_0_0_10));
   INV_X1 i_0_0_22 (.A(n_0_0_11), .ZN(n_0_11));
   AOI22_X1 i_0_0_23 (.A1(RAM_DATA_RD2[11]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[11]), .ZN(n_0_0_11));
   INV_X1 i_0_0_24 (.A(n_0_0_12), .ZN(n_0_12));
   AOI22_X1 i_0_0_25 (.A1(RAM_DATA_RD2[12]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[12]), .ZN(n_0_0_12));
   INV_X1 i_0_0_26 (.A(n_0_0_13), .ZN(n_0_13));
   AOI22_X1 i_0_0_27 (.A1(RAM_DATA_RD2[13]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[13]), .ZN(n_0_0_13));
   INV_X1 i_0_0_28 (.A(n_0_0_14), .ZN(n_0_14));
   AOI22_X1 i_0_0_29 (.A1(RAM_DATA_RD2[14]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[14]), .ZN(n_0_0_14));
   INV_X1 i_0_0_30 (.A(n_0_0_15), .ZN(n_0_15));
   AOI22_X1 i_0_0_31 (.A1(RAM_DATA_RD2[15]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[15]), .ZN(n_0_0_15));
   INV_X1 i_0_0_32 (.A(n_0_0_16), .ZN(n_0_16));
   AOI22_X1 i_0_0_33 (.A1(RAM_DATA_RD2[16]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[16]), .ZN(n_0_0_16));
   INV_X1 i_0_0_34 (.A(n_0_0_17), .ZN(n_0_17));
   AOI22_X1 i_0_0_35 (.A1(RAM_DATA_RD2[17]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[17]), .ZN(n_0_0_17));
   INV_X1 i_0_0_36 (.A(n_0_0_18), .ZN(n_0_18));
   AOI22_X1 i_0_0_37 (.A1(RAM_DATA_RD2[18]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[18]), .ZN(n_0_0_18));
   INV_X1 i_0_0_38 (.A(n_0_0_19), .ZN(n_0_19));
   AOI22_X1 i_0_0_39 (.A1(RAM_DATA_RD2[19]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[19]), .ZN(n_0_0_19));
   INV_X1 i_0_0_40 (.A(n_0_0_20), .ZN(n_0_20));
   AOI22_X1 i_0_0_41 (.A1(RAM_DATA_RD2[20]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[20]), .ZN(n_0_0_20));
   INV_X1 i_0_0_42 (.A(n_0_0_21), .ZN(n_0_21));
   AOI22_X1 i_0_0_43 (.A1(RAM_DATA_RD2[21]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[21]), .ZN(n_0_0_21));
   INV_X1 i_0_0_44 (.A(n_0_0_22), .ZN(n_0_22));
   AOI22_X1 i_0_0_45 (.A1(RAM_DATA_RD2[22]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[22]), .ZN(n_0_0_22));
   INV_X1 i_0_0_46 (.A(n_0_0_23), .ZN(n_0_23));
   AOI22_X1 i_0_0_47 (.A1(RAM_DATA_RD2[23]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[23]), .ZN(n_0_0_23));
   INV_X1 i_0_0_48 (.A(n_0_0_24), .ZN(n_0_24));
   AOI22_X1 i_0_0_49 (.A1(RAM_DATA_RD2[24]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[24]), .ZN(n_0_0_24));
   INV_X1 i_0_0_50 (.A(n_0_0_25), .ZN(n_0_25));
   AOI22_X1 i_0_0_51 (.A1(RAM_DATA_RD2[25]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[25]), .ZN(n_0_0_25));
   INV_X1 i_0_0_52 (.A(n_0_0_26), .ZN(n_0_26));
   AOI22_X1 i_0_0_53 (.A1(RAM_DATA_RD2[26]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[26]), .ZN(n_0_0_26));
   INV_X1 i_0_0_54 (.A(n_0_0_27), .ZN(n_0_27));
   AOI22_X1 i_0_0_55 (.A1(RAM_DATA_RD2[27]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[27]), .ZN(n_0_0_27));
   INV_X1 i_0_0_56 (.A(n_0_0_28), .ZN(n_0_28));
   AOI22_X1 i_0_0_57 (.A1(RAM_DATA_RD2[28]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[28]), .ZN(n_0_0_28));
   INV_X1 i_0_0_58 (.A(n_0_0_29), .ZN(n_0_29));
   AOI22_X1 i_0_0_59 (.A1(RAM_DATA_RD2[29]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[29]), .ZN(n_0_0_29));
   INV_X1 i_0_0_60 (.A(n_0_0_30), .ZN(n_0_30));
   AOI22_X1 i_0_0_61 (.A1(RAM_DATA_RD2[30]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[30]), .ZN(n_0_0_30));
   INV_X1 i_0_0_62 (.A(n_0_0_31), .ZN(n_0_31));
   AOI22_X1 i_0_0_63 (.A1(RAM_DATA_RD2[31]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[31]), .ZN(n_0_0_31));
   INV_X1 i_0_0_64 (.A(n_0_0_32), .ZN(n_0_32));
   AOI22_X1 i_0_0_65 (.A1(RAM_DATA_RD2[32]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[32]), .ZN(n_0_0_32));
   INV_X1 i_0_0_66 (.A(n_0_0_33), .ZN(n_0_33));
   AOI22_X1 i_0_0_67 (.A1(RAM_DATA_RD2[33]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[33]), .ZN(n_0_0_33));
   INV_X1 i_0_0_68 (.A(n_0_0_34), .ZN(n_0_34));
   AOI22_X1 i_0_0_69 (.A1(RAM_DATA_RD2[34]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[34]), .ZN(n_0_0_34));
   INV_X1 i_0_0_70 (.A(n_0_0_35), .ZN(n_0_35));
   AOI22_X1 i_0_0_71 (.A1(RAM_DATA_RD2[35]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[35]), .ZN(n_0_0_35));
   INV_X1 i_0_0_72 (.A(n_0_0_36), .ZN(n_0_36));
   AOI22_X1 i_0_0_73 (.A1(RAM_DATA_RD2[36]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[36]), .ZN(n_0_0_36));
   INV_X1 i_0_0_74 (.A(n_0_0_37), .ZN(n_0_37));
   AOI22_X1 i_0_0_75 (.A1(RAM_DATA_RD2[37]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[37]), .ZN(n_0_0_37));
   INV_X1 i_0_0_76 (.A(n_0_0_38), .ZN(n_0_38));
   AOI22_X1 i_0_0_77 (.A1(RAM_DATA_RD2[38]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[38]), .ZN(n_0_0_38));
   INV_X1 i_0_0_78 (.A(n_0_0_39), .ZN(n_0_39));
   AOI22_X1 i_0_0_79 (.A1(RAM_DATA_RD2[39]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[39]), .ZN(n_0_0_39));
   INV_X1 i_0_0_80 (.A(n_0_0_40), .ZN(n_0_40));
   AOI22_X1 i_0_0_81 (.A1(RAM_DATA_RD2[40]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[40]), .ZN(n_0_0_40));
   INV_X1 i_0_0_82 (.A(n_0_0_41), .ZN(n_0_41));
   AOI22_X1 i_0_0_83 (.A1(RAM_DATA_RD2[41]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[41]), .ZN(n_0_0_41));
   INV_X1 i_0_0_84 (.A(n_0_0_42), .ZN(n_0_42));
   AOI22_X1 i_0_0_85 (.A1(RAM_DATA_RD2[42]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[42]), .ZN(n_0_0_42));
   INV_X1 i_0_0_86 (.A(n_0_0_43), .ZN(n_0_43));
   AOI22_X1 i_0_0_87 (.A1(RAM_DATA_RD2[43]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[43]), .ZN(n_0_0_43));
   INV_X1 i_0_0_88 (.A(n_0_0_44), .ZN(n_0_44));
   AOI22_X1 i_0_0_89 (.A1(RAM_DATA_RD2[44]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[44]), .ZN(n_0_0_44));
   INV_X1 i_0_0_90 (.A(n_0_0_45), .ZN(n_0_45));
   AOI22_X1 i_0_0_91 (.A1(RAM_DATA_RD2[45]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[45]), .ZN(n_0_0_45));
   INV_X1 i_0_0_92 (.A(n_0_0_46), .ZN(n_0_46));
   AOI22_X1 i_0_0_93 (.A1(RAM_DATA_RD2[46]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[46]), .ZN(n_0_0_46));
   INV_X1 i_0_0_94 (.A(n_0_0_47), .ZN(n_0_47));
   AOI22_X1 i_0_0_95 (.A1(RAM_DATA_RD2[47]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[47]), .ZN(n_0_0_47));
   INV_X1 i_0_0_96 (.A(n_0_0_48), .ZN(n_0_48));
   AOI22_X1 i_0_0_97 (.A1(RAM_DATA_RD2[48]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[48]), .ZN(n_0_0_48));
   INV_X1 i_0_0_98 (.A(n_0_0_49), .ZN(n_0_49));
   AOI22_X1 i_0_0_99 (.A1(RAM_DATA_RD2[49]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[49]), .ZN(n_0_0_49));
   INV_X1 i_0_0_100 (.A(n_0_0_50), .ZN(n_0_50));
   AOI22_X1 i_0_0_101 (.A1(RAM_DATA_RD2[50]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[50]), .ZN(n_0_0_50));
   INV_X1 i_0_0_102 (.A(n_0_0_51), .ZN(n_0_51));
   AOI22_X1 i_0_0_103 (.A1(RAM_DATA_RD2[51]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[51]), .ZN(n_0_0_51));
   INV_X1 i_0_0_104 (.A(n_0_0_52), .ZN(n_0_52));
   AOI22_X1 i_0_0_105 (.A1(RAM_DATA_RD2[52]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[52]), .ZN(n_0_0_52));
   INV_X1 i_0_0_106 (.A(n_0_0_53), .ZN(n_0_53));
   AOI22_X1 i_0_0_107 (.A1(RAM_DATA_RD2[53]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[53]), .ZN(n_0_0_53));
   INV_X1 i_0_0_108 (.A(n_0_0_54), .ZN(n_0_54));
   AOI22_X1 i_0_0_109 (.A1(RAM_DATA_RD2[54]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[54]), .ZN(n_0_0_54));
   INV_X1 i_0_0_110 (.A(n_0_0_55), .ZN(n_0_55));
   AOI22_X1 i_0_0_111 (.A1(RAM_DATA_RD2[55]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[55]), .ZN(n_0_0_55));
   INV_X1 i_0_0_112 (.A(n_0_0_56), .ZN(n_0_56));
   AOI22_X1 i_0_0_113 (.A1(RAM_DATA_RD2[56]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[56]), .ZN(n_0_0_56));
   INV_X1 i_0_0_114 (.A(n_0_0_57), .ZN(n_0_57));
   AOI22_X1 i_0_0_115 (.A1(RAM_DATA_RD2[57]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[57]), .ZN(n_0_0_57));
   INV_X1 i_0_0_116 (.A(n_0_0_58), .ZN(n_0_58));
   AOI22_X1 i_0_0_117 (.A1(RAM_DATA_RD2[58]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[58]), .ZN(n_0_0_58));
   INV_X1 i_0_0_118 (.A(n_0_0_59), .ZN(n_0_59));
   AOI22_X1 i_0_0_119 (.A1(RAM_DATA_RD2[59]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[59]), .ZN(n_0_0_59));
   INV_X1 i_0_0_120 (.A(n_0_0_60), .ZN(n_0_60));
   AOI22_X1 i_0_0_121 (.A1(RAM_DATA_RD2[60]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[60]), .ZN(n_0_0_60));
   INV_X1 i_0_0_122 (.A(n_0_0_61), .ZN(n_0_61));
   AOI22_X1 i_0_0_123 (.A1(RAM_DATA_RD2[61]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[61]), .ZN(n_0_0_61));
   INV_X1 i_0_0_124 (.A(n_0_0_62), .ZN(n_0_62));
   AOI22_X1 i_0_0_125 (.A1(RAM_DATA_RD2[62]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[62]), .ZN(n_0_0_62));
   INV_X1 i_0_0_126 (.A(n_0_0_63), .ZN(n_0_63));
   AOI22_X1 i_0_0_127 (.A1(RAM_DATA_RD2[63]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(m_val[63]), .ZN(n_0_0_63));
   INV_X1 i_0_0_128 (.A(n_0_0_64), .ZN(n_0_64));
   AOI22_X1 i_0_0_129 (.A1(RAM_DATA_RD1[0]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[0]), .ZN(n_0_0_64));
   INV_X1 i_0_0_130 (.A(n_0_0_65), .ZN(n_0_65));
   AOI22_X1 i_0_0_131 (.A1(RAM_DATA_RD1[1]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[1]), .ZN(n_0_0_65));
   INV_X1 i_0_0_132 (.A(n_0_0_66), .ZN(n_0_66));
   AOI22_X1 i_0_0_133 (.A1(RAM_DATA_RD1[2]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[2]), .ZN(n_0_0_66));
   INV_X1 i_0_0_134 (.A(n_0_0_67), .ZN(n_0_67));
   AOI22_X1 i_0_0_135 (.A1(RAM_DATA_RD1[3]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[3]), .ZN(n_0_0_67));
   INV_X1 i_0_0_136 (.A(n_0_0_68), .ZN(n_0_68));
   AOI22_X1 i_0_0_137 (.A1(RAM_DATA_RD1[4]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[4]), .ZN(n_0_0_68));
   INV_X1 i_0_0_138 (.A(n_0_0_69), .ZN(n_0_69));
   AOI22_X1 i_0_0_139 (.A1(RAM_DATA_RD1[5]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[5]), .ZN(n_0_0_69));
   INV_X1 i_0_0_140 (.A(n_0_0_70), .ZN(n_0_70));
   AOI22_X1 i_0_0_141 (.A1(RAM_DATA_RD1[6]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[6]), .ZN(n_0_0_70));
   INV_X1 i_0_0_142 (.A(n_0_0_71), .ZN(n_0_71));
   AOI22_X1 i_0_0_143 (.A1(RAM_DATA_RD1[7]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[7]), .ZN(n_0_0_71));
   INV_X1 i_0_0_144 (.A(n_0_0_72), .ZN(n_0_72));
   AOI22_X1 i_0_0_145 (.A1(RAM_DATA_RD1[8]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[8]), .ZN(n_0_0_72));
   INV_X1 i_0_0_146 (.A(n_0_0_73), .ZN(n_0_73));
   AOI22_X1 i_0_0_147 (.A1(RAM_DATA_RD1[9]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[9]), .ZN(n_0_0_73));
   INV_X1 i_0_0_148 (.A(n_0_0_74), .ZN(n_0_74));
   AOI22_X1 i_0_0_149 (.A1(RAM_DATA_RD1[10]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[10]), .ZN(n_0_0_74));
   INV_X1 i_0_0_150 (.A(n_0_0_75), .ZN(n_0_75));
   AOI22_X1 i_0_0_151 (.A1(RAM_DATA_RD1[11]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[11]), .ZN(n_0_0_75));
   INV_X1 i_0_0_152 (.A(n_0_0_76), .ZN(n_0_76));
   AOI22_X1 i_0_0_153 (.A1(RAM_DATA_RD1[12]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[12]), .ZN(n_0_0_76));
   INV_X1 i_0_0_154 (.A(n_0_0_77), .ZN(n_0_77));
   AOI22_X1 i_0_0_155 (.A1(RAM_DATA_RD1[13]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[13]), .ZN(n_0_0_77));
   INV_X1 i_0_0_156 (.A(n_0_0_78), .ZN(n_0_78));
   AOI22_X1 i_0_0_157 (.A1(RAM_DATA_RD1[14]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[14]), .ZN(n_0_0_78));
   INV_X1 i_0_0_158 (.A(n_0_0_79), .ZN(n_0_79));
   AOI22_X1 i_0_0_159 (.A1(RAM_DATA_RD1[15]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[15]), .ZN(n_0_0_79));
   INV_X1 i_0_0_160 (.A(n_0_0_80), .ZN(n_0_80));
   AOI22_X1 i_0_0_161 (.A1(RAM_DATA_RD1[16]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[16]), .ZN(n_0_0_80));
   INV_X1 i_0_0_162 (.A(n_0_0_81), .ZN(n_0_81));
   AOI22_X1 i_0_0_163 (.A1(RAM_DATA_RD1[17]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[17]), .ZN(n_0_0_81));
   INV_X1 i_0_0_164 (.A(n_0_0_82), .ZN(n_0_82));
   AOI22_X1 i_0_0_165 (.A1(RAM_DATA_RD1[18]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[18]), .ZN(n_0_0_82));
   INV_X1 i_0_0_166 (.A(n_0_0_83), .ZN(n_0_83));
   AOI22_X1 i_0_0_167 (.A1(RAM_DATA_RD1[19]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[19]), .ZN(n_0_0_83));
   INV_X1 i_0_0_168 (.A(n_0_0_84), .ZN(n_0_84));
   AOI22_X1 i_0_0_169 (.A1(RAM_DATA_RD1[20]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[20]), .ZN(n_0_0_84));
   INV_X1 i_0_0_170 (.A(n_0_0_85), .ZN(n_0_85));
   AOI22_X1 i_0_0_171 (.A1(RAM_DATA_RD1[21]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[21]), .ZN(n_0_0_85));
   INV_X1 i_0_0_172 (.A(n_0_0_86), .ZN(n_0_86));
   AOI22_X1 i_0_0_173 (.A1(RAM_DATA_RD1[22]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[22]), .ZN(n_0_0_86));
   INV_X1 i_0_0_174 (.A(n_0_0_87), .ZN(n_0_87));
   AOI22_X1 i_0_0_175 (.A1(RAM_DATA_RD1[23]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[23]), .ZN(n_0_0_87));
   INV_X1 i_0_0_176 (.A(n_0_0_88), .ZN(n_0_88));
   AOI22_X1 i_0_0_177 (.A1(RAM_DATA_RD1[24]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[24]), .ZN(n_0_0_88));
   INV_X1 i_0_0_178 (.A(n_0_0_89), .ZN(n_0_89));
   AOI22_X1 i_0_0_179 (.A1(RAM_DATA_RD1[25]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[25]), .ZN(n_0_0_89));
   INV_X1 i_0_0_180 (.A(n_0_0_90), .ZN(n_0_90));
   AOI22_X1 i_0_0_181 (.A1(RAM_DATA_RD1[26]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[26]), .ZN(n_0_0_90));
   INV_X1 i_0_0_182 (.A(n_0_0_91), .ZN(n_0_91));
   AOI22_X1 i_0_0_183 (.A1(RAM_DATA_RD1[27]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[27]), .ZN(n_0_0_91));
   INV_X1 i_0_0_184 (.A(n_0_0_92), .ZN(n_0_92));
   AOI22_X1 i_0_0_185 (.A1(RAM_DATA_RD1[28]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[28]), .ZN(n_0_0_92));
   INV_X1 i_0_0_186 (.A(n_0_0_93), .ZN(n_0_93));
   AOI22_X1 i_0_0_187 (.A1(RAM_DATA_RD1[29]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[29]), .ZN(n_0_0_93));
   INV_X1 i_0_0_188 (.A(n_0_0_94), .ZN(n_0_94));
   AOI22_X1 i_0_0_189 (.A1(RAM_DATA_RD1[30]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[30]), .ZN(n_0_0_94));
   INV_X1 i_0_0_190 (.A(n_0_0_95), .ZN(n_0_95));
   AOI22_X1 i_0_0_191 (.A1(RAM_DATA_RD1[31]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[31]), .ZN(n_0_0_95));
   INV_X1 i_0_0_192 (.A(n_0_0_96), .ZN(n_0_96));
   AOI22_X1 i_0_0_193 (.A1(RAM_DATA_RD1[32]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[32]), .ZN(n_0_0_96));
   INV_X1 i_0_0_194 (.A(n_0_0_97), .ZN(n_0_97));
   AOI22_X1 i_0_0_195 (.A1(RAM_DATA_RD1[33]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[33]), .ZN(n_0_0_97));
   INV_X1 i_0_0_196 (.A(n_0_0_98), .ZN(n_0_98));
   AOI22_X1 i_0_0_197 (.A1(RAM_DATA_RD1[34]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[34]), .ZN(n_0_0_98));
   INV_X1 i_0_0_198 (.A(n_0_0_99), .ZN(n_0_99));
   AOI22_X1 i_0_0_199 (.A1(RAM_DATA_RD1[35]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[35]), .ZN(n_0_0_99));
   INV_X1 i_0_0_200 (.A(n_0_0_100), .ZN(n_0_100));
   AOI22_X1 i_0_0_201 (.A1(RAM_DATA_RD1[36]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[36]), .ZN(n_0_0_100));
   INV_X1 i_0_0_202 (.A(n_0_0_101), .ZN(n_0_101));
   AOI22_X1 i_0_0_203 (.A1(RAM_DATA_RD1[37]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[37]), .ZN(n_0_0_101));
   INV_X1 i_0_0_204 (.A(n_0_0_102), .ZN(n_0_102));
   AOI22_X1 i_0_0_205 (.A1(RAM_DATA_RD1[38]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[38]), .ZN(n_0_0_102));
   INV_X1 i_0_0_206 (.A(n_0_0_103), .ZN(n_0_103));
   AOI22_X1 i_0_0_207 (.A1(RAM_DATA_RD1[39]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[39]), .ZN(n_0_0_103));
   INV_X1 i_0_0_208 (.A(n_0_0_104), .ZN(n_0_104));
   AOI22_X1 i_0_0_209 (.A1(RAM_DATA_RD1[40]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[40]), .ZN(n_0_0_104));
   INV_X1 i_0_0_210 (.A(n_0_0_105), .ZN(n_0_105));
   AOI22_X1 i_0_0_211 (.A1(RAM_DATA_RD1[41]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[41]), .ZN(n_0_0_105));
   INV_X1 i_0_0_212 (.A(n_0_0_106), .ZN(n_0_106));
   AOI22_X1 i_0_0_213 (.A1(RAM_DATA_RD1[42]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[42]), .ZN(n_0_0_106));
   INV_X1 i_0_0_214 (.A(n_0_0_107), .ZN(n_0_107));
   AOI22_X1 i_0_0_215 (.A1(RAM_DATA_RD1[43]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[43]), .ZN(n_0_0_107));
   INV_X1 i_0_0_216 (.A(n_0_0_108), .ZN(n_0_108));
   AOI22_X1 i_0_0_217 (.A1(RAM_DATA_RD1[44]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[44]), .ZN(n_0_0_108));
   INV_X1 i_0_0_218 (.A(n_0_0_109), .ZN(n_0_109));
   AOI22_X1 i_0_0_219 (.A1(RAM_DATA_RD1[45]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[45]), .ZN(n_0_0_109));
   INV_X1 i_0_0_220 (.A(n_0_0_110), .ZN(n_0_110));
   AOI22_X1 i_0_0_221 (.A1(RAM_DATA_RD1[46]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[46]), .ZN(n_0_0_110));
   INV_X1 i_0_0_222 (.A(n_0_0_111), .ZN(n_0_111));
   AOI22_X1 i_0_0_223 (.A1(RAM_DATA_RD1[47]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[47]), .ZN(n_0_0_111));
   INV_X1 i_0_0_224 (.A(n_0_0_112), .ZN(n_0_112));
   AOI22_X1 i_0_0_225 (.A1(RAM_DATA_RD1[48]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[48]), .ZN(n_0_0_112));
   INV_X1 i_0_0_226 (.A(n_0_0_113), .ZN(n_0_113));
   AOI22_X1 i_0_0_227 (.A1(RAM_DATA_RD1[49]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[49]), .ZN(n_0_0_113));
   INV_X1 i_0_0_228 (.A(n_0_0_114), .ZN(n_0_114));
   AOI22_X1 i_0_0_229 (.A1(RAM_DATA_RD1[50]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[50]), .ZN(n_0_0_114));
   INV_X1 i_0_0_230 (.A(n_0_0_115), .ZN(n_0_115));
   AOI22_X1 i_0_0_231 (.A1(RAM_DATA_RD1[51]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[51]), .ZN(n_0_0_115));
   INV_X1 i_0_0_232 (.A(n_0_0_116), .ZN(n_0_116));
   AOI22_X1 i_0_0_233 (.A1(RAM_DATA_RD1[52]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[52]), .ZN(n_0_0_116));
   INV_X1 i_0_0_234 (.A(n_0_0_117), .ZN(n_0_117));
   AOI22_X1 i_0_0_235 (.A1(RAM_DATA_RD1[53]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[53]), .ZN(n_0_0_117));
   INV_X1 i_0_0_236 (.A(n_0_0_118), .ZN(n_0_118));
   AOI22_X1 i_0_0_237 (.A1(RAM_DATA_RD1[54]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[54]), .ZN(n_0_0_118));
   INV_X1 i_0_0_238 (.A(n_0_0_119), .ZN(n_0_119));
   AOI22_X1 i_0_0_239 (.A1(RAM_DATA_RD1[55]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[55]), .ZN(n_0_0_119));
   INV_X1 i_0_0_240 (.A(n_0_0_120), .ZN(n_0_120));
   AOI22_X1 i_0_0_241 (.A1(RAM_DATA_RD1[56]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[56]), .ZN(n_0_0_120));
   INV_X1 i_0_0_242 (.A(n_0_0_121), .ZN(n_0_121));
   AOI22_X1 i_0_0_243 (.A1(RAM_DATA_RD1[57]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[57]), .ZN(n_0_0_121));
   INV_X1 i_0_0_244 (.A(n_0_0_122), .ZN(n_0_122));
   AOI22_X1 i_0_0_245 (.A1(RAM_DATA_RD1[58]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[58]), .ZN(n_0_0_122));
   INV_X1 i_0_0_246 (.A(n_0_0_123), .ZN(n_0_123));
   AOI22_X1 i_0_0_247 (.A1(RAM_DATA_RD1[59]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[59]), .ZN(n_0_0_123));
   INV_X1 i_0_0_248 (.A(n_0_0_124), .ZN(n_0_124));
   AOI22_X1 i_0_0_249 (.A1(RAM_DATA_RD1[60]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[60]), .ZN(n_0_0_124));
   INV_X1 i_0_0_250 (.A(n_0_0_125), .ZN(n_0_125));
   AOI22_X1 i_0_0_251 (.A1(RAM_DATA_RD1[61]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[61]), .ZN(n_0_0_125));
   INV_X1 i_0_0_252 (.A(n_0_0_126), .ZN(n_0_126));
   AOI22_X1 i_0_0_253 (.A1(RAM_DATA_RD1[62]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[62]), .ZN(n_0_0_126));
   INV_X1 i_0_0_254 (.A(n_0_0_127), .ZN(n_0_127));
   AOI22_X1 i_0_0_255 (.A1(RAM_DATA_RD1[63]), .A2(n_0_0_497), .B1(n_0_0_128), 
      .B2(n_val[63]), .ZN(n_0_0_127));
   AOI21_X1 i_0_0_256 (.A(RST), .B1(n_0_0_281), .B2(n_0_0_499), .ZN(n_0_0_128));
   AND2_X1 i_0_0_257 (.A1(n_0_0_321), .A2(n_0_0_129), .ZN(n_0_128));
   OAI21_X1 i_0_0_258 (.A(n_0_0_130), .B1(n_0_0_139), .B2(n_0_0_322), .ZN(
      n_0_0_129));
   OAI21_X1 i_0_0_259 (.A(Final_Calc_Enable), .B1(n_0_0_219), .B2(n_0_0_322), 
      .ZN(n_0_0_130));
   OAI21_X1 i_0_0_260 (.A(n_0_0_226), .B1(n_0_0_131), .B2(RST), .ZN(n_0_129));
   OAI21_X1 i_0_0_261 (.A(Matrix_Multiplication2_Enable), .B1(n_0_0_608), 
      .B2(n_0_0_322), .ZN(n_0_0_131));
   INV_X1 i_0_0_262 (.A(n_0_0_132), .ZN(n_0_130));
   AOI22_X1 i_0_0_263 (.A1(Interpolate_DONE), .A2(n_0_0_475), .B1(n_0_0_133), 
      .B2(Matrix_Multiplication1_Enable), .ZN(n_0_0_132));
   AOI21_X1 i_0_0_264 (.A(RST), .B1(n_0_0_255), .B2(INT), .ZN(n_0_0_133));
   AOI21_X1 i_0_0_265 (.A(RST), .B1(n_0_0_327), .B2(n_0_0_134), .ZN(n_0_131));
   NAND2_X1 i_0_0_266 (.A1(n_0_0_219), .A2(counter[0]), .ZN(n_0_0_134));
   INV_X1 i_0_0_267 (.A(n_0_0_135), .ZN(n_0_132));
   AOI21_X1 i_0_0_268 (.A(n_0_0_446), .B1(n_0_0_136), .B2(n_0_0_219), .ZN(
      n_0_0_135));
   NOR2_X1 i_0_0_269 (.A1(n_0_0_301), .A2(RST), .ZN(n_0_0_136));
   OAI22_X1 i_0_0_270 (.A1(RST), .A2(n_0_0_137), .B1(n_0_0_184), .B2(n_0_0_553), 
      .ZN(n_0_133));
   AOI21_X1 i_0_0_271 (.A(n_0_0_138), .B1(n_0_0_228), .B2(n_0_0_255), .ZN(
      n_0_0_137));
   NAND3_X1 i_0_0_272 (.A1(n_0_0_139), .A2(n_0_0_299), .A3(n_0_0_181), .ZN(
      n_0_0_138));
   NAND4_X1 i_0_0_273 (.A1(n_0_0_152), .A2(n_0_0_542), .A3(n_0_0_140), .A4(
      n_0_0_165), .ZN(n_0_0_139));
   NOR3_X1 i_0_0_274 (.A1(n_0_0_148), .A2(n_0_0_143), .A3(n_0_0_141), .ZN(
      n_0_0_140));
   NAND4_X1 i_0_0_275 (.A1(n_0_0_158), .A2(n_0_0_597), .A3(n_0_0_609), .A4(
      n_0_0_176), .ZN(n_0_0_141));
   NAND4_X1 i_0_0_277 (.A1(n_0_0_147), .A2(n_0_0_144), .A3(n_0_0_154), .A4(
      n_0_0_153), .ZN(n_0_0_143));
   NOR3_X1 i_0_0_278 (.A1(n_0_0_145), .A2(n_0_0_167), .A3(n_0_0_150), .ZN(
      n_0_0_144));
   NAND3_X1 i_0_0_279 (.A1(n_0_0_174), .A2(n_0_0_596), .A3(n_0_0_541), .ZN(
      n_0_0_145));
   XOR2_X1 i_0_0_281 (.A(n_val[4]), .B(n_0_0_178), .Z(n_0_0_147));
   XNOR2_X1 i_0_0_282 (.A(n_val[10]), .B(n_0_0_170), .ZN(n_0_0_148));
   XNOR2_X1 i_0_0_284 (.A(n_val[3]), .B(n_0_0_171), .ZN(n_0_0_150));
   XNOR2_X1 i_0_0_285 (.A(n_val[5]), .B(n_0_0_156), .ZN(n_0_0_151));
   XOR2_X1 i_0_0_286 (.A(n_val[0]), .B(n_0_0_162), .Z(n_0_0_152));
   XOR2_X1 i_0_0_287 (.A(n_val[9]), .B(n_0_0_169), .Z(n_0_0_153));
   XOR2_X1 i_0_0_288 (.A(n_val[12]), .B(n_0_0_155), .Z(n_0_0_154));
   AOI22_X1 i_0_0_289 (.A1(MATRIX_CNT[12]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[12]), .ZN(n_0_0_155));
   AOI22_X1 i_0_0_290 (.A1(MATRIX_CNT[5]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[5]), .ZN(n_0_0_156));
   XOR2_X1 i_0_0_292 (.A(n_val[8]), .B(n_0_0_159), .Z(n_0_0_158));
   AOI22_X1 i_0_0_293 (.A1(MATRIX_CNT[8]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[8]), .ZN(n_0_0_159));
   AOI22_X1 i_0_0_296 (.A1(MATRIX_CNT[0]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[0]), .ZN(n_0_0_162));
   XNOR2_X1 i_0_0_297 (.A(n_val[2]), .B(n_0_0_164), .ZN(n_0_0_163));
   AOI22_X1 i_0_0_298 (.A1(MATRIX_CNT[2]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[2]), .ZN(n_0_0_164));
   XOR2_X1 i_0_0_299 (.A(n_val[1]), .B(n_0_0_166), .Z(n_0_0_165));
   AOI22_X1 i_0_0_300 (.A1(MATRIX_CNT[1]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[1]), .ZN(n_0_0_166));
   XNOR2_X1 i_0_0_301 (.A(n_val[6]), .B(n_0_0_168), .ZN(n_0_0_167));
   AOI22_X1 i_0_0_302 (.A1(MATRIX_CNT[6]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[6]), .ZN(n_0_0_168));
   AOI22_X1 i_0_0_303 (.A1(MATRIX_CNT[9]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[9]), .ZN(n_0_0_169));
   AOI22_X1 i_0_0_304 (.A1(MATRIX_CNT[10]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[10]), .ZN(n_0_0_170));
   AOI22_X1 i_0_0_305 (.A1(MATRIX_CNT[3]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[3]), .ZN(n_0_0_171));
   XOR2_X1 i_0_0_308 (.A(n_val[11]), .B(n_0_0_175), .Z(n_0_0_174));
   AOI22_X1 i_0_0_309 (.A1(MATRIX_CNT[11]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[11]), .ZN(n_0_0_175));
   XOR2_X1 i_0_0_310 (.A(n_val[7]), .B(n_0_0_177), .Z(n_0_0_176));
   AOI22_X1 i_0_0_311 (.A1(MATRIX_CNT[7]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[7]), .ZN(n_0_0_177));
   AOI22_X1 i_0_0_312 (.A1(MATRIX_CNT[4]), .A2(n_0_0_180), .B1(n_0_0_179), 
      .B2(NEW_MATRIX_CNT[4]), .ZN(n_0_0_178));
   NOR2_X1 i_0_0_313 (.A1(Matrix_Multiplication2_Enable), .A2(n_0_0_565), 
      .ZN(n_0_0_179));
   NOR2_X1 i_0_0_314 (.A1(n_0_0_566), .A2(Matrix_Multiplication2_Enable), 
      .ZN(n_0_0_180));
   NAND2_X1 i_0_0_315 (.A1(Interpolate_DONE), .A2(n_0_0_476), .ZN(n_0_0_181));
   OAI211_X1 i_0_0_316 (.A(n_0_0_496), .B(n_0_0_513), .C1(n_0_0_227), .C2(
      n_0_0_498), .ZN(n_0_134));
   NAND2_X1 i_0_0_317 (.A1(n_0_0_226), .A2(n_0_0_182), .ZN(n_0_135));
   NAND3_X1 i_0_0_318 (.A1(n_0_0_183), .A2(n_0_0_231), .A3(n_0_0_283), .ZN(
      n_0_0_182));
   NAND2_X1 i_0_0_319 (.A1(next[0]), .A2(n_0_0_184), .ZN(n_0_0_183));
   AND4_X1 i_0_0_320 (.A1(n_0_0_185), .A2(n_0_0_196), .A3(n_0_0_205), .A4(
      n_0_0_195), .ZN(n_0_0_184));
   NOR4_X1 i_0_0_321 (.A1(n_0_0_188), .A2(n_0_0_203), .A3(n_0_0_193), .A4(
      n_0_0_186), .ZN(n_0_0_185));
   OAI211_X1 i_0_0_322 (.A(n_0_0_187), .B(n_0_0_541), .C1(n_0_0_202), .C2(
      n_val[11]), .ZN(n_0_0_186));
   AOI221_X1 i_0_0_323 (.A(n_0_0_199), .B1(n_0_0_222), .B2(n_val[6]), .C1(
      n_val[11]), .C2(n_0_0_202), .ZN(n_0_0_187));
   OR4_X1 i_0_0_324 (.A1(n_0_0_191), .A2(n_0_0_211), .A3(n_val[13]), .A4(
      n_0_0_189), .ZN(n_0_0_188));
   OAI211_X1 i_0_0_325 (.A(n_0_0_190), .B(n_0_0_604), .C1(n_val[1]), .C2(
      n_0_0_208), .ZN(n_0_0_189));
   AOI22_X1 i_0_0_326 (.A1(n_val[2]), .A2(n_0_0_213), .B1(n_0_0_208), .B2(
      n_val[1]), .ZN(n_0_0_190));
   OAI211_X1 i_0_0_327 (.A(n_0_0_192), .B(n_0_0_209), .C1(n_0_0_214), .C2(
      n_val[5]), .ZN(n_0_0_191));
   AOI211_X1 i_0_0_328 (.A(n_0_0_574), .B(n_0_0_221), .C1(n_0_0_207), .C2(
      n_val[9]), .ZN(n_0_0_192));
   OAI21_X1 i_0_0_329 (.A(n_0_0_194), .B1(n_0_0_207), .B2(n_val[9]), .ZN(
      n_0_0_193));
   AOI21_X1 i_0_0_330 (.A(n_0_0_540), .B1(n_0_0_214), .B2(n_val[5]), .ZN(
      n_0_0_194));
   XOR2_X1 i_0_0_331 (.A(n_val[3]), .B(n_0_0_215), .Z(n_0_0_195));
   XOR2_X1 i_0_0_332 (.A(n_val[8]), .B(n_0_0_217), .Z(n_0_0_196));
   XNOR2_X1 i_0_0_335 (.A(n_val[12]), .B(n_0_0_218), .ZN(n_0_0_199));
   AOI22_X1 i_0_0_338 (.A1(VECTOR_CNT[11]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[11]), .ZN(n_0_0_202));
   XNOR2_X1 i_0_0_339 (.A(n_val[0]), .B(n_0_0_204), .ZN(n_0_0_203));
   AOI22_X1 i_0_0_340 (.A1(VECTOR_CNT[0]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[0]), .ZN(n_0_0_204));
   XOR2_X1 i_0_0_341 (.A(n_val[4]), .B(n_0_0_206), .Z(n_0_0_205));
   AOI22_X1 i_0_0_342 (.A1(VECTOR_CNT[4]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[4]), .ZN(n_0_0_206));
   AOI22_X1 i_0_0_343 (.A1(VECTOR_CNT[9]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[9]), .ZN(n_0_0_207));
   AOI22_X1 i_0_0_344 (.A1(VECTOR_CNT[1]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[1]), .ZN(n_0_0_208));
   XOR2_X1 i_0_0_345 (.A(n_val[10]), .B(n_0_0_210), .Z(n_0_0_209));
   AOI22_X1 i_0_0_346 (.A1(VECTOR_CNT[10]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[10]), .ZN(n_0_0_210));
   XNOR2_X1 i_0_0_347 (.A(n_val[7]), .B(n_0_0_212), .ZN(n_0_0_211));
   AOI22_X1 i_0_0_348 (.A1(VECTOR_CNT[7]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[7]), .ZN(n_0_0_212));
   AOI22_X1 i_0_0_349 (.A1(VECTOR_CNT[2]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[2]), .ZN(n_0_0_213));
   AOI22_X1 i_0_0_350 (.A1(VECTOR_CNT[5]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[5]), .ZN(n_0_0_214));
   AOI22_X1 i_0_0_351 (.A1(VECTOR_CNT[3]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[3]), .ZN(n_0_0_215));
   AOI22_X1 i_0_0_353 (.A1(VECTOR_CNT[8]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[8]), .ZN(n_0_0_217));
   AOI22_X1 i_0_0_354 (.A1(VECTOR_CNT[12]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[12]), .ZN(n_0_0_218));
   NOR2_X1 i_0_0_357 (.A1(n_val[6]), .A2(n_0_0_222), .ZN(n_0_0_221));
   AOI22_X1 i_0_0_358 (.A1(VECTOR_CNT[6]), .A2(n_0_0_225), .B1(n_0_0_223), 
      .B2(NEW_VECTOR_CNT[6]), .ZN(n_0_0_222));
   NOR2_X1 i_0_0_359 (.A1(Final_Calc_Enable), .A2(n_0_0_224), .ZN(n_0_0_223));
   NOR2_X1 i_0_0_360 (.A1(n_0_0_558), .A2(n_0_0_216), .ZN(n_0_0_224));
   NOR2_X1 i_0_0_361 (.A1(n_0_0_546), .A2(Final_Calc_Enable), .ZN(n_0_0_225));
   NAND3_X1 i_0_0_362 (.A1(n_0_0_255), .A2(n_0_0_231), .A3(n_0_0_227), .ZN(
      n_0_0_226));
   INV_X1 i_0_0_363 (.A(n_0_0_228), .ZN(n_0_0_227));
   OR4_X1 i_0_0_364 (.A1(n_0_0_242), .A2(n_0_0_241), .A3(n_0_0_235), .A4(
      n_0_0_229), .ZN(n_0_0_228));
   NAND4_X1 i_0_0_365 (.A1(n_0_0_234), .A2(n_0_0_514), .A3(n_0_0_230), .A4(
      n_0_0_252), .ZN(n_0_0_229));
   AOI221_X1 i_0_0_366 (.A(n_0_0_515), .B1(n_0_0_259), .B2(n_val[3]), .C1(
      n_val[9]), .C2(n_0_0_260), .ZN(n_0_0_230));
   OAI22_X1 i_0_0_369 (.A1(n_val[1]), .A2(n_0_0_261), .B1(n_0_0_256), .B2(
      n_val[0]), .ZN(n_0_0_233));
   AOI211_X1 i_0_0_370 (.A(n_0_0_574), .B(n_0_0_247), .C1(n_0_0_243), .C2(
      n_val[6]), .ZN(n_0_0_234));
   OAI211_X1 i_0_0_371 (.A(n_0_0_240), .B(n_0_0_236), .C1(n_val[3]), .C2(
      n_0_0_259), .ZN(n_0_0_235));
   AOI211_X1 i_0_0_372 (.A(n_val[14]), .B(n_0_0_237), .C1(n_val[1]), .C2(
      n_0_0_261), .ZN(n_0_0_236));
   OAI221_X1 i_0_0_373 (.A(n_0_0_238), .B1(n_0_0_243), .B2(n_val[6]), .C1(
      n_val[10]), .C2(n_0_0_254), .ZN(n_0_0_237));
   AOI22_X1 i_0_0_374 (.A1(n_val[12]), .A2(n_0_0_264), .B1(n_0_0_257), .B2(
      n_val[2]), .ZN(n_0_0_238));
   AOI221_X1 i_0_0_376 (.A(n_0_0_244), .B1(n_0_0_256), .B2(n_val[0]), .C1(
      n_val[4]), .C2(n_0_0_258), .ZN(n_0_0_240));
   OAI211_X1 i_0_0_377 (.A(n_0_0_262), .B(n_0_0_596), .C1(n_0_0_257), .C2(
      n_val[2]), .ZN(n_0_0_241));
   OAI221_X1 i_0_0_378 (.A(n_0_0_245), .B1(n_0_0_258), .B2(n_val[4]), .C1(
      n_val[9]), .C2(n_0_0_260), .ZN(n_0_0_242));
   AOI22_X1 i_0_0_379 (.A1(MATRIX_CNT[6]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[6]), .ZN(n_0_0_243));
   NOR2_X1 i_0_0_380 (.A1(n_val[7]), .A2(n_0_0_263), .ZN(n_0_0_244));
   XOR2_X1 i_0_0_381 (.A(n_val[5]), .B(n_0_0_246), .Z(n_0_0_245));
   AOI22_X1 i_0_0_382 (.A1(MATRIX_CNT[5]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[5]), .ZN(n_0_0_246));
   XNOR2_X1 i_0_0_383 (.A(n_val[11]), .B(n_0_0_248), .ZN(n_0_0_247));
   AOI22_X1 i_0_0_384 (.A1(MATRIX_CNT[11]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[11]), .ZN(n_0_0_248));
   XOR2_X1 i_0_0_388 (.A(n_val[8]), .B(n_0_0_253), .Z(n_0_0_252));
   AOI22_X1 i_0_0_389 (.A1(MATRIX_CNT[8]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[8]), .ZN(n_0_0_253));
   AOI22_X1 i_0_0_390 (.A1(MATRIX_CNT[10]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[10]), .ZN(n_0_0_254));
   AOI22_X1 i_0_0_392 (.A1(MATRIX_CNT[0]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[0]), .ZN(n_0_0_256));
   AOI22_X1 i_0_0_393 (.A1(MATRIX_CNT[2]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[2]), .ZN(n_0_0_257));
   AOI22_X1 i_0_0_394 (.A1(MATRIX_CNT[4]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[4]), .ZN(n_0_0_258));
   AOI22_X1 i_0_0_395 (.A1(MATRIX_CNT[3]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[3]), .ZN(n_0_0_259));
   AOI22_X1 i_0_0_396 (.A1(MATRIX_CNT[9]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[9]), .ZN(n_0_0_260));
   AOI22_X1 i_0_0_397 (.A1(MATRIX_CNT[1]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[1]), .ZN(n_0_0_261));
   NAND2_X1 i_0_0_398 (.A1(n_val[7]), .A2(n_0_0_263), .ZN(n_0_0_262));
   AOI22_X1 i_0_0_399 (.A1(MATRIX_CNT[7]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[7]), .ZN(n_0_0_263));
   AOI22_X1 i_0_0_400 (.A1(MATRIX_CNT[12]), .A2(n_0_0_266), .B1(n_0_0_265), 
      .B2(NEW_MATRIX_CNT[12]), .ZN(n_0_0_264));
   NOR2_X1 i_0_0_401 (.A1(Matrix_Multiplication1_Enable), .A2(n_0_0_565), 
      .ZN(n_0_0_265));
   NOR2_X1 i_0_0_402 (.A1(n_0_0_566), .A2(Matrix_Multiplication1_Enable), 
      .ZN(n_0_0_266));
   OAI21_X1 i_0_0_403 (.A(n_0_0_267), .B1(n_0_0_513), .B2(Interpolate_DONE), 
      .ZN(n_0_137));
   NAND2_X1 i_0_0_404 (.A1(n_0_0_474), .A2(Interpolate_Enable), .ZN(n_0_0_267));
   NAND2_X1 i_0_0_405 (.A1(n_0_0_416), .A2(n_0_0_268), .ZN(n_0_138));
   AOI22_X1 i_0_0_406 (.A1(n_0_0_284), .A2(NEW_MATRIX_ADD[0]), .B1(MATRIX_ADD[0]), 
      .B2(n_0_0_544), .ZN(n_0_0_268));
   NAND2_X1 i_0_0_407 (.A1(n_0_0_419), .A2(n_0_0_269), .ZN(n_0_139));
   AOI22_X1 i_0_0_408 (.A1(n_0_0_284), .A2(NEW_MATRIX_ADD[1]), .B1(MATRIX_ADD[1]), 
      .B2(n_0_0_544), .ZN(n_0_0_269));
   NAND2_X1 i_0_0_409 (.A1(n_0_0_417), .A2(n_0_0_270), .ZN(n_0_140));
   AOI22_X1 i_0_0_410 (.A1(n_0_0_284), .A2(NEW_MATRIX_ADD[2]), .B1(MATRIX_ADD[2]), 
      .B2(n_0_0_544), .ZN(n_0_0_270));
   NAND2_X1 i_0_0_411 (.A1(n_0_0_418), .A2(n_0_0_271), .ZN(n_0_141));
   AOI22_X1 i_0_0_412 (.A1(n_0_0_284), .A2(NEW_MATRIX_ADD[3]), .B1(MATRIX_ADD[3]), 
      .B2(n_0_0_544), .ZN(n_0_0_271));
   INV_X1 i_0_0_413 (.A(n_0_0_272), .ZN(n_0_142));
   AOI22_X1 i_0_0_414 (.A1(n_0_0_284), .A2(NEW_MATRIX_ADD[4]), .B1(MATRIX_ADD[4]), 
      .B2(n_0_0_544), .ZN(n_0_0_272));
   NAND2_X1 i_0_0_415 (.A1(n_0_0_273), .A2(n_0_0_399), .ZN(n_0_143));
   AOI22_X1 i_0_0_416 (.A1(n_0_0_284), .A2(NEW_MATRIX_ADD[5]), .B1(MATRIX_ADD[5]), 
      .B2(n_0_0_544), .ZN(n_0_0_273));
   NAND2_X1 i_0_0_417 (.A1(n_0_0_418), .A2(n_0_0_274), .ZN(n_0_144));
   AOI22_X1 i_0_0_418 (.A1(n_0_0_284), .A2(NEW_MATRIX_ADD[6]), .B1(MATRIX_ADD[6]), 
      .B2(n_0_0_544), .ZN(n_0_0_274));
   NAND2_X1 i_0_0_419 (.A1(n_0_0_418), .A2(n_0_0_275), .ZN(n_0_145));
   AOI22_X1 i_0_0_420 (.A1(n_0_0_284), .A2(NEW_MATRIX_ADD[7]), .B1(MATRIX_ADD[7]), 
      .B2(n_0_0_544), .ZN(n_0_0_275));
   INV_X1 i_0_0_421 (.A(n_0_0_276), .ZN(n_0_146));
   AOI221_X1 i_0_0_422 (.A(n_0_0_421), .B1(n_0_0_544), .B2(MATRIX_ADD[8]), 
      .C1(n_0_0_284), .C2(NEW_MATRIX_ADD[8]), .ZN(n_0_0_276));
   INV_X1 i_0_0_423 (.A(n_0_0_277), .ZN(n_0_147));
   AOI22_X1 i_0_0_424 (.A1(n_0_0_284), .A2(NEW_MATRIX_ADD[9]), .B1(MATRIX_ADD[9]), 
      .B2(n_0_0_544), .ZN(n_0_0_277));
   NAND2_X1 i_0_0_425 (.A1(n_0_0_278), .A2(n_0_0_399), .ZN(n_0_148));
   AOI22_X1 i_0_0_426 (.A1(n_0_0_284), .A2(NEW_MATRIX_ADD[10]), .B1(
      MATRIX_ADD[10]), .B2(n_0_0_544), .ZN(n_0_0_278));
   INV_X1 i_0_0_427 (.A(n_0_0_279), .ZN(n_0_149));
   AOI221_X1 i_0_0_428 (.A(n_0_0_421), .B1(n_0_0_544), .B2(MATRIX_ADD[11]), 
      .C1(n_0_0_284), .C2(NEW_MATRIX_ADD[11]), .ZN(n_0_0_279));
   NAND2_X1 i_0_0_429 (.A1(n_0_0_280), .A2(n_0_0_399), .ZN(n_0_150));
   AOI22_X1 i_0_0_430 (.A1(n_0_0_284), .A2(NEW_MATRIX_ADD[12]), .B1(
      MATRIX_ADD[12]), .B2(n_0_0_544), .ZN(n_0_0_280));
   OAI21_X1 i_0_0_437 (.A(n_0_0_285), .B1(n_0_0_551), .B2(Final_Calc_Enable), 
      .ZN(n_0_0_284));
   AOI21_X1 i_0_0_438 (.A(n_0_0_428), .B1(n_0_0_546), .B2(n_0_0_557), .ZN(
      n_0_0_285));
   NAND2_X1 i_0_0_439 (.A1(n_0_0_286), .A2(n_0_0_399), .ZN(n_0_154));
   AOI22_X1 i_0_0_440 (.A1(NEW_VECTOR2_ADD[0]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[0]), .ZN(n_0_0_286));
   NAND2_X1 i_0_0_441 (.A1(n_0_0_287), .A2(n_0_0_399), .ZN(n_0_155));
   AOI22_X1 i_0_0_442 (.A1(NEW_VECTOR2_ADD[1]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[1]), .ZN(n_0_0_287));
   NAND2_X1 i_0_0_443 (.A1(n_0_0_288), .A2(n_0_0_399), .ZN(n_0_156));
   AOI22_X1 i_0_0_444 (.A1(NEW_VECTOR2_ADD[2]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[2]), .ZN(n_0_0_288));
   INV_X1 i_0_0_445 (.A(n_0_0_289), .ZN(n_0_157));
   AOI22_X1 i_0_0_446 (.A1(NEW_VECTOR2_ADD[3]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[3]), .ZN(n_0_0_289));
   NAND2_X1 i_0_0_447 (.A1(n_0_0_290), .A2(n_0_0_399), .ZN(n_0_158));
   AOI22_X1 i_0_0_448 (.A1(NEW_VECTOR2_ADD[4]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[4]), .ZN(n_0_0_290));
   INV_X1 i_0_0_449 (.A(n_0_0_291), .ZN(n_0_159));
   AOI22_X1 i_0_0_450 (.A1(NEW_VECTOR2_ADD[5]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[5]), .ZN(n_0_0_291));
   NAND2_X1 i_0_0_451 (.A1(n_0_0_292), .A2(n_0_0_399), .ZN(n_0_160));
   AOI22_X1 i_0_0_452 (.A1(NEW_VECTOR2_ADD[6]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[6]), .ZN(n_0_0_292));
   INV_X1 i_0_0_453 (.A(n_0_0_293), .ZN(n_0_161));
   AOI22_X1 i_0_0_454 (.A1(NEW_VECTOR2_ADD[7]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[7]), .ZN(n_0_0_293));
   INV_X1 i_0_0_455 (.A(n_0_0_294), .ZN(n_0_162));
   AOI22_X1 i_0_0_456 (.A1(NEW_VECTOR2_ADD[8]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[8]), .ZN(n_0_0_294));
   INV_X1 i_0_0_457 (.A(n_0_0_295), .ZN(n_0_163));
   AOI22_X1 i_0_0_458 (.A1(NEW_VECTOR2_ADD[9]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[9]), .ZN(n_0_0_295));
   NAND2_X1 i_0_0_459 (.A1(n_0_0_296), .A2(n_0_0_399), .ZN(n_0_164));
   AOI22_X1 i_0_0_460 (.A1(NEW_VECTOR2_ADD[10]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[10]), .ZN(n_0_0_296));
   INV_X1 i_0_0_461 (.A(n_0_0_297), .ZN(n_0_165));
   AOI22_X1 i_0_0_462 (.A1(NEW_VECTOR2_ADD[11]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[11]), .ZN(n_0_0_297));
   NAND2_X1 i_0_0_463 (.A1(n_0_0_298), .A2(n_0_0_399), .ZN(n_0_166));
   AOI22_X1 i_0_0_464 (.A1(NEW_VECTOR2_ADD[12]), .A2(n_0_0_550), .B1(n_0_0_302), 
      .B2(VECTOR2_ADD[12]), .ZN(n_0_0_298));
   NOR2_X1 i_0_0_471 (.A1(n_0_0_216), .A2(n_0_0_303), .ZN(n_0_0_302));
   OAI21_X1 i_0_0_472 (.A(n_0_0_321), .B1(n_0_0_219), .B2(n_0_0_555), .ZN(
      n_0_0_303));
   NAND2_X1 i_0_0_473 (.A1(n_0_0_318), .A2(n_0_0_304), .ZN(n_0_170));
   AOI22_X1 i_0_0_474 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[0]), .B1(VECTOR_ADD[0]), 
      .B2(n_0_0_324), .ZN(n_0_0_304));
   NAND2_X1 i_0_0_475 (.A1(n_0_0_309), .A2(n_0_0_305), .ZN(n_0_171));
   AOI22_X1 i_0_0_476 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[1]), .B1(VECTOR_ADD[1]), 
      .B2(n_0_0_324), .ZN(n_0_0_305));
   NAND2_X1 i_0_0_477 (.A1(n_0_0_319), .A2(n_0_0_306), .ZN(n_0_172));
   AOI22_X1 i_0_0_478 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[2]), .B1(VECTOR_ADD[2]), 
      .B2(n_0_0_324), .ZN(n_0_0_306));
   NAND2_X1 i_0_0_479 (.A1(n_0_0_320), .A2(n_0_0_307), .ZN(n_0_173));
   AOI22_X1 i_0_0_480 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[3]), .B1(VECTOR_ADD[3]), 
      .B2(n_0_0_324), .ZN(n_0_0_307));
   NAND2_X1 i_0_0_481 (.A1(n_0_0_309), .A2(n_0_0_308), .ZN(n_0_174));
   AOI22_X1 i_0_0_482 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[4]), .B1(VECTOR_ADD[4]), 
      .B2(n_0_0_324), .ZN(n_0_0_308));
   NOR3_X1 i_0_0_483 (.A1(n_0_0_520), .A2(n_0_0_422), .A3(n_0_0_420), .ZN(
      n_0_0_309));
   NAND2_X1 i_0_0_484 (.A1(n_0_0_310), .A2(n_0_0_399), .ZN(n_0_175));
   AOI22_X1 i_0_0_485 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[5]), .B1(VECTOR_ADD[5]), 
      .B2(n_0_0_324), .ZN(n_0_0_310));
   NAND2_X1 i_0_0_486 (.A1(n_0_0_319), .A2(n_0_0_311), .ZN(n_0_176));
   AOI22_X1 i_0_0_487 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[6]), .B1(VECTOR_ADD[6]), 
      .B2(n_0_0_324), .ZN(n_0_0_311));
   NAND2_X1 i_0_0_488 (.A1(n_0_0_320), .A2(n_0_0_312), .ZN(n_0_177));
   AOI22_X1 i_0_0_489 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[7]), .B1(VECTOR_ADD[7]), 
      .B2(n_0_0_324), .ZN(n_0_0_312));
   INV_X1 i_0_0_490 (.A(n_0_0_313), .ZN(n_0_178));
   AOI22_X1 i_0_0_491 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[8]), .B1(VECTOR_ADD[8]), 
      .B2(n_0_0_324), .ZN(n_0_0_313));
   INV_X1 i_0_0_492 (.A(n_0_0_314), .ZN(n_0_179));
   AOI22_X1 i_0_0_493 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[9]), .B1(VECTOR_ADD[9]), 
      .B2(n_0_0_324), .ZN(n_0_0_314));
   NAND2_X1 i_0_0_494 (.A1(n_0_0_318), .A2(n_0_0_315), .ZN(n_0_180));
   AOI22_X1 i_0_0_495 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[10]), .B1(
      VECTOR_ADD[10]), .B2(n_0_0_324), .ZN(n_0_0_315));
   INV_X1 i_0_0_496 (.A(n_0_0_316), .ZN(n_0_181));
   AOI22_X1 i_0_0_497 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[11]), .B1(
      VECTOR_ADD[11]), .B2(n_0_0_324), .ZN(n_0_0_316));
   NAND2_X1 i_0_0_498 (.A1(n_0_0_318), .A2(n_0_0_317), .ZN(n_0_182));
   AOI22_X1 i_0_0_499 (.A1(n_0_0_326), .A2(NEW_VECTOR_ADD[12]), .B1(
      VECTOR_ADD[12]), .B2(n_0_0_324), .ZN(n_0_0_317));
   AND2_X1 i_0_0_500 (.A1(n_0_0_320), .A2(n_0_0_319), .ZN(n_0_0_318));
   NOR2_X1 i_0_0_501 (.A1(n_0_0_520), .A2(n_0_0_420), .ZN(n_0_0_319));
   NOR3_X1 i_0_0_502 (.A1(n_0_0_518), .A2(n_0_0_422), .A3(n_0_0_421), .ZN(
      n_0_0_320));
   AOI211_X1 i_0_0_509 (.A(RST), .B(n_0_0_255), .C1(n_0_0_325), .C2(n_0_0_283), 
      .ZN(n_0_0_324));
   OAI211_X1 i_0_0_510 (.A(n_0_0_555), .B(next[0]), .C1(counter[1]), .C2(
      counter[0]), .ZN(n_0_0_325));
   OAI21_X1 i_0_0_511 (.A(n_0_0_556), .B1(n_0_0_554), .B2(n_0_0_327), .ZN(
      n_0_0_326));
   OR3_X1 i_0_0_512 (.A1(n_0_0_219), .A2(counter[0]), .A3(counter[1]), .ZN(
      n_0_0_327));
   NAND4_X1 i_0_0_513 (.A1(n_0_0_416), .A2(n_0_0_330), .A3(n_0_0_329), .A4(
      n_0_0_328), .ZN(n_0_186));
   NAND2_X1 i_0_0_514 (.A1(NEW_MATRIX_ADD[0]), .A2(n_0_0_357), .ZN(n_0_0_328));
   NAND2_X1 i_0_0_515 (.A1(n_0_0_354), .A2(RAM_ADD_RD1[0]), .ZN(n_0_0_329));
   AOI221_X1 i_0_0_516 (.A(n_0_0_475), .B1(n_0_0_360), .B2(VECTOR2_ADD[0]), 
      .C1(n_0_0_359), .C2(VECTOR_ADD[0]), .ZN(n_0_0_330));
   NAND3_X1 i_0_0_517 (.A1(n_0_0_416), .A2(n_0_0_332), .A3(n_0_0_331), .ZN(
      n_0_187));
   AOI22_X1 i_0_0_518 (.A1(VECTOR_ADD[1]), .A2(n_0_0_359), .B1(n_0_0_357), 
      .B2(NEW_MATRIX_ADD[1]), .ZN(n_0_0_331));
   AOI22_X1 i_0_0_519 (.A1(n_0_0_354), .A2(RAM_ADD_RD1[1]), .B1(VECTOR2_ADD[1]), 
      .B2(n_0_0_360), .ZN(n_0_0_332));
   NAND3_X1 i_0_0_520 (.A1(n_0_0_417), .A2(n_0_0_334), .A3(n_0_0_333), .ZN(
      n_0_188));
   AOI22_X1 i_0_0_521 (.A1(n_0_0_354), .A2(RAM_ADD_RD1[2]), .B1(VECTOR2_ADD[2]), 
      .B2(n_0_0_360), .ZN(n_0_0_333));
   AOI22_X1 i_0_0_522 (.A1(VECTOR_ADD[2]), .A2(n_0_0_359), .B1(n_0_0_357), 
      .B2(NEW_MATRIX_ADD[2]), .ZN(n_0_0_334));
   NAND3_X1 i_0_0_523 (.A1(n_0_0_336), .A2(n_0_0_335), .A3(n_0_0_456), .ZN(
      n_0_189));
   AOI22_X1 i_0_0_524 (.A1(VECTOR_ADD[3]), .A2(n_0_0_359), .B1(n_0_0_357), 
      .B2(NEW_MATRIX_ADD[3]), .ZN(n_0_0_335));
   AOI22_X1 i_0_0_525 (.A1(n_0_0_354), .A2(RAM_ADD_RD1[3]), .B1(VECTOR2_ADD[3]), 
      .B2(n_0_0_360), .ZN(n_0_0_336));
   NAND2_X1 i_0_0_526 (.A1(n_0_0_338), .A2(n_0_0_337), .ZN(n_0_190));
   AOI22_X1 i_0_0_527 (.A1(n_0_0_354), .A2(RAM_ADD_RD1[4]), .B1(
      NEW_MATRIX_ADD[4]), .B2(n_0_0_357), .ZN(n_0_0_337));
   AOI221_X1 i_0_0_528 (.A(n_0_0_361), .B1(n_0_0_360), .B2(VECTOR2_ADD[4]), 
      .C1(n_0_0_359), .C2(VECTOR_ADD[4]), .ZN(n_0_0_338));
   NAND2_X1 i_0_0_529 (.A1(n_0_0_340), .A2(n_0_0_339), .ZN(n_0_191));
   AOI22_X1 i_0_0_530 (.A1(VECTOR2_ADD[5]), .A2(n_0_0_360), .B1(n_0_0_357), 
      .B2(NEW_MATRIX_ADD[5]), .ZN(n_0_0_339));
   AOI22_X1 i_0_0_531 (.A1(n_0_0_354), .A2(RAM_ADD_RD1[5]), .B1(VECTOR_ADD[5]), 
      .B2(n_0_0_359), .ZN(n_0_0_340));
   NAND3_X1 i_0_0_532 (.A1(n_0_0_341), .A2(n_0_0_456), .A3(n_0_0_342), .ZN(
      n_0_192));
   AOI221_X1 i_0_0_533 (.A(n_0_0_361), .B1(n_0_0_359), .B2(VECTOR_ADD[6]), 
      .C1(n_0_0_357), .C2(NEW_MATRIX_ADD[6]), .ZN(n_0_0_341));
   AOI22_X1 i_0_0_534 (.A1(n_0_0_354), .A2(RAM_ADD_RD1[6]), .B1(VECTOR2_ADD[6]), 
      .B2(n_0_0_360), .ZN(n_0_0_342));
   NAND3_X1 i_0_0_535 (.A1(n_0_0_344), .A2(n_0_0_343), .A3(n_0_0_456), .ZN(
      n_0_193));
   AOI22_X1 i_0_0_536 (.A1(VECTOR_ADD[7]), .A2(n_0_0_359), .B1(n_0_0_357), 
      .B2(NEW_MATRIX_ADD[7]), .ZN(n_0_0_343));
   AOI22_X1 i_0_0_537 (.A1(n_0_0_354), .A2(RAM_ADD_RD1[7]), .B1(VECTOR2_ADD[7]), 
      .B2(n_0_0_360), .ZN(n_0_0_344));
   NAND3_X1 i_0_0_538 (.A1(n_0_0_345), .A2(n_0_0_513), .A3(n_0_0_346), .ZN(
      n_0_194));
   AOI221_X1 i_0_0_539 (.A(n_0_0_421), .B1(n_0_0_359), .B2(VECTOR_ADD[8]), 
      .C1(n_0_0_354), .C2(RAM_ADD_RD1[8]), .ZN(n_0_0_345));
   AOI22_X1 i_0_0_540 (.A1(VECTOR2_ADD[8]), .A2(n_0_0_360), .B1(n_0_0_357), 
      .B2(NEW_MATRIX_ADD[8]), .ZN(n_0_0_346));
   NAND2_X1 i_0_0_541 (.A1(n_0_0_348), .A2(n_0_0_347), .ZN(n_0_195));
   AOI22_X1 i_0_0_542 (.A1(VECTOR2_ADD[9]), .A2(n_0_0_360), .B1(n_0_0_357), 
      .B2(NEW_MATRIX_ADD[9]), .ZN(n_0_0_347));
   AOI22_X1 i_0_0_543 (.A1(n_0_0_354), .A2(RAM_ADD_RD1[9]), .B1(VECTOR_ADD[9]), 
      .B2(n_0_0_359), .ZN(n_0_0_348));
   NAND2_X1 i_0_0_544 (.A1(n_0_0_350), .A2(n_0_0_349), .ZN(n_0_196));
   AOI22_X1 i_0_0_545 (.A1(n_0_0_354), .A2(RAM_ADD_RD1[10]), .B1(
      NEW_MATRIX_ADD[10]), .B2(n_0_0_357), .ZN(n_0_0_349));
   AOI221_X1 i_0_0_546 (.A(n_0_0_361), .B1(n_0_0_360), .B2(VECTOR2_ADD[10]), 
      .C1(n_0_0_359), .C2(VECTOR_ADD[10]), .ZN(n_0_0_350));
   NAND3_X1 i_0_0_547 (.A1(n_0_0_352), .A2(n_0_0_351), .A3(n_0_0_456), .ZN(
      n_0_197));
   AOI22_X1 i_0_0_548 (.A1(VECTOR_ADD[11]), .A2(n_0_0_359), .B1(n_0_0_357), 
      .B2(NEW_MATRIX_ADD[11]), .ZN(n_0_0_351));
   AOI22_X1 i_0_0_549 (.A1(n_0_0_354), .A2(RAM_ADD_RD1[11]), .B1(VECTOR2_ADD[11]), 
      .B2(n_0_0_360), .ZN(n_0_0_352));
   NAND2_X1 i_0_0_550 (.A1(n_0_0_358), .A2(n_0_0_353), .ZN(n_0_198));
   AOI22_X1 i_0_0_551 (.A1(n_0_0_354), .A2(RAM_ADD_RD1[12]), .B1(
      NEW_MATRIX_ADD[12]), .B2(n_0_0_357), .ZN(n_0_0_353));
   OAI21_X1 i_0_0_552 (.A(n_0_0_496), .B1(n_0_0_356), .B2(n_0_0_355), .ZN(
      n_0_0_354));
   OAI21_X1 i_0_0_553 (.A(n_0_0_231), .B1(n_0_0_397), .B2(next[2]), .ZN(
      n_0_0_355));
   AOI221_X1 i_0_0_554 (.A(next[1]), .B1(n_0_0_398), .B2(Back), .C1(n_0_0_427), 
      .C2(counter[1]), .ZN(n_0_0_356));
   AND2_X1 i_0_0_555 (.A1(n_0_0_429), .A2(n_0_0_231), .ZN(n_0_0_357));
   AOI221_X1 i_0_0_556 (.A(n_0_0_361), .B1(n_0_0_360), .B2(VECTOR2_ADD[12]), 
      .C1(n_0_0_359), .C2(VECTOR_ADD[12]), .ZN(n_0_0_358));
   NOR2_X1 i_0_0_557 (.A1(n_0_0_449), .A2(n_0_0_425), .ZN(n_0_0_359));
   NOR3_X1 i_0_0_558 (.A1(n_0_0_425), .A2(counter[0]), .A3(counter[1]), .ZN(
      n_0_0_360));
   NAND2_X1 i_0_0_559 (.A1(n_0_0_513), .A2(n_0_0_399), .ZN(n_0_0_361));
   NAND2_X1 i_0_0_560 (.A1(n_0_0_378), .A2(n_0_0_362), .ZN(n_0_199));
   AOI21_X1 i_0_0_561 (.A(n_0_0_363), .B1(n_0_0_383), .B2(NEW_VECTOR_ADD[0]), 
      .ZN(n_0_0_362));
   OAI21_X1 i_0_0_562 (.A(n_0_0_364), .B1(n_0_0_299), .B2(RST), .ZN(n_0_0_363));
   AOI22_X1 i_0_0_563 (.A1(RAM_ADD_RD2[0]), .A2(n_0_0_239), .B1(n_0_0_426), 
      .B2(MATRIX_ADD[0]), .ZN(n_0_0_364));
   NAND2_X1 i_0_0_564 (.A1(n_0_0_382), .A2(n_0_0_365), .ZN(n_0_200));
   AOI222_X1 i_0_0_565 (.A1(MATRIX_ADD[1]), .A2(n_0_0_426), .B1(n_0_0_383), 
      .B2(NEW_VECTOR_ADD[1]), .C1(RAM_ADD_RD2[1]), .C2(n_0_0_239), .ZN(n_0_0_365));
   NAND2_X1 i_0_0_566 (.A1(n_0_0_379), .A2(n_0_0_366), .ZN(n_0_201));
   AOI222_X1 i_0_0_567 (.A1(MATRIX_ADD[2]), .A2(n_0_0_426), .B1(n_0_0_383), 
      .B2(NEW_VECTOR_ADD[2]), .C1(RAM_ADD_RD2[2]), .C2(n_0_0_239), .ZN(n_0_0_366));
   NAND2_X1 i_0_0_568 (.A1(n_0_0_380), .A2(n_0_0_367), .ZN(n_0_202));
   AOI222_X1 i_0_0_569 (.A1(MATRIX_ADD[3]), .A2(n_0_0_426), .B1(n_0_0_383), 
      .B2(NEW_VECTOR_ADD[3]), .C1(RAM_ADD_RD2[3]), .C2(n_0_0_239), .ZN(n_0_0_367));
   NAND2_X1 i_0_0_570 (.A1(n_0_0_382), .A2(n_0_0_368), .ZN(n_0_203));
   AOI222_X1 i_0_0_571 (.A1(MATRIX_ADD[4]), .A2(n_0_0_426), .B1(n_0_0_383), 
      .B2(NEW_VECTOR_ADD[4]), .C1(RAM_ADD_RD2[4]), .C2(n_0_0_239), .ZN(n_0_0_368));
   NAND3_X1 i_0_0_572 (.A1(n_0_0_399), .A2(n_0_0_370), .A3(n_0_0_369), .ZN(
      n_0_204));
   AOI22_X1 i_0_0_573 (.A1(RAM_ADD_RD2[5]), .A2(n_0_0_239), .B1(n_0_0_426), 
      .B2(MATRIX_ADD[5]), .ZN(n_0_0_369));
   NAND2_X1 i_0_0_574 (.A1(NEW_VECTOR_ADD[5]), .A2(n_0_0_383), .ZN(n_0_0_370));
   NAND2_X1 i_0_0_575 (.A1(n_0_0_379), .A2(n_0_0_371), .ZN(n_0_205));
   AOI222_X1 i_0_0_576 (.A1(MATRIX_ADD[6]), .A2(n_0_0_426), .B1(n_0_0_383), 
      .B2(NEW_VECTOR_ADD[6]), .C1(RAM_ADD_RD2[6]), .C2(n_0_0_239), .ZN(n_0_0_371));
   NAND2_X1 i_0_0_577 (.A1(n_0_0_380), .A2(n_0_0_372), .ZN(n_0_206));
   AOI222_X1 i_0_0_578 (.A1(MATRIX_ADD[7]), .A2(n_0_0_426), .B1(n_0_0_383), 
      .B2(NEW_VECTOR_ADD[7]), .C1(RAM_ADD_RD2[7]), .C2(n_0_0_239), .ZN(n_0_0_372));
   INV_X1 i_0_0_579 (.A(n_0_0_373), .ZN(n_0_207));
   AOI222_X1 i_0_0_580 (.A1(MATRIX_ADD[8]), .A2(n_0_0_426), .B1(n_0_0_383), 
      .B2(NEW_VECTOR_ADD[8]), .C1(RAM_ADD_RD2[8]), .C2(n_0_0_239), .ZN(n_0_0_373));
   INV_X1 i_0_0_581 (.A(n_0_0_374), .ZN(n_0_208));
   AOI222_X1 i_0_0_582 (.A1(MATRIX_ADD[9]), .A2(n_0_0_426), .B1(n_0_0_383), 
      .B2(NEW_VECTOR_ADD[9]), .C1(RAM_ADD_RD2[9]), .C2(n_0_0_239), .ZN(n_0_0_374));
   NAND2_X1 i_0_0_583 (.A1(n_0_0_378), .A2(n_0_0_375), .ZN(n_0_209));
   AOI222_X1 i_0_0_584 (.A1(MATRIX_ADD[10]), .A2(n_0_0_426), .B1(n_0_0_383), 
      .B2(NEW_VECTOR_ADD[10]), .C1(RAM_ADD_RD2[10]), .C2(n_0_0_239), .ZN(
      n_0_0_375));
   INV_X1 i_0_0_585 (.A(n_0_0_376), .ZN(n_0_210));
   AOI222_X1 i_0_0_586 (.A1(MATRIX_ADD[11]), .A2(n_0_0_426), .B1(n_0_0_383), 
      .B2(NEW_VECTOR_ADD[11]), .C1(RAM_ADD_RD2[11]), .C2(n_0_0_239), .ZN(
      n_0_0_376));
   NAND2_X1 i_0_0_587 (.A1(n_0_0_378), .A2(n_0_0_377), .ZN(n_0_211));
   AOI222_X1 i_0_0_588 (.A1(MATRIX_ADD[12]), .A2(n_0_0_426), .B1(n_0_0_383), 
      .B2(NEW_VECTOR_ADD[12]), .C1(RAM_ADD_RD2[12]), .C2(n_0_0_239), .ZN(
      n_0_0_377));
   AND2_X1 i_0_0_589 (.A1(n_0_0_382), .A2(n_0_0_380), .ZN(n_0_0_378));
   AND2_X1 i_0_0_590 (.A1(n_0_0_382), .A2(n_0_0_399), .ZN(n_0_0_379));
   NOR2_X1 i_0_0_591 (.A1(n_0_0_422), .A2(n_0_0_381), .ZN(n_0_0_380));
   NOR3_X1 i_0_0_592 (.A1(n_0_0_561), .A2(n_0_0_498), .A3(n_0_0_397), .ZN(
      n_0_0_381));
   AOI21_X1 i_0_0_593 (.A(n_0_0_420), .B1(n_0_0_520), .B2(INT), .ZN(n_0_0_382));
   NOR3_X1 i_0_0_594 (.A1(n_0_0_560), .A2(n_0_0_322), .A3(RST), .ZN(n_0_0_383));
   NAND2_X1 i_0_0_595 (.A1(n_0_0_416), .A2(n_0_0_384), .ZN(n_0_212));
   AOI22_X1 i_0_0_596 (.A1(n_0_0_400), .A2(NEW_RESULT_ADD[0]), .B1(n_0_0_401), 
      .B2(RESULT_ADD[0]), .ZN(n_0_0_384));
   NAND2_X1 i_0_0_597 (.A1(n_0_0_418), .A2(n_0_0_385), .ZN(n_0_213));
   AOI22_X1 i_0_0_598 (.A1(n_0_0_400), .A2(NEW_RESULT_ADD[1]), .B1(n_0_0_401), 
      .B2(RESULT_ADD[1]), .ZN(n_0_0_385));
   NAND2_X1 i_0_0_599 (.A1(n_0_0_417), .A2(n_0_0_386), .ZN(n_0_214));
   AOI22_X1 i_0_0_600 (.A1(n_0_0_400), .A2(NEW_RESULT_ADD[2]), .B1(n_0_0_401), 
      .B2(RESULT_ADD[2]), .ZN(n_0_0_386));
   NAND2_X1 i_0_0_601 (.A1(n_0_0_416), .A2(n_0_0_387), .ZN(n_0_215));
   AOI22_X1 i_0_0_602 (.A1(n_0_0_400), .A2(NEW_RESULT_ADD[3]), .B1(n_0_0_401), 
      .B2(RESULT_ADD[3]), .ZN(n_0_0_387));
   NAND2_X1 i_0_0_603 (.A1(n_0_0_418), .A2(n_0_0_388), .ZN(n_0_216));
   AOI22_X1 i_0_0_604 (.A1(n_0_0_400), .A2(NEW_RESULT_ADD[4]), .B1(n_0_0_401), 
      .B2(RESULT_ADD[4]), .ZN(n_0_0_388));
   NAND2_X1 i_0_0_605 (.A1(n_0_0_419), .A2(n_0_0_389), .ZN(n_0_217));
   AOI22_X1 i_0_0_606 (.A1(n_0_0_400), .A2(NEW_RESULT_ADD[5]), .B1(n_0_0_401), 
      .B2(RESULT_ADD[5]), .ZN(n_0_0_389));
   INV_X1 i_0_0_607 (.A(n_0_0_390), .ZN(n_0_218));
   AOI221_X1 i_0_0_608 (.A(n_0_0_420), .B1(n_0_0_401), .B2(RESULT_ADD[6]), 
      .C1(n_0_0_400), .C2(NEW_RESULT_ADD[6]), .ZN(n_0_0_390));
   NAND2_X1 i_0_0_609 (.A1(n_0_0_419), .A2(n_0_0_391), .ZN(n_0_219));
   AOI22_X1 i_0_0_610 (.A1(n_0_0_400), .A2(NEW_RESULT_ADD[7]), .B1(n_0_0_401), 
      .B2(RESULT_ADD[7]), .ZN(n_0_0_391));
   NAND2_X1 i_0_0_611 (.A1(n_0_0_392), .A2(n_0_0_399), .ZN(n_0_220));
   AOI22_X1 i_0_0_612 (.A1(n_0_0_400), .A2(NEW_RESULT_ADD[8]), .B1(n_0_0_401), 
      .B2(RESULT_ADD[8]), .ZN(n_0_0_392));
   INV_X1 i_0_0_613 (.A(n_0_0_393), .ZN(n_0_221));
   AOI22_X1 i_0_0_614 (.A1(n_0_0_400), .A2(NEW_RESULT_ADD[9]), .B1(n_0_0_401), 
      .B2(RESULT_ADD[9]), .ZN(n_0_0_393));
   NAND2_X1 i_0_0_615 (.A1(n_0_0_416), .A2(n_0_0_394), .ZN(n_0_222));
   AOI22_X1 i_0_0_616 (.A1(n_0_0_400), .A2(NEW_RESULT_ADD[10]), .B1(n_0_0_401), 
      .B2(RESULT_ADD[10]), .ZN(n_0_0_394));
   INV_X1 i_0_0_617 (.A(n_0_0_395), .ZN(n_0_223));
   AOI22_X1 i_0_0_618 (.A1(n_0_0_400), .A2(NEW_RESULT_ADD[11]), .B1(n_0_0_401), 
      .B2(RESULT_ADD[11]), .ZN(n_0_0_395));
   NAND2_X1 i_0_0_619 (.A1(n_0_0_416), .A2(n_0_0_396), .ZN(n_0_224));
   AOI22_X1 i_0_0_620 (.A1(n_0_0_400), .A2(NEW_RESULT_ADD[12]), .B1(n_0_0_401), 
      .B2(RESULT_ADD[12]), .ZN(n_0_0_396));
   NAND3_X1 i_0_0_627 (.A1(n_0_0_549), .A2(n_0_0_519), .A3(n_0_0_517), .ZN(
      n_0_0_400));
   OAI211_X1 i_0_0_628 (.A(n_0_0_543), .B(n_0_0_525), .C1(n_0_0_402), .C2(RST), 
      .ZN(n_0_0_401));
   NAND2_X1 i_0_0_629 (.A1(next[1]), .A2(n_0_0_523), .ZN(n_0_0_402));
   NAND2_X1 i_0_0_630 (.A1(n_0_0_416), .A2(n_0_0_403), .ZN(n_0_228));
   AOI22_X1 i_0_0_631 (.A1(n_0_0_423), .A2(RESULT_ADD[0]), .B1(RAM_ADD_WR[0]), 
      .B2(n_0_0_249), .ZN(n_0_0_403));
   NAND2_X1 i_0_0_632 (.A1(n_0_0_418), .A2(n_0_0_404), .ZN(n_0_229));
   AOI22_X1 i_0_0_633 (.A1(n_0_0_423), .A2(RESULT_ADD[1]), .B1(RAM_ADD_WR[1]), 
      .B2(n_0_0_249), .ZN(n_0_0_404));
   NAND2_X1 i_0_0_634 (.A1(n_0_0_417), .A2(n_0_0_405), .ZN(n_0_230));
   AOI22_X1 i_0_0_635 (.A1(n_0_0_423), .A2(RESULT_ADD[2]), .B1(RAM_ADD_WR[2]), 
      .B2(n_0_0_249), .ZN(n_0_0_405));
   NAND2_X1 i_0_0_636 (.A1(n_0_0_416), .A2(n_0_0_406), .ZN(n_0_231));
   AOI22_X1 i_0_0_637 (.A1(n_0_0_423), .A2(RESULT_ADD[3]), .B1(RAM_ADD_WR[3]), 
      .B2(n_0_0_249), .ZN(n_0_0_406));
   NAND2_X1 i_0_0_638 (.A1(n_0_0_418), .A2(n_0_0_407), .ZN(n_0_232));
   AOI22_X1 i_0_0_639 (.A1(n_0_0_423), .A2(RESULT_ADD[4]), .B1(RAM_ADD_WR[4]), 
      .B2(n_0_0_249), .ZN(n_0_0_407));
   NAND2_X1 i_0_0_640 (.A1(n_0_0_419), .A2(n_0_0_408), .ZN(n_0_233));
   AOI22_X1 i_0_0_641 (.A1(n_0_0_423), .A2(RESULT_ADD[5]), .B1(RAM_ADD_WR[5]), 
      .B2(n_0_0_249), .ZN(n_0_0_408));
   INV_X1 i_0_0_642 (.A(n_0_0_409), .ZN(n_0_234));
   AOI221_X1 i_0_0_643 (.A(n_0_0_420), .B1(n_0_0_249), .B2(RAM_ADD_WR[6]), 
      .C1(n_0_0_423), .C2(RESULT_ADD[6]), .ZN(n_0_0_409));
   NAND2_X1 i_0_0_644 (.A1(n_0_0_419), .A2(n_0_0_410), .ZN(n_0_235));
   AOI22_X1 i_0_0_645 (.A1(n_0_0_423), .A2(RESULT_ADD[7]), .B1(RAM_ADD_WR[7]), 
      .B2(n_0_0_249), .ZN(n_0_0_410));
   NAND2_X1 i_0_0_646 (.A1(n_0_0_411), .A2(n_0_0_399), .ZN(n_0_236));
   AOI22_X1 i_0_0_647 (.A1(n_0_0_423), .A2(RESULT_ADD[8]), .B1(RAM_ADD_WR[8]), 
      .B2(n_0_0_249), .ZN(n_0_0_411));
   INV_X1 i_0_0_648 (.A(n_0_0_412), .ZN(n_0_237));
   AOI22_X1 i_0_0_649 (.A1(n_0_0_423), .A2(RESULT_ADD[9]), .B1(RAM_ADD_WR[9]), 
      .B2(n_0_0_249), .ZN(n_0_0_412));
   NAND2_X1 i_0_0_650 (.A1(n_0_0_416), .A2(n_0_0_413), .ZN(n_0_238));
   AOI22_X1 i_0_0_651 (.A1(n_0_0_423), .A2(RESULT_ADD[10]), .B1(RAM_ADD_WR[10]), 
      .B2(n_0_0_249), .ZN(n_0_0_413));
   INV_X1 i_0_0_652 (.A(n_0_0_414), .ZN(n_0_239));
   AOI22_X1 i_0_0_653 (.A1(n_0_0_423), .A2(RESULT_ADD[11]), .B1(RAM_ADD_WR[11]), 
      .B2(n_0_0_249), .ZN(n_0_0_414));
   NAND2_X1 i_0_0_654 (.A1(n_0_0_416), .A2(n_0_0_415), .ZN(n_0_240));
   AOI22_X1 i_0_0_655 (.A1(n_0_0_423), .A2(RESULT_ADD[12]), .B1(RAM_ADD_WR[12]), 
      .B2(n_0_0_249), .ZN(n_0_0_415));
   NOR3_X1 i_0_0_656 (.A1(n_0_0_422), .A2(n_0_0_421), .A3(n_0_0_420), .ZN(
      n_0_0_416));
   NOR2_X1 i_0_0_657 (.A1(n_0_0_422), .A2(n_0_0_420), .ZN(n_0_0_417));
   NOR2_X1 i_0_0_658 (.A1(n_0_0_422), .A2(n_0_0_421), .ZN(n_0_0_418));
   NOR2_X1 i_0_0_659 (.A1(n_0_0_421), .A2(n_0_0_420), .ZN(n_0_0_419));
   NOR3_X1 i_0_0_660 (.A1(n_0_0_608), .A2(n_0_0_526), .A3(RST), .ZN(n_0_0_420));
   AND3_X1 i_0_0_661 (.A1(Matrix_Multiplication1_Enable), .A2(n_0_0_255), 
      .A3(n_0_0_231), .ZN(n_0_0_421));
   NOR2_X1 i_0_0_662 (.A1(n_0_0_555), .A2(n_0_0_553), .ZN(n_0_0_422));
   OR3_X1 i_0_0_663 (.A1(n_0_0_428), .A2(n_0_0_426), .A3(n_0_0_424), .ZN(
      n_0_0_423));
   NOR3_X1 i_0_0_664 (.A1(INT), .A2(RST), .A3(n_0_0_250), .ZN(n_0_0_424));
   INV_X1 i_0_0_665 (.A(n_0_0_426), .ZN(n_0_0_425));
   AND3_X1 i_0_0_666 (.A1(n_0_0_283), .A2(n_0_0_231), .A3(n_0_0_427), .ZN(
      n_0_0_426));
   NOR2_X1 i_0_0_667 (.A1(n_0_0_323), .A2(Final_Calc_Enable), .ZN(n_0_0_427));
   AND2_X1 i_0_0_668 (.A1(n_0_0_321), .A2(n_0_0_429), .ZN(n_0_0_428));
   OAI22_X1 i_0_0_669 (.A1(Matrix_Multiplication1_Enable), .A2(n_0_0_251), 
      .B1(n_0_0_608), .B2(Matrix_Multiplication2_Enable), .ZN(n_0_0_429));
   INV_X1 i_0_0_670 (.A(n_0_0_430), .ZN(n_0_241));
   AOI222_X1 i_0_0_671 (.A1(n_0_0_450), .A2(NEW_Element_Result[0]), .B1(
      RAM_DATA_RD1[0]), .B2(n_0_0_446), .C1(Element_Result[0]), .C2(n_0_0_447), 
      .ZN(n_0_0_430));
   INV_X1 i_0_0_672 (.A(n_0_0_431), .ZN(n_0_242));
   AOI222_X1 i_0_0_673 (.A1(n_0_0_450), .A2(NEW_Element_Result[1]), .B1(
      RAM_DATA_RD1[1]), .B2(n_0_0_446), .C1(Element_Result[1]), .C2(n_0_0_447), 
      .ZN(n_0_0_431));
   INV_X1 i_0_0_674 (.A(n_0_0_432), .ZN(n_0_243));
   AOI222_X1 i_0_0_675 (.A1(n_0_0_450), .A2(NEW_Element_Result[2]), .B1(
      RAM_DATA_RD1[2]), .B2(n_0_0_446), .C1(Element_Result[2]), .C2(n_0_0_447), 
      .ZN(n_0_0_432));
   INV_X1 i_0_0_676 (.A(n_0_0_433), .ZN(n_0_244));
   AOI222_X1 i_0_0_677 (.A1(n_0_0_450), .A2(NEW_Element_Result[3]), .B1(
      RAM_DATA_RD1[3]), .B2(n_0_0_446), .C1(Element_Result[3]), .C2(n_0_0_447), 
      .ZN(n_0_0_433));
   INV_X1 i_0_0_678 (.A(n_0_0_434), .ZN(n_0_245));
   AOI222_X1 i_0_0_679 (.A1(n_0_0_450), .A2(NEW_Element_Result[4]), .B1(
      RAM_DATA_RD1[4]), .B2(n_0_0_446), .C1(Element_Result[4]), .C2(n_0_0_447), 
      .ZN(n_0_0_434));
   INV_X1 i_0_0_680 (.A(n_0_0_435), .ZN(n_0_246));
   AOI222_X1 i_0_0_681 (.A1(n_0_0_450), .A2(NEW_Element_Result[5]), .B1(
      RAM_DATA_RD1[5]), .B2(n_0_0_446), .C1(Element_Result[5]), .C2(n_0_0_447), 
      .ZN(n_0_0_435));
   INV_X1 i_0_0_682 (.A(n_0_0_436), .ZN(n_0_247));
   AOI222_X1 i_0_0_683 (.A1(n_0_0_450), .A2(NEW_Element_Result[6]), .B1(
      RAM_DATA_RD1[6]), .B2(n_0_0_446), .C1(Element_Result[6]), .C2(n_0_0_447), 
      .ZN(n_0_0_436));
   INV_X1 i_0_0_684 (.A(n_0_0_437), .ZN(n_0_248));
   AOI222_X1 i_0_0_685 (.A1(n_0_0_450), .A2(NEW_Element_Result[7]), .B1(
      RAM_DATA_RD1[7]), .B2(n_0_0_446), .C1(Element_Result[7]), .C2(n_0_0_447), 
      .ZN(n_0_0_437));
   INV_X1 i_0_0_686 (.A(n_0_0_438), .ZN(n_0_249));
   AOI222_X1 i_0_0_687 (.A1(n_0_0_450), .A2(NEW_Element_Result[8]), .B1(
      RAM_DATA_RD1[8]), .B2(n_0_0_446), .C1(Element_Result[8]), .C2(n_0_0_447), 
      .ZN(n_0_0_438));
   INV_X1 i_0_0_688 (.A(n_0_0_439), .ZN(n_0_250));
   AOI222_X1 i_0_0_689 (.A1(n_0_0_450), .A2(NEW_Element_Result[9]), .B1(
      RAM_DATA_RD1[9]), .B2(n_0_0_446), .C1(Element_Result[9]), .C2(n_0_0_447), 
      .ZN(n_0_0_439));
   INV_X1 i_0_0_690 (.A(n_0_0_440), .ZN(n_0_251));
   AOI222_X1 i_0_0_691 (.A1(n_0_0_450), .A2(NEW_Element_Result[10]), .B1(
      RAM_DATA_RD1[10]), .B2(n_0_0_446), .C1(Element_Result[10]), .C2(n_0_0_447), 
      .ZN(n_0_0_440));
   INV_X1 i_0_0_696 (.A(n_0_0_443), .ZN(n_0_254));
   AOI222_X1 i_0_0_697 (.A1(n_0_0_450), .A2(NEW_Element_Result[13]), .B1(
      RAM_DATA_RD1[13]), .B2(n_0_0_446), .C1(Element_Result[13]), .C2(n_0_0_447), 
      .ZN(n_0_0_443));
   INV_X1 i_0_0_698 (.A(n_0_0_444), .ZN(n_0_255));
   AOI222_X1 i_0_0_699 (.A1(n_0_0_450), .A2(NEW_Element_Result[14]), .B1(
      RAM_DATA_RD1[14]), .B2(n_0_0_446), .C1(Element_Result[14]), .C2(n_0_0_447), 
      .ZN(n_0_0_444));
   INV_X1 i_0_0_700 (.A(n_0_0_445), .ZN(n_0_256));
   AOI222_X1 i_0_0_701 (.A1(n_0_0_450), .A2(NEW_Element_Result[15]), .B1(
      RAM_DATA_RD1[15]), .B2(n_0_0_446), .C1(Element_Result[15]), .C2(n_0_0_447), 
      .ZN(n_0_0_445));
   AOI21_X1 i_0_0_704 (.A(n_0_0_282), .B1(n_0_0_449), .B2(next[0]), .ZN(
      n_0_0_448));
   NAND2_X1 i_0_0_705 (.A1(n_0_0_301), .A2(counter[0]), .ZN(n_0_0_449));
   OAI21_X1 i_0_0_707 (.A(n_0_0_559), .B1(n_0_0_455), .B2(n_0_0_452), .ZN(
      n_0_0_451));
   NAND2_X1 i_0_0_708 (.A1(n_0_0_454), .A2(n_0_0_453), .ZN(n_0_0_452));
   NOR4_X1 i_0_0_709 (.A1(NEW_VECTOR_CNT[7]), .A2(NEW_VECTOR_CNT[6]), .A3(
      NEW_VECTOR_CNT[5]), .A4(NEW_VECTOR_CNT[4]), .ZN(n_0_0_453));
   NOR4_X1 i_0_0_710 (.A1(NEW_VECTOR_CNT[3]), .A2(NEW_VECTOR_CNT[2]), .A3(
      NEW_VECTOR_CNT[1]), .A4(NEW_VECTOR_CNT[0]), .ZN(n_0_0_454));
   NAND2_X1 i_0_0_711 (.A1(n_0_0_457), .A2(n_0_0_629), .ZN(n_0_0_455));
   NOR4_X1 i_0_0_713 (.A1(NEW_VECTOR_CNT[11]), .A2(NEW_VECTOR_CNT[10]), .A3(
      NEW_VECTOR_CNT[9]), .A4(NEW_VECTOR_CNT[8]), .ZN(n_0_0_457));
   INV_X1 i_0_0_714 (.A(n_0_0_458), .ZN(n_0_257));
   AOI22_X1 i_0_0_715 (.A1(RAM_DATA_RD1[0]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_15), .ZN(n_0_0_458));
   INV_X1 i_0_0_716 (.A(n_0_0_459), .ZN(n_0_258));
   AOI22_X1 i_0_0_717 (.A1(RAM_DATA_RD1[1]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_14), .ZN(n_0_0_459));
   INV_X1 i_0_0_718 (.A(n_0_0_460), .ZN(n_0_259));
   AOI22_X1 i_0_0_719 (.A1(RAM_DATA_RD1[2]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_13), .ZN(n_0_0_460));
   INV_X1 i_0_0_720 (.A(n_0_0_461), .ZN(n_0_260));
   AOI22_X1 i_0_0_721 (.A1(RAM_DATA_RD1[3]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_12), .ZN(n_0_0_461));
   INV_X1 i_0_0_722 (.A(n_0_0_462), .ZN(n_0_261));
   AOI22_X1 i_0_0_723 (.A1(RAM_DATA_RD1[4]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_11), .ZN(n_0_0_462));
   INV_X1 i_0_0_724 (.A(n_0_0_463), .ZN(n_0_262));
   AOI22_X1 i_0_0_725 (.A1(RAM_DATA_RD1[5]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_10), .ZN(n_0_0_463));
   INV_X1 i_0_0_726 (.A(n_0_0_464), .ZN(n_0_263));
   AOI22_X1 i_0_0_727 (.A1(RAM_DATA_RD1[6]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_9), .ZN(n_0_0_464));
   INV_X1 i_0_0_728 (.A(n_0_0_465), .ZN(n_0_264));
   AOI22_X1 i_0_0_729 (.A1(RAM_DATA_RD1[7]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_8), .ZN(n_0_0_465));
   INV_X1 i_0_0_730 (.A(n_0_0_466), .ZN(n_0_265));
   AOI22_X1 i_0_0_731 (.A1(RAM_DATA_RD1[8]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_7), .ZN(n_0_0_466));
   INV_X1 i_0_0_732 (.A(n_0_0_467), .ZN(n_0_266));
   AOI22_X1 i_0_0_733 (.A1(RAM_DATA_RD1[9]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_6), .ZN(n_0_0_467));
   INV_X1 i_0_0_734 (.A(n_0_0_468), .ZN(n_0_267));
   AOI22_X1 i_0_0_735 (.A1(RAM_DATA_RD1[10]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_5), .ZN(n_0_0_468));
   INV_X1 i_0_0_736 (.A(n_0_0_469), .ZN(n_0_268));
   AOI22_X1 i_0_0_737 (.A1(RAM_DATA_RD1[11]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_4), .ZN(n_0_0_469));
   INV_X1 i_0_0_738 (.A(n_0_0_470), .ZN(n_0_269));
   AOI22_X1 i_0_0_739 (.A1(RAM_DATA_RD1[12]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_3), .ZN(n_0_0_470));
   INV_X1 i_0_0_740 (.A(n_0_0_471), .ZN(n_0_270));
   AOI22_X1 i_0_0_741 (.A1(RAM_DATA_RD1[13]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_2), .ZN(n_0_0_471));
   INV_X1 i_0_0_742 (.A(n_0_0_472), .ZN(n_0_271));
   AOI22_X1 i_0_0_743 (.A1(RAM_DATA_RD1[14]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_1), .ZN(n_0_0_472));
   INV_X1 i_0_0_744 (.A(n_0_0_473), .ZN(n_0_272));
   AOI22_X1 i_0_0_745 (.A1(RAM_DATA_RD1[15]), .A2(n_0_0_475), .B1(n_0_0_474), 
      .B2(n_0), .ZN(n_0_0_473));
   AOI21_X1 i_0_0_746 (.A(RST), .B1(n_0_0_476), .B2(INT), .ZN(n_0_0_474));
   AND2_X1 i_0_0_747 (.A1(n_0_0_231), .A2(n_0_0_476), .ZN(n_0_0_475));
   NOR3_X1 i_0_0_748 (.A1(n_0_0_397), .A2(next[0]), .A3(next[2]), .ZN(n_0_0_476));
   INV_X1 i_0_0_749 (.A(n_0_0_477), .ZN(n_0_273));
   AOI222_X1 i_0_0_750 (.A1(FINAL_RESULT[0]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[0]), .C1(n_0_0_494), .C2(NEW_Element_Result[0]), .ZN(
      n_0_0_477));
   INV_X1 i_0_0_751 (.A(n_0_0_478), .ZN(n_0_274));
   AOI222_X1 i_0_0_752 (.A1(FINAL_RESULT[1]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[1]), .C1(n_0_0_494), .C2(NEW_Element_Result[1]), .ZN(
      n_0_0_478));
   INV_X1 i_0_0_753 (.A(n_0_0_479), .ZN(n_0_275));
   AOI222_X1 i_0_0_754 (.A1(FINAL_RESULT[2]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[2]), .C1(n_0_0_494), .C2(NEW_Element_Result[2]), .ZN(
      n_0_0_479));
   INV_X1 i_0_0_755 (.A(n_0_0_480), .ZN(n_0_276));
   AOI222_X1 i_0_0_756 (.A1(FINAL_RESULT[3]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[3]), .C1(n_0_0_494), .C2(NEW_Element_Result[3]), .ZN(
      n_0_0_480));
   INV_X1 i_0_0_757 (.A(n_0_0_481), .ZN(n_0_277));
   AOI222_X1 i_0_0_758 (.A1(FINAL_RESULT[4]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[4]), .C1(n_0_0_494), .C2(NEW_Element_Result[4]), .ZN(
      n_0_0_481));
   INV_X1 i_0_0_759 (.A(n_0_0_482), .ZN(n_0_278));
   AOI222_X1 i_0_0_760 (.A1(FINAL_RESULT[5]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[5]), .C1(n_0_0_494), .C2(NEW_Element_Result[5]), .ZN(
      n_0_0_482));
   INV_X1 i_0_0_761 (.A(n_0_0_483), .ZN(n_0_279));
   AOI222_X1 i_0_0_762 (.A1(FINAL_RESULT[6]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[6]), .C1(n_0_0_494), .C2(NEW_Element_Result[6]), .ZN(
      n_0_0_483));
   INV_X1 i_0_0_763 (.A(n_0_0_484), .ZN(n_0_280));
   AOI222_X1 i_0_0_764 (.A1(FINAL_RESULT[7]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[7]), .C1(n_0_0_494), .C2(NEW_Element_Result[7]), .ZN(
      n_0_0_484));
   INV_X1 i_0_0_765 (.A(n_0_0_485), .ZN(n_0_281));
   AOI222_X1 i_0_0_766 (.A1(FINAL_RESULT[8]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[8]), .C1(n_0_0_494), .C2(NEW_Element_Result[8]), .ZN(
      n_0_0_485));
   INV_X1 i_0_0_767 (.A(n_0_0_486), .ZN(n_0_282));
   AOI222_X1 i_0_0_768 (.A1(FINAL_RESULT[9]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[9]), .C1(n_0_0_494), .C2(NEW_Element_Result[9]), .ZN(
      n_0_0_486));
   INV_X1 i_0_0_769 (.A(n_0_0_487), .ZN(n_0_283));
   AOI222_X1 i_0_0_770 (.A1(FINAL_RESULT[10]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[10]), .C1(n_0_0_494), .C2(NEW_Element_Result[10]), 
      .ZN(n_0_0_487));
   INV_X1 i_0_0_775 (.A(n_0_0_490), .ZN(n_0_286));
   AOI222_X1 i_0_0_776 (.A1(FINAL_RESULT[13]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[13]), .C1(n_0_0_494), .C2(NEW_Element_Result[13]), 
      .ZN(n_0_0_490));
   INV_X1 i_0_0_777 (.A(n_0_0_491), .ZN(n_0_287));
   AOI222_X1 i_0_0_778 (.A1(FINAL_RESULT[14]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[14]), .C1(n_0_0_494), .C2(NEW_Element_Result[14]), 
      .ZN(n_0_0_491));
   INV_X1 i_0_0_779 (.A(n_0_0_492), .ZN(n_0_288));
   AOI222_X1 i_0_0_780 (.A1(FINAL_RESULT[15]), .A2(n_0_0_552), .B1(n_0_0_545), 
      .B2(RAM_DATA_WR[15]), .C1(n_0_0_494), .C2(NEW_Element_Result[15]), 
      .ZN(n_0_0_492));
   INV_X1 i_0_0_781 (.A(n_0_0_494), .ZN(n_0_0_493));
   NOR4_X1 i_0_0_783 (.A1(n_0_0_495), .A2(next[0]), .A3(next[1]), .A4(next[2]), 
      .ZN(n_0_289));
   NAND2_X1 i_0_0_784 (.A1(n_0_0_496), .A2(n_0_0_495), .ZN(n_0_290));
   NAND2_X1 i_0_0_785 (.A1(Back), .A2(n_0_0_231), .ZN(n_0_0_495));
   NAND3_X1 i_0_0_786 (.A1(n_0_0_281), .A2(n_0_0_231), .A3(n_0_0_397), .ZN(
      n_0_0_496));
   NOR2_X1 i_0_0_787 (.A1(n_0_0_498), .A2(next[1]), .ZN(n_0_0_497));
   NAND2_X1 i_0_0_788 (.A1(n_0_0_281), .A2(n_0_0_231), .ZN(n_0_0_498));
   NOR2_X1 i_0_0_789 (.A1(n_0_0_322), .A2(next[1]), .ZN(n_0_0_499));
   INV_X1 i_0_0_790 (.A(n_0_0_500), .ZN(n_0_291));
   AOI22_X1 i_0_0_791 (.A1(MATRIX_CNT[0]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[0]), .ZN(n_0_0_500));
   INV_X1 i_0_0_792 (.A(n_0_0_501), .ZN(n_0_292));
   AOI22_X1 i_0_0_793 (.A1(MATRIX_CNT[1]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[1]), .ZN(n_0_0_501));
   INV_X1 i_0_0_794 (.A(n_0_0_502), .ZN(n_0_293));
   AOI22_X1 i_0_0_795 (.A1(MATRIX_CNT[2]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[2]), .ZN(n_0_0_502));
   INV_X1 i_0_0_796 (.A(n_0_0_503), .ZN(n_0_294));
   AOI22_X1 i_0_0_797 (.A1(MATRIX_CNT[3]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[3]), .ZN(n_0_0_503));
   INV_X1 i_0_0_798 (.A(n_0_0_504), .ZN(n_0_295));
   AOI22_X1 i_0_0_799 (.A1(MATRIX_CNT[4]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[4]), .ZN(n_0_0_504));
   INV_X1 i_0_0_800 (.A(n_0_0_505), .ZN(n_0_296));
   AOI22_X1 i_0_0_801 (.A1(MATRIX_CNT[5]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[5]), .ZN(n_0_0_505));
   INV_X1 i_0_0_802 (.A(n_0_0_506), .ZN(n_0_297));
   AOI22_X1 i_0_0_803 (.A1(MATRIX_CNT[6]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[6]), .ZN(n_0_0_506));
   INV_X1 i_0_0_804 (.A(n_0_0_507), .ZN(n_0_298));
   AOI22_X1 i_0_0_805 (.A1(MATRIX_CNT[7]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[7]), .ZN(n_0_0_507));
   INV_X1 i_0_0_806 (.A(n_0_0_508), .ZN(n_0_299));
   AOI22_X1 i_0_0_807 (.A1(MATRIX_CNT[8]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[8]), .ZN(n_0_0_508));
   INV_X1 i_0_0_808 (.A(n_0_0_509), .ZN(n_0_300));
   AOI22_X1 i_0_0_809 (.A1(MATRIX_CNT[9]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[9]), .ZN(n_0_0_509));
   INV_X1 i_0_0_810 (.A(n_0_0_510), .ZN(n_0_301));
   AOI22_X1 i_0_0_811 (.A1(MATRIX_CNT[10]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[10]), .ZN(n_0_0_510));
   INV_X1 i_0_0_812 (.A(n_0_0_511), .ZN(n_0_302));
   AOI22_X1 i_0_0_813 (.A1(MATRIX_CNT[11]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[11]), .ZN(n_0_0_511));
   INV_X1 i_0_0_814 (.A(n_0_0_512), .ZN(n_0_303));
   AOI22_X1 i_0_0_815 (.A1(MATRIX_CNT[12]), .A2(n_0_0_521), .B1(n_0_0_516), 
      .B2(NEW_MATRIX_CNT[12]), .ZN(n_0_0_512));
   NAND2_X1 i_0_0_822 (.A1(n_0_0_519), .A2(n_0_0_517), .ZN(n_0_0_516));
   NAND2_X1 i_0_0_823 (.A1(n_0_0_518), .A2(n_0_0_524), .ZN(n_0_0_517));
   NOR2_X1 i_0_0_824 (.A1(n_0_0_610), .A2(RST), .ZN(n_0_0_518));
   NAND2_X1 i_0_0_825 (.A1(n_0_0_520), .A2(n_0_0_526), .ZN(n_0_0_519));
   NOR2_X1 i_0_0_826 (.A1(n_0_0_567), .A2(RST), .ZN(n_0_0_520));
   OAI21_X1 i_0_0_827 (.A(n_0_0_525), .B1(n_0_0_522), .B2(RST), .ZN(n_0_0_521));
   OAI21_X1 i_0_0_828 (.A(n_0_0_608), .B1(n_0_0_523), .B2(n_0_0_251), .ZN(
      n_0_0_522));
   AND2_X1 i_0_0_829 (.A1(n_0_0_612), .A2(n_0_0_524), .ZN(n_0_0_523));
   NAND2_X1 i_0_0_830 (.A1(INT), .A2(Matrix_Multiplication1_Enable), .ZN(
      n_0_0_524));
   NAND4_X1 i_0_0_831 (.A1(n_0_0_323), .A2(n_0_0_321), .A3(n_0_0_568), .A4(
      n_0_0_526), .ZN(n_0_0_525));
   NAND2_X1 i_0_0_832 (.A1(INT), .A2(Matrix_Multiplication2_Enable), .ZN(
      n_0_0_526));
   INV_X1 i_0_0_833 (.A(n_0_0_527), .ZN(n_0_151));
   AOI22_X1 i_0_0_834 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[0]), .B1(VECTOR_CNT[0]), 
      .B2(n_0_0_544), .ZN(n_0_0_527));
   INV_X1 i_0_0_835 (.A(n_0_0_528), .ZN(n_0_152));
   AOI22_X1 i_0_0_836 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[1]), .B1(VECTOR_CNT[1]), 
      .B2(n_0_0_544), .ZN(n_0_0_528));
   INV_X1 i_0_0_837 (.A(n_0_0_529), .ZN(n_0_153));
   AOI22_X1 i_0_0_838 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[2]), .B1(VECTOR_CNT[2]), 
      .B2(n_0_0_544), .ZN(n_0_0_529));
   INV_X1 i_0_0_839 (.A(n_0_0_530), .ZN(n_0_167));
   AOI22_X1 i_0_0_840 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[3]), .B1(VECTOR_CNT[3]), 
      .B2(n_0_0_544), .ZN(n_0_0_530));
   INV_X1 i_0_0_841 (.A(n_0_0_531), .ZN(n_0_168));
   AOI22_X1 i_0_0_842 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[4]), .B1(VECTOR_CNT[4]), 
      .B2(n_0_0_544), .ZN(n_0_0_531));
   INV_X1 i_0_0_843 (.A(n_0_0_532), .ZN(n_0_169));
   AOI22_X1 i_0_0_844 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[5]), .B1(VECTOR_CNT[5]), 
      .B2(n_0_0_544), .ZN(n_0_0_532));
   INV_X1 i_0_0_845 (.A(n_0_0_533), .ZN(n_0_183));
   AOI22_X1 i_0_0_846 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[6]), .B1(VECTOR_CNT[6]), 
      .B2(n_0_0_544), .ZN(n_0_0_533));
   INV_X1 i_0_0_847 (.A(n_0_0_534), .ZN(n_0_184));
   AOI22_X1 i_0_0_848 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[7]), .B1(VECTOR_CNT[7]), 
      .B2(n_0_0_544), .ZN(n_0_0_534));
   INV_X1 i_0_0_849 (.A(n_0_0_535), .ZN(n_0_185));
   AOI22_X1 i_0_0_850 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[8]), .B1(VECTOR_CNT[8]), 
      .B2(n_0_0_544), .ZN(n_0_0_535));
   INV_X1 i_0_0_851 (.A(n_0_0_536), .ZN(n_0_225));
   AOI22_X1 i_0_0_852 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[9]), .B1(VECTOR_CNT[9]), 
      .B2(n_0_0_544), .ZN(n_0_0_536));
   INV_X1 i_0_0_853 (.A(n_0_0_537), .ZN(n_0_226));
   AOI22_X1 i_0_0_854 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[10]), .B1(
      VECTOR_CNT[10]), .B2(n_0_0_544), .ZN(n_0_0_537));
   INV_X1 i_0_0_855 (.A(n_0_0_538), .ZN(n_0_227));
   AOI22_X1 i_0_0_856 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[11]), .B1(
      VECTOR_CNT[11]), .B2(n_0_0_544), .ZN(n_0_0_538));
   INV_X1 i_0_0_857 (.A(n_0_0_539), .ZN(n_0_304));
   AOI22_X1 i_0_0_858 (.A1(n_0_0_548), .A2(NEW_VECTOR_CNT[12]), .B1(
      VECTOR_CNT[12]), .B2(n_0_0_544), .ZN(n_0_0_539));
   INV_X1 i_0_0_865 (.A(n_0_0_544), .ZN(n_0_0_543));
   NOR3_X1 i_0_0_866 (.A1(RST), .A2(n_0_0_547), .A3(n_0_0_546), .ZN(n_0_0_544));
   OAI211_X1 i_0_0_868 (.A(n_0_0_251), .B(n_0_0_608), .C1(n_0_0_220), .C2(
      counter[0]), .ZN(n_0_0_546));
   NOR2_X1 i_0_0_869 (.A1(n_0_0_250), .A2(n_0_0_555), .ZN(n_0_0_547));
   NAND2_X1 i_0_0_870 (.A1(n_0_0_556), .A2(n_0_0_549), .ZN(n_0_0_548));
   INV_X1 i_0_0_871 (.A(n_0_0_550), .ZN(n_0_0_549));
   AND2_X1 i_0_0_872 (.A1(n_0_0_552), .A2(n_0_0_555), .ZN(n_0_0_550));
   INV_X1 i_0_0_873 (.A(n_0_0_552), .ZN(n_0_0_551));
   NAND3_X1 i_0_0_875 (.A1(next[0]), .A2(n_0_0_283), .A3(n_0_0_321), .ZN(
      n_0_0_553));
   NAND2_X1 i_0_0_876 (.A1(n_0_0_321), .A2(n_0_0_555), .ZN(n_0_0_554));
   NAND2_X1 i_0_0_877 (.A1(INT), .A2(Final_Calc_Enable), .ZN(n_0_0_555));
   AOI21_X1 i_0_0_878 (.A(n_0_0_559), .B1(n_0_0_558), .B2(n_0_0_557), .ZN(
      n_0_0_556));
   NOR2_X1 i_0_0_879 (.A1(INT), .A2(RST), .ZN(n_0_0_557));
   OAI21_X1 i_0_0_880 (.A(n_0_0_563), .B1(n_0_0_611), .B2(n_0_0_251), .ZN(
      n_0_0_558));
   NOR2_X1 i_0_0_881 (.A1(RST), .A2(n_0_0_560), .ZN(n_0_0_559));
   AOI21_X1 i_0_0_882 (.A(n_0_0_562), .B1(n_0_0_561), .B2(n_0_0_255), .ZN(
      n_0_0_560));
   NOR2_X1 i_0_0_883 (.A1(Matrix_Multiplication1_Enable), .A2(n_0_0_611), 
      .ZN(n_0_0_561));
   NOR2_X1 i_0_0_884 (.A1(n_0_0_563), .A2(Matrix_Multiplication2_Enable), 
      .ZN(n_0_0_562));
   NAND2_X1 i_0_0_885 (.A1(n_0_0_568), .A2(n_0_0_609), .ZN(n_0_0_563));
   NAND2_X1 i_0_0_886 (.A1(n_0_0_232), .A2(n_0_0_564), .ZN(n_0_305));
   OAI21_X1 i_0_0_887 (.A(n_0_0_231), .B1(n_0_0_566), .B2(n_0_0_216), .ZN(
      n_0_0_564));
   INV_X1 i_0_0_888 (.A(n_0_0_566), .ZN(n_0_0_565));
   NAND2_X1 i_0_0_889 (.A1(n_0_0_610), .A2(n_0_0_567), .ZN(n_0_0_566));
   OR2_X1 i_0_0_890 (.A1(n_0_0_608), .A2(n_0_0_568), .ZN(n_0_0_567));
   NAND3_X1 i_0_0_891 (.A1(n_0_0_573), .A2(n_0_0_572), .A3(n_0_0_569), .ZN(
      n_0_0_568));
   NOR4_X1 i_0_0_892 (.A1(n_0_0_601), .A2(n_0_0_574), .A3(n_0_0_571), .A4(
      n_0_0_570), .ZN(n_0_0_569));
   NAND4_X1 i_0_0_893 (.A1(n_0_0_605), .A2(n_0_0_604), .A3(n_0_0_603), .A4(
      n_0_0_602), .ZN(n_0_0_570));
   NAND3_X1 i_0_0_894 (.A1(n_0_0_600), .A2(n_0_0_596), .A3(n_0_0_592), .ZN(
      n_0_0_571));
   NOR4_X1 i_0_0_895 (.A1(n_0_0_599), .A2(n_0_0_598), .A3(n_0_0_595), .A4(
      n_0_0_593), .ZN(n_0_0_572));
   NOR4_X1 i_0_0_896 (.A1(n_0_0_607), .A2(n_0_0_606), .A3(n_val[15]), .A4(
      n_0_0_594), .ZN(n_0_0_573));
   NAND4_X1 i_0_0_897 (.A1(n_0_0_588), .A2(n_0_0_587), .A3(n_0_0_586), .A4(
      n_0_0_575), .ZN(n_0_0_574));
   NOR2_X1 i_0_0_898 (.A1(n_0_0_581), .A2(n_0_0_576), .ZN(n_0_0_575));
   NAND4_X1 i_0_0_899 (.A1(n_0_0_580), .A2(n_0_0_579), .A3(n_0_0_578), .A4(
      n_0_0_577), .ZN(n_0_0_576));
   NOR4_X1 i_0_0_900 (.A1(n_val[51]), .A2(n_val[50]), .A3(n_val[49]), .A4(
      n_val[48]), .ZN(n_0_0_577));
   NOR4_X1 i_0_0_901 (.A1(n_val[55]), .A2(n_val[54]), .A3(n_val[53]), .A4(
      n_val[52]), .ZN(n_0_0_578));
   NOR4_X1 i_0_0_902 (.A1(n_val[63]), .A2(n_val[62]), .A3(n_val[61]), .A4(
      n_val[60]), .ZN(n_0_0_579));
   NOR4_X1 i_0_0_903 (.A1(n_val[59]), .A2(n_val[58]), .A3(n_val[57]), .A4(
      n_val[56]), .ZN(n_0_0_580));
   NAND4_X1 i_0_0_904 (.A1(n_0_0_585), .A2(n_0_0_584), .A3(n_0_0_583), .A4(
      n_0_0_582), .ZN(n_0_0_581));
   NOR4_X1 i_0_0_905 (.A1(n_val[39]), .A2(n_val[38]), .A3(n_val[37]), .A4(
      n_val[36]), .ZN(n_0_0_582));
   NOR4_X1 i_0_0_906 (.A1(n_val[35]), .A2(n_val[34]), .A3(n_val[33]), .A4(
      n_val[32]), .ZN(n_0_0_583));
   NOR4_X1 i_0_0_907 (.A1(n_val[43]), .A2(n_val[42]), .A3(n_val[41]), .A4(
      n_val[40]), .ZN(n_0_0_584));
   NOR4_X1 i_0_0_908 (.A1(n_val[47]), .A2(n_val[46]), .A3(n_val[45]), .A4(
      n_val[44]), .ZN(n_0_0_585));
   NOR4_X1 i_0_0_909 (.A1(n_val[23]), .A2(n_val[22]), .A3(n_val[21]), .A4(
      n_val[20]), .ZN(n_0_0_586));
   NOR4_X1 i_0_0_910 (.A1(n_val[19]), .A2(n_val[18]), .A3(n_val[17]), .A4(
      n_val[16]), .ZN(n_0_0_587));
   AND3_X1 i_0_0_911 (.A1(n_0_0_591), .A2(n_0_0_590), .A3(n_0_0_589), .ZN(
      n_0_0_588));
   NOR4_X1 i_0_0_912 (.A1(n_val[31]), .A2(n_val[30]), .A3(n_val[29]), .A4(
      n_val[28]), .ZN(n_0_0_589));
   NOR2_X1 i_0_0_913 (.A1(n_val[27]), .A2(n_val[24]), .ZN(n_0_0_590));
   NOR2_X1 i_0_0_914 (.A1(n_val[26]), .A2(n_val[25]), .ZN(n_0_0_591));
   XNOR2_X1 i_0_0_915 (.A(n_val[12]), .B(NEW_VECTOR_CNT[12]), .ZN(n_0_0_592));
   XOR2_X1 i_0_0_916 (.A(n_val[7]), .B(NEW_VECTOR_CNT[7]), .Z(n_0_0_593));
   XOR2_X1 i_0_0_917 (.A(n_val[8]), .B(NEW_VECTOR_CNT[8]), .Z(n_0_0_594));
   XOR2_X1 i_0_0_918 (.A(n_val[5]), .B(NEW_VECTOR_CNT[5]), .Z(n_0_0_595));
   XOR2_X1 i_0_0_921 (.A(n_val[11]), .B(NEW_VECTOR_CNT[11]), .Z(n_0_0_598));
   XOR2_X1 i_0_0_922 (.A(n_val[2]), .B(NEW_VECTOR_CNT[2]), .Z(n_0_0_599));
   XNOR2_X1 i_0_0_923 (.A(n_val[10]), .B(NEW_VECTOR_CNT[10]), .ZN(n_0_0_600));
   XOR2_X1 i_0_0_924 (.A(n_val[3]), .B(NEW_VECTOR_CNT[3]), .Z(n_0_0_601));
   XNOR2_X1 i_0_0_925 (.A(n_val[1]), .B(NEW_VECTOR_CNT[1]), .ZN(n_0_0_602));
   XNOR2_X1 i_0_0_926 (.A(n_val[4]), .B(NEW_VECTOR_CNT[4]), .ZN(n_0_0_603));
   XNOR2_X1 i_0_0_928 (.A(n_val[6]), .B(NEW_VECTOR_CNT[6]), .ZN(n_0_0_605));
   XOR2_X1 i_0_0_929 (.A(n_val[9]), .B(NEW_VECTOR_CNT[9]), .Z(n_0_0_606));
   XOR2_X1 i_0_0_930 (.A(n_val[0]), .B(NEW_VECTOR_CNT[0]), .Z(n_0_0_607));
   NAND2_X1 i_0_0_931 (.A1(n_0_0_283), .A2(n_0_0_323), .ZN(n_0_0_608));
   NOR2_X1 i_0_0_932 (.A1(n_0_0_282), .A2(next[0]), .ZN(n_0_0_609));
   NAND2_X1 i_0_0_933 (.A1(n_0_0_255), .A2(n_0_0_611), .ZN(n_0_0_610));
   INV_X1 i_0_0_934 (.A(n_0_0_612), .ZN(n_0_0_611));
   NAND4_X1 i_0_0_935 (.A1(n_0_0_619), .A2(n_0_0_618), .A3(n_0_0_617), .A4(
      n_0_0_613), .ZN(n_0_0_612));
   NOR3_X1 i_0_0_936 (.A1(n_0_0_616), .A2(n_0_0_615), .A3(n_0_0_614), .ZN(
      n_0_0_613));
   NAND4_X1 i_0_0_937 (.A1(n_0_0_634), .A2(n_0_0_628), .A3(n_0_0_627), .A4(
      n_0_0_201), .ZN(n_0_0_614));
   NAND4_X1 i_0_0_938 (.A1(n_0_0_633), .A2(n_0_0_631), .A3(n_0_0_630), .A4(
      n_0_0_623), .ZN(n_0_0_615));
   NAND4_X1 i_0_0_939 (.A1(n_0_0_157), .A2(n_0_0_142), .A3(n_0_0_637), .A4(
      n_0_0_636), .ZN(n_0_0_616));
   AND4_X1 i_0_0_940 (.A1(n_0_0_635), .A2(n_0_0_625), .A3(n_0_0_624), .A4(
      n_0_0_622), .ZN(n_0_0_617));
   NOR4_X1 i_0_0_941 (.A1(n_0_0_200), .A2(n_0_0_197), .A3(n_0_0_160), .A4(
      m_val[15]), .ZN(n_0_0_618));
   NOR4_X1 i_0_0_942 (.A1(n_0_0_632), .A2(n_0_0_621), .A3(n_0_0_620), .A4(
      n_0_0_198), .ZN(n_0_0_619));
   NAND3_X1 i_0_0_943 (.A1(n_0_0_161), .A2(n_0_0_638), .A3(n_0_0_626), .ZN(
      n_0_0_620));
   XOR2_X1 i_0_0_944 (.A(NEW_VECTOR_CNT[4]), .B(m_val[4]), .Z(n_0_0_621));
   NOR4_X1 i_0_0_945 (.A1(m_val[63]), .A2(m_val[62]), .A3(m_val[61]), .A4(
      m_val[60]), .ZN(n_0_0_622));
   XNOR2_X1 i_0_0_947 (.A(NEW_VECTOR_CNT[7]), .B(m_val[7]), .ZN(n_0_0_624));
   NOR4_X1 i_0_0_948 (.A1(m_val[51]), .A2(m_val[50]), .A3(m_val[49]), .A4(
      m_val[48]), .ZN(n_0_0_625));
   NOR4_X1 i_0_0_949 (.A1(m_val[47]), .A2(m_val[46]), .A3(m_val[45]), .A4(
      m_val[44]), .ZN(n_0_0_626));
   NOR4_X1 i_0_0_950 (.A1(m_val[59]), .A2(m_val[58]), .A3(m_val[57]), .A4(
      m_val[56]), .ZN(n_0_0_627));
   NOR4_X1 i_0_0_951 (.A1(m_val[55]), .A2(m_val[54]), .A3(m_val[53]), .A4(
      m_val[52]), .ZN(n_0_0_628));
   XNOR2_X1 i_0_0_953 (.A(NEW_VECTOR_CNT[0]), .B(m_val[0]), .ZN(n_0_0_630));
   XNOR2_X1 i_0_0_954 (.A(NEW_VECTOR_CNT[9]), .B(m_val[9]), .ZN(n_0_0_631));
   XOR2_X1 i_0_0_955 (.A(NEW_VECTOR_CNT[11]), .B(m_val[11]), .Z(n_0_0_632));
   XNOR2_X1 i_0_0_956 (.A(NEW_VECTOR_CNT[3]), .B(m_val[3]), .ZN(n_0_0_633));
   XNOR2_X1 i_0_0_957 (.A(NEW_VECTOR_CNT[10]), .B(m_val[10]), .ZN(n_0_0_634));
   XNOR2_X1 i_0_0_959 (.A(NEW_VECTOR_CNT[8]), .B(m_val[8]), .ZN(n_0_0_636));
   NOR4_X1 i_0_0_960 (.A1(m_val[31]), .A2(m_val[30]), .A3(m_val[29]), .A4(
      m_val[28]), .ZN(n_0_0_637));
   NOR4_X1 i_0_0_961 (.A1(m_val[35]), .A2(m_val[34]), .A3(m_val[33]), .A4(
      m_val[32]), .ZN(n_0_0_638));
   NOR4_X1 i_0_0_962 (.A1(n_0_0_149), .A2(n_0_0_146), .A3(m_val[43]), .A4(
      m_val[42]), .ZN(n_0_0_142));
   OR2_X1 i_0_0_963 (.A1(m_val[41]), .A2(m_val[40]), .ZN(n_0_0_146));
   OR4_X1 i_0_0_964 (.A1(m_val[39]), .A2(m_val[38]), .A3(m_val[37]), .A4(
      m_val[36]), .ZN(n_0_0_149));
   NOR4_X1 i_0_0_965 (.A1(m_val[19]), .A2(m_val[18]), .A3(m_val[17]), .A4(
      m_val[16]), .ZN(n_0_0_157));
   XOR2_X1 i_0_0_966 (.A(NEW_VECTOR_CNT[2]), .B(m_val[2]), .Z(n_0_0_160));
   NOR4_X1 i_0_0_967 (.A1(n_0_0_172), .A2(m_val[20]), .A3(m_val[21]), .A4(
      n_0_0_173), .ZN(n_0_0_161));
   OR4_X1 i_0_0_968 (.A1(m_val[27]), .A2(m_val[26]), .A3(m_val[25]), .A4(
      m_val[24]), .ZN(n_0_0_172));
   OR2_X1 i_0_0_969 (.A1(m_val[23]), .A2(m_val[22]), .ZN(n_0_0_173));
   XOR2_X1 i_0_0_970 (.A(NEW_VECTOR_CNT[12]), .B(m_val[12]), .Z(n_0_0_197));
   XOR2_X1 i_0_0_971 (.A(NEW_VECTOR_CNT[5]), .B(m_val[5]), .Z(n_0_0_198));
   XOR2_X1 i_0_0_972 (.A(NEW_VECTOR_CNT[1]), .B(m_val[1]), .Z(n_0_0_200));
   XNOR2_X1 i_0_0_973 (.A(NEW_VECTOR_CNT[6]), .B(m_val[6]), .ZN(n_0_0_201));
   NOR3_X1 i_0_0_974 (.A1(n_0_0_301), .A2(n_0_0_219), .A3(counter[0]), .ZN(
      n_0_0_216));
   NAND2_X1 i_0_0_975 (.A1(next[0]), .A2(n_0_0_283), .ZN(n_0_0_219));
   NAND2_X1 i_0_0_976 (.A1(counter[1]), .A2(n_0_0_283), .ZN(n_0_0_220));
   NOR2_X1 i_0_0_977 (.A1(n_0_0_322), .A2(RST), .ZN(n_0_0_231));
   NAND2_X1 i_0_0_978 (.A1(RAM_ENABLE_WR), .A2(n_0_0_239), .ZN(n_0_0_232));
   AND2_X1 i_0_0_979 (.A1(n_0_0_299), .A2(n_0_0_249), .ZN(n_0_0_239));
   NOR3_X1 i_0_0_980 (.A1(RST), .A2(n_0_0_283), .A3(n_0_0_255), .ZN(n_0_0_249));
   NOR2_X1 i_0_0_981 (.A1(n_0_0_283), .A2(n_0_0_255), .ZN(n_0_0_250));
   NAND2_X1 i_0_0_982 (.A1(next[1]), .A2(n_0_0_281), .ZN(n_0_0_251));
   NOR3_X1 i_0_0_983 (.A1(n_0_0_397), .A2(n_0_0_323), .A3(next[2]), .ZN(
      n_0_0_255));
   NOR2_X1 i_0_0_984 (.A1(n_0_0_323), .A2(next[2]), .ZN(n_0_0_281));
   NAND2_X1 i_0_0_985 (.A1(n_0_0_397), .A2(next[2]), .ZN(n_0_0_282));
   NOR2_X1 i_0_0_986 (.A1(n_0_0_398), .A2(next[1]), .ZN(n_0_0_283));
   NOR2_X1 i_0_0_987 (.A1(n_0_0_300), .A2(n_0_0_322), .ZN(n_0_0_299));
   NOR4_X1 i_0_0_988 (.A1(next[2]), .A2(next[1]), .A3(next[0]), .A4(Back), 
      .ZN(n_0_0_300));
   INV_X1 i_0_0_989 (.A(CLK), .ZN(n_0_136));
   INV_X1 i_0_0_990 (.A(counter[1]), .ZN(n_0_0_301));
   INV_X1 i_0_0_992 (.A(INT), .ZN(n_0_0_322));
   INV_X1 i_0_0_993 (.A(next[0]), .ZN(n_0_0_323));
   INV_X1 i_0_0_994 (.A(next[1]), .ZN(n_0_0_397));
   INV_X1 i_0_0_995 (.A(next[2]), .ZN(n_0_0_398));
   INV_X1 i_0_0_996 (.A(n_0_0_422), .ZN(n_0_0_399));
   INV_X1 i_0_0_997 (.A(n_0_0_421), .ZN(n_0_0_456));
   INV_X1 i_0_0_998 (.A(n_0_0_475), .ZN(n_0_0_513));
   INV_X1 i_0_0_276 (.A(m_val[14]), .ZN(n_0_0_635));
   INV_X1 i_0_0_280 (.A(m_val[13]), .ZN(n_0_0_623));
   INV_X1 i_0_0_283 (.A(n_val[13]), .ZN(n_0_0_596));
   INV_X1 i_0_0_291 (.A(n_val[14]), .ZN(n_0_0_604));
   AOI211_X1 i_0_0_294 (.A(n_0_0_233), .B(n_val[15]), .C1(n_0_0_254), .C2(
      n_val[10]), .ZN(n_0_0_514));
   NOR2_X1 i_0_0_295 (.A1(n_val[12]), .A2(n_0_0_264), .ZN(n_0_0_515));
   NOR2_X1 i_0_0_306 (.A1(n_0_0_213), .A2(n_val[2]), .ZN(n_0_0_540));
   INV_X1 i_0_0_307 (.A(n_val[15]), .ZN(n_0_0_541));
   INV_X1 i_0_0_333 (.A(n_0_0_163), .ZN(n_0_0_542));
   NOR3_X1 i_0_0_334 (.A1(n_0_0_151), .A2(n_val[14]), .A3(n_0_0_574), .ZN(
      n_0_0_597));
   INV_X1 i_0_0_336 (.A(NEW_VECTOR_CNT[12]), .ZN(n_0_0_629));
   INV_X1 i_0_0_337 (.A(RST), .ZN(n_0_0_321));
   OAI21_X1 i_0_0_352 (.A(n_0_0_441), .B1(n_0_0_641), .B2(n_0_0_442), .ZN(
      n_0_252));
   AOI22_X1 i_0_0_355 (.A1(RAM_DATA_RD1[11]), .A2(n_0_0_446), .B1(
      Element_Result[11]), .B2(n_0_0_447), .ZN(n_0_0_441));
   INV_X1 i_0_0_356 (.A(n_0_0_450), .ZN(n_0_0_442));
   NAND2_X1 i_0_0_367 (.A1(n_0_0_489), .A2(n_0_0_488), .ZN(n_0_253));
   AOI22_X1 i_0_0_368 (.A1(RAM_DATA_RD1[12]), .A2(n_0_0_446), .B1(
      Element_Result[12]), .B2(n_0_0_447), .ZN(n_0_0_488));
   NOR3_X1 i_0_0_375 (.A1(n_0_0_255), .A2(RST), .A3(n_0_0_448), .ZN(n_0_0_447));
   NOR2_X1 i_0_0_385 (.A1(n_0_0_553), .A2(n_0_0_449), .ZN(n_0_0_446));
   NAND2_X1 i_0_0_386 (.A1(NEW_Element_Result[12]), .A2(n_0_0_450), .ZN(
      n_0_0_489));
   OAI21_X1 i_0_0_387 (.A(n_0_0_451), .B1(INT), .B2(n_0_0_493), .ZN(n_0_0_450));
   OAI21_X1 i_0_0_391 (.A(n_0_0_639), .B1(n_0_0_641), .B2(n_0_0_640), .ZN(
      n_0_284));
   AOI22_X1 i_0_0_431 (.A1(FINAL_RESULT[11]), .A2(n_0_0_552), .B1(
      RAM_DATA_WR[11]), .B2(n_0_0_545), .ZN(n_0_0_639));
   INV_X1 i_0_0_432 (.A(n_0_0_494), .ZN(n_0_0_640));
   INV_X1 i_0_0_433 (.A(NEW_Element_Result[11]), .ZN(n_0_0_641));
   NAND2_X1 i_0_0_434 (.A1(n_0_0_645), .A2(n_0_0_642), .ZN(n_0_285));
   AOI21_X1 i_0_0_435 (.A(n_0_0_643), .B1(FINAL_RESULT[12]), .B2(n_0_0_552), 
      .ZN(n_0_0_642));
   NOR3_X1 i_0_0_436 (.A1(n_0_0_553), .A2(counter[0]), .A3(n_0_0_301), .ZN(
      n_0_0_552));
   INV_X1 i_0_0_465 (.A(n_0_0_644), .ZN(n_0_0_643));
   NAND2_X1 i_0_0_466 (.A1(n_0_0_545), .A2(RAM_DATA_WR[12]), .ZN(n_0_0_644));
   NOR2_X1 i_0_0_467 (.A1(n_0_0_546), .A2(RST), .ZN(n_0_0_545));
   NAND2_X1 i_0_0_468 (.A1(NEW_Element_Result[12]), .A2(n_0_0_494), .ZN(
      n_0_0_645));
   AOI21_X1 i_0_0_469 (.A(RST), .B1(n_0_0_608), .B2(n_0_0_251), .ZN(n_0_0_494));
   add_sub_cla__0_1293 ELEMENT_adder (.sub(), .in1(Element_Result), .in2(
      Multiplication_Result), .cin(), .out(NEW_Element_Result), .cout(), 
      .invalid());
endmodule
