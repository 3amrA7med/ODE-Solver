/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 21:04:59 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2522491783 */

module carry_lookahead_adder_4bit__4_800(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_9;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_14;
   wire n_0_15;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_4;
   wire n_0_5;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_16;

   XNOR2_X1 i_0_1 (.A(cin), .B(n_0_7), .ZN(sum[0]));
   XNOR2_X1 i_0_0 (.A(n_0_6), .B(n_0_0), .ZN(sum[1]));
   XNOR2_X1 i_0_2 (.A(in1[1]), .B(in0[1]), .ZN(n_0_0));
   XOR2_X1 i_0_3 (.A(n_0_9), .B(n_0_3), .Z(sum[2]));
   XNOR2_X1 i_0_4 (.A(n_0_13), .B(n_0_1), .ZN(sum[3]));
   NAND2_X1 i_0_5 (.A1(n_0_11), .A2(n_0_5), .ZN(n_0_9));
   INV_X1 i_0_6 (.A(n_0_2), .ZN(n_0_1));
   OAI21_X1 i_0_7 (.A(n_0_5), .B1(n_0_3), .B2(n_0_12), .ZN(n_0_2));
   OAI21_X1 i_0_8 (.A(n_0_17), .B1(in1[1]), .B2(in0[1]), .ZN(n_0_3));
   NOR2_X1 i_0_9 (.A1(n_0_18), .A2(n_0_19), .ZN(n_0_6));
   XNOR2_X1 i_0_13 (.A(in1[0]), .B(in0[0]), .ZN(n_0_7));
   AOI21_X1 i_0_10 (.A(n_0_16), .B1(n_0_10), .B2(n_0_8), .ZN(cout));
   AOI21_X1 i_0_11 (.A(n_0_4), .B1(n_0_14), .B2(n_0_17), .ZN(n_0_8));
   NOR2_X1 i_0_12 (.A1(n_0_12), .A2(n_0_15), .ZN(n_0_14));
   NOR2_X1 i_0_14 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_15));
   OAI21_X1 i_0_15 (.A(n_0_20), .B1(n_0_19), .B2(n_0_18), .ZN(n_0_17));
   AOI21_X1 i_0_16 (.A(cin), .B1(in1[0]), .B2(in0[0]), .ZN(n_0_18));
   NOR2_X1 i_0_17 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_19));
   NAND2_X1 i_0_18 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_20));
   INV_X1 i_0_19 (.A(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_20 (.A1(in0[2]), .A2(in1[2]), .ZN(n_0_5));
   NAND2_X1 i_0_21 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_12), .ZN(n_0_11));
   NOR2_X1 i_0_23 (.A1(in0[2]), .A2(in1[2]), .ZN(n_0_12));
   AOI21_X1 i_0_24 (.A(n_0_16), .B1(in1[3]), .B2(in0[3]), .ZN(n_0_13));
   NOR2_X1 i_0_25 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_16));
endmodule

module carry_lookahead_adder_4bit__4_791(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_10;
   wire n_0_11;
   wire n_0_7;
   wire n_0_1;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_8;
   wire n_0_9;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;

   XNOR2_X1 i_0_1 (.A(cin), .B(n_0_7), .ZN(sum[0]));
   XNOR2_X1 i_0_0 (.A(n_0_10), .B(n_0_1), .ZN(sum[3]));
   NOR2_X1 i_0_2 (.A1(n_0_14), .A2(n_0_11), .ZN(n_0_10));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(n_0_11));
   NAND2_X1 i_0_8 (.A1(n_0_8), .A2(n_0_4), .ZN(n_0_7));
   NAND2_X1 i_0_4 (.A1(n_0_12), .A2(n_0_13), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_0));
   NAND2_X1 i_0_6 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_2));
   NAND2_X1 i_0_7 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_3));
   NAND2_X1 i_0_9 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_4), .ZN(n_0_5));
   NOR2_X1 i_0_11 (.A1(n_0_5), .A2(cin), .ZN(n_0_6));
   OR2_X1 i_0_12 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_8));
   OAI21_X1 i_0_13 (.A(n_0_8), .B1(in1[1]), .B2(in0[1]), .ZN(n_0_9));
   OAI211_X1 i_0_14 (.A(n_0_2), .B(n_0_3), .C1(n_0_6), .C2(n_0_9), .ZN(n_0_12));
   OR2_X1 i_0_15 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_13));
   NOR2_X1 i_0_16 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_14));
   INV_X1 i_0_17 (.A(n_0_14), .ZN(n_0_15));
   NAND3_X1 i_0_18 (.A1(n_0_12), .A2(n_0_13), .A3(n_0_15), .ZN(n_0_16));
   NAND2_X1 i_0_19 (.A1(n_0_16), .A2(n_0_0), .ZN(cout));
   XNOR2_X1 i_0_20 (.A(n_0_18), .B(n_0_17), .ZN(sum[1]));
   XOR2_X1 i_0_21 (.A(in1[1]), .B(in0[1]), .Z(n_0_17));
   OAI21_X1 i_0_22 (.A(n_0_8), .B1(cin), .B2(n_0_5), .ZN(n_0_18));
   XNOR2_X1 i_0_23 (.A(n_0_20), .B(n_0_19), .ZN(sum[2]));
   OAI21_X1 i_0_24 (.A(n_0_3), .B1(n_0_6), .B2(n_0_9), .ZN(n_0_19));
   NAND2_X1 i_0_25 (.A1(n_0_13), .A2(n_0_2), .ZN(n_0_20));
endmodule

module carry_lookahead_adder_4bit__4_782(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_3;
   wire n_0_9;
   wire n_0_5;
   wire n_0_14;
   wire n_0_1;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_0;
   wire n_0_2;
   wire n_0_4;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_19;
   wire n_0_20;

   XOR2_X1 i_0_0 (.A(n_0_9), .B(n_0_3), .Z(sum[2]));
   XNOR2_X1 i_0_1 (.A(n_0_13), .B(n_0_1), .ZN(sum[3]));
   INV_X1 i_0_2 (.A(n_0_14), .ZN(n_0_3));
   NAND2_X1 i_0_3 (.A1(n_0_2), .A2(n_0_5), .ZN(n_0_9));
   NAND2_X1 i_0_4 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_5));
   NAND2_X1 i_0_5 (.A1(n_0_17), .A2(n_0_0), .ZN(n_0_14));
   NAND2_X1 i_0_6 (.A1(n_0_16), .A2(n_0_2), .ZN(n_0_1));
   NAND2_X1 i_0_7 (.A1(n_0_15), .A2(n_0_19), .ZN(cout));
   NAND3_X1 i_0_8 (.A1(n_0_16), .A2(n_0_4), .A3(n_0_2), .ZN(n_0_15));
   NAND3_X1 i_0_9 (.A1(n_0_17), .A2(n_0_5), .A3(n_0_0), .ZN(n_0_16));
   OAI211_X1 i_0_10 (.A(n_0_8), .B(n_0_18), .C1(cin), .C2(n_0_12), .ZN(n_0_17));
   OR2_X1 i_0_11 (.A1(in0[1]), .A2(in1[1]), .ZN(n_0_18));
   NAND2_X1 i_0_12 (.A1(in0[1]), .A2(in1[1]), .ZN(n_0_0));
   OR2_X1 i_0_13 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_2));
   INV_X1 i_0_14 (.A(n_0_20), .ZN(n_0_4));
   XNOR2_X1 i_0_15 (.A(cin), .B(n_0_6), .ZN(sum[0]));
   NAND2_X1 i_0_16 (.A1(n_0_8), .A2(n_0_7), .ZN(n_0_6));
   NAND2_X1 i_0_17 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_7));
   OR2_X1 i_0_18 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_8));
   XNOR2_X1 i_0_19 (.A(n_0_11), .B(n_0_10), .ZN(sum[1]));
   XOR2_X1 i_0_20 (.A(in1[1]), .B(in0[1]), .Z(n_0_10));
   OAI21_X1 i_0_21 (.A(n_0_8), .B1(n_0_12), .B2(cin), .ZN(n_0_11));
   INV_X1 i_0_22 (.A(n_0_7), .ZN(n_0_12));
   AOI21_X1 i_0_23 (.A(n_0_20), .B1(in1[3]), .B2(in0[3]), .ZN(n_0_13));
   NAND2_X1 i_0_24 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_19));
   NOR2_X1 i_0_25 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_20));
endmodule

module carry_lookahead_adder_4bit__4_773(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;

   AOI21_X1 i_0_0 (.A(n_0_15), .B1(n_0_13), .B2(n_0_14), .ZN(cout));
   XNOR2_X1 i_0_1 (.A(cin), .B(n_0_0), .ZN(sum[0]));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_1));
   OR2_X1 i_0_4 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_2));
   XNOR2_X1 i_0_5 (.A(n_0_4), .B(n_0_3), .ZN(sum[1]));
   XOR2_X1 i_0_6 (.A(in1[1]), .B(in0[1]), .Z(n_0_3));
   OAI21_X1 i_0_7 (.A(n_0_2), .B1(n_0_5), .B2(cin), .ZN(n_0_4));
   INV_X1 i_0_8 (.A(n_0_1), .ZN(n_0_5));
   XNOR2_X1 i_0_9 (.A(n_0_7), .B(n_0_6), .ZN(sum[2]));
   NAND2_X1 i_0_10 (.A1(n_0_11), .A2(n_0_10), .ZN(n_0_6));
   AOI21_X1 i_0_11 (.A(n_0_9), .B1(n_0_4), .B2(n_0_8), .ZN(n_0_7));
   NAND2_X1 i_0_12 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_8));
   NOR2_X1 i_0_13 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_9));
   NAND2_X1 i_0_14 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_10));
   OR2_X1 i_0_15 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_11));
   XNOR2_X1 i_0_16 (.A(n_0_13), .B(n_0_12), .ZN(sum[3]));
   AOI21_X1 i_0_17 (.A(n_0_15), .B1(in1[3]), .B2(in0[3]), .ZN(n_0_12));
   OAI21_X1 i_0_18 (.A(n_0_11), .B1(n_0_16), .B2(n_0_7), .ZN(n_0_13));
   NAND2_X1 i_0_19 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_14));
   NOR2_X1 i_0_20 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_15));
   INV_X1 i_0_21 (.A(n_0_10), .ZN(n_0_16));
endmodule

module carry_lookahead_adder_4bit__4_764(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_7;
   wire n_0_8;
   wire n_0_2;
   wire n_0_5;
   wire n_0_10;
   wire n_0_3;
   wire n_0_4;
   wire n_0_6;
   wire n_0_9;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;

   MUX2_X1 i_0_0 (.A(n_0_18), .B(n_0_24), .S(n_0_2), .Z(v));
   XNOR2_X1 i_0_1 (.A(in1[0]), .B(n_0_0), .ZN(sum[0]));
   XNOR2_X1 i_0_2 (.A(in0[0]), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_3 (.A(n_0_8), .B(n_0_1), .ZN(sum[2]));
   OAI21_X1 i_0_4 (.A(n_0_7), .B1(n_0_9), .B2(n_0_4), .ZN(n_0_1));
   NAND2_X1 i_0_5 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_7));
   NAND2_X1 i_0_6 (.A1(n_0_15), .A2(n_0_14), .ZN(n_0_8));
   INV_X1 i_0_7 (.A(n_0_10), .ZN(n_0_2));
   NAND2_X1 i_0_8 (.A1(n_0_5), .A2(n_0_23), .ZN(sum[3]));
   NAND2_X1 i_0_9 (.A1(n_0_10), .A2(n_0_3), .ZN(n_0_5));
   NAND2_X1 i_0_10 (.A1(n_0_17), .A2(n_0_22), .ZN(n_0_10));
   NAND2_X1 i_0_11 (.A1(n_0_20), .A2(n_0_19), .ZN(n_0_3));
   XOR2_X1 i_0_12 (.A(n_0_9), .B(n_0_4), .Z(sum[1]));
   INV_X1 i_0_13 (.A(n_0_6), .ZN(n_0_4));
   XOR2_X1 i_0_14 (.A(in0[1]), .B(in1[1]), .Z(n_0_6));
   NAND2_X1 i_0_15 (.A1(n_0_12), .A2(n_0_11), .ZN(n_0_9));
   OR2_X1 i_0_16 (.A1(cin), .A2(in0[0]), .ZN(n_0_11));
   INV_X1 i_0_17 (.A(n_0_13), .ZN(n_0_12));
   AOI21_X1 i_0_18 (.A(in1[0]), .B1(cin), .B2(in0[0]), .ZN(n_0_13));
   NAND2_X1 i_0_19 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_14));
   OR2_X1 i_0_20 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_15));
   AND2_X1 i_0_21 (.A1(n_0_15), .A2(n_0_14), .ZN(n_0_16));
   NAND4_X1 i_0_22 (.A1(n_0_16), .A2(n_0_6), .A3(n_0_12), .A4(n_0_11), .ZN(
      n_0_17));
   NOR2_X1 i_0_23 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_18));
   INV_X1 i_0_24 (.A(n_0_18), .ZN(n_0_19));
   NAND2_X1 i_0_25 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_20));
   NAND3_X1 i_0_26 (.A1(n_0_15), .A2(in0[1]), .A3(in1[1]), .ZN(n_0_21));
   AND2_X1 i_0_27 (.A1(n_0_21), .A2(n_0_14), .ZN(n_0_22));
   NAND4_X1 i_0_28 (.A1(n_0_17), .A2(n_0_22), .A3(n_0_19), .A4(n_0_20), .ZN(
      n_0_23));
   INV_X1 i_0_29 (.A(n_0_20), .ZN(n_0_24));
endmodule

module carry_lookahead_adder_20bit__4_801(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [19:0]in0;
   input [19:0]in1;
   input cin;
   output [19:0]sum;
   output cout;
   output v;

   wire c1;
   wire c2;
   wire c3;
   wire c4;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_0;

   carry_lookahead_adder_4bit__4_800 cla0 (.in0({in0[3], in0[2], in0[1], in0[0]}), 
      .in1({n_18, n_17, n_16, n_19}), .cin(sub), .sum({sum[3], sum[2], sum[1], 
      sum[0]}), .cout(c1), .v());
   carry_lookahead_adder_4bit__4_791 cla1 (.in0({in0[7], in0[6], in0[5], in0[4]}), 
      .in1({n_15, n_14, n_13, n_12}), .cin(c1), .sum({sum[7], sum[6], sum[5], 
      sum[4]}), .cout(c2), .v());
   carry_lookahead_adder_4bit__4_782 cla2 (.in0({in0[11], in0[10], in0[9], 
      in0[8]}), .in1({n_11, n_10, n_9, n_8}), .cin(c2), .sum({sum[11], sum[10], 
      sum[9], sum[8]}), .cout(c3), .v());
   carry_lookahead_adder_4bit__4_773 cla3 (.in0({in0[15], in0[14], in0[13], 
      in0[12]}), .in1({n_7, n_6, n_5, n_4}), .cin(c3), .sum({sum[15], sum[14], 
      sum[13], sum[12]}), .cout(c4), .v());
   carry_lookahead_adder_4bit__4_764 cla4 (.in0({in0[19], in0[18], in0[17], 
      in0[16]}), .in1({n_3, n_2, n_1, n_0}), .cin(c4), .sum({sum[19], sum[18], 
      sum[17], sum[16]}), .cout(), .v(v));
   XOR2_X1 i_0_0 (.A(in1[16]), .B(sub), .Z(n_0));
   XOR2_X1 i_0_1 (.A(sub), .B(in1[17]), .Z(n_1));
   XOR2_X1 i_0_2 (.A(sub), .B(in1[18]), .Z(n_2));
   XOR2_X1 i_0_3 (.A(sub), .B(in1[19]), .Z(n_3));
   XOR2_X1 i_0_4 (.A(in1[12]), .B(sub), .Z(n_4));
   XOR2_X1 i_0_5 (.A(sub), .B(in1[13]), .Z(n_5));
   XOR2_X1 i_0_6 (.A(sub), .B(in1[14]), .Z(n_6));
   XOR2_X1 i_0_7 (.A(sub), .B(in1[15]), .Z(n_7));
   XOR2_X1 i_0_8 (.A(in1[8]), .B(sub), .Z(n_8));
   XOR2_X1 i_0_9 (.A(sub), .B(in1[9]), .Z(n_9));
   XOR2_X1 i_0_10 (.A(sub), .B(in1[10]), .Z(n_10));
   XOR2_X1 i_0_11 (.A(sub), .B(in1[11]), .Z(n_11));
   XOR2_X1 i_0_12 (.A(in1[4]), .B(sub), .Z(n_12));
   XOR2_X1 i_0_13 (.A(sub), .B(in1[5]), .Z(n_13));
   XOR2_X1 i_0_14 (.A(sub), .B(in1[6]), .Z(n_14));
   XOR2_X1 i_0_15 (.A(sub), .B(in1[7]), .Z(n_15));
   XNOR2_X1 i_0_18 (.A(in1[1]), .B(n_0_2), .ZN(n_16));
   XNOR2_X1 i_0_19 (.A(in1[2]), .B(n_0_2), .ZN(n_17));
   NAND2_X1 i_0_16 (.A1(n_0_3), .A2(n_0_1), .ZN(n_18));
   NAND2_X1 i_0_17 (.A1(in1[3]), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_20 (.A(sub), .ZN(n_0_2));
   NAND2_X1 i_0_21 (.A1(n_0_0), .A2(sub), .ZN(n_0_3));
   INV_X1 i_0_22 (.A(in1[3]), .ZN(n_0_0));
   XOR2_X1 i_0_23 (.A(in1[0]), .B(sub), .Z(n_19));
endmodule

module add_sub_cla__4_802(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   wire v;
   wire [19:0]tempOut;
   wire n_0_7;
   wire n_0_8;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_9;
   wire n_1_0;
   wire [19:0]tempIn11;
   wire n_1_5;
   wire n_1_12;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;
   wire n_1_28;
   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_52;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire [19:0]tempIn22;
   wire n_1_87;
   wire n_1_88;
   wire n_1_89;
   wire n_1_90;
   wire n_1_91;
   wire n_1_92;
   wire n_1_93;
   wire n_1_94;
   wire n_1_95;
   wire n_1_96;
   wire n_1_97;
   wire n_1_98;
   wire n_1_99;
   wire n_1_102;
   wire n_1_105;
   wire n_1_106;
   wire n_1_107;
   wire n_1_108;
   wire n_1_109;
   wire n_1_112;
   wire n_1_113;
   wire n_1_114;
   wire n_1_123;
   wire n_1_124;
   wire n_1_148;
   wire n_1_151;
   wire n_1_156;
   wire n_1_157;
   wire n_1_158;
   wire n_1_159;
   wire n_1_15;
   wire n_1_6;
   wire n_1_72;
   wire n_1_73;
   wire n_1_13;
   wire n_1_74;
   wire n_1_75;
   wire n_1_138;
   wire n_1_139;
   wire n_1_140;
   wire n_1_141;
   wire n_1_161;
   wire n_1_162;
   wire n_1_163;
   wire n_1_116;
   wire n_1_167;
   wire n_1_168;
   wire n_1_170;
   wire n_1_171;
   wire n_1_172;
   wire n_1_173;
   wire n_1_174;
   wire n_1_175;
   wire n_1_176;
   wire n_1_177;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_14;
   wire n_1_16;
   wire n_1_17;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_40;
   wire n_1_41;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;
   wire n_1_60;
   wire n_1_61;
   wire n_1_62;
   wire n_1_63;
   wire n_1_64;
   wire n_1_65;
   wire n_1_66;
   wire n_1_67;
   wire n_1_68;
   wire n_1_69;
   wire n_1_70;
   wire n_1_71;
   wire n_1_76;
   wire n_1_77;
   wire n_1_78;
   wire n_1_79;
   wire n_1_80;
   wire n_1_81;
   wire n_1_82;
   wire n_1_83;
   wire n_1_84;
   wire n_1_85;
   wire n_1_86;
   wire n_1_100;
   wire n_1_101;
   wire n_1_103;
   wire n_1_104;
   wire n_1_110;
   wire n_1_111;
   wire n_1_115;
   wire n_1_117;
   wire n_1_118;
   wire n_1_119;
   wire n_1_120;
   wire n_1_121;
   wire n_1_122;
   wire n_1_125;
   wire n_1_126;
   wire n_1_127;
   wire n_1_128;
   wire n_1_129;
   wire n_1_130;
   wire n_1_131;
   wire n_1_132;
   wire n_1_133;
   wire n_1_134;
   wire n_1_135;
   wire n_1_136;
   wire n_1_137;
   wire n_1_142;
   wire n_1_143;
   wire n_1_144;
   wire n_1_145;
   wire n_1_146;
   wire n_1_147;
   wire n_1_149;
   wire n_1_150;
   wire n_1_152;
   wire n_1_153;
   wire n_1_154;
   wire n_1_155;
   wire n_1_160;
   wire n_1_164;
   wire n_1_165;
   wire n_1_166;
   wire n_1_169;
   wire n_1_178;
   wire n_1_179;
   wire n_1_180;
   wire n_1_181;
   wire n_1_182;
   wire n_1_183;
   wire n_1_184;
   wire n_1_185;
   wire n_1_186;
   wire n_1_187;
   wire n_1_188;
   wire n_1_189;
   wire n_1_190;
   wire n_1_191;

   carry_lookahead_adder_20bit__4_801 cs0 (.sub(sub), .in0({in1[12], 
      tempIn11[18], tempIn11[17], tempIn11[16], tempIn11[15], tempIn11[14], 
      tempIn11[13], tempIn11[12], tempIn11[11], tempIn11[10], tempIn11[9], 
      tempIn11[8], tempIn11[7], tempIn11[6], tempIn11[5], tempIn11[4], 
      tempIn11[3], tempIn11[2], tempIn11[1], tempIn11[0]}), .in1({in2[12], 
      tempIn22[18], tempIn22[17], tempIn22[16], tempIn22[15], tempIn22[14], 
      tempIn22[13], tempIn22[12], tempIn22[11], tempIn22[10], tempIn22[9], 
      tempIn22[8], tempIn22[7], tempIn22[6], tempIn22[5], tempIn22[4], 
      tempIn22[3], tempIn22[2], tempIn22[1], tempIn22[0]}), .cin(), .sum({
      tempOut[19], tempOut[18], tempOut[17], tempOut[16], tempOut[15], 
      tempOut[14], tempOut[13], out[12], out[11], out[10], out[9], out[8], 
      out[7], out[6], out[5], out[4], out[3], out[2], out[1], out[0]}), .cout(), 
      .v(v));
   INV_X1 i_0_0 (.A(tempOut[18]), .ZN(n_0_7));
   INV_X1 i_0_1 (.A(tempOut[19]), .ZN(n_0_8));
   NAND2_X1 i_0_2 (.A1(n_0_0), .A2(n_0_3), .ZN(invalid));
   NAND2_X1 i_0_3 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND3_X1 i_0_4 (.A1(n_0_4), .A2(n_0_7), .A3(n_0_8), .ZN(n_0_1));
   NAND4_X1 i_0_5 (.A1(tempOut[18]), .A2(tempOut[19]), .A3(tempOut[16]), 
      .A4(n_0_9), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(v), .ZN(n_0_3));
   NOR3_X1 i_0_7 (.A1(tempOut[16]), .A2(n_0_5), .A3(tempOut[17]), .ZN(n_0_4));
   OR4_X1 i_0_8 (.A1(tempOut[15]), .A2(tempOut[13]), .A3(out[12]), .A4(
      tempOut[14]), .ZN(n_0_5));
   AND4_X1 i_0_9 (.A1(tempOut[15]), .A2(tempOut[13]), .A3(out[12]), .A4(
      tempOut[14]), .ZN(n_0_6));
   AND2_X1 i_0_10 (.A1(n_0_6), .A2(tempOut[17]), .ZN(n_0_9));
   OAI21_X1 i_1_0 (.A(n_1_0), .B1(n_1_19), .B2(n_1_2), .ZN(out[13]));
   NAND2_X1 i_1_1 (.A1(in1[13]), .A2(n_1_2), .ZN(n_1_0));
   NAND2_X1 i_1_4 (.A1(n_1_41), .A2(n_1_20), .ZN(out[15]));
   OAI21_X1 i_1_2 (.A(n_1_5), .B1(n_1_63), .B2(n_1_6), .ZN(tempIn11[3]));
   AOI22_X1 i_1_3 (.A1(in1[3]), .A2(n_1_49), .B1(n_1_79), .B2(n_1_120), .ZN(
      n_1_5));
   OAI21_X1 i_1_5 (.A(n_1_12), .B1(n_1_80), .B2(n_1_15), .ZN(tempIn11[6]));
   AOI22_X1 i_1_6 (.A1(in1[6]), .A2(n_1_49), .B1(n_1_77), .B2(n_1_13), .ZN(
      n_1_12));
   AOI222_X1 i_1_7 (.A1(n_1_156), .A2(n_1_49), .B1(n_1_79), .B2(n_1_21), 
      .C1(n_1_77), .C2(n_1_126), .ZN(tempIn11[8]));
   AOI222_X1 i_1_8 (.A1(n_1_157), .A2(n_1_49), .B1(n_1_79), .B2(n_1_24), 
      .C1(n_1_77), .C2(n_1_21), .ZN(tempIn11[9]));
   AOI221_X1 i_1_9 (.A(n_1_22), .B1(in1[6]), .B2(n_1_122), .C1(in1[8]), .C2(
      n_1_84), .ZN(n_1_21));
   INV_X1 i_1_10 (.A(n_1_23), .ZN(n_1_22));
   AOI22_X1 i_1_11 (.A1(in1[4]), .A2(n_1_134), .B1(in1[2]), .B2(n_1_131), 
      .ZN(n_1_23));
   AOI222_X1 i_1_12 (.A1(n_1_158), .A2(n_1_49), .B1(n_1_79), .B2(n_1_27), 
      .C1(n_1_77), .C2(n_1_24), .ZN(tempIn11[10]));
   AOI221_X1 i_1_13 (.A(n_1_25), .B1(in1[7]), .B2(n_1_122), .C1(in1[9]), 
      .C2(n_1_84), .ZN(n_1_24));
   INV_X1 i_1_14 (.A(n_1_26), .ZN(n_1_25));
   AOI22_X1 i_1_15 (.A1(in1[5]), .A2(n_1_134), .B1(in1[3]), .B2(n_1_131), 
      .ZN(n_1_26));
   AOI222_X1 i_1_16 (.A1(n_1_159), .A2(n_1_49), .B1(n_1_77), .B2(n_1_27), 
      .C1(n_1_79), .C2(n_1_31), .ZN(tempIn11[11]));
   AOI221_X1 i_1_17 (.A(n_1_28), .B1(in1[8]), .B2(n_1_122), .C1(in1[4]), 
      .C2(n_1_131), .ZN(n_1_27));
   INV_X1 i_1_18 (.A(n_1_29), .ZN(n_1_28));
   AOI22_X1 i_1_19 (.A1(in1[10]), .A2(n_1_84), .B1(in1[6]), .B2(n_1_134), 
      .ZN(n_1_29));
   OAI21_X1 i_1_20 (.A(n_1_30), .B1(n_1_63), .B2(n_1_31), .ZN(tempIn11[12]));
   AOI21_X1 i_1_21 (.A(n_1_43), .B1(n_1_79), .B2(n_1_35), .ZN(n_1_30));
   AOI221_X1 i_1_22 (.A(n_1_32), .B1(in1[9]), .B2(n_1_122), .C1(in1[11]), 
      .C2(n_1_84), .ZN(n_1_31));
   INV_X1 i_1_23 (.A(n_1_33), .ZN(n_1_32));
   AOI22_X1 i_1_24 (.A1(in1[5]), .A2(n_1_131), .B1(in1[7]), .B2(n_1_134), 
      .ZN(n_1_33));
   INV_X1 i_1_25 (.A(n_1_34), .ZN(tempIn11[13]));
   AOI221_X1 i_1_26 (.A(n_1_43), .B1(n_1_79), .B2(n_1_38), .C1(n_1_77), .C2(
      n_1_35), .ZN(n_1_34));
   AOI221_X1 i_1_27 (.A(n_1_36), .B1(n_1_85), .B2(n_1_48), .C1(n_1_156), 
      .C2(n_1_134), .ZN(n_1_35));
   OAI33_X1 i_1_28 (.A1(n_1_100), .A2(n_1_85), .A3(in1[6]), .B1(n_1_101), 
      .B2(n_1_85), .B3(in1[10]), .ZN(n_1_36));
   INV_X1 i_1_29 (.A(n_1_37), .ZN(tempIn11[14]));
   AOI221_X1 i_1_30 (.A(n_1_43), .B1(n_1_77), .B2(n_1_38), .C1(n_1_79), .C2(
      n_1_44), .ZN(n_1_37));
   AOI221_X1 i_1_31 (.A(n_1_39), .B1(n_1_85), .B2(n_1_48), .C1(n_1_133), 
      .C2(n_1_131), .ZN(n_1_38));
   OAI33_X1 i_1_32 (.A1(n_1_101), .A2(n_1_85), .A3(in1[11]), .B1(n_1_100), 
      .B2(n_1_86), .B3(in1[9]), .ZN(n_1_39));
   INV_X1 i_1_33 (.A(n_1_42), .ZN(tempIn11[15]));
   AOI221_X1 i_1_34 (.A(n_1_43), .B1(n_1_79), .B2(n_1_47), .C1(n_1_77), .C2(
      n_1_44), .ZN(n_1_42));
   AND2_X1 i_1_35 (.A1(in1[12]), .A2(n_1_49), .ZN(n_1_43));
   AOI221_X1 i_1_36 (.A(n_1_48), .B1(n_1_158), .B2(n_1_134), .C1(n_1_156), 
      .C2(n_1_131), .ZN(n_1_44));
   AOI221_X1 i_1_37 (.A(n_1_45), .B1(n_1_158), .B2(n_1_52), .C1(n_1_77), 
      .C2(n_1_46), .ZN(tempIn11[16]));
   NOR3_X1 i_1_38 (.A1(in1[12]), .A2(n_1_77), .A3(n_1_52), .ZN(n_1_45));
   INV_X1 i_1_39 (.A(n_1_47), .ZN(n_1_46));
   AOI221_X1 i_1_40 (.A(n_1_48), .B1(n_1_157), .B2(n_1_131), .C1(n_1_159), 
      .C2(n_1_134), .ZN(n_1_47));
   NOR2_X1 i_1_41 (.A1(in1[12]), .A2(n_1_101), .ZN(n_1_48));
   AOI221_X1 i_1_42 (.A(n_1_56), .B1(n_1_159), .B2(n_1_52), .C1(n_1_158), 
      .C2(n_1_58), .ZN(tempIn11[17]));
   NOR3_X1 i_1_43 (.A1(n_1_100), .A2(n_1_85), .A3(n_1_80), .ZN(n_1_52));
   AOI21_X1 i_1_44 (.A(in1[12]), .B1(n_1_3), .B2(n_1_131), .ZN(n_1_56));
   OAI21_X1 i_1_45 (.A(n_1_57), .B1(n_1_159), .B2(n_1_59), .ZN(tempIn11[18]));
   NAND2_X1 i_1_46 (.A1(in1[12]), .A2(n_1_59), .ZN(n_1_57));
   INV_X1 i_1_47 (.A(n_1_59), .ZN(n_1_58));
   NAND3_X1 i_1_48 (.A1(n_1_3), .A2(n_1_131), .A3(n_1_62), .ZN(n_1_59));
   AOI222_X1 i_1_49 (.A1(n_1_148), .A2(n_1_3), .B1(n_1_116), .B2(n_1_179), 
      .C1(n_1_169), .C2(n_1_87), .ZN(tempIn22[9]));
   AOI222_X1 i_1_50 (.A1(n_1_190), .A2(n_1_3), .B1(n_1_169), .B2(n_1_89), 
      .C1(n_1_116), .C2(n_1_87), .ZN(tempIn22[10]));
   AOI221_X1 i_1_51 (.A(n_1_88), .B1(in2[3]), .B2(n_1_70), .C1(in2[5]), .C2(
      n_1_186), .ZN(n_1_87));
   OAI22_X1 i_1_52 (.A1(n_1_148), .A2(n_1_146), .B1(n_1_184), .B2(n_1_145), 
      .ZN(n_1_88));
   AOI222_X1 i_1_53 (.A1(n_1_191), .A2(n_1_3), .B1(n_1_116), .B2(n_1_89), 
      .C1(n_1_169), .C2(n_1_92), .ZN(tempIn22[11]));
   AOI221_X1 i_1_54 (.A(n_1_90), .B1(in2[4]), .B2(n_1_70), .C1(in2[6]), .C2(
      n_1_186), .ZN(n_1_89));
   OAI22_X1 i_1_55 (.A1(n_1_190), .A2(n_1_146), .B1(n_1_185), .B2(n_1_145), 
      .ZN(n_1_90));
   OAI21_X1 i_1_56 (.A(n_1_91), .B1(n_1_160), .B2(n_1_92), .ZN(tempIn22[12]));
   AOI21_X1 i_1_57 (.A(n_1_106), .B1(n_1_169), .B2(n_1_95), .ZN(n_1_91));
   AOI221_X1 i_1_58 (.A(n_1_93), .B1(in2[5]), .B2(n_1_70), .C1(in2[7]), .C2(
      n_1_186), .ZN(n_1_92));
   OAI22_X1 i_1_59 (.A1(n_1_148), .A2(n_1_145), .B1(n_1_191), .B2(n_1_146), 
      .ZN(n_1_93));
   INV_X1 i_1_60 (.A(n_1_94), .ZN(tempIn22[13]));
   AOI221_X1 i_1_61 (.A(n_1_106), .B1(n_1_169), .B2(n_1_98), .C1(n_1_116), 
      .C2(n_1_95), .ZN(n_1_94));
   AOI221_X1 i_1_62 (.A(n_1_96), .B1(n_1_65), .B2(n_1_114), .C1(n_1_185), 
      .C2(n_1_186), .ZN(n_1_95));
   OAI33_X1 i_1_63 (.A1(n_1_65), .A2(n_1_149), .A3(in2[6]), .B1(n_1_65), 
      .B2(n_1_68), .B3(in2[10]), .ZN(n_1_96));
   INV_X1 i_1_64 (.A(n_1_97), .ZN(tempIn22[14]));
   AOI221_X1 i_1_65 (.A(n_1_106), .B1(n_1_116), .B2(n_1_98), .C1(n_1_169), 
      .C2(n_1_107), .ZN(n_1_97));
   AOI221_X1 i_1_66 (.A(n_1_99), .B1(n_1_184), .B2(n_1_70), .C1(n_1_65), 
      .C2(n_1_114), .ZN(n_1_98));
   OAI21_X1 i_1_67 (.A(n_1_102), .B1(in2[11]), .B2(n_1_145), .ZN(n_1_99));
   NAND2_X1 i_1_68 (.A1(n_1_148), .A2(n_1_186), .ZN(n_1_102));
   INV_X1 i_1_69 (.A(n_1_105), .ZN(tempIn22[15]));
   AOI221_X1 i_1_70 (.A(n_1_106), .B1(n_1_113), .B2(n_1_169), .C1(n_1_116), 
      .C2(n_1_107), .ZN(n_1_105));
   NOR2_X1 i_1_71 (.A1(n_1_151), .A2(n_1_2), .ZN(n_1_106));
   AOI221_X1 i_1_72 (.A(n_1_114), .B1(n_1_190), .B2(n_1_186), .C1(n_1_185), 
      .C2(n_1_70), .ZN(n_1_107));
   AOI221_X1 i_1_73 (.A(n_1_108), .B1(n_1_151), .B2(n_1_109), .C1(n_1_116), 
      .C2(n_1_112), .ZN(tempIn22[16]));
   NOR4_X1 i_1_74 (.A1(n_1_65), .A2(n_1_149), .A3(n_1_178), .A4(in2[10]), 
      .ZN(n_1_108));
   AOI21_X1 i_1_75 (.A(n_1_116), .B1(n_1_70), .B2(n_1_169), .ZN(n_1_109));
   INV_X1 i_1_76 (.A(n_1_113), .ZN(n_1_112));
   AOI221_X1 i_1_77 (.A(n_1_114), .B1(n_1_148), .B2(n_1_70), .C1(n_1_191), 
      .C2(n_1_186), .ZN(n_1_113));
   NOR2_X1 i_1_78 (.A1(in2[12]), .A2(n_1_68), .ZN(n_1_114));
   AOI21_X1 i_1_163 (.A(n_1_123), .B1(n_1_151), .B2(n_1_124), .ZN(tempIn22[18]));
   NOR2_X1 i_1_164 (.A1(in2[11]), .A2(n_1_124), .ZN(n_1_123));
   NAND2_X1 i_1_165 (.A1(n_1_189), .A2(n_1_62), .ZN(n_1_124));
   INV_X1 i_1_79 (.A(in2[9]), .ZN(n_1_148));
   INV_X1 i_1_80 (.A(in2[12]), .ZN(n_1_151));
   INV_X1 i_1_81 (.A(in1[8]), .ZN(n_1_156));
   INV_X1 i_1_82 (.A(in1[9]), .ZN(n_1_157));
   INV_X1 i_1_83 (.A(in1[10]), .ZN(n_1_158));
   INV_X1 i_1_84 (.A(in1[11]), .ZN(n_1_159));
   INV_X1 i_1_85 (.A(n_1_128), .ZN(n_1_15));
   INV_X1 i_1_86 (.A(n_1_81), .ZN(n_1_6));
   OAI211_X1 i_1_87 (.A(n_1_72), .B(n_1_78), .C1(n_1_111), .C2(n_1_50), .ZN(
      tempIn11[2]));
   NAND2_X1 i_1_88 (.A1(n_1_71), .A2(in1[1]), .ZN(n_1_72));
   OAI221_X1 i_1_89 (.A(n_1_73), .B1(n_1_132), .B2(n_1_50), .C1(n_1_117), 
      .C2(n_1_63), .ZN(tempIn11[5]));
   NAND2_X1 i_1_90 (.A1(n_1_13), .A2(n_1_79), .ZN(n_1_73));
   OAI211_X1 i_1_91 (.A(n_1_75), .B(n_1_74), .C1(n_1_83), .C2(n_1_132), .ZN(
      n_1_13));
   NAND2_X1 i_1_92 (.A1(n_1_122), .A2(in1[3]), .ZN(n_1_74));
   NAND2_X1 i_1_93 (.A1(n_1_134), .A2(in1[1]), .ZN(n_1_75));
   OAI21_X1 i_1_94 (.A(n_1_138), .B1(n_1_150), .B2(n_1_2), .ZN(tempIn22[1]));
   NAND3_X1 i_1_95 (.A1(n_1_140), .A2(n_1_116), .A3(in2[0]), .ZN(n_1_138));
   OAI221_X1 i_1_96 (.A(n_1_139), .B1(n_1_152), .B2(n_1_2), .C1(n_1_162), 
      .C2(n_1_178), .ZN(tempIn22[2]));
   NAND3_X1 i_1_97 (.A1(n_1_140), .A2(n_1_116), .A3(in2[1]), .ZN(n_1_139));
   INV_X1 i_1_98 (.A(n_1_146), .ZN(n_1_140));
   INV_X1 i_1_99 (.A(n_1_141), .ZN(tempIn22[3]));
   OAI221_X1 i_1_100 (.A(n_1_161), .B1(in2[3]), .B2(n_1_2), .C1(n_1_178), 
      .C2(n_1_144), .ZN(n_1_141));
   OAI211_X1 i_1_101 (.A(n_1_162), .B(n_1_116), .C1(n_1_152), .C2(n_1_146), 
      .ZN(n_1_161));
   NAND3_X1 i_1_102 (.A1(n_1_149), .A2(in2[0]), .A3(n_1_66), .ZN(n_1_162));
   OAI221_X1 i_1_103 (.A(n_1_163), .B1(n_1_182), .B2(n_1_2), .C1(n_1_178), 
      .C2(n_1_167), .ZN(tempIn22[5]));
   OAI21_X1 i_1_104 (.A(n_1_116), .B1(n_1_142), .B2(n_1_137), .ZN(n_1_163));
   INV_X1 i_1_105 (.A(n_1_160), .ZN(n_1_116));
   OAI211_X1 i_1_106 (.A(n_1_171), .B(n_1_170), .C1(n_1_160), .C2(n_1_167), 
      .ZN(tempIn22[6]));
   AOI21_X1 i_1_107 (.A(n_1_168), .B1(n_1_186), .B2(in2[1]), .ZN(n_1_167));
   OAI22_X1 i_1_108 (.A1(n_1_182), .A2(n_1_146), .B1(n_1_145), .B2(n_1_153), 
      .ZN(n_1_168));
   NAND2_X1 i_1_109 (.A1(n_1_3), .A2(in2[6]), .ZN(n_1_170));
   NAND2_X1 i_1_110 (.A1(n_1_174), .A2(n_1_169), .ZN(n_1_171));
   INV_X1 i_1_111 (.A(n_1_172), .ZN(tempIn22[7]));
   OAI211_X1 i_1_112 (.A(n_1_177), .B(n_1_173), .C1(n_1_174), .C2(n_1_160), 
      .ZN(n_1_172));
   NAND2_X1 i_1_113 (.A1(n_1_3), .A2(n_1_184), .ZN(n_1_173));
   OAI21_X1 i_1_114 (.A(n_1_175), .B1(n_1_152), .B2(n_1_143), .ZN(n_1_174));
   AOI21_X1 i_1_115 (.A(n_1_176), .B1(n_1_70), .B2(in2[0]), .ZN(n_1_175));
   OAI22_X1 i_1_116 (.A1(n_1_183), .A2(n_1_146), .B1(n_1_145), .B2(n_1_154), 
      .ZN(n_1_176));
   NAND3_X1 i_1_117 (.A1(n_1_165), .A2(n_1_164), .A3(n_1_169), .ZN(n_1_177));
   INV_X1 i_1_118 (.A(n_1_1), .ZN(out[14]));
   OAI22_X1 i_1_119 (.A1(in2[14]), .A2(n_1_2), .B1(in1[14]), .B2(n_1_3), 
      .ZN(n_1_1));
   INV_X1 i_1_120 (.A(n_1_3), .ZN(n_1_2));
   OAI21_X1 i_1_121 (.A(n_1_18), .B1(n_1_8), .B2(n_1_7), .ZN(n_1_3));
   INV_X1 i_1_122 (.A(n_1_7), .ZN(n_1_4));
   NOR2_X1 i_1_123 (.A1(n_1_41), .A2(in2[15]), .ZN(n_1_7));
   INV_X1 i_1_124 (.A(n_1_9), .ZN(n_1_8));
   OAI21_X1 i_1_125 (.A(n_1_17), .B1(n_1_14), .B2(n_1_11), .ZN(n_1_9));
   INV_X1 i_1_126 (.A(n_1_11), .ZN(n_1_10));
   NOR2_X1 i_1_127 (.A1(n_1_40), .A2(in2[14]), .ZN(n_1_11));
   INV_X1 i_1_128 (.A(n_1_16), .ZN(n_1_14));
   NAND2_X1 i_1_129 (.A1(in1[13]), .A2(n_1_19), .ZN(n_1_16));
   NAND2_X1 i_1_130 (.A1(n_1_40), .A2(in2[14]), .ZN(n_1_17));
   NAND2_X1 i_1_131 (.A1(n_1_41), .A2(in2[15]), .ZN(n_1_18));
   INV_X1 i_1_132 (.A(in2[13]), .ZN(n_1_19));
   INV_X1 i_1_133 (.A(in2[15]), .ZN(n_1_20));
   INV_X1 i_1_134 (.A(in1[14]), .ZN(n_1_40));
   INV_X1 i_1_135 (.A(in1[15]), .ZN(n_1_41));
   AND2_X1 i_1_136 (.A1(in1[0]), .A2(n_1_49), .ZN(tempIn11[0]));
   INV_X1 i_1_137 (.A(n_1_50), .ZN(n_1_49));
   AOI21_X1 i_1_138 (.A(n_1_55), .B1(n_1_18), .B2(n_1_51), .ZN(n_1_50));
   OAI21_X1 i_1_139 (.A(n_1_10), .B1(n_1_60), .B2(n_1_54), .ZN(n_1_51));
   INV_X1 i_1_140 (.A(n_1_54), .ZN(n_1_53));
   NOR2_X1 i_1_141 (.A1(in1[13]), .A2(n_1_61), .ZN(n_1_54));
   INV_X1 i_1_142 (.A(n_1_4), .ZN(n_1_55));
   INV_X1 i_1_143 (.A(n_1_17), .ZN(n_1_60));
   INV_X1 i_1_144 (.A(in2[13]), .ZN(n_1_61));
   NAND2_X1 i_1_145 (.A1(n_1_53), .A2(n_1_16), .ZN(n_1_62));
   NAND2_X1 i_1_146 (.A1(n_1_62), .A2(n_1_50), .ZN(n_1_63));
   NAND2_X1 i_1_147 (.A1(n_1_17), .A2(n_1_10), .ZN(n_1_64));
   XNOR2_X1 i_1_148 (.A(n_1_64), .B(n_1_54), .ZN(n_1_65));
   INV_X1 i_1_149 (.A(n_1_65), .ZN(n_1_66));
   NAND2_X1 i_1_150 (.A1(n_1_18), .A2(n_1_4), .ZN(n_1_67));
   XNOR2_X1 i_1_151 (.A(n_1_67), .B(n_1_51), .ZN(n_1_68));
   NAND2_X1 i_1_152 (.A1(n_1_66), .A2(n_1_68), .ZN(n_1_69));
   INV_X1 i_1_153 (.A(n_1_69), .ZN(n_1_70));
   NOR2_X1 i_1_154 (.A1(n_1_69), .A2(n_1_63), .ZN(n_1_71));
   AOI22_X1 i_1_155 (.A1(n_1_71), .A2(in1[0]), .B1(in1[1]), .B2(n_1_49), 
      .ZN(n_1_76));
   INV_X1 i_1_156 (.A(n_1_76), .ZN(tempIn11[1]));
   INV_X1 i_1_157 (.A(n_1_63), .ZN(n_1_77));
   NAND2_X1 i_1_158 (.A1(n_1_81), .A2(n_1_79), .ZN(n_1_78));
   INV_X1 i_1_159 (.A(n_1_80), .ZN(n_1_79));
   NAND2_X1 i_1_160 (.A1(n_1_104), .A2(n_1_50), .ZN(n_1_80));
   OAI22_X1 i_1_161 (.A1(n_1_111), .A2(n_1_83), .B1(n_1_110), .B2(n_1_82), 
      .ZN(n_1_81));
   NAND2_X1 i_1_162 (.A1(n_1_100), .A2(n_1_86), .ZN(n_1_82));
   INV_X1 i_1_166 (.A(n_1_84), .ZN(n_1_83));
   NOR2_X1 i_1_167 (.A1(n_1_101), .A2(n_1_86), .ZN(n_1_84));
   INV_X1 i_1_168 (.A(n_1_86), .ZN(n_1_85));
   XOR2_X1 i_1_169 (.A(n_1_64), .B(n_1_14), .Z(n_1_86));
   INV_X1 i_1_170 (.A(n_1_101), .ZN(n_1_100));
   AOI21_X1 i_1_171 (.A(n_1_103), .B1(n_1_8), .B2(n_1_67), .ZN(n_1_101));
   AND3_X1 i_1_172 (.A1(n_1_18), .A2(n_1_4), .A3(n_1_9), .ZN(n_1_103));
   INV_X1 i_1_173 (.A(n_1_62), .ZN(n_1_104));
   INV_X1 i_1_174 (.A(in1[0]), .ZN(n_1_110));
   INV_X1 i_1_175 (.A(in1[2]), .ZN(n_1_111));
   OAI21_X1 i_1_176 (.A(n_1_115), .B1(n_1_80), .B2(n_1_117), .ZN(tempIn11[4]));
   AOI22_X1 i_1_177 (.A1(n_1_77), .A2(n_1_120), .B1(in1[4]), .B2(n_1_49), 
      .ZN(n_1_115));
   AOI21_X1 i_1_178 (.A(n_1_118), .B1(in1[4]), .B2(n_1_84), .ZN(n_1_117));
   OAI22_X1 i_1_179 (.A1(n_1_110), .A2(n_1_119), .B1(n_1_82), .B2(n_1_111), 
      .ZN(n_1_118));
   NAND2_X1 i_1_180 (.A1(n_1_101), .A2(n_1_85), .ZN(n_1_119));
   INV_X1 i_1_181 (.A(n_1_121), .ZN(n_1_120));
   AOI22_X1 i_1_182 (.A1(in1[3]), .A2(n_1_84), .B1(n_1_122), .B2(in1[1]), 
      .ZN(n_1_121));
   INV_X1 i_1_183 (.A(n_1_82), .ZN(n_1_122));
   AOI21_X1 i_1_184 (.A(n_1_125), .B1(n_1_79), .B2(n_1_126), .ZN(tempIn11[7]));
   OAI22_X1 i_1_185 (.A1(n_1_63), .A2(n_1_128), .B1(in1[7]), .B2(n_1_50), 
      .ZN(n_1_125));
   AOI221_X1 i_1_186 (.A(n_1_127), .B1(in1[1]), .B2(n_1_131), .C1(n_1_134), 
      .C2(in1[3]), .ZN(n_1_126));
   OAI22_X1 i_1_187 (.A1(n_1_132), .A2(n_1_82), .B1(n_1_133), .B2(n_1_83), 
      .ZN(n_1_127));
   NAND2_X1 i_1_188 (.A1(n_1_130), .A2(n_1_129), .ZN(n_1_128));
   AOI222_X1 i_1_189 (.A1(in1[0]), .A2(n_1_131), .B1(n_1_134), .B2(in1[2]), 
      .C1(in1[6]), .C2(n_1_84), .ZN(n_1_129));
   NAND2_X1 i_1_190 (.A1(in1[4]), .A2(n_1_122), .ZN(n_1_130));
   AND2_X1 i_1_191 (.A1(n_1_101), .A2(n_1_86), .ZN(n_1_131));
   INV_X1 i_1_192 (.A(in1[5]), .ZN(n_1_132));
   INV_X1 i_1_193 (.A(in1[7]), .ZN(n_1_133));
   INV_X1 i_1_194 (.A(n_1_119), .ZN(n_1_134));
   AND2_X1 i_1_195 (.A1(n_1_3), .A2(in2[0]), .ZN(tempIn22[0]));
   OAI211_X1 i_1_196 (.A(n_1_135), .B(n_1_136), .C1(n_1_154), .C2(n_1_147), 
      .ZN(tempIn22[4]));
   NAND3_X1 i_1_197 (.A1(n_1_2), .A2(n_1_62), .A3(n_1_144), .ZN(n_1_135));
   OAI211_X1 i_1_198 (.A(n_1_2), .B(n_1_104), .C1(n_1_142), .C2(n_1_137), 
      .ZN(n_1_136));
   OAI22_X1 i_1_199 (.A1(n_1_152), .A2(n_1_145), .B1(n_1_154), .B2(n_1_146), 
      .ZN(n_1_137));
   AND3_X1 i_1_200 (.A1(n_1_68), .A2(n_1_65), .A3(in2[0]), .ZN(n_1_142));
   NAND2_X1 i_1_201 (.A1(n_1_68), .A2(n_1_65), .ZN(n_1_143));
   OAI22_X1 i_1_202 (.A1(n_1_150), .A2(n_1_145), .B1(n_1_153), .B2(n_1_146), 
      .ZN(n_1_144));
   NAND2_X1 i_1_203 (.A1(n_1_149), .A2(n_1_66), .ZN(n_1_145));
   NAND2_X1 i_1_204 (.A1(n_1_149), .A2(n_1_65), .ZN(n_1_146));
   INV_X1 i_1_205 (.A(n_1_3), .ZN(n_1_147));
   INV_X1 i_1_206 (.A(n_1_68), .ZN(n_1_149));
   INV_X1 i_1_207 (.A(in2[1]), .ZN(n_1_150));
   INV_X1 i_1_208 (.A(in2[2]), .ZN(n_1_152));
   INV_X1 i_1_209 (.A(in2[3]), .ZN(n_1_153));
   INV_X1 i_1_210 (.A(in2[4]), .ZN(n_1_154));
   AOI221_X1 i_1_211 (.A(n_1_155), .B1(n_1_179), .B2(n_1_169), .C1(n_1_185), 
      .C2(n_1_3), .ZN(tempIn22[8]));
   AND4_X1 i_1_212 (.A1(n_1_2), .A2(n_1_62), .A3(n_1_165), .A4(n_1_164), 
      .ZN(n_1_155));
   NAND2_X1 i_1_213 (.A1(n_1_2), .A2(n_1_62), .ZN(n_1_160));
   NAND2_X1 i_1_214 (.A1(in2[1]), .A2(n_1_70), .ZN(n_1_164));
   AOI21_X1 i_1_215 (.A(n_1_166), .B1(n_1_186), .B2(in2[3]), .ZN(n_1_165));
   OAI22_X1 i_1_216 (.A1(n_1_182), .A2(n_1_145), .B1(n_1_184), .B2(n_1_146), 
      .ZN(n_1_166));
   INV_X1 i_1_217 (.A(n_1_178), .ZN(n_1_169));
   NAND2_X1 i_1_218 (.A1(n_1_2), .A2(n_1_104), .ZN(n_1_178));
   NOR2_X1 i_1_219 (.A1(n_1_181), .A2(n_1_180), .ZN(n_1_179));
   OAI22_X1 i_1_220 (.A1(n_1_69), .A2(n_1_152), .B1(n_1_143), .B2(n_1_154), 
      .ZN(n_1_180));
   OAI22_X1 i_1_221 (.A1(n_1_183), .A2(n_1_145), .B1(n_1_185), .B2(n_1_146), 
      .ZN(n_1_181));
   INV_X1 i_1_222 (.A(in2[5]), .ZN(n_1_182));
   INV_X1 i_1_223 (.A(in2[6]), .ZN(n_1_183));
   INV_X1 i_1_224 (.A(in2[7]), .ZN(n_1_184));
   INV_X1 i_1_225 (.A(in2[8]), .ZN(n_1_185));
   INV_X1 i_1_226 (.A(n_1_143), .ZN(n_1_186));
   INV_X1 i_1_227 (.A(n_1_187), .ZN(tempIn22[17]));
   OAI21_X1 i_1_228 (.A(n_1_188), .B1(in2[12]), .B2(n_1_189), .ZN(n_1_187));
   OAI221_X1 i_1_229 (.A(n_1_189), .B1(n_1_190), .B2(n_1_104), .C1(n_1_191), 
      .C2(n_1_62), .ZN(n_1_188));
   AND2_X1 i_1_230 (.A1(n_1_7), .A2(n_1_70), .ZN(n_1_189));
   INV_X1 i_1_231 (.A(in2[10]), .ZN(n_1_190));
   INV_X1 i_1_232 (.A(in2[11]), .ZN(n_1_191));
endmodule

module carry_lookahead_adder_4bit__4_711(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_0;
   wire n_0_1;
   wire n_0_6;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;

   XNOR2_X1 i_0_0 (.A(n_0_6), .B(n_0_0), .ZN(sum[1]));
   XNOR2_X1 i_0_1 (.A(in1[1]), .B(in0[1]), .ZN(n_0_0));
   AOI22_X1 i_0_2 (.A1(n_0_16), .A2(n_0_12), .B1(in1[3]), .B2(in0[3]), .ZN(n_0_1));
   NOR2_X1 i_0_3 (.A1(n_0_1), .A2(n_0_17), .ZN(cout));
   BUF_X1 i_0_4 (.A(n_0_10), .Z(n_0_6));
   XOR2_X1 i_0_5 (.A(cin), .B(n_0_2), .Z(sum[0]));
   AOI21_X1 i_0_6 (.A(n_0_4), .B1(in1[0]), .B2(in0[0]), .ZN(n_0_2));
   NAND2_X1 i_0_7 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_3));
   NOR2_X1 i_0_8 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_4));
   XNOR2_X1 i_0_9 (.A(n_0_7), .B(n_0_5), .ZN(sum[2]));
   NAND2_X1 i_0_10 (.A1(n_0_9), .A2(n_0_8), .ZN(n_0_5));
   NAND2_X1 i_0_11 (.A1(n_0_12), .A2(n_0_11), .ZN(n_0_7));
   NAND2_X1 i_0_12 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_8));
   OAI21_X1 i_0_13 (.A(n_0_10), .B1(in1[1]), .B2(in0[1]), .ZN(n_0_9));
   OAI21_X1 i_0_14 (.A(n_0_3), .B1(n_0_13), .B2(n_0_4), .ZN(n_0_10));
   NAND2_X1 i_0_15 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_11));
   OR2_X1 i_0_16 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_12));
   INV_X1 i_0_17 (.A(cin), .ZN(n_0_13));
   XNOR2_X1 i_0_18 (.A(n_0_15), .B(n_0_14), .ZN(sum[3]));
   NAND2_X1 i_0_19 (.A1(n_0_12), .A2(n_0_16), .ZN(n_0_14));
   AOI21_X1 i_0_20 (.A(n_0_17), .B1(in1[3]), .B2(in0[3]), .ZN(n_0_15));
   NAND3_X1 i_0_21 (.A1(n_0_11), .A2(n_0_8), .A3(n_0_9), .ZN(n_0_16));
   NOR2_X1 i_0_22 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_17));
endmodule

module carry_lookahead_adder_4bit__4_720(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_10;
   wire n_0_11;
   wire n_0_7;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_8;
   wire n_0_9;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;

   XNOR2_X1 i_0_0 (.A(cin), .B(n_0_7), .ZN(sum[0]));
   XNOR2_X1 i_0_1 (.A(n_0_10), .B(n_0_1), .ZN(sum[3]));
   NOR2_X1 i_0_2 (.A1(n_0_13), .A2(n_0_11), .ZN(n_0_10));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(n_0_11));
   NAND2_X1 i_0_4 (.A1(n_0_6), .A2(n_0_8), .ZN(n_0_7));
   AOI21_X1 i_0_5 (.A(n_0_13), .B1(n_0_1), .B2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_0));
   NAND2_X1 i_0_7 (.A1(n_0_3), .A2(n_0_2), .ZN(n_0_1));
   OAI211_X1 i_0_8 (.A(n_0_9), .B(n_0_12), .C1(n_0_5), .C2(n_0_4), .ZN(n_0_2));
   OR2_X1 i_0_9 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_3));
   NOR2_X1 i_0_10 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_4));
   AOI22_X1 i_0_11 (.A1(in1[0]), .A2(in0[0]), .B1(cin), .B2(n_0_6), .ZN(n_0_5));
   OR2_X1 i_0_12 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_6));
   NAND2_X1 i_0_13 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_8));
   NAND2_X1 i_0_14 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_9));
   NAND2_X1 i_0_15 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_12));
   NOR2_X1 i_0_16 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_13));
   XNOR2_X1 i_0_17 (.A(n_0_5), .B(n_0_14), .ZN(sum[1]));
   XOR2_X1 i_0_18 (.A(in1[1]), .B(in0[1]), .Z(n_0_14));
   XNOR2_X1 i_0_19 (.A(n_0_16), .B(n_0_15), .ZN(sum[2]));
   OAI21_X1 i_0_20 (.A(n_0_9), .B1(n_0_5), .B2(n_0_4), .ZN(n_0_15));
   NAND2_X1 i_0_21 (.A1(n_0_3), .A2(n_0_12), .ZN(n_0_16));
endmodule

module carry_lookahead_adder_4bit__4_729(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_10;
   wire n_0_11;
   wire n_0_7;
   wire n_0_13;
   wire n_0_15;
   wire n_0_1;
   wire n_0_12;
   wire n_0_18;
   wire n_0_0;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_8;
   wire n_0_9;
   wire n_0_14;
   wire n_0_16;
   wire n_0_17;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;

   XNOR2_X1 i_0_0 (.A(cin), .B(n_0_7), .ZN(sum[0]));
   XNOR2_X1 i_0_1 (.A(n_0_10), .B(n_0_1), .ZN(sum[3]));
   NOR2_X1 i_0_2 (.A1(n_0_13), .A2(n_0_11), .ZN(n_0_10));
   INV_X1 i_0_3 (.A(n_0_12), .ZN(n_0_11));
   NAND2_X1 i_0_4 (.A1(n_0_15), .A2(n_0_4), .ZN(n_0_7));
   BUF_X1 i_0_5 (.A(n_0_20), .Z(n_0_13));
   BUF_X1 i_0_6 (.A(n_0_3), .Z(n_0_15));
   BUF_X1 i_0_7 (.A(n_0_18), .Z(n_0_1));
   BUF_X1 i_0_8 (.A(n_0_0), .Z(n_0_12));
   OAI21_X1 i_0_9 (.A(n_0_25), .B1(n_0_16), .B2(n_0_19), .ZN(n_0_18));
   NAND2_X1 i_0_10 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_0));
   NOR2_X1 i_0_11 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_2));
   OR2_X1 i_0_12 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_3));
   NAND2_X1 i_0_13 (.A1(in1[0]), .A2(in0[0]), .ZN(n_0_4));
   INV_X1 i_0_14 (.A(n_0_4), .ZN(n_0_5));
   OAI21_X1 i_0_15 (.A(n_0_3), .B1(n_0_5), .B2(cin), .ZN(n_0_6));
   NOR2_X1 i_0_16 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_8));
   INV_X1 i_0_17 (.A(in1[1]), .ZN(n_0_9));
   INV_X1 i_0_18 (.A(in0[1]), .ZN(n_0_14));
   OAI22_X1 i_0_19 (.A1(n_0_6), .A2(n_0_8), .B1(n_0_9), .B2(n_0_14), .ZN(n_0_16));
   NAND2_X1 i_0_20 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_17));
   INV_X1 i_0_21 (.A(n_0_17), .ZN(n_0_19));
   NOR2_X1 i_0_22 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_20));
   INV_X1 i_0_23 (.A(n_0_20), .ZN(n_0_21));
   OAI21_X1 i_0_24 (.A(n_0_21), .B1(n_0_16), .B2(n_0_19), .ZN(n_0_22));
   OAI21_X1 i_0_25 (.A(n_0_0), .B1(n_0_22), .B2(n_0_2), .ZN(cout));
   XNOR2_X1 i_0_26 (.A(n_0_6), .B(n_0_23), .ZN(sum[1]));
   XOR2_X1 i_0_27 (.A(in1[1]), .B(in0[1]), .Z(n_0_23));
   XNOR2_X1 i_0_28 (.A(n_0_16), .B(n_0_24), .ZN(sum[2]));
   NAND2_X1 i_0_29 (.A1(n_0_25), .A2(n_0_17), .ZN(n_0_24));
   INV_X1 i_0_30 (.A(n_0_2), .ZN(n_0_25));
endmodule

module carry_lookahead_adder_4bit__4_738(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_7;
   wire n_0_3;
   wire n_0_1;
   wire n_0_4;
   wire n_0_5;
   wire n_0_8;
   wire n_0_16;
   wire n_0_0;
   wire n_0_2;
   wire n_0_6;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;

   XNOR2_X1 i_0_0 (.A(cin), .B(n_0_7), .ZN(sum[0]));
   XNOR2_X1 i_0_1 (.A(n_0_13), .B(n_0_1), .ZN(sum[3]));
   NAND2_X1 i_0_2 (.A1(n_0_6), .A2(n_0_9), .ZN(n_0_7));
   NAND2_X1 i_0_3 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_3));
   AOI21_X1 i_0_4 (.A(n_0_15), .B1(n_0_1), .B2(n_0_14), .ZN(cout));
   OAI21_X1 i_0_5 (.A(n_0_2), .B1(n_0_5), .B2(n_0_4), .ZN(n_0_1));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(n_0_4));
   XNOR2_X1 i_0_7 (.A(n_0_5), .B(n_0_0), .ZN(sum[2]));
   AOI21_X1 i_0_8 (.A(n_0_16), .B1(n_0_11), .B2(n_0_8), .ZN(n_0_5));
   NAND2_X1 i_0_9 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_8));
   NOR2_X1 i_0_10 (.A1(in1[1]), .A2(in0[1]), .ZN(n_0_16));
   NAND2_X1 i_0_11 (.A1(n_0_2), .A2(n_0_3), .ZN(n_0_0));
   OR2_X1 i_0_12 (.A1(in0[2]), .A2(in1[2]), .ZN(n_0_2));
   OR2_X1 i_0_13 (.A1(in0[0]), .A2(in1[0]), .ZN(n_0_6));
   NAND2_X1 i_0_14 (.A1(in0[0]), .A2(in1[0]), .ZN(n_0_9));
   INV_X1 i_0_15 (.A(n_0_9), .ZN(n_0_10));
   OAI21_X1 i_0_16 (.A(n_0_6), .B1(n_0_10), .B2(cin), .ZN(n_0_11));
   XNOR2_X1 i_0_17 (.A(in0[1]), .B(in1[1]), .ZN(n_0_12));
   XOR2_X1 i_0_18 (.A(n_0_11), .B(n_0_12), .Z(sum[1]));
   AOI21_X1 i_0_19 (.A(n_0_15), .B1(in1[3]), .B2(in0[3]), .ZN(n_0_13));
   NAND2_X1 i_0_20 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_14));
   NOR2_X1 i_0_21 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_15));
endmodule

module carry_lookahead_adder_4bit(in0, in1, cin, sum, cout, v);
   input [3:0]in0;
   input [3:0]in1;
   input cin;
   output [3:0]sum;
   output cout;
   output v;

   wire n_0_4;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_32;

   OAI211_X1 i_0_0 (.A(in1[1]), .B(in0[1]), .C1(in0[2]), .C2(in1[2]), .ZN(n_0_4));
   NOR2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(v));
   AOI21_X1 i_0_2 (.A(n_0_32), .B1(n_0_26), .B2(n_0_27), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(n_0_1));
   NAND3_X1 i_0_4 (.A1(n_0_26), .A2(n_0_10), .A3(n_0_27), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(n_0_5), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_11), .A2(n_0_7), .ZN(n_0_6));
   OR2_X1 i_0_8 (.A1(in1[2]), .A2(in0[2]), .ZN(n_0_7));
   INV_X1 i_0_9 (.A(n_0_21), .ZN(n_0_11));
   XNOR2_X1 i_0_10 (.A(n_0_12), .B(in1[0]), .ZN(sum[0]));
   XNOR2_X1 i_0_11 (.A(cin), .B(in0[0]), .ZN(n_0_12));
   AND2_X1 i_0_12 (.A1(n_0_19), .A2(n_0_13), .ZN(sum[1]));
   NAND3_X1 i_0_13 (.A1(n_0_30), .A2(n_0_31), .A3(n_0_21), .ZN(n_0_13));
   INV_X1 i_0_14 (.A(n_0_14), .ZN(sum[2]));
   NAND2_X1 i_0_15 (.A1(n_0_15), .A2(n_0_18), .ZN(n_0_14));
   OAI21_X1 i_0_16 (.A(n_0_17), .B1(n_0_20), .B2(n_0_16), .ZN(n_0_15));
   INV_X1 i_0_17 (.A(n_0_22), .ZN(n_0_16));
   INV_X1 i_0_18 (.A(n_0_23), .ZN(n_0_17));
   NAND3_X1 i_0_19 (.A1(n_0_19), .A2(n_0_23), .A3(n_0_22), .ZN(n_0_18));
   INV_X1 i_0_20 (.A(n_0_20), .ZN(n_0_19));
   AOI21_X1 i_0_21 (.A(n_0_21), .B1(n_0_30), .B2(n_0_31), .ZN(n_0_20));
   XNOR2_X1 i_0_22 (.A(in0[1]), .B(in1[1]), .ZN(n_0_21));
   NAND2_X1 i_0_23 (.A1(in0[1]), .A2(in1[1]), .ZN(n_0_22));
   NAND2_X1 i_0_24 (.A1(n_0_7), .A2(n_0_5), .ZN(n_0_23));
   INV_X1 i_0_25 (.A(n_0_24), .ZN(sum[3]));
   NAND2_X1 i_0_26 (.A1(n_0_28), .A2(n_0_25), .ZN(n_0_24));
   NAND3_X1 i_0_27 (.A1(n_0_26), .A2(n_0_27), .A3(n_0_8), .ZN(n_0_25));
   INV_X1 i_0_28 (.A(n_0_29), .ZN(n_0_26));
   INV_X1 i_0_29 (.A(n_0_3), .ZN(n_0_27));
   OAI21_X1 i_0_30 (.A(n_0_9), .B1(n_0_29), .B2(n_0_3), .ZN(n_0_28));
   AOI21_X1 i_0_31 (.A(n_0_6), .B1(n_0_30), .B2(n_0_31), .ZN(n_0_29));
   OAI21_X1 i_0_32 (.A(in1[0]), .B1(cin), .B2(in0[0]), .ZN(n_0_30));
   NAND2_X1 i_0_33 (.A1(cin), .A2(in0[0]), .ZN(n_0_31));
   INV_X1 i_0_34 (.A(n_0_9), .ZN(n_0_8));
   AOI21_X1 i_0_35 (.A(n_0_32), .B1(in1[3]), .B2(in0[3]), .ZN(n_0_9));
   NAND2_X1 i_0_36 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_10));
   NOR2_X1 i_0_37 (.A1(in1[3]), .A2(in0[3]), .ZN(n_0_32));
endmodule

module carry_lookahead_adder_20bit(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [19:0]in0;
   input [19:0]in1;
   input cin;
   output [19:0]sum;
   output cout;
   output v;

   wire c1;
   wire c2;
   wire c3;
   wire c4;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   carry_lookahead_adder_4bit__4_711 cla0 (.in0({in0[3], in0[2], in0[1], in0[0]}), 
      .in1({n_18, n_17, n_16, n_15}), .cin(sub), .sum({sum[3], sum[2], sum[1], 
      sum[0]}), .cout(c1), .v());
   carry_lookahead_adder_4bit__4_720 cla1 (.in0({in0[7], in0[6], in0[5], in0[4]}), 
      .in1({n_14, n_13, n_12, n_19}), .cin(c1), .sum({sum[7], sum[6], sum[5], 
      sum[4]}), .cout(c2), .v());
   carry_lookahead_adder_4bit__4_729 cla2 (.in0({in0[11], in0[10], in0[9], 
      in0[8]}), .in1({n_11, n_10, n_9, n_8}), .cin(c2), .sum({sum[11], sum[10], 
      sum[9], sum[8]}), .cout(c3), .v());
   carry_lookahead_adder_4bit__4_738 cla3 (.in0({in0[15], in0[14], in0[13], 
      in0[12]}), .in1({n_7, n_6, n_5, n_4}), .cin(c3), .sum({sum[15], sum[14], 
      sum[13], sum[12]}), .cout(c4), .v());
   carry_lookahead_adder_4bit cla4 (.in0({in0[19], in0[18], in0[17], in0[16]}), 
      .in1({n_3, n_2, n_1, n_0}), .cin(c4), .sum({sum[19], sum[18], sum[17], 
      sum[16]}), .cout(), .v(v));
   XOR2_X1 i_0_0 (.A(in1[16]), .B(sub), .Z(n_0));
   XOR2_X1 i_0_1 (.A(sub), .B(in1[17]), .Z(n_1));
   XOR2_X1 i_0_2 (.A(sub), .B(in1[18]), .Z(n_2));
   XOR2_X1 i_0_3 (.A(sub), .B(in1[19]), .Z(n_3));
   XOR2_X1 i_0_4 (.A(in1[12]), .B(sub), .Z(n_4));
   XOR2_X1 i_0_5 (.A(sub), .B(in1[13]), .Z(n_5));
   XOR2_X1 i_0_6 (.A(sub), .B(in1[14]), .Z(n_6));
   XOR2_X1 i_0_7 (.A(sub), .B(in1[15]), .Z(n_7));
   XOR2_X1 i_0_8 (.A(in1[8]), .B(sub), .Z(n_8));
   XOR2_X1 i_0_9 (.A(sub), .B(in1[9]), .Z(n_9));
   XOR2_X1 i_0_10 (.A(sub), .B(in1[10]), .Z(n_10));
   XOR2_X1 i_0_11 (.A(sub), .B(in1[11]), .Z(n_11));
   XOR2_X1 i_0_13 (.A(sub), .B(in1[5]), .Z(n_12));
   XOR2_X1 i_0_14 (.A(sub), .B(in1[6]), .Z(n_13));
   XOR2_X1 i_0_15 (.A(sub), .B(in1[7]), .Z(n_14));
   XNOR2_X1 i_0_12 (.A(in1[0]), .B(n_0_3), .ZN(n_15));
   XNOR2_X1 i_0_16 (.A(in1[1]), .B(n_0_3), .ZN(n_16));
   XNOR2_X1 i_0_17 (.A(in1[2]), .B(n_0_3), .ZN(n_17));
   NAND2_X1 i_0_18 (.A1(n_0_1), .A2(n_0_0), .ZN(n_18));
   NAND2_X1 i_0_19 (.A1(in1[3]), .A2(n_0_3), .ZN(n_0_0));
   NAND2_X1 i_0_20 (.A1(n_0_2), .A2(sub), .ZN(n_0_1));
   INV_X1 i_0_21 (.A(in1[3]), .ZN(n_0_2));
   XNOR2_X1 i_0_22 (.A(in1[4]), .B(n_0_3), .ZN(n_19));
   INV_X1 i_0_23 (.A(sub), .ZN(n_0_3));
endmodule

module add_sub_cla(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   wire v;
   wire [19:0]tempOut;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_1_1;
   wire [19:0]tempIn11;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;
   wire n_1_28;
   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_52;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire [19:0]tempIn22;
   wire n_1_81;
   wire n_1_82;
   wire n_1_83;
   wire n_1_84;
   wire n_1_85;
   wire n_1_86;
   wire n_1_87;
   wire n_1_88;
   wire n_1_89;
   wire n_1_90;
   wire n_1_91;
   wire n_1_92;
   wire n_1_93;
   wire n_1_94;
   wire n_1_95;
   wire n_1_96;
   wire n_1_97;
   wire n_1_98;
   wire n_1_99;
   wire n_1_102;
   wire n_1_105;
   wire n_1_106;
   wire n_1_107;
   wire n_1_108;
   wire n_1_109;
   wire n_1_112;
   wire n_1_113;
   wire n_1_114;
   wire n_1_123;
   wire n_1_124;
   wire n_1_146;
   wire n_1_147;
   wire n_1_148;
   wire n_1_151;
   wire n_1_155;
   wire n_1_156;
   wire n_1_157;
   wire n_1_158;
   wire n_1_159;
   wire n_1_153;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_78;
   wire n_1_63;
   wire n_1_65;
   wire n_1_66;
   wire n_1_67;
   wire n_1_69;
   wire n_1_70;
   wire n_1_110;
   wire n_1_73;
   wire n_1_74;
   wire n_1_15;
   wire n_1_75;
   wire n_1_76;
   wire n_1_77;
   wire n_1_79;
   wire n_1_80;
   wire n_1_120;
   wire n_1_127;
   wire n_1_133;
   wire n_1_134;
   wire n_1_135;
   wire n_1_136;
   wire n_1_138;
   wire n_1_139;
   wire n_1_140;
   wire n_1_141;
   wire n_1_142;
   wire n_1_144;
   wire n_1_145;
   wire n_1_161;
   wire n_1_162;
   wire n_1_163;
   wire n_1_164;
   wire n_1_165;
   wire n_1_55;
   wire n_1_166;
   wire n_1_167;
   wire n_1_168;
   wire n_1_40;
   wire n_1_169;
   wire n_1_170;
   wire n_1_60;
   wire n_1_171;
   wire n_1_172;
   wire n_1_54;
   wire n_1_174;
   wire n_1_175;
   wire n_1_176;
   wire n_1_49;
   wire n_1_177;
   wire n_1_178;
   wire n_1_41;
   wire n_1_179;
   wire n_1_62;
   wire n_1_180;
   wire n_1_61;
   wire n_1_64;
   wire n_1_181;
   wire n_1_182;
   wire n_1_183;
   wire n_1_184;
   wire n_1_51;
   wire n_1_50;
   wire n_1_186;
   wire n_1_187;
   wire n_1_188;
   wire n_1_189;
   wire n_1_190;
   wire n_1_191;
   wire n_1_192;
   wire n_1_193;
   wire n_1_111;
   wire n_1_194;
   wire n_1_116;
   wire n_1_117;
   wire n_1_200;
   wire n_1_103;
   wire n_1_0;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_16;
   wire n_1_17;
   wire n_1_53;
   wire n_1_68;
   wire n_1_71;
   wire n_1_72;
   wire n_1_100;
   wire n_1_101;
   wire n_1_104;
   wire n_1_115;
   wire n_1_118;
   wire n_1_119;
   wire n_1_121;
   wire n_1_122;
   wire n_1_125;
   wire n_1_126;
   wire n_1_128;
   wire n_1_129;
   wire n_1_130;
   wire n_1_131;
   wire n_1_132;
   wire n_1_137;
   wire n_1_143;
   wire n_1_149;
   wire n_1_150;
   wire n_1_152;
   wire n_1_154;
   wire n_1_160;
   wire n_1_173;
   wire n_1_185;
   wire n_1_195;
   wire n_1_196;
   wire n_1_197;
   wire n_1_198;
   wire n_1_199;
   wire n_1_201;
   wire n_1_202;
   wire n_1_203;
   wire n_1_204;
   wire n_1_205;
   wire n_1_206;
   wire n_1_207;
   wire n_1_208;
   wire n_1_209;
   wire n_1_210;
   wire n_1_211;

   carry_lookahead_adder_20bit cs0 (.sub(sub), .in0({in1[12], tempIn11[18], 
      tempIn11[17], tempIn11[16], tempIn11[15], tempIn11[14], tempIn11[13], 
      tempIn11[12], tempIn11[11], tempIn11[10], tempIn11[9], tempIn11[8], 
      tempIn11[7], tempIn11[6], tempIn11[5], tempIn11[4], tempIn11[3], 
      tempIn11[2], tempIn11[1], tempIn11[0]}), .in1({in2[12], tempIn22[18], 
      tempIn22[17], tempIn22[16], tempIn22[15], tempIn22[14], tempIn22[13], 
      tempIn22[12], tempIn22[11], tempIn22[10], tempIn22[9], tempIn22[8], 
      tempIn22[7], tempIn22[6], tempIn22[5], tempIn22[4], tempIn22[3], 
      tempIn22[2], tempIn22[1], tempIn22[0]}), .cin(), .sum({tempOut[19], 
      tempOut[18], tempOut[17], tempOut[16], tempOut[15], tempOut[14], 
      tempOut[13], out[12], out[11], out[10], out[9], out[8], out[7], out[6], 
      out[5], out[4], out[3], out[2], out[1], out[0]}), .cout(), .v(v));
   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_10), .ZN(invalid));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_9), .ZN(n_0_0));
   NAND3_X1 i_0_2 (.A1(n_0_8), .A2(n_0_7), .A3(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_3), .ZN(n_0_2));
   NAND3_X1 i_0_4 (.A1(n_0_5), .A2(n_0_6), .A3(n_0_4), .ZN(n_0_3));
   NOR4_X1 i_0_5 (.A1(tempOut[15]), .A2(tempOut[14]), .A3(tempOut[13]), .A4(
      out[12]), .ZN(n_0_4));
   INV_X1 i_0_6 (.A(tempOut[16]), .ZN(n_0_5));
   INV_X1 i_0_7 (.A(tempOut[17]), .ZN(n_0_6));
   INV_X1 i_0_8 (.A(tempOut[18]), .ZN(n_0_7));
   INV_X1 i_0_9 (.A(tempOut[19]), .ZN(n_0_8));
   NAND3_X1 i_0_10 (.A1(tempOut[19]), .A2(tempOut[18]), .A3(n_0_11), .ZN(n_0_9));
   INV_X1 i_0_11 (.A(v), .ZN(n_0_10));
   NOR2_X1 i_0_12 (.A1(n_0_13), .A2(n_0_12), .ZN(n_0_11));
   NAND4_X1 i_0_13 (.A1(tempOut[17]), .A2(tempOut[16]), .A3(tempOut[15]), 
      .A4(out[12]), .ZN(n_0_12));
   NAND2_X1 i_0_14 (.A1(tempOut[14]), .A2(tempOut[13]), .ZN(n_0_13));
   OAI21_X1 i_1_0 (.A(n_1_1), .B1(n_1_153), .B2(n_1_104), .ZN(out[14]));
   NAND2_X1 i_1_1 (.A1(in1[14]), .A2(n_1_104), .ZN(n_1_1));
   NAND2_X1 i_1_4 (.A1(n_1_0), .A2(n_1_71), .ZN(out[15]));
   AND2_X1 i_1_2 (.A1(in1[0]), .A2(n_1_55), .ZN(tempIn11[0]));
   AOI222_X1 i_1_3 (.A1(n_1_155), .A2(n_1_55), .B1(n_1_54), .B2(n_1_18), 
      .C1(n_1_51), .C2(n_1_15), .ZN(tempIn11[7]));
   AOI222_X1 i_1_5 (.A1(n_1_156), .A2(n_1_55), .B1(n_1_54), .B2(n_1_21), 
      .C1(n_1_51), .C2(n_1_18), .ZN(tempIn11[8]));
   AOI221_X1 i_1_6 (.A(n_1_19), .B1(in1[5]), .B2(n_1_40), .C1(in1[7]), .C2(
      n_1_41), .ZN(n_1_18));
   INV_X1 i_1_7 (.A(n_1_20), .ZN(n_1_19));
   AOI22_X1 i_1_8 (.A1(in1[3]), .A2(n_1_49), .B1(in1[1]), .B2(n_1_60), .ZN(
      n_1_20));
   AOI222_X1 i_1_33 (.A1(n_1_157), .A2(n_1_55), .B1(n_1_54), .B2(n_1_24), 
      .C1(n_1_51), .C2(n_1_21), .ZN(tempIn11[9]));
   AOI221_X1 i_1_9 (.A(n_1_22), .B1(in1[6]), .B2(n_1_40), .C1(in1[8]), .C2(
      n_1_41), .ZN(n_1_21));
   INV_X1 i_1_10 (.A(n_1_23), .ZN(n_1_22));
   AOI22_X1 i_1_11 (.A1(in1[4]), .A2(n_1_49), .B1(in1[2]), .B2(n_1_60), .ZN(
      n_1_23));
   AOI222_X1 i_1_12 (.A1(n_1_158), .A2(n_1_55), .B1(n_1_54), .B2(n_1_27), 
      .C1(n_1_51), .C2(n_1_24), .ZN(tempIn11[10]));
   AOI221_X1 i_1_13 (.A(n_1_25), .B1(in1[7]), .B2(n_1_40), .C1(in1[9]), .C2(
      n_1_41), .ZN(n_1_24));
   INV_X1 i_1_14 (.A(n_1_26), .ZN(n_1_25));
   AOI22_X1 i_1_15 (.A1(in1[5]), .A2(n_1_49), .B1(in1[3]), .B2(n_1_60), .ZN(
      n_1_26));
   AOI222_X1 i_1_41 (.A1(n_1_159), .A2(n_1_55), .B1(n_1_51), .B2(n_1_27), 
      .C1(n_1_54), .C2(n_1_31), .ZN(tempIn11[11]));
   AOI221_X1 i_1_16 (.A(n_1_28), .B1(in1[8]), .B2(n_1_40), .C1(in1[4]), .C2(
      n_1_60), .ZN(n_1_27));
   INV_X1 i_1_17 (.A(n_1_29), .ZN(n_1_28));
   AOI22_X1 i_1_18 (.A1(in1[10]), .A2(n_1_41), .B1(in1[6]), .B2(n_1_49), 
      .ZN(n_1_29));
   OAI21_X1 i_1_45 (.A(n_1_30), .B1(n_1_50), .B2(n_1_31), .ZN(tempIn11[12]));
   AOI21_X1 i_1_46 (.A(n_1_43), .B1(n_1_54), .B2(n_1_35), .ZN(n_1_30));
   AOI221_X1 i_1_47 (.A(n_1_32), .B1(in1[9]), .B2(n_1_40), .C1(in1[11]), 
      .C2(n_1_41), .ZN(n_1_31));
   INV_X1 i_1_48 (.A(n_1_33), .ZN(n_1_32));
   AOI22_X1 i_1_49 (.A1(in1[5]), .A2(n_1_60), .B1(in1[7]), .B2(n_1_49), .ZN(
      n_1_33));
   INV_X1 i_1_50 (.A(n_1_34), .ZN(tempIn11[13]));
   AOI221_X1 i_1_51 (.A(n_1_43), .B1(n_1_54), .B2(n_1_38), .C1(n_1_51), .C2(
      n_1_35), .ZN(n_1_34));
   AOI221_X1 i_1_52 (.A(n_1_36), .B1(n_1_62), .B2(n_1_48), .C1(n_1_156), 
      .C2(n_1_49), .ZN(n_1_35));
   OAI33_X1 i_1_53 (.A1(n_1_64), .A2(n_1_62), .A3(in1[6]), .B1(n_1_63), .B2(
      n_1_62), .B3(in1[10]), .ZN(n_1_36));
   INV_X1 i_1_54 (.A(n_1_37), .ZN(tempIn11[14]));
   AOI221_X1 i_1_55 (.A(n_1_43), .B1(n_1_51), .B2(n_1_38), .C1(n_1_54), .C2(
      n_1_44), .ZN(n_1_37));
   AOI221_X1 i_1_56 (.A(n_1_39), .B1(n_1_62), .B2(n_1_48), .C1(n_1_155), 
      .C2(n_1_60), .ZN(n_1_38));
   OAI33_X1 i_1_57 (.A1(n_1_63), .A2(n_1_62), .A3(in1[11]), .B1(n_1_64), 
      .B2(n_1_61), .B3(in1[9]), .ZN(n_1_39));
   INV_X1 i_1_60 (.A(n_1_42), .ZN(tempIn11[15]));
   AOI221_X1 i_1_61 (.A(n_1_43), .B1(n_1_54), .B2(n_1_47), .C1(n_1_51), .C2(
      n_1_44), .ZN(n_1_42));
   AND2_X1 i_1_62 (.A1(in1[12]), .A2(n_1_55), .ZN(n_1_43));
   AOI221_X1 i_1_63 (.A(n_1_48), .B1(n_1_158), .B2(n_1_49), .C1(n_1_156), 
      .C2(n_1_60), .ZN(n_1_44));
   AOI221_X1 i_1_64 (.A(n_1_45), .B1(n_1_158), .B2(n_1_52), .C1(n_1_51), 
      .C2(n_1_46), .ZN(tempIn11[16]));
   NOR3_X1 i_1_65 (.A1(in1[12]), .A2(n_1_51), .A3(n_1_52), .ZN(n_1_45));
   INV_X1 i_1_66 (.A(n_1_47), .ZN(n_1_46));
   AOI221_X1 i_1_67 (.A(n_1_48), .B1(n_1_157), .B2(n_1_60), .C1(n_1_159), 
      .C2(n_1_49), .ZN(n_1_47));
   NOR2_X1 i_1_68 (.A1(in1[12]), .A2(n_1_63), .ZN(n_1_48));
   AOI221_X1 i_1_72 (.A(n_1_56), .B1(n_1_159), .B2(n_1_52), .C1(n_1_158), 
      .C2(n_1_58), .ZN(tempIn11[17]));
   NOR3_X1 i_1_19 (.A1(n_1_64), .A2(n_1_62), .A3(n_1_118), .ZN(n_1_52));
   AOI21_X1 i_1_20 (.A(in1[12]), .B1(n_1_101), .B2(n_1_60), .ZN(n_1_56));
   OAI21_X1 i_1_21 (.A(n_1_57), .B1(n_1_159), .B2(n_1_59), .ZN(tempIn11[18]));
   NAND2_X1 i_1_22 (.A1(in1[12]), .A2(n_1_59), .ZN(n_1_57));
   INV_X1 i_1_23 (.A(n_1_59), .ZN(n_1_58));
   NAND3_X1 i_1_25 (.A1(n_1_101), .A2(n_1_60), .A3(n_1_119), .ZN(n_1_59));
   AOI222_X1 i_1_26 (.A1(n_1_146), .A2(n_1_101), .B1(n_1_116), .B2(n_1_78), 
      .C1(n_1_110), .C2(n_1_81), .ZN(tempIn22[7]));
   AOI222_X1 i_1_27 (.A1(n_1_147), .A2(n_1_101), .B1(n_1_110), .B2(n_1_84), 
      .C1(n_1_116), .C2(n_1_81), .ZN(tempIn22[8]));
   AOI221_X1 i_1_28 (.A(n_1_82), .B1(in2[1]), .B2(n_1_206), .C1(in2[3]), 
      .C2(n_1_195), .ZN(n_1_81));
   OAI21_X1 i_1_29 (.A(n_1_83), .B1(n_1_146), .B2(n_1_202), .ZN(n_1_82));
   NAND2_X1 i_1_30 (.A1(in2[5]), .A2(n_1_132), .ZN(n_1_83));
   AOI222_X1 i_1_31 (.A1(n_1_148), .A2(n_1_101), .B1(n_1_116), .B2(n_1_84), 
      .C1(n_1_110), .C2(n_1_87), .ZN(tempIn22[9]));
   AOI221_X1 i_1_32 (.A(n_1_85), .B1(in2[8]), .B2(n_1_103), .C1(in2[2]), 
      .C2(n_1_206), .ZN(n_1_84));
   INV_X1 i_1_34 (.A(n_1_86), .ZN(n_1_85));
   AOI22_X1 i_1_35 (.A1(in2[6]), .A2(n_1_132), .B1(in2[4]), .B2(n_1_195), 
      .ZN(n_1_86));
   AOI222_X1 i_1_36 (.A1(n_1_210), .A2(n_1_101), .B1(n_1_110), .B2(n_1_89), 
      .C1(n_1_116), .C2(n_1_87), .ZN(tempIn22[10]));
   AOI221_X1 i_1_37 (.A(n_1_88), .B1(in2[3]), .B2(n_1_206), .C1(in2[5]), 
      .C2(n_1_195), .ZN(n_1_87));
   OAI22_X1 i_1_38 (.A1(n_1_148), .A2(n_1_202), .B1(n_1_146), .B2(n_1_137), 
      .ZN(n_1_88));
   AOI222_X1 i_1_39 (.A1(n_1_211), .A2(n_1_101), .B1(n_1_116), .B2(n_1_89), 
      .C1(n_1_110), .C2(n_1_92), .ZN(tempIn22[11]));
   AOI221_X1 i_1_40 (.A(n_1_90), .B1(in2[4]), .B2(n_1_206), .C1(in2[6]), 
      .C2(n_1_195), .ZN(n_1_89));
   OAI22_X1 i_1_42 (.A1(n_1_210), .A2(n_1_202), .B1(n_1_147), .B2(n_1_137), 
      .ZN(n_1_90));
   OAI21_X1 i_1_43 (.A(n_1_91), .B1(n_1_117), .B2(n_1_92), .ZN(tempIn22[12]));
   AOI21_X1 i_1_44 (.A(n_1_106), .B1(n_1_110), .B2(n_1_95), .ZN(n_1_91));
   AOI221_X1 i_1_58 (.A(n_1_93), .B1(in2[5]), .B2(n_1_206), .C1(in2[7]), 
      .C2(n_1_195), .ZN(n_1_92));
   OAI22_X1 i_1_59 (.A1(n_1_148), .A2(n_1_137), .B1(n_1_211), .B2(n_1_202), 
      .ZN(n_1_93));
   INV_X1 i_1_69 (.A(n_1_94), .ZN(tempIn22[13]));
   AOI221_X1 i_1_70 (.A(n_1_106), .B1(n_1_110), .B2(n_1_98), .C1(n_1_116), 
      .C2(n_1_95), .ZN(n_1_94));
   AOI221_X1 i_1_71 (.A(n_1_96), .B1(n_1_196), .B2(n_1_114), .C1(n_1_147), 
      .C2(n_1_195), .ZN(n_1_95));
   OAI33_X1 i_1_73 (.A1(n_1_196), .A2(n_1_150), .A3(in2[6]), .B1(n_1_196), 
      .B2(n_1_197), .B3(in2[10]), .ZN(n_1_96));
   INV_X1 i_1_74 (.A(n_1_97), .ZN(tempIn22[14]));
   AOI221_X1 i_1_75 (.A(n_1_106), .B1(n_1_116), .B2(n_1_98), .C1(n_1_110), 
      .C2(n_1_107), .ZN(n_1_97));
   AOI221_X1 i_1_76 (.A(n_1_99), .B1(n_1_146), .B2(n_1_206), .C1(n_1_196), 
      .C2(n_1_114), .ZN(n_1_98));
   OAI21_X1 i_1_77 (.A(n_1_102), .B1(in2[11]), .B2(n_1_137), .ZN(n_1_99));
   NAND2_X1 i_1_78 (.A1(n_1_148), .A2(n_1_195), .ZN(n_1_102));
   INV_X1 i_1_79 (.A(n_1_105), .ZN(tempIn22[15]));
   AOI221_X1 i_1_80 (.A(n_1_106), .B1(n_1_113), .B2(n_1_110), .C1(n_1_116), 
      .C2(n_1_107), .ZN(n_1_105));
   NOR2_X1 i_1_81 (.A1(n_1_151), .A2(n_1_104), .ZN(n_1_106));
   AOI221_X1 i_1_82 (.A(n_1_114), .B1(n_1_210), .B2(n_1_195), .C1(n_1_147), 
      .C2(n_1_206), .ZN(n_1_107));
   AOI221_X1 i_1_83 (.A(n_1_108), .B1(n_1_151), .B2(n_1_109), .C1(n_1_116), 
      .C2(n_1_112), .ZN(tempIn22[16]));
   NOR4_X1 i_1_84 (.A1(n_1_196), .A2(n_1_150), .A3(n_1_111), .A4(in2[10]), 
      .ZN(n_1_108));
   AOI21_X1 i_1_85 (.A(n_1_116), .B1(n_1_206), .B2(n_1_110), .ZN(n_1_109));
   INV_X1 i_1_86 (.A(n_1_113), .ZN(n_1_112));
   AOI221_X1 i_1_87 (.A(n_1_114), .B1(n_1_148), .B2(n_1_206), .C1(n_1_211), 
      .C2(n_1_195), .ZN(n_1_113));
   NOR2_X1 i_1_88 (.A1(in2[12]), .A2(n_1_197), .ZN(n_1_114));
   AOI21_X1 i_1_89 (.A(n_1_123), .B1(n_1_151), .B2(n_1_124), .ZN(tempIn22[18]));
   NOR2_X1 i_1_90 (.A1(in2[11]), .A2(n_1_124), .ZN(n_1_123));
   NAND2_X1 i_1_91 (.A1(n_1_209), .A2(n_1_119), .ZN(n_1_124));
   INV_X1 i_1_92 (.A(in2[7]), .ZN(n_1_146));
   INV_X1 i_1_93 (.A(in2[8]), .ZN(n_1_147));
   INV_X1 i_1_94 (.A(in2[9]), .ZN(n_1_148));
   INV_X1 i_1_95 (.A(in2[12]), .ZN(n_1_151));
   INV_X1 i_1_96 (.A(in1[7]), .ZN(n_1_155));
   INV_X1 i_1_97 (.A(in1[8]), .ZN(n_1_156));
   INV_X1 i_1_198 (.A(in1[9]), .ZN(n_1_157));
   INV_X1 i_1_98 (.A(in1[10]), .ZN(n_1_158));
   INV_X1 i_1_99 (.A(in1[11]), .ZN(n_1_159));
   INV_X1 i_1_100 (.A(in2[14]), .ZN(n_1_153));
   NAND3_X1 i_1_101 (.A1(n_1_4), .A2(n_1_3), .A3(n_1_2), .ZN(tempIn22[4]));
   NAND2_X1 i_1_102 (.A1(n_1_101), .A2(in2[4]), .ZN(n_1_2));
   NAND3_X1 i_1_103 (.A1(n_1_104), .A2(n_1_204), .A3(n_1_7), .ZN(n_1_3));
   NAND3_X1 i_1_104 (.A1(n_1_104), .A2(n_1_119), .A3(n_1_191), .ZN(n_1_4));
   NAND3_X1 i_1_105 (.A1(n_1_198), .A2(n_1_6), .A3(n_1_5), .ZN(tempIn22[5]));
   NAND2_X1 i_1_106 (.A1(n_1_101), .A2(in2[5]), .ZN(n_1_5));
   NAND3_X1 i_1_107 (.A1(n_1_104), .A2(n_1_119), .A3(n_1_7), .ZN(n_1_6));
   NAND3_X1 i_1_108 (.A1(n_1_185), .A2(n_1_9), .A3(n_1_8), .ZN(n_1_7));
   NAND2_X1 i_1_109 (.A1(n_1_132), .A2(in2[2]), .ZN(n_1_8));
   NAND2_X1 i_1_110 (.A1(n_1_103), .A2(in2[4]), .ZN(n_1_9));
   INV_X1 i_1_111 (.A(n_1_66), .ZN(n_1_78));
   INV_X1 i_1_24 (.A(n_1_64), .ZN(n_1_63));
   OAI22_X1 i_1_112 (.A1(n_1_74), .A2(n_1_135), .B1(n_1_140), .B2(n_1_121), 
      .ZN(tempIn11[1]));
   NAND2_X1 i_1_113 (.A1(n_1_73), .A2(n_1_65), .ZN(tempIn22[6]));
   AOI22_X1 i_1_114 (.A1(n_1_66), .A2(n_1_110), .B1(in2[6]), .B2(n_1_101), 
      .ZN(n_1_65));
   NAND4_X1 i_1_115 (.A1(n_1_205), .A2(n_1_67), .A3(n_1_70), .A4(n_1_69), 
      .ZN(n_1_66));
   NAND2_X1 i_1_116 (.A1(n_1_195), .A2(in2[2]), .ZN(n_1_67));
   NAND2_X1 i_1_117 (.A1(n_1_132), .A2(in2[4]), .ZN(n_1_69));
   NAND2_X1 i_1_118 (.A1(n_1_103), .A2(in2[6]), .ZN(n_1_70));
   INV_X1 i_1_119 (.A(n_1_111), .ZN(n_1_110));
   NAND2_X1 i_1_120 (.A1(n_1_199), .A2(n_1_116), .ZN(n_1_73));
   NAND2_X1 i_1_121 (.A1(n_1_206), .A2(n_1_51), .ZN(n_1_74));
   INV_X1 i_1_122 (.A(n_1_167), .ZN(n_1_15));
   NAND2_X1 i_1_123 (.A1(n_1_80), .A2(n_1_75), .ZN(tempIn11[2]));
   INV_X1 i_1_124 (.A(n_1_76), .ZN(n_1_75));
   OAI21_X1 i_1_125 (.A(n_1_77), .B1(n_1_79), .B2(n_1_118), .ZN(n_1_76));
   NAND2_X1 i_1_126 (.A1(n_1_55), .A2(in1[2]), .ZN(n_1_77));
   INV_X1 i_1_127 (.A(n_1_133), .ZN(n_1_79));
   NAND3_X1 i_1_128 (.A1(n_1_206), .A2(in1[1]), .A3(n_1_51), .ZN(n_1_80));
   OAI211_X1 i_1_129 (.A(n_1_120), .B(n_1_127), .C1(n_1_184), .C2(n_1_121), 
      .ZN(tempIn11[3]));
   NAND2_X1 i_1_130 (.A1(n_1_139), .A2(n_1_54), .ZN(n_1_120));
   NAND2_X1 i_1_131 (.A1(n_1_133), .A2(n_1_51), .ZN(n_1_127));
   OAI21_X1 i_1_132 (.A(n_1_134), .B1(n_1_180), .B2(n_1_135), .ZN(n_1_133));
   NAND3_X1 i_1_133 (.A1(n_1_64), .A2(n_1_62), .A3(in1[2]), .ZN(n_1_134));
   INV_X1 i_1_134 (.A(in1[0]), .ZN(n_1_135));
   OAI211_X1 i_1_135 (.A(n_1_138), .B(n_1_136), .C1(n_1_141), .C2(n_1_118), 
      .ZN(tempIn11[4]));
   NAND2_X1 i_1_136 (.A1(n_1_55), .A2(in1[4]), .ZN(n_1_136));
   NAND2_X1 i_1_137 (.A1(n_1_139), .A2(n_1_51), .ZN(n_1_138));
   OAI22_X1 i_1_138 (.A1(n_1_184), .A2(n_1_179), .B1(n_1_180), .B2(n_1_140), 
      .ZN(n_1_139));
   INV_X1 i_1_139 (.A(in1[1]), .ZN(n_1_140));
   INV_X1 i_1_140 (.A(n_1_161), .ZN(n_1_141));
   NAND3_X1 i_1_141 (.A1(n_1_144), .A2(n_1_145), .A3(n_1_142), .ZN(tempIn11[5]));
   NAND2_X1 i_1_142 (.A1(n_1_55), .A2(in1[5]), .ZN(n_1_142));
   NAND2_X1 i_1_143 (.A1(n_1_175), .A2(n_1_54), .ZN(n_1_144));
   NAND2_X1 i_1_144 (.A1(n_1_161), .A2(n_1_51), .ZN(n_1_145));
   OAI211_X1 i_1_145 (.A(n_1_163), .B(n_1_162), .C1(n_1_164), .C2(n_1_179), 
      .ZN(n_1_161));
   NAND2_X1 i_1_146 (.A1(n_1_49), .A2(in1[0]), .ZN(n_1_162));
   NAND2_X1 i_1_147 (.A1(n_1_40), .A2(in1[2]), .ZN(n_1_163));
   INV_X1 i_1_148 (.A(in1[4]), .ZN(n_1_164));
   NAND3_X1 i_1_149 (.A1(n_1_166), .A2(n_1_174), .A3(n_1_165), .ZN(tempIn11[6]));
   NAND2_X1 i_1_150 (.A1(n_1_55), .A2(in1[6]), .ZN(n_1_165));
   INV_X1 i_1_151 (.A(n_1_121), .ZN(n_1_55));
   NAND2_X1 i_1_152 (.A1(n_1_167), .A2(n_1_54), .ZN(n_1_166));
   NAND4_X1 i_1_153 (.A1(n_1_169), .A2(n_1_168), .A3(n_1_172), .A4(n_1_170), 
      .ZN(n_1_167));
   NAND2_X1 i_1_154 (.A1(n_1_40), .A2(in1[4]), .ZN(n_1_168));
   INV_X1 i_1_155 (.A(n_1_180), .ZN(n_1_40));
   NAND2_X1 i_1_156 (.A1(n_1_41), .A2(in1[6]), .ZN(n_1_169));
   NAND2_X1 i_1_157 (.A1(n_1_60), .A2(in1[0]), .ZN(n_1_170));
   INV_X1 i_1_158 (.A(n_1_171), .ZN(n_1_60));
   NAND2_X1 i_1_159 (.A1(n_1_181), .A2(n_1_61), .ZN(n_1_171));
   NAND2_X1 i_1_160 (.A1(n_1_49), .A2(in1[2]), .ZN(n_1_172));
   INV_X1 i_1_161 (.A(n_1_118), .ZN(n_1_54));
   NAND2_X1 i_1_162 (.A1(n_1_175), .A2(n_1_51), .ZN(n_1_174));
   OAI211_X1 i_1_163 (.A(n_1_178), .B(n_1_176), .C1(n_1_184), .C2(n_1_180), 
      .ZN(n_1_175));
   NAND2_X1 i_1_164 (.A1(n_1_49), .A2(in1[1]), .ZN(n_1_176));
   INV_X1 i_1_165 (.A(n_1_177), .ZN(n_1_49));
   NAND2_X1 i_1_166 (.A1(n_1_62), .A2(n_1_181), .ZN(n_1_177));
   NAND2_X1 i_1_167 (.A1(n_1_41), .A2(in1[5]), .ZN(n_1_178));
   INV_X1 i_1_168 (.A(n_1_179), .ZN(n_1_41));
   NAND2_X1 i_1_169 (.A1(n_1_64), .A2(n_1_62), .ZN(n_1_179));
   INV_X1 i_1_170 (.A(n_1_61), .ZN(n_1_62));
   NAND2_X1 i_1_171 (.A1(n_1_64), .A2(n_1_61), .ZN(n_1_180));
   XNOR2_X1 i_1_172 (.A(n_1_149), .B(n_1_16), .ZN(n_1_61));
   INV_X1 i_1_173 (.A(n_1_181), .ZN(n_1_64));
   NAND2_X1 i_1_174 (.A1(n_1_183), .A2(n_1_182), .ZN(n_1_181));
   NAND2_X1 i_1_175 (.A1(n_1_68), .A2(n_1_173), .ZN(n_1_182));
   NAND2_X1 i_1_176 (.A1(n_1_53), .A2(n_1_160), .ZN(n_1_183));
   INV_X1 i_1_177 (.A(in1[3]), .ZN(n_1_184));
   INV_X1 i_1_178 (.A(n_1_50), .ZN(n_1_51));
   NAND2_X1 i_1_179 (.A1(n_1_121), .A2(n_1_119), .ZN(n_1_50));
   OAI21_X1 i_1_180 (.A(n_1_186), .B1(n_1_192), .B2(n_1_104), .ZN(tempIn22[1]));
   NAND2_X1 i_1_181 (.A1(n_1_188), .A2(in2[0]), .ZN(n_1_186));
   OAI21_X1 i_1_182 (.A(n_1_187), .B1(n_1_131), .B2(n_1_111), .ZN(tempIn22[2]));
   AOI22_X1 i_1_183 (.A1(n_1_188), .A2(in2[1]), .B1(in2[2]), .B2(n_1_101), 
      .ZN(n_1_187));
   NOR2_X1 i_1_184 (.A1(n_1_202), .A2(n_1_117), .ZN(n_1_188));
   INV_X1 i_1_185 (.A(n_1_189), .ZN(tempIn22[3]));
   OAI211_X1 i_1_186 (.A(n_1_194), .B(n_1_190), .C1(n_1_111), .C2(n_1_191), 
      .ZN(n_1_189));
   NAND2_X1 i_1_187 (.A1(n_1_101), .A2(n_1_193), .ZN(n_1_190));
   OAI22_X1 i_1_188 (.A1(n_1_193), .A2(n_1_202), .B1(n_1_137), .B2(n_1_192), 
      .ZN(n_1_191));
   INV_X1 i_1_189 (.A(in2[1]), .ZN(n_1_192));
   INV_X1 i_1_190 (.A(in2[3]), .ZN(n_1_193));
   NAND2_X1 i_1_191 (.A1(n_1_204), .A2(n_1_104), .ZN(n_1_111));
   NAND3_X1 i_1_192 (.A1(n_1_131), .A2(n_1_200), .A3(n_1_116), .ZN(n_1_194));
   INV_X1 i_1_193 (.A(n_1_117), .ZN(n_1_116));
   NAND2_X1 i_1_194 (.A1(n_1_104), .A2(n_1_119), .ZN(n_1_117));
   NAND2_X1 i_1_195 (.A1(n_1_103), .A2(in2[2]), .ZN(n_1_200));
   INV_X1 i_1_196 (.A(n_1_202), .ZN(n_1_103));
   INV_X1 i_1_197 (.A(in1[15]), .ZN(n_1_0));
   NAND2_X1 i_1_199 (.A1(n_1_0), .A2(in2[15]), .ZN(n_1_10));
   INV_X1 i_1_200 (.A(in2[14]), .ZN(n_1_11));
   OR2_X1 i_1_201 (.A1(n_1_11), .A2(in1[14]), .ZN(n_1_12));
   NAND2_X1 i_1_202 (.A1(n_1_11), .A2(in1[14]), .ZN(n_1_13));
   INV_X1 i_1_203 (.A(in2[13]), .ZN(n_1_14));
   NAND2_X1 i_1_204 (.A1(n_1_14), .A2(in1[13]), .ZN(n_1_16));
   INV_X1 i_1_205 (.A(n_1_12), .ZN(n_1_17));
   OAI21_X1 i_1_206 (.A(n_1_13), .B1(n_1_16), .B2(n_1_17), .ZN(n_1_53));
   INV_X1 i_1_207 (.A(n_1_53), .ZN(n_1_68));
   INV_X1 i_1_208 (.A(in2[15]), .ZN(n_1_71));
   NAND2_X1 i_1_209 (.A1(n_1_71), .A2(in1[15]), .ZN(n_1_72));
   INV_X1 i_1_210 (.A(n_1_72), .ZN(n_1_100));
   OAI21_X1 i_1_211 (.A(n_1_10), .B1(n_1_53), .B2(n_1_100), .ZN(n_1_101));
   INV_X1 i_1_212 (.A(n_1_101), .ZN(n_1_104));
   INV_X1 i_1_213 (.A(in1[13]), .ZN(n_1_115));
   AOI22_X1 i_1_214 (.A1(n_1_115), .A2(n_1_104), .B1(n_1_101), .B2(n_1_14), 
      .ZN(out[13]));
   NAND3_X1 i_1_215 (.A1(n_1_16), .A2(n_1_125), .A3(n_1_121), .ZN(n_1_118));
   NAND2_X1 i_1_216 (.A1(n_1_16), .A2(n_1_125), .ZN(n_1_119));
   AOI21_X1 i_1_217 (.A(n_1_130), .B1(n_1_10), .B2(n_1_122), .ZN(n_1_121));
   OAI21_X1 i_1_218 (.A(n_1_13), .B1(n_1_129), .B2(n_1_126), .ZN(n_1_122));
   INV_X1 i_1_219 (.A(n_1_126), .ZN(n_1_125));
   NOR2_X1 i_1_220 (.A1(in1[13]), .A2(n_1_128), .ZN(n_1_126));
   INV_X1 i_1_221 (.A(in2[13]), .ZN(n_1_128));
   INV_X1 i_1_222 (.A(n_1_12), .ZN(n_1_129));
   INV_X1 i_1_223 (.A(n_1_72), .ZN(n_1_130));
   AND2_X1 i_1_224 (.A1(n_1_101), .A2(in2[0]), .ZN(tempIn22[0]));
   NAND2_X1 i_1_225 (.A1(in2[0]), .A2(n_1_132), .ZN(n_1_131));
   INV_X1 i_1_226 (.A(n_1_137), .ZN(n_1_132));
   NAND2_X1 i_1_227 (.A1(n_1_150), .A2(n_1_143), .ZN(n_1_137));
   XNOR2_X1 i_1_228 (.A(n_1_125), .B(n_1_149), .ZN(n_1_143));
   NAND2_X1 i_1_229 (.A1(n_1_13), .A2(n_1_12), .ZN(n_1_149));
   OAI22_X1 i_1_230 (.A1(n_1_173), .A2(n_1_152), .B1(n_1_122), .B2(n_1_160), 
      .ZN(n_1_150));
   INV_X1 i_1_231 (.A(n_1_154), .ZN(n_1_152));
   OAI21_X1 i_1_232 (.A(n_1_13), .B1(n_1_129), .B2(n_1_126), .ZN(n_1_154));
   INV_X1 i_1_233 (.A(n_1_173), .ZN(n_1_160));
   NAND2_X1 i_1_234 (.A1(n_1_10), .A2(n_1_72), .ZN(n_1_173));
   NAND2_X1 i_1_235 (.A1(in2[0]), .A2(n_1_195), .ZN(n_1_185));
   NOR2_X1 i_1_236 (.A1(n_1_150), .A2(n_1_143), .ZN(n_1_195));
   INV_X1 i_1_237 (.A(n_1_143), .ZN(n_1_196));
   INV_X1 i_1_238 (.A(n_1_150), .ZN(n_1_197));
   NAND3_X1 i_1_239 (.A1(n_1_204), .A2(n_1_104), .A3(n_1_199), .ZN(n_1_198));
   OAI21_X1 i_1_240 (.A(n_1_201), .B1(n_1_203), .B2(n_1_202), .ZN(n_1_199));
   AOI22_X1 i_1_241 (.A1(n_1_195), .A2(in2[1]), .B1(in2[3]), .B2(n_1_132), 
      .ZN(n_1_201));
   NAND2_X1 i_1_242 (.A1(n_1_150), .A2(n_1_196), .ZN(n_1_202));
   INV_X1 i_1_243 (.A(in2[5]), .ZN(n_1_203));
   INV_X1 i_1_244 (.A(n_1_119), .ZN(n_1_204));
   NAND2_X1 i_1_245 (.A1(in2[0]), .A2(n_1_206), .ZN(n_1_205));
   AND2_X1 i_1_246 (.A1(n_1_197), .A2(n_1_143), .ZN(n_1_206));
   INV_X1 i_1_247 (.A(n_1_207), .ZN(tempIn22[17]));
   OAI21_X1 i_1_248 (.A(n_1_208), .B1(in2[12]), .B2(n_1_209), .ZN(n_1_207));
   OAI221_X1 i_1_249 (.A(n_1_209), .B1(n_1_210), .B2(n_1_204), .C1(n_1_211), 
      .C2(n_1_119), .ZN(n_1_208));
   AND2_X1 i_1_250 (.A1(n_1_130), .A2(n_1_206), .ZN(n_1_209));
   INV_X1 i_1_251 (.A(in2[10]), .ZN(n_1_210));
   INV_X1 i_1_252 (.A(in2[11]), .ZN(n_1_211));
endmodule

module full_adder__4_338(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_334(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_339(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_338 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_334 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_328(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
endmodule

module ripple_adder_2bit__4_329(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   full_adder__4_328 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout());
endmodule

module full_adder__4_319(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in0), .B(in1), .ZN(sum));
endmodule

module ripple_adder_2bit__4_320(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   full_adder__4_319 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout());
endmodule

module mux2X1__4_311(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_330(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire [1:0]s0;
   wire [1:0]s1;

   ripple_adder_2bit__4_329 ra0 (.in0({uc_0, in0[0]}), .in1({uc_1, in1[0]}), 
      .cin(), .sum({uc_2, s0[0]}), .cout());
   ripple_adder_2bit__4_320 ra1 (.in0({uc_3, in0[0]}), .in1({uc_4, in1[0]}), 
      .cin(), .sum({uc_5, s1[0]}), .cout());
   mux2X1__4_311 ms0 (.in0({uc_6, s0[0]}), .in1({uc_7, s1[0]}), .sel(cin), 
      .out({uc_8, sum[0]}));
endmodule

module carry_select_adder_16bit__4_340(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [15:0]in0;
   input [15:0]in1;
   input cin;
   output [15:0]sum;
   output cout;
   output v;

   wire c;

   ripple_adder_2bit__4_339 ra0 (.in0({in0[1], in0[0]}), .in1({n_1, n_0}), .cin(), 
      .sum({sum[1], sum[0]}), .cout(c));
   carry_select_adder_2bit__4_330 csa0 (.in0({uc_0, in0[2]}), .in1({uc_1, n_2}), 
      .cin(c), .sum({uc_2, sum[2]}), .cout());
   INV_X1 i_10 (.A(in1[0]), .ZN(n_0));
   INV_X1 i_11 (.A(in1[1]), .ZN(n_1));
   INV_X1 i_12 (.A(in1[2]), .ZN(n_2));
endmodule

module full_adder__4_519(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_515(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_520(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_519 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_515 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_509(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_505(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_510(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_509 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_505 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_500(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_496(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_501(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_500 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_496 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module mux2X1__4_492(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module mux2X1__parameterized0__4_490(in0, in1, sel, out);
   input [0:0]in0;
   input [0:0]in1;
   input sel;
   output [0:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_511(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;
   wire [1:0]s0;
   wire c1;
   wire [1:0]s1;

   ripple_adder_2bit__4_510 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), 
      .cout(c0));
   ripple_adder_2bit__4_501 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), 
      .cout(c1));
   mux2X1__4_492 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
   mux2X1__parameterized0__4_490 mc0 (.in0(c0), .in1(c1), .sel(cin), .out(cout));
endmodule

module full_adder__4_486(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_482(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_487(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_486 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_482 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_477(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_473(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_478(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_477 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_473 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module mux2X1__4_469(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module mux2X1__parameterized0__4_467(in0, in1, sel, out);
   input [0:0]in0;
   input [0:0]in1;
   input sel;
   output [0:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_488(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;
   wire [1:0]s0;
   wire c1;
   wire [1:0]s1;

   ripple_adder_2bit__4_487 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), 
      .cout(c0));
   ripple_adder_2bit__4_478 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), 
      .cout(c1));
   mux2X1__4_469 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
   mux2X1__parameterized0__4_467 mc0 (.in0(c0), .in1(c1), .sel(cin), .out(cout));
endmodule

module full_adder__4_463(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_459(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_464(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_463 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_459 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_454(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_450(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_455(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_454 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_450 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module mux2X1__4_446(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module mux2X1__parameterized0__4_444(in0, in1, sel, out);
   input [0:0]in0;
   input [0:0]in1;
   input sel;
   output [0:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_465(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;
   wire [1:0]s0;
   wire c1;
   wire [1:0]s1;

   ripple_adder_2bit__4_464 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), 
      .cout(c0));
   ripple_adder_2bit__4_455 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), 
      .cout(c1));
   mux2X1__4_446 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
   mux2X1__parameterized0__4_444 mc0 (.in0(c0), .in1(c1), .sel(cin), .out(cout));
endmodule

module full_adder__4_440(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_436(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_441(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_440 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_436 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_431(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_427(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_432(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_431 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_427 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module mux2X1__4_423(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module mux2X1__parameterized0__4_421(in0, in1, sel, out);
   input [0:0]in0;
   input [0:0]in1;
   input sel;
   output [0:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_442(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;
   wire [1:0]s0;
   wire c1;
   wire [1:0]s1;

   ripple_adder_2bit__4_441 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), 
      .cout(c0));
   ripple_adder_2bit__4_432 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), 
      .cout(c1));
   mux2X1__4_423 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
   mux2X1__parameterized0__4_421 mc0 (.in0(c0), .in1(c1), .sel(cin), .out(cout));
endmodule

module full_adder__4_417(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_413(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_418(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_417 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_413 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_408(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_404(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_409(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_408 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_404 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module mux2X1__4_400(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module mux2X1__parameterized0__4_398(in0, in1, sel, out);
   input [0:0]in0;
   input [0:0]in1;
   input sel;
   output [0:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_419(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;
   wire [1:0]s0;
   wire c1;
   wire [1:0]s1;

   ripple_adder_2bit__4_418 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), 
      .cout(c0));
   ripple_adder_2bit__4_409 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), 
      .cout(c1));
   mux2X1__4_400 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
   mux2X1__parameterized0__4_398 mc0 (.in0(c0), .in1(c1), .sel(cin), .out(cout));
endmodule

module full_adder__4_394(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_390(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_395(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_394 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_390 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_385(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_381(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_386(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_385 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_381 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module mux2X1__4_377(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module mux2X1__parameterized0__4_375(in0, in1, sel, out);
   input [0:0]in0;
   input [0:0]in1;
   input sel;
   output [0:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_396(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;
   wire [1:0]s0;
   wire c1;
   wire [1:0]s1;

   ripple_adder_2bit__4_395 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), 
      .cout(c0));
   ripple_adder_2bit__4_386 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), 
      .cout(c1));
   mux2X1__4_377 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
   mux2X1__parameterized0__4_375 mc0 (.in0(c0), .in1(c1), .sel(cin), .out(cout));
endmodule

module full_adder__4_371(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_367(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(cin), .Z(sum));
endmodule

module ripple_adder_2bit__4_372(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_371 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_367 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout());
endmodule

module full_adder__4_362(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_358(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(cin), .Z(sum));
endmodule

module ripple_adder_2bit__4_363(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_362 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_358 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout());
endmodule

module mux2X1__4_354(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module carry_select_adder_2bit__4_373(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire [1:0]s0;
   wire [1:0]s1;

   ripple_adder_2bit__4_372 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), .cout());
   ripple_adder_2bit__4_363 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), .cout());
   mux2X1__4_354 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
endmodule

module carry_select_adder_16bit__4_521(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [15:0]in0;
   input [15:0]in1;
   input cin;
   output [15:0]sum;
   output cout;
   output v;

   wire c;

   ripple_adder_2bit__4_520 ra0 (.in0({in0[1], in0[0]}), .in1({in1[1], in1[0]}), 
      .cin(), .sum({sum[1], sum[0]}), .cout(c));
   carry_select_adder_2bit__4_511 csa0 (.in0({in0[3], in0[2]}), .in1({in1[3], 
      in1[2]}), .cin(c), .sum({sum[3], sum[2]}), .cout(n_0));
   carry_select_adder_2bit__4_488 csa1 (.in0({in0[5], in0[4]}), .in1({in1[5], 
      in1[4]}), .cin(n_0), .sum({sum[5], sum[4]}), .cout(n_1));
   carry_select_adder_2bit__4_465 csa2 (.in0({in0[7], in0[6]}), .in1({in1[7], 
      in1[6]}), .cin(n_1), .sum({sum[7], sum[6]}), .cout(n_2));
   carry_select_adder_2bit__4_442 csa3 (.in0({in0[9], in0[8]}), .in1({in1[9], 
      in1[8]}), .cin(n_2), .sum({sum[9], sum[8]}), .cout(n_3));
   carry_select_adder_2bit__4_419 csa4 (.in0({in0[11], in0[10]}), .in1({in1[11], 
      in1[10]}), .cin(n_3), .sum({sum[11], sum[10]}), .cout(n_4));
   carry_select_adder_2bit__4_396 csa5 (.in0({in0[13], in0[12]}), .in1({in1[13], 
      in1[12]}), .cin(n_4), .sum({sum[13], sum[12]}), .cout(n_5));
   carry_select_adder_2bit__4_373 csa6 (.in0({in0[15], in0[14]}), .in1({in1[15], 
      in1[14]}), .cin(n_5), .sum({sum[15], sum[14]}), .cout());
endmodule

module full_adder__4_700(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_696(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_701(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_700 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_696 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_690(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_686(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_691(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_690 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_686 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_681(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_677(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_682(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_681 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_677 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module mux2X1__4_673(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module mux2X1__parameterized0__4_671(in0, in1, sel, out);
   input [0:0]in0;
   input [0:0]in1;
   input sel;
   output [0:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_692(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;
   wire [1:0]s0;
   wire c1;
   wire [1:0]s1;

   ripple_adder_2bit__4_691 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), 
      .cout(c0));
   ripple_adder_2bit__4_682 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), 
      .cout(c1));
   mux2X1__4_673 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
   mux2X1__parameterized0__4_671 mc0 (.in0(c0), .in1(c1), .sel(cin), .out(cout));
endmodule

module full_adder__4_667(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_663(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_668(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_667 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_663 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_658(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_654(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_659(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_658 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_654 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module mux2X1__4_650(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module mux2X1__parameterized0__4_648(in0, in1, sel, out);
   input [0:0]in0;
   input [0:0]in1;
   input sel;
   output [0:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_669(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;
   wire [1:0]s0;
   wire c1;
   wire [1:0]s1;

   ripple_adder_2bit__4_668 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), 
      .cout(c0));
   ripple_adder_2bit__4_659 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), 
      .cout(c1));
   mux2X1__4_650 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
   mux2X1__parameterized0__4_648 mc0 (.in0(c0), .in1(c1), .sel(cin), .out(cout));
endmodule

module full_adder__4_644(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_640(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_645(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_644 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_640 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_635(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_631(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_636(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_635 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_631 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module mux2X1__4_627(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module mux2X1__parameterized0__4_625(in0, in1, sel, out);
   input [0:0]in0;
   input [0:0]in1;
   input sel;
   output [0:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_646(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;
   wire [1:0]s0;
   wire c1;
   wire [1:0]s1;

   ripple_adder_2bit__4_645 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), 
      .cout(c0));
   ripple_adder_2bit__4_636 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), 
      .cout(c1));
   mux2X1__4_627 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
   mux2X1__parameterized0__4_625 mc0 (.in0(c0), .in1(c1), .sel(cin), .out(cout));
endmodule

module full_adder__4_621(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_617(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_622(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_621 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_617 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_612(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_608(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_613(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_612 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_608 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module mux2X1__4_604(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module mux2X1__parameterized0__4_602(in0, in1, sel, out);
   input [0:0]in0;
   input [0:0]in1;
   input sel;
   output [0:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_623(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;
   wire [1:0]s0;
   wire c1;
   wire [1:0]s1;

   ripple_adder_2bit__4_622 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), 
      .cout(c0));
   ripple_adder_2bit__4_613 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), 
      .cout(c1));
   mux2X1__4_604 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
   mux2X1__parameterized0__4_602 mc0 (.in0(c0), .in1(c1), .sel(cin), .out(cout));
endmodule

module full_adder__4_598(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_594(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_599(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_598 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_594 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_589(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_585(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_590(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_589 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_585 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module mux2X1__4_581(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module mux2X1__parameterized0__4_579(in0, in1, sel, out);
   input [0:0]in0;
   input [0:0]in1;
   input sel;
   output [0:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_600(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;
   wire [1:0]s0;
   wire c1;
   wire [1:0]s1;

   ripple_adder_2bit__4_599 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), 
      .cout(c0));
   ripple_adder_2bit__4_590 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), 
      .cout(c1));
   mux2X1__4_581 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
   mux2X1__parameterized0__4_579 mc0 (.in0(c0), .in1(c1), .sel(cin), .out(cout));
endmodule

module full_adder__4_575(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_571(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_576(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_575 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_571 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module full_adder__4_566(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_562(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit__4_567(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_566 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_562 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout(cout));
endmodule

module mux2X1__4_558(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module mux2X1__parameterized0__4_556(in0, in1, sel, out);
   input [0:0]in0;
   input [0:0]in1;
   input sel;
   output [0:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_577(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;
   wire [1:0]s0;
   wire c1;
   wire [1:0]s1;

   ripple_adder_2bit__4_576 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), 
      .cout(c0));
   ripple_adder_2bit__4_567 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), 
      .cout(c1));
   mux2X1__4_558 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
   mux2X1__parameterized0__4_556 mc0 (.in0(c0), .in1(c1), .sel(cin), .out(cout));
endmodule

module full_adder__4_552(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
   AND2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_548(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(cin), .Z(sum));
endmodule

module ripple_adder_2bit__4_553(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_552 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_548 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout());
endmodule

module full_adder__4_543(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder__4_539(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(cin), .Z(sum));
endmodule

module ripple_adder_2bit__4_544(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_543 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder__4_539 fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), 
      .cout());
endmodule

module mux2X1__4_535(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
   MUX2_X1 i_0_1 (.A(in0[1]), .B(in1[1]), .S(sel), .Z(out[1]));
endmodule

module carry_select_adder_2bit__4_554(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire [1:0]s0;
   wire [1:0]s1;

   ripple_adder_2bit__4_553 ra0 (.in0(in0), .in1(in1), .cin(), .sum(s0), .cout());
   ripple_adder_2bit__4_544 ra1 (.in0(in0), .in1(in1), .cin(), .sum(s1), .cout());
   mux2X1__4_535 ms0 (.in0(s0), .in1(s1), .sel(cin), .out(sum));
endmodule

module carry_select_adder_16bit__4_702(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [15:0]in0;
   input [15:0]in1;
   input cin;
   output [15:0]sum;
   output cout;
   output v;

   wire c;

   ripple_adder_2bit__4_701 ra0 (.in0({in0[1], in0[0]}), .in1({in1[1], in1[0]}), 
      .cin(), .sum({sum[1], sum[0]}), .cout(c));
   carry_select_adder_2bit__4_692 csa0 (.in0({in0[3], in0[2]}), .in1({in1[3], 
      in1[2]}), .cin(c), .sum({sum[3], sum[2]}), .cout(n_0));
   carry_select_adder_2bit__4_669 csa1 (.in0({in0[5], in0[4]}), .in1({in1[5], 
      in1[4]}), .cin(n_0), .sum({sum[5], sum[4]}), .cout(n_1));
   carry_select_adder_2bit__4_646 csa2 (.in0({in0[7], in0[6]}), .in1({in1[7], 
      in1[6]}), .cin(n_1), .sum({sum[7], sum[6]}), .cout(n_2));
   carry_select_adder_2bit__4_623 csa3 (.in0({in0[9], in0[8]}), .in1({in1[9], 
      in1[8]}), .cin(n_2), .sum({sum[9], sum[8]}), .cout(n_3));
   carry_select_adder_2bit__4_600 csa4 (.in0({in0[11], in0[10]}), .in1({in1[11], 
      in1[10]}), .cin(n_3), .sum({sum[11], sum[10]}), .cout(n_4));
   carry_select_adder_2bit__4_577 csa5 (.in0({in0[13], in0[12]}), .in1({in1[13], 
      in1[12]}), .cin(n_4), .sum({sum[13], sum[12]}), .cout(n_5));
   carry_select_adder_2bit__4_554 csa6 (.in0({in0[15], in0[14]}), .in1({in1[15], 
      in1[14]}), .cin(n_5), .sum({sum[15], sum[14]}), .cout());
endmodule

module full_adder__4_3(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in1), .B(in0), .ZN(sum));
   OR2_X1 i_0_1 (.A1(in1), .A2(in0), .ZN(cout));
endmodule

module full_adder(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(sum));
   AOI22_X1 i_0_2 (.A1(in0), .A2(in1), .B1(cin), .B2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module ripple_adder_2bit(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire c0;

   full_adder__4_3 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), 
      .cout(c0));
   full_adder fa1 (.in0(in0[1]), .in1(in1[1]), .cin(c0), .sum(sum[1]), .cout(
      cout));
endmodule

module full_adder__4_42(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XOR2_X1 i_0_0 (.A(in0), .B(in1), .Z(sum));
endmodule

module ripple_adder_2bit__4_43(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   full_adder__4_42 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), .cout());
endmodule

module full_adder__4_33(in0, in1, cin, sum, cout);
   input in0;
   input in1;
   input cin;
   output sum;
   output cout;

   XNOR2_X1 i_0_0 (.A(in0), .B(in1), .ZN(sum));
endmodule

module ripple_adder_2bit__4_34(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   full_adder__4_33 fa0 (.in0(in0[0]), .in1(in1[0]), .cin(), .sum(sum[0]), .cout());
endmodule

module mux2X1__4_25(in0, in1, sel, out);
   input [1:0]in0;
   input [1:0]in1;
   input sel;
   output [1:0]out;

   MUX2_X1 i_0_0 (.A(in0[0]), .B(in1[0]), .S(sel), .Z(out[0]));
endmodule

module carry_select_adder_2bit__4_44(in0, in1, cin, sum, cout);
   input [1:0]in0;
   input [1:0]in1;
   input cin;
   output [1:0]sum;
   output cout;

   wire [1:0]s0;
   wire [1:0]s1;

   ripple_adder_2bit__4_43 ra0 (.in0({uc_0, in0[0]}), .in1({uc_1, in1[0]}), 
      .cin(), .sum({uc_2, s0[0]}), .cout());
   ripple_adder_2bit__4_34 ra1 (.in0({uc_3, in0[0]}), .in1({uc_4, in1[0]}), 
      .cin(), .sum({uc_5, s1[0]}), .cout());
   mux2X1__4_25 ms0 (.in0({uc_6, s0[0]}), .in1({uc_7, s1[0]}), .sel(cin), 
      .out({uc_8, sum[0]}));
endmodule

module carry_select_adder_16bit(sub, in0, in1, cin, sum, cout, v);
   input sub;
   input [15:0]in0;
   input [15:0]in1;
   input cin;
   output [15:0]sum;
   output cout;
   output v;

   wire c;

   ripple_adder_2bit ra0 (.in0({in0[1], in0[0]}), .in1({n_1, n_0}), .cin(), 
      .sum({sum[1], sum[0]}), .cout(c));
   carry_select_adder_2bit__4_44 csa0 (.in0({uc_0, in0[2]}), .in1({uc_1, n_2}), 
      .cin(c), .sum({uc_2, sum[2]}), .cout());
   INV_X1 i_10 (.A(in1[0]), .ZN(n_0));
   INV_X1 i_11 (.A(in1[1]), .ZN(n_1));
   INV_X1 i_12 (.A(in1[2]), .ZN(n_2));
endmodule

module Division_CSA(reset, clk, dividend, divisor, Q, ready, overFlow, 
      divideByZero);
   input reset;
   input clk;
   input [15:0]dividend;
   input [15:0]divisor;
   output [15:0]Q;
   output ready;
   output overFlow;
   output divideByZero;

   wire [15:0]sum3;
   wire [15:0]sum2;
   wire [15:0]negated_second_operand_number;
   wire [15:0]second_operand_number;
   wire [4:0]number_of_bits_in_dividend;
   wire sign;
   wire n_0_0__0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_90;
   wire n_0_91;
   wire n_0_93;
   wire n_0_97;
   wire n_0_98;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_141;
   wire n_0_142;
   wire n_0_147;
   wire n_0_148;
   wire n_0_152;
   wire n_0_153;
   wire n_0_157;
   wire n_0_158;
   wire n_0_162;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_50;
   wire n_0_160;
   wire n_0_161;
   wire n_0_154;
   wire n_0_146;
   wire n_0_145;
   wire n_0_138;
   wire n_0_100;
   wire n_0_99;
   wire n_0_0__1;
   wire n_0_51;
   wire n_0_52;
   wire n_0_89;
   wire n_0_92;
   wire n_0_95;
   wire n_0_164;
   wire n_0_165;
   wire n_0_96;
   wire n_0_159;
   wire n_0_150;
   wire n_0_151;
   wire n_0_101;
   wire n_0_134;
   wire n_0_135;
   wire n_0_166;
   wire n_0_167;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_163;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_155;
   wire n_0_156;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_149;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_143;
   wire n_0_144;
   wire n_0_332;
   wire n_0_139;
   wire n_0_140;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_137;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_53;
   wire n_0_342;
   wire n_0_136;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_83;
   wire n_0_82;
   wire n_0_60;
   wire n_0_347;
   wire n_0_94;
   wire n_0_348;
   wire n_0_88;
   wire n_0_349;
   wire n_0_87;

   carry_select_adder_16bit__4_340 csa0 (.sub(), .in0({uc_0, uc_1, uc_2, uc_3, 
      uc_4, uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, dividend[15], 
      dividend[14], dividend[13]}), .in1({uc_13, uc_14, uc_15, uc_16, uc_17, 
      uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, divisor[15], 
      divisor[14], divisor[13]}), .cin(), .sum({uc_26, uc_27, uc_28, uc_29, 
      uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, n_8, n_7, 
      n_5}), .cout(), .v());
   carry_select_adder_16bit__4_521 csa3 (.sub(), .in0({n_12, n_13, n_14, n_15, 
      n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_2}), 
      .in1({second_operand_number[15], second_operand_number[14], 
      second_operand_number[13], second_operand_number[12], 
      second_operand_number[11], second_operand_number[10], 
      second_operand_number[9], second_operand_number[8], 
      second_operand_number[7], second_operand_number[6], 
      second_operand_number[5], second_operand_number[4], 
      second_operand_number[3], second_operand_number[2], 
      second_operand_number[1], negated_second_operand_number[0]}), .cin(), 
      .sum(sum3), .cout(), .v());
   carry_select_adder_16bit__4_702 csa2 (.sub(), .in0({n_12, n_13, n_14, n_15, 
      n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_2}), 
      .in1(negated_second_operand_number), .cin(), .sum(sum2), .cout(), .v());
   carry_select_adder_16bit csa1 (.sub(), .in0({uc_39, uc_40, uc_41, uc_42, 
      uc_43, uc_44, uc_45, uc_46, uc_47, uc_48, uc_49, uc_50, uc_51, divisor[15], 
      divisor[14], divisor[13]}), .in1({uc_52, uc_53, uc_54, uc_55, uc_56, uc_57, 
      uc_58, uc_59, uc_60, uc_61, uc_62, uc_63, uc_64, dividend[15], 
      dividend[14], dividend[13]}), .cin(), .sum({uc_65, uc_66, uc_67, uc_68, 
      uc_69, uc_70, uc_71, uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, n_11, n_10, 
      n_9}), .cout(), .v());
   DFF_X1 divideByZero_reg (.D(n_116), .CK(n_6), .Q(divideByZero), .QN());
   DFF_X1 overFlow_reg (.D(n_133), .CK(clk), .Q(overFlow), .QN());
   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_96), .SE(1'b0), .GCK(n_0));
   DFF_X1 \Q_reg[14]  (.D(n_0_0__1), .CK(n_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_55), .CK(n_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_54), .CK(n_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_53), .CK(n_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_52), .CK(n_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_51), .CK(n_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_50), .CK(n_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_49), .CK(n_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_48), .CK(n_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_47), .CK(n_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_46), .CK(n_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_45), .CK(n_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_44), .CK(n_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_43), .CK(n_0), .Q(Q[0]), .QN());
   CLKGATETST_X1 clk_gate_A_reg (.CK(clk), .E(n_94), .SE(1'b0), .GCK(n_1));
   DFF_X1 \A_reg[31]  (.D(n_93), .CK(n_1), .Q(n_12), .QN());
   DFF_X1 \A_reg[30]  (.D(n_92), .CK(n_1), .Q(n_13), .QN());
   DFF_X1 \A_reg[29]  (.D(n_91), .CK(n_1), .Q(n_14), .QN());
   DFF_X1 \A_reg[28]  (.D(n_90), .CK(n_1), .Q(n_15), .QN());
   DFF_X1 \A_reg[27]  (.D(n_89), .CK(n_1), .Q(n_16), .QN());
   DFF_X1 \A_reg[26]  (.D(n_88), .CK(n_1), .Q(n_17), .QN());
   DFF_X1 \A_reg[25]  (.D(n_87), .CK(n_1), .Q(n_18), .QN());
   DFF_X1 \A_reg[24]  (.D(n_86), .CK(n_1), .Q(n_19), .QN());
   DFF_X1 \A_reg[23]  (.D(n_85), .CK(n_1), .Q(n_20), .QN());
   DFF_X1 \A_reg[22]  (.D(n_84), .CK(n_1), .Q(n_21), .QN());
   DFF_X1 \A_reg[21]  (.D(n_83), .CK(n_1), .Q(n_22), .QN());
   DFF_X1 \A_reg[20]  (.D(n_82), .CK(n_1), .Q(n_23), .QN());
   DFF_X1 \A_reg[19]  (.D(n_81), .CK(n_1), .Q(n_24), .QN());
   DFF_X1 \A_reg[18]  (.D(n_80), .CK(n_1), .Q(n_25), .QN());
   DFF_X1 \A_reg[17]  (.D(n_79), .CK(n_1), .Q(n_26), .QN());
   DFF_X1 \A_reg[16]  (.D(n_78), .CK(n_1), .Q(n_2), .QN());
   CLKGATETST_X1 clk_gate_A_reg__15 (.CK(clk), .E(n_95), .SE(1'b0), .GCK(n_3));
   DFF_X1 \A_reg[15]  (.D(n_77), .CK(n_3), .Q(n_27), .QN());
   DFF_X1 \A_reg[14]  (.D(n_76), .CK(n_3), .Q(n_28), .QN());
   DFF_X1 \A_reg[13]  (.D(n_75), .CK(n_3), .Q(n_29), .QN());
   DFF_X1 \A_reg[12]  (.D(n_74), .CK(n_3), .Q(n_30), .QN());
   DFF_X1 \A_reg[11]  (.D(n_73), .CK(n_3), .Q(n_31), .QN());
   DFF_X1 \A_reg[10]  (.D(n_72), .CK(n_3), .Q(n_32), .QN());
   DFF_X1 \A_reg[9]  (.D(n_71), .CK(n_3), .Q(n_33), .QN());
   DFF_X1 \A_reg[8]  (.D(n_70), .CK(n_3), .Q(n_34), .QN());
   DFF_X1 \A_reg[7]  (.D(n_69), .CK(n_3), .Q(n_35), .QN());
   DFF_X1 \A_reg[6]  (.D(n_68), .CK(n_3), .Q(n_36), .QN());
   DFF_X1 \A_reg[5]  (.D(n_67), .CK(n_3), .Q(n_37), .QN());
   DFF_X1 \A_reg[4]  (.D(n_66), .CK(n_3), .Q(n_38), .QN());
   DFF_X1 \A_reg[3]  (.D(n_65), .CK(n_3), .Q(n_39), .QN());
   DFF_X1 \A_reg[2]  (.D(n_64), .CK(n_3), .Q(n_40), .QN());
   DFF_X1 \A_reg[1]  (.D(n_63), .CK(n_3), .Q(n_41), .QN());
   DFF_X1 \A_reg[0]  (.D(n_62), .CK(n_3), .Q(n_42), .QN());
   DFF_X1 \negated_second_operand_number_reg[15]  (.D(n_125), .CK(n_6), .Q(
      negated_second_operand_number[15]), .QN());
   DFF_X1 \negated_second_operand_number_reg[14]  (.D(n_114), .CK(n_6), .Q(
      negated_second_operand_number[14]), .QN());
   DFF_X1 \negated_second_operand_number_reg[13]  (.D(n_113), .CK(n_6), .Q(
      negated_second_operand_number[13]), .QN());
   DFF_X1 \negated_second_operand_number_reg[12]  (.D(n_112), .CK(n_6), .Q(
      negated_second_operand_number[12]), .QN());
   DFF_X1 \negated_second_operand_number_reg[11]  (.D(n_111), .CK(n_6), .Q(
      negated_second_operand_number[11]), .QN());
   DFF_X1 \negated_second_operand_number_reg[10]  (.D(n_110), .CK(n_6), .Q(
      negated_second_operand_number[10]), .QN());
   DFF_X1 \negated_second_operand_number_reg[9]  (.D(n_109), .CK(n_6), .Q(
      negated_second_operand_number[9]), .QN());
   DFF_X1 \negated_second_operand_number_reg[8]  (.D(n_108), .CK(n_6), .Q(
      negated_second_operand_number[8]), .QN());
   DFF_X1 \negated_second_operand_number_reg[7]  (.D(n_107), .CK(n_6), .Q(
      negated_second_operand_number[7]), .QN());
   DFF_X1 \negated_second_operand_number_reg[6]  (.D(n_106), .CK(n_6), .Q(
      negated_second_operand_number[6]), .QN());
   DFF_X1 \negated_second_operand_number_reg[5]  (.D(n_105), .CK(n_6), .Q(
      negated_second_operand_number[5]), .QN());
   DFF_X1 \negated_second_operand_number_reg[4]  (.D(n_104), .CK(n_6), .Q(
      negated_second_operand_number[4]), .QN());
   DFF_X1 \negated_second_operand_number_reg[3]  (.D(n_103), .CK(n_6), .Q(
      negated_second_operand_number[3]), .QN());
   DFF_X1 \negated_second_operand_number_reg[2]  (.D(n_102), .CK(n_6), .Q(
      negated_second_operand_number[2]), .QN());
   DFF_X1 \negated_second_operand_number_reg[1]  (.D(n_100), .CK(n_6), .Q(
      negated_second_operand_number[1]), .QN());
   DFF_X1 \second_operand_number_reg[15]  (.D(n_126), .CK(n_6), .Q(
      second_operand_number[15]), .QN());
   DFF_X1 \second_operand_number_reg[14]  (.D(n_124), .CK(n_6), .Q(
      second_operand_number[14]), .QN());
   DFF_X1 \second_operand_number_reg[13]  (.D(n_123), .CK(n_6), .Q(
      second_operand_number[13]), .QN());
   DFF_X1 \second_operand_number_reg[12]  (.D(n_127), .CK(n_6), .Q(
      second_operand_number[12]), .QN());
   DFF_X1 \second_operand_number_reg[11]  (.D(n_128), .CK(n_6), .Q(
      second_operand_number[11]), .QN());
   DFF_X1 \second_operand_number_reg[10]  (.D(n_129), .CK(n_6), .Q(
      second_operand_number[10]), .QN());
   DFF_X1 \second_operand_number_reg[9]  (.D(n_122), .CK(n_6), .Q(
      second_operand_number[9]), .QN());
   DFF_X1 \second_operand_number_reg[8]  (.D(n_130), .CK(n_6), .Q(
      second_operand_number[8]), .QN());
   DFF_X1 \second_operand_number_reg[7]  (.D(n_131), .CK(n_6), .Q(
      second_operand_number[7]), .QN());
   DFF_X1 \second_operand_number_reg[6]  (.D(n_121), .CK(n_6), .Q(
      second_operand_number[6]), .QN());
   DFF_X1 \second_operand_number_reg[5]  (.D(n_132), .CK(n_6), .Q(
      second_operand_number[5]), .QN());
   DFF_X1 \second_operand_number_reg[4]  (.D(n_120), .CK(n_6), .Q(
      second_operand_number[4]), .QN());
   DFF_X1 \second_operand_number_reg[3]  (.D(n_119), .CK(n_6), .Q(
      second_operand_number[3]), .QN());
   DFF_X1 \second_operand_number_reg[2]  (.D(n_101), .CK(n_6), .Q(
      second_operand_number[2]), .QN());
   DFF_X1 \second_operand_number_reg[1]  (.D(n_118), .CK(n_6), .Q(
      second_operand_number[1]), .QN());
   DFF_X1 ready_reg (.D(n_134), .CK(clk), .Q(ready), .QN());
   CLKGATETST_X1 clk_gate_number_of_bits_in_dividend_reg (.CK(clk), .E(n_61), 
      .SE(1'b0), .GCK(n_4));
   DFF_X1 \number_of_bits_in_dividend_reg[4]  (.D(n_115), .CK(n_4), .Q(
      number_of_bits_in_dividend[4]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[3]  (.D(n_60), .CK(n_4), .Q(
      number_of_bits_in_dividend[3]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[2]  (.D(n_59), .CK(n_4), .Q(
      number_of_bits_in_dividend[2]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[1]  (.D(n_58), .CK(n_4), .Q(
      number_of_bits_in_dividend[1]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[0]  (.D(n_57), .CK(n_4), .Q(
      number_of_bits_in_dividend[0]), .QN());
   DFF_X1 sign_reg (.D(n_56), .CK(n_6), .Q(sign), .QN());
   CLKGATETST_X1 clk_gate_divideByZero_reg (.CK(clk), .E(reset), .SE(1'b0), 
      .GCK(n_6));
   DFF_X1 \negated_second_operand_number_reg[0]  (.D(n_117), .CK(n_6), .Q(
      negated_second_operand_number[0]), .QN());
   INV_X1 i_0_1 (.A(n_42), .ZN(n_0_0__0));
   NOR2_X1 i_0_2 (.A1(n_0_0__0), .A2(reset), .ZN(n_43));
   NAND2_X1 i_0_3 (.A1(sign), .A2(n_42), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_41), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_1), .A2(n_0_2), .ZN(n_0_3));
   OAI21_X1 i_0_6 (.A(n_0_3), .B1(n_0_2), .B2(n_0_1), .ZN(n_0_4));
   NOR2_X1 i_0_7 (.A1(n_0_4), .A2(reset), .ZN(n_44));
   NAND2_X1 i_0_8 (.A1(n_0_3), .A2(sign), .ZN(n_0_5));
   XOR2_X1 i_0_9 (.A(n_0_5), .B(n_40), .Z(n_0_6));
   NOR2_X1 i_0_10 (.A1(n_0_6), .A2(reset), .ZN(n_45));
   INV_X1 i_0_11 (.A(sign), .ZN(n_0_7));
   INV_X1 i_0_12 (.A(n_40), .ZN(n_0_8));
   AOI21_X1 i_0_13 (.A(n_0_7), .B1(n_0_5), .B2(n_0_8), .ZN(n_0_9));
   XNOR2_X1 i_0_14 (.A(n_0_9), .B(n_39), .ZN(n_0_10));
   NOR2_X1 i_0_15 (.A1(n_0_10), .A2(reset), .ZN(n_46));
   OAI21_X1 i_0_16 (.A(sign), .B1(n_0_9), .B2(n_39), .ZN(n_0_11));
   XOR2_X1 i_0_17 (.A(n_0_11), .B(n_38), .Z(n_0_12));
   NOR2_X1 i_0_18 (.A1(n_0_12), .A2(reset), .ZN(n_47));
   INV_X1 i_0_19 (.A(n_38), .ZN(n_0_13));
   AOI21_X1 i_0_20 (.A(n_0_7), .B1(n_0_11), .B2(n_0_13), .ZN(n_0_14));
   XNOR2_X1 i_0_21 (.A(n_0_14), .B(n_37), .ZN(n_0_15));
   NOR2_X1 i_0_22 (.A1(n_0_15), .A2(reset), .ZN(n_48));
   OAI21_X1 i_0_23 (.A(sign), .B1(n_0_14), .B2(n_37), .ZN(n_0_16));
   XOR2_X1 i_0_24 (.A(n_0_16), .B(n_36), .Z(n_0_17));
   NOR2_X1 i_0_25 (.A1(n_0_17), .A2(reset), .ZN(n_49));
   INV_X1 i_0_26 (.A(n_36), .ZN(n_0_18));
   AOI21_X1 i_0_27 (.A(n_0_7), .B1(n_0_16), .B2(n_0_18), .ZN(n_0_19));
   XNOR2_X1 i_0_28 (.A(n_0_19), .B(n_35), .ZN(n_0_20));
   NOR2_X1 i_0_29 (.A1(n_0_20), .A2(reset), .ZN(n_50));
   OAI21_X1 i_0_30 (.A(sign), .B1(n_0_19), .B2(n_35), .ZN(n_0_21));
   XOR2_X1 i_0_31 (.A(n_0_21), .B(n_34), .Z(n_0_22));
   NOR2_X1 i_0_32 (.A1(n_0_22), .A2(reset), .ZN(n_51));
   INV_X1 i_0_33 (.A(n_34), .ZN(n_0_23));
   AOI21_X1 i_0_34 (.A(n_0_7), .B1(n_0_21), .B2(n_0_23), .ZN(n_0_24));
   XNOR2_X1 i_0_35 (.A(n_0_24), .B(n_33), .ZN(n_0_25));
   NOR2_X1 i_0_36 (.A1(n_0_25), .A2(reset), .ZN(n_52));
   OAI21_X1 i_0_37 (.A(sign), .B1(n_0_24), .B2(n_33), .ZN(n_0_26));
   XOR2_X1 i_0_38 (.A(n_0_26), .B(n_32), .Z(n_0_27));
   NOR2_X1 i_0_39 (.A1(n_0_27), .A2(reset), .ZN(n_53));
   INV_X1 i_0_40 (.A(n_32), .ZN(n_0_28));
   AOI21_X1 i_0_41 (.A(n_0_7), .B1(n_0_26), .B2(n_0_28), .ZN(n_0_29));
   XNOR2_X1 i_0_42 (.A(n_0_29), .B(n_31), .ZN(n_0_30));
   NOR2_X1 i_0_43 (.A1(n_0_30), .A2(reset), .ZN(n_54));
   OAI21_X1 i_0_44 (.A(sign), .B1(n_0_29), .B2(n_31), .ZN(n_0_31));
   XOR2_X1 i_0_45 (.A(n_0_31), .B(n_30), .Z(n_0_32));
   NOR2_X1 i_0_46 (.A1(n_0_32), .A2(reset), .ZN(n_55));
   INV_X1 i_0_47 (.A(dividend[12]), .ZN(n_0_33));
   INV_X1 i_0_48 (.A(divisor[12]), .ZN(n_0_34));
   OAI22_X1 i_0_49 (.A1(n_0_33), .A2(divisor[12]), .B1(n_0_34), .B2(dividend[12]), 
      .ZN(n_56));
   NAND2_X1 i_0_50 (.A1(n_0_0__1), .A2(number_of_bits_in_dividend[0]), .ZN(n_57));
   NOR2_X1 i_0_51 (.A1(number_of_bits_in_dividend[1]), .A2(
      number_of_bits_in_dividend[0]), .ZN(n_0_35));
   INV_X1 i_0_52 (.A(n_0_35), .ZN(n_0_36));
   AOI21_X1 i_0_53 (.A(reset), .B1(number_of_bits_in_dividend[1]), .B2(
      number_of_bits_in_dividend[0]), .ZN(n_0_37));
   NAND2_X1 i_0_54 (.A1(n_0_36), .A2(n_0_37), .ZN(n_58));
   NOR3_X1 i_0_55 (.A1(number_of_bits_in_dividend[1]), .A2(
      number_of_bits_in_dividend[0]), .A3(number_of_bits_in_dividend[2]), 
      .ZN(n_0_38));
   INV_X1 i_0_56 (.A(n_0_38), .ZN(n_0_39));
   INV_X1 i_0_57 (.A(number_of_bits_in_dividend[2]), .ZN(n_0_40));
   OAI211_X1 i_0_58 (.A(n_0_39), .B(n_0_0__1), .C1(n_0_35), .C2(n_0_40), 
      .ZN(n_59));
   INV_X1 i_0_59 (.A(number_of_bits_in_dividend[3]), .ZN(n_0_41));
   NAND2_X1 i_0_60 (.A1(n_0_38), .A2(n_0_41), .ZN(n_0_42));
   OAI211_X1 i_0_61 (.A(n_0_42), .B(n_0_0__1), .C1(n_0_38), .C2(n_0_41), 
      .ZN(n_60));
   INV_X1 i_0_62 (.A(dividend[15]), .ZN(n_0_43));
   INV_X1 i_0_63 (.A(dividend[14]), .ZN(n_0_44));
   AOI22_X1 i_0_64 (.A1(n_0_43), .A2(divisor[15]), .B1(n_0_44), .B2(divisor[14]), 
      .ZN(n_0_45));
   INV_X1 i_0_65 (.A(dividend[13]), .ZN(n_0_46));
   OAI22_X1 i_0_66 (.A1(n_0_44), .A2(divisor[14]), .B1(n_0_46), .B2(divisor[13]), 
      .ZN(n_0_47));
   INV_X1 i_0_67 (.A(divisor[15]), .ZN(n_0_48));
   AOI22_X1 i_0_68 (.A1(n_0_45), .A2(n_0_47), .B1(n_0_48), .B2(dividend[15]), 
      .ZN(n_0_49));
   OR2_X1 i_0_73 (.A1(divisor[1]), .A2(divisor[0]), .ZN(n_0_54));
   OR3_X1 i_0_74 (.A1(n_0_54), .A2(divisor[2]), .A3(divisor[3]), .ZN(n_0_55));
   OR4_X1 i_0_75 (.A1(n_0_55), .A2(divisor[5]), .A3(divisor[6]), .A4(divisor[4]), 
      .ZN(n_0_56));
   OR3_X1 i_0_76 (.A1(n_0_56), .A2(divisor[7]), .A3(divisor[8]), .ZN(n_0_57));
   OAI21_X1 i_0_77 (.A(divisor[12]), .B1(n_0_57), .B2(divisor[9]), .ZN(n_0_58));
   XNOR2_X1 i_0_78 (.A(n_0_58), .B(divisor[10]), .ZN(n_0_59));
   OR2_X1 i_0_80 (.A1(n_0_55), .A2(divisor[4]), .ZN(n_0_61));
   OAI21_X1 i_0_81 (.A(divisor[12]), .B1(n_0_61), .B2(divisor[5]), .ZN(n_0_62));
   XNOR2_X1 i_0_82 (.A(n_0_62), .B(divisor[6]), .ZN(n_0_63));
   AOI22_X1 i_0_83 (.A1(n_0_59), .A2(n_0_60), .B1(n_0_63), .B2(n_8), .ZN(n_0_64));
   OAI21_X1 i_0_84 (.A(divisor[12]), .B1(n_0_56), .B2(divisor[7]), .ZN(n_0_65));
   XNOR2_X1 i_0_85 (.A(n_0_65), .B(divisor[8]), .ZN(n_0_66));
   NOR3_X1 i_0_86 (.A1(n_0_57), .A2(divisor[9]), .A3(divisor[10]), .ZN(n_0_67));
   INV_X1 i_0_87 (.A(divisor[11]), .ZN(n_0_68));
   NAND3_X1 i_0_88 (.A1(n_0_67), .A2(n_0_68), .A3(divisor[12]), .ZN(n_0_69));
   INV_X1 i_0_89 (.A(n_0_69), .ZN(n_0_70));
   OAI22_X1 i_0_90 (.A1(n_0_66), .A2(n_0_60), .B1(n_0_70), .B2(n_8), .ZN(n_0_71));
   INV_X1 i_0_91 (.A(n_7), .ZN(n_0_72));
   AOI22_X1 i_0_92 (.A1(n_0_64), .A2(n_7), .B1(n_0_71), .B2(n_0_72), .ZN(n_0_73));
   INV_X1 i_0_93 (.A(n_0_73), .ZN(n_0_74));
   NAND2_X1 i_0_94 (.A1(n_0_56), .A2(divisor[12]), .ZN(n_0_75));
   XNOR2_X1 i_0_95 (.A(n_0_75), .B(divisor[7]), .ZN(n_0_76));
   INV_X1 i_0_96 (.A(n_0_76), .ZN(n_0_77));
   NAND2_X1 i_0_97 (.A1(n_0_57), .A2(divisor[12]), .ZN(n_0_78));
   XNOR2_X1 i_0_98 (.A(n_0_78), .B(divisor[9]), .ZN(n_0_79));
   INV_X1 i_0_99 (.A(n_0_79), .ZN(n_0_80));
   AOI221_X1 i_0_100 (.A(n_0_60), .B1(n_0_77), .B2(n_7), .C1(n_0_80), .C2(n_0_72), 
      .ZN(n_0_81));
   NOR2_X1 i_0_103 (.A1(n_0_67), .A2(n_0_34), .ZN(n_0_84));
   XOR2_X1 i_0_104 (.A(n_0_84), .B(divisor[11]), .Z(n_0_85));
   AOI21_X1 i_0_105 (.A(n_0_81), .B1(n_0_83), .B2(n_0_85), .ZN(n_0_86));
   NAND2_X1 i_0_110 (.A1(divisor[12]), .A2(divisor[0]), .ZN(n_0_90));
   XNOR2_X1 i_0_111 (.A(n_0_90), .B(divisor[1]), .ZN(n_0_91));
   NAND2_X1 i_0_115 (.A1(n_0_54), .A2(divisor[12]), .ZN(n_0_93));
   OAI21_X1 i_0_119 (.A(divisor[12]), .B1(n_0_54), .B2(divisor[2]), .ZN(n_0_97));
   XNOR2_X1 i_0_120 (.A(n_0_97), .B(divisor[3]), .ZN(n_0_98));
   NAND2_X1 i_0_125 (.A1(n_0_55), .A2(divisor[12]), .ZN(n_0_102));
   XNOR2_X1 i_0_126 (.A(n_0_102), .B(divisor[4]), .ZN(n_0_103));
   AOI22_X1 i_0_127 (.A1(n_0_103), .A2(n_0_60), .B1(divisor[0]), .B2(n_8), 
      .ZN(n_0_104));
   INV_X1 i_0_128 (.A(n_0_94), .ZN(n_0_105));
   OAI22_X1 i_0_129 (.A1(n_0_104), .A2(n_7), .B1(n_0_105), .B2(n_0_82), .ZN(
      n_0_106));
   NAND2_X1 i_0_130 (.A1(n_0_61), .A2(divisor[12]), .ZN(n_0_107));
   XNOR2_X1 i_0_131 (.A(n_0_107), .B(divisor[5]), .ZN(n_0_108));
   OAI22_X1 i_0_132 (.A1(n_0_108), .A2(n_8), .B1(n_0_60), .B2(n_0_91), .ZN(
      n_0_109));
   OAI22_X1 i_0_133 (.A1(n_0_109), .A2(n_7), .B1(n_0_82), .B2(n_0_99), .ZN(
      n_0_110));
   OAI221_X1 i_0_134 (.A(n_0_88), .B1(n_0_87), .B2(n_0_106), .C1(n_0_110), 
      .C2(n_5), .ZN(n_0_111));
   INV_X1 i_0_135 (.A(n_0_108), .ZN(n_0_112));
   OAI22_X1 i_0_137 (.A1(n_0_76), .A2(n_8), .B1(n_0_98), .B2(n_0_60), .ZN(
      n_0_113));
   OAI22_X1 i_0_138 (.A1(n_0_113), .A2(n_7), .B1(n_0_109), .B2(n_0_72), .ZN(
      n_0_114));
   OAI22_X1 i_0_139 (.A1(n_0_63), .A2(n_8), .B1(n_0_94), .B2(n_0_60), .ZN(
      n_0_115));
   AOI22_X1 i_0_140 (.A1(n_0_115), .A2(n_0_72), .B1(n_0_104), .B2(n_7), .ZN(
      n_0_116));
   OAI221_X1 i_0_141 (.A(n_0_88), .B1(n_0_114), .B2(n_5), .C1(n_0_116), .C2(
      n_0_87), .ZN(n_0_117));
   AOI22_X1 i_0_143 (.A1(n_0_66), .A2(n_0_60), .B1(n_0_103), .B2(n_8), .ZN(
      n_0_118));
   OAI22_X1 i_0_144 (.A1(n_0_118), .A2(n_7), .B1(n_0_115), .B2(n_0_72), .ZN(
      n_0_119));
   AOI22_X1 i_0_145 (.A1(n_0_79), .A2(n_0_60), .B1(n_0_108), .B2(n_8), .ZN(
      n_0_120));
   OAI22_X1 i_0_146 (.A1(n_0_120), .A2(n_7), .B1(n_0_113), .B2(n_0_72), .ZN(
      n_0_121));
   AOI221_X1 i_0_147 (.A(n_0_53), .B1(n_0_119), .B2(n_5), .C1(n_0_121), .C2(
      n_0_87), .ZN(n_0_122));
   AOI22_X1 i_0_149 (.A1(n_0_64), .A2(n_0_72), .B1(n_0_118), .B2(n_7), .ZN(
      n_0_123));
   OAI221_X1 i_0_150 (.A(n_0_72), .B1(n_0_76), .B2(n_0_60), .C1(n_0_85), 
      .C2(n_8), .ZN(n_0_124));
   OAI21_X1 i_0_151 (.A(n_0_124), .B1(n_0_72), .B2(n_0_120), .ZN(n_0_125));
   OAI221_X1 i_0_152 (.A(n_0_88), .B1(n_0_87), .B2(n_0_123), .C1(n_0_125), 
      .C2(n_5), .ZN(n_0_126));
   INV_X1 i_0_153 (.A(n_0_85), .ZN(n_0_127));
   AOI21_X1 i_0_155 (.A(n_7), .B1(n_0_59), .B2(n_8), .ZN(n_0_128));
   AOI21_X1 i_0_156 (.A(n_0_128), .B1(n_7), .B2(n_0_71), .ZN(n_0_129));
   OAI21_X1 i_0_157 (.A(n_0_88), .B1(n_0_129), .B2(n_5), .ZN(n_0_130));
   NAND2_X1 i_0_159 (.A1(n_0_129), .A2(n_5), .ZN(n_0_131));
   AOI21_X1 i_0_160 (.A(n_5), .B1(n_0_80), .B2(n_7), .ZN(n_0_132));
   OAI211_X1 i_0_161 (.A(n_0_132), .B(n_8), .C1(n_0_85), .C2(n_7), .ZN(n_0_133));
   OAI221_X1 i_0_170 (.A(n_0_88), .B1(n_0_100), .B2(n_0_87), .C1(n_0_106), 
      .C2(n_5), .ZN(n_0_141));
   INV_X1 i_0_171 (.A(n_0_103), .ZN(n_0_142));
   OAI22_X1 i_0_177 (.A1(n_0_116), .A2(n_5), .B1(n_0_110), .B2(n_0_87), .ZN(
      n_0_147));
   INV_X1 i_0_178 (.A(n_0_63), .ZN(n_0_148));
   OAI221_X1 i_0_183 (.A(n_0_88), .B1(n_0_114), .B2(n_0_87), .C1(n_0_119), 
      .C2(n_5), .ZN(n_0_152));
   INV_X1 i_0_184 (.A(n_0_66), .ZN(n_0_153));
   OAI221_X1 i_0_189 (.A(n_0_88), .B1(n_0_121), .B2(n_0_87), .C1(n_0_123), 
      .C2(n_5), .ZN(n_0_157));
   INV_X1 i_0_190 (.A(n_0_59), .ZN(n_0_158));
   OAI221_X1 i_0_195 (.A(n_0_88), .B1(n_5), .B2(n_0_73), .C1(n_0_125), .C2(
      n_0_87), .ZN(n_0_162));
   AND3_X1 i_0_204 (.A1(number_of_bits_in_dividend[1]), .A2(
      number_of_bits_in_dividend[0]), .A3(number_of_bits_in_dividend[3]), 
      .ZN(n_0_168));
   AND3_X1 i_0_205 (.A1(n_0_168), .A2(number_of_bits_in_dividend[4]), .A3(
      number_of_bits_in_dividend[2]), .ZN(n_0_169));
   AND2_X1 i_0_206 (.A1(n_0_169), .A2(n_0_0__1), .ZN(n_0_170));
   INV_X1 i_0_207 (.A(n_0_170), .ZN(n_61));
   NOR2_X1 i_0_208 (.A1(n_0_169), .A2(reset), .ZN(n_0_171));
   INV_X1 i_0_209 (.A(n_0_171), .ZN(n_0_172));
   NOR2_X1 i_0_210 (.A1(n_0_172), .A2(n_12), .ZN(n_0_173));
   INV_X1 i_0_211 (.A(n_0_173), .ZN(n_0_174));
   NOR2_X1 i_0_212 (.A1(n_0_174), .A2(sum2[15]), .ZN(n_0_175));
   NOR2_X1 i_0_213 (.A1(n_61), .A2(ready), .ZN(n_0_176));
   NOR4_X1 i_0_214 (.A1(n_30), .A2(n_29), .A3(n_28), .A4(n_27), .ZN(n_0_177));
   NAND2_X1 i_0_215 (.A1(n_0_176), .A2(n_0_177), .ZN(n_0_178));
   INV_X1 i_0_216 (.A(n_0_178), .ZN(n_0_179));
   AOI21_X1 i_0_217 (.A(n_0_175), .B1(n_0_179), .B2(n_42), .ZN(n_0_180));
   NAND2_X1 i_0_218 (.A1(n_0_171), .A2(n_12), .ZN(n_0_181));
   OAI21_X1 i_0_219 (.A(n_0_180), .B1(sum3[15]), .B2(n_0_181), .ZN(n_62));
   OAI22_X1 i_0_220 (.A1(n_0_178), .A2(n_0_4), .B1(n_0_172), .B2(n_0_0__0), 
      .ZN(n_63));
   OAI22_X1 i_0_221 (.A1(n_0_178), .A2(n_0_6), .B1(n_0_2), .B2(n_0_172), 
      .ZN(n_64));
   OAI22_X1 i_0_222 (.A1(n_0_178), .A2(n_0_10), .B1(n_0_172), .B2(n_0_8), 
      .ZN(n_65));
   NOR2_X1 i_0_223 (.A1(n_11), .A2(n_10), .ZN(n_0_182));
   INV_X1 i_0_224 (.A(n_0_182), .ZN(n_0_183));
   OAI21_X1 i_0_225 (.A(n_0_49), .B1(n_9), .B2(n_0_183), .ZN(n_0_184));
   NAND3_X1 i_0_226 (.A1(n_0_184), .A2(dividend[0]), .A3(reset), .ZN(n_0_185));
   INV_X1 i_0_227 (.A(n_39), .ZN(n_0_186));
   OAI221_X1 i_0_228 (.A(n_0_185), .B1(n_0_186), .B2(n_0_172), .C1(n_0_12), 
      .C2(n_0_178), .ZN(n_66));
   NAND2_X1 i_0_229 (.A1(dividend[0]), .A2(dividend[12]), .ZN(n_0_187));
   XNOR2_X1 i_0_230 (.A(n_0_187), .B(dividend[1]), .ZN(n_0_188));
   INV_X1 i_0_231 (.A(dividend[0]), .ZN(n_0_189));
   INV_X1 i_0_232 (.A(n_9), .ZN(n_0_190));
   NOR3_X1 i_0_233 (.A1(n_0_183), .A2(n_0_189), .A3(n_0_190), .ZN(n_0_191));
   AOI22_X1 i_0_234 (.A1(n_0_184), .A2(n_0_188), .B1(n_0_49), .B2(n_0_191), 
      .ZN(n_0_192));
   OAI222_X1 i_0_235 (.A1(n_0_15), .A2(n_0_178), .B1(n_0_192), .B2(n_0_0__1), 
      .C1(n_0_13), .C2(n_0_172), .ZN(n_67));
   INV_X1 i_0_236 (.A(n_0_184), .ZN(n_0_193));
   INV_X1 i_0_237 (.A(n_0_188), .ZN(n_0_194));
   OR2_X1 i_0_238 (.A1(dividend[1]), .A2(dividend[0]), .ZN(n_0_195));
   NAND2_X1 i_0_239 (.A1(n_0_195), .A2(dividend[12]), .ZN(n_0_196));
   XNOR2_X1 i_0_240 (.A(n_0_196), .B(dividend[2]), .ZN(n_0_197));
   INV_X1 i_0_241 (.A(n_0_197), .ZN(n_0_198));
   INV_X1 i_0_242 (.A(n_10), .ZN(n_0_199));
   AOI22_X1 i_0_243 (.A1(n_0_198), .A2(n_0_199), .B1(n_0_189), .B2(n_10), 
      .ZN(n_0_200));
   INV_X1 i_0_244 (.A(n_11), .ZN(n_0_201));
   NAND2_X1 i_0_245 (.A1(n_0_200), .A2(n_0_201), .ZN(n_0_202));
   OAI221_X1 i_0_246 (.A(n_0_193), .B1(n_0_194), .B2(n_0_183), .C1(n_0_202), 
      .C2(n_9), .ZN(n_0_203));
   OAI211_X1 i_0_247 (.A(n_0_203), .B(reset), .C1(n_0_193), .C2(n_0_197), 
      .ZN(n_0_204));
   INV_X1 i_0_248 (.A(n_37), .ZN(n_0_205));
   OAI221_X1 i_0_249 (.A(n_0_204), .B1(n_0_205), .B2(n_0_172), .C1(n_0_178), 
      .C2(n_0_17), .ZN(n_68));
   OAI21_X1 i_0_250 (.A(dividend[12]), .B1(n_0_195), .B2(dividend[2]), .ZN(
      n_0_206));
   XNOR2_X1 i_0_251 (.A(n_0_206), .B(dividend[3]), .ZN(n_0_207));
   NAND2_X1 i_0_252 (.A1(n_0_201), .A2(n_10), .ZN(n_0_208));
   INV_X1 i_0_253 (.A(n_0_208), .ZN(n_0_209));
   AOI22_X1 i_0_254 (.A1(n_0_207), .A2(n_0_182), .B1(n_0_209), .B2(n_0_188), 
      .ZN(n_0_210));
   OAI221_X1 i_0_255 (.A(n_0_193), .B1(n_9), .B2(n_0_210), .C1(n_0_202), 
      .C2(n_0_190), .ZN(n_0_211));
   OAI211_X1 i_0_256 (.A(n_0_211), .B(reset), .C1(n_0_193), .C2(n_0_207), 
      .ZN(n_0_212));
   OAI221_X1 i_0_257 (.A(n_0_212), .B1(n_0_18), .B2(n_0_172), .C1(n_0_178), 
      .C2(n_0_20), .ZN(n_69));
   OR4_X1 i_0_258 (.A1(dividend[1]), .A2(dividend[0]), .A3(dividend[2]), 
      .A4(dividend[3]), .ZN(n_0_213));
   NAND2_X1 i_0_259 (.A1(n_0_213), .A2(dividend[12]), .ZN(n_0_214));
   XNOR2_X1 i_0_260 (.A(n_0_214), .B(dividend[4]), .ZN(n_0_215));
   INV_X1 i_0_261 (.A(n_0_215), .ZN(n_0_216));
   OAI22_X1 i_0_262 (.A1(n_0_216), .A2(n_0_183), .B1(n_0_198), .B2(n_0_208), 
      .ZN(n_0_217));
   NOR2_X1 i_0_263 (.A1(n_0_201), .A2(n_10), .ZN(n_0_218));
   AOI21_X1 i_0_264 (.A(n_0_217), .B1(dividend[0]), .B2(n_0_218), .ZN(n_0_219));
   OAI221_X1 i_0_265 (.A(n_0_193), .B1(n_0_210), .B2(n_0_190), .C1(n_0_219), 
      .C2(n_9), .ZN(n_0_220));
   OAI211_X1 i_0_266 (.A(n_0_220), .B(reset), .C1(n_0_193), .C2(n_0_215), 
      .ZN(n_0_221));
   INV_X1 i_0_267 (.A(n_35), .ZN(n_0_222));
   OAI221_X1 i_0_268 (.A(n_0_221), .B1(n_0_222), .B2(n_0_172), .C1(n_0_22), 
      .C2(n_0_178), .ZN(n_70));
   OAI21_X1 i_0_269 (.A(dividend[12]), .B1(n_0_213), .B2(dividend[4]), .ZN(
      n_0_223));
   XNOR2_X1 i_0_270 (.A(n_0_223), .B(dividend[5]), .ZN(n_0_224));
   INV_X1 i_0_271 (.A(n_0_224), .ZN(n_0_225));
   OAI22_X1 i_0_272 (.A1(n_0_225), .A2(n_11), .B1(n_0_194), .B2(n_0_201), 
      .ZN(n_0_226));
   AOI22_X1 i_0_273 (.A1(n_0_226), .A2(n_0_199), .B1(n_0_209), .B2(n_0_207), 
      .ZN(n_0_227));
   AOI22_X1 i_0_274 (.A1(n_0_227), .A2(n_0_190), .B1(n_0_219), .B2(n_9), 
      .ZN(n_0_228));
   OAI221_X1 i_0_275 (.A(reset), .B1(n_0_224), .B2(n_0_193), .C1(n_0_228), 
      .C2(n_0_184), .ZN(n_0_229));
   OAI221_X1 i_0_276 (.A(n_0_229), .B1(n_0_23), .B2(n_0_172), .C1(n_0_25), 
      .C2(n_0_178), .ZN(n_71));
   OR3_X1 i_0_277 (.A1(n_0_213), .A2(dividend[4]), .A3(dividend[5]), .ZN(n_0_230));
   NAND2_X1 i_0_278 (.A1(n_0_230), .A2(dividend[12]), .ZN(n_0_231));
   XNOR2_X1 i_0_279 (.A(n_0_231), .B(dividend[6]), .ZN(n_0_232));
   OAI222_X1 i_0_280 (.A1(n_0_232), .A2(n_0_183), .B1(n_0_200), .B2(n_0_201), 
      .C1(n_0_208), .C2(n_0_215), .ZN(n_0_233));
   OAI221_X1 i_0_281 (.A(n_0_193), .B1(n_0_190), .B2(n_0_227), .C1(n_0_233), 
      .C2(n_9), .ZN(n_0_234));
   OAI211_X1 i_0_282 (.A(n_0_234), .B(reset), .C1(n_0_193), .C2(n_0_232), 
      .ZN(n_0_235));
   INV_X1 i_0_283 (.A(n_33), .ZN(n_0_236));
   OAI221_X1 i_0_284 (.A(n_0_235), .B1(n_0_236), .B2(n_0_172), .C1(n_0_27), 
      .C2(n_0_178), .ZN(n_72));
   OR2_X1 i_0_285 (.A1(n_0_230), .A2(dividend[6]), .ZN(n_0_237));
   NAND2_X1 i_0_286 (.A1(n_0_237), .A2(dividend[12]), .ZN(n_0_238));
   XNOR2_X1 i_0_287 (.A(n_0_238), .B(dividend[7]), .ZN(n_0_239));
   AOI22_X1 i_0_288 (.A1(n_0_239), .A2(n_0_201), .B1(n_11), .B2(n_0_207), 
      .ZN(n_0_240));
   INV_X1 i_0_289 (.A(n_0_240), .ZN(n_0_241));
   OAI22_X1 i_0_290 (.A1(n_0_241), .A2(n_10), .B1(n_0_226), .B2(n_0_199), 
      .ZN(n_0_242));
   AOI22_X1 i_0_291 (.A1(n_0_233), .A2(n_9), .B1(n_0_242), .B2(n_0_190), 
      .ZN(n_0_243));
   OAI221_X1 i_0_292 (.A(reset), .B1(n_0_239), .B2(n_0_193), .C1(n_0_243), 
      .C2(n_0_184), .ZN(n_0_244));
   OAI221_X1 i_0_293 (.A(n_0_244), .B1(n_0_28), .B2(n_0_172), .C1(n_0_30), 
      .C2(n_0_178), .ZN(n_73));
   OAI221_X1 i_0_294 (.A(n_10), .B1(n_0_197), .B2(n_0_201), .C1(n_0_232), 
      .C2(n_11), .ZN(n_0_245));
   OAI21_X1 i_0_295 (.A(dividend[12]), .B1(n_0_237), .B2(dividend[7]), .ZN(
      n_0_246));
   XNOR2_X1 i_0_296 (.A(n_0_246), .B(dividend[8]), .ZN(n_0_247));
   OAI22_X1 i_0_297 (.A1(n_0_247), .A2(n_11), .B1(n_0_215), .B2(n_0_201), 
      .ZN(n_0_248));
   OAI21_X1 i_0_298 (.A(n_0_245), .B1(n_10), .B2(n_0_248), .ZN(n_0_249));
   INV_X1 i_0_299 (.A(n_0_249), .ZN(n_0_250));
   OAI221_X1 i_0_300 (.A(n_0_193), .B1(n_0_190), .B2(n_0_242), .C1(n_0_250), 
      .C2(n_9), .ZN(n_0_251));
   OAI211_X1 i_0_301 (.A(n_0_251), .B(reset), .C1(n_0_193), .C2(n_0_247), 
      .ZN(n_0_252));
   INV_X1 i_0_302 (.A(n_31), .ZN(n_0_253));
   OAI221_X1 i_0_303 (.A(n_0_252), .B1(n_0_253), .B2(n_0_172), .C1(n_0_32), 
      .C2(n_0_178), .ZN(n_74));
   OR4_X1 i_0_304 (.A1(n_0_230), .A2(dividend[6]), .A3(dividend[7]), .A4(
      dividend[8]), .ZN(n_0_254));
   NAND2_X1 i_0_305 (.A1(n_0_254), .A2(dividend[12]), .ZN(n_0_255));
   XNOR2_X1 i_0_306 (.A(n_0_255), .B(dividend[9]), .ZN(n_0_256));
   OAI22_X1 i_0_307 (.A1(n_0_256), .A2(n_11), .B1(n_0_224), .B2(n_0_201), 
      .ZN(n_0_257));
   AOI22_X1 i_0_308 (.A1(n_0_257), .A2(n_0_199), .B1(n_0_240), .B2(n_10), 
      .ZN(n_0_258));
   OAI221_X1 i_0_309 (.A(n_0_193), .B1(n_0_258), .B2(n_9), .C1(n_0_249), 
      .C2(n_0_190), .ZN(n_0_259));
   INV_X1 i_0_310 (.A(n_0_256), .ZN(n_0_260));
   OAI21_X1 i_0_311 (.A(n_0_259), .B1(n_0_193), .B2(n_0_260), .ZN(n_0_261));
   AOI22_X1 i_0_312 (.A1(n_0_261), .A2(reset), .B1(n_30), .B2(n_0_171), .ZN(
      n_0_262));
   NAND2_X1 i_0_313 (.A1(n_0_262), .A2(n_0_178), .ZN(n_75));
   INV_X1 i_0_314 (.A(n_29), .ZN(n_0_263));
   OAI21_X1 i_0_315 (.A(dividend[12]), .B1(n_0_254), .B2(dividend[9]), .ZN(
      n_0_264));
   XNOR2_X1 i_0_316 (.A(n_0_264), .B(dividend[10]), .ZN(n_0_265));
   AOI22_X1 i_0_317 (.A1(n_0_265), .A2(n_0_201), .B1(n_0_232), .B2(n_11), 
      .ZN(n_0_266));
   OAI22_X1 i_0_318 (.A1(n_0_266), .A2(n_10), .B1(n_0_248), .B2(n_0_199), 
      .ZN(n_0_267));
   AOI221_X1 i_0_319 (.A(n_0_184), .B1(n_0_258), .B2(n_9), .C1(n_0_267), 
      .C2(n_0_190), .ZN(n_0_268));
   OAI21_X1 i_0_320 (.A(reset), .B1(n_0_265), .B2(n_0_193), .ZN(n_0_269));
   OAI221_X1 i_0_321 (.A(n_0_178), .B1(n_0_172), .B2(n_0_263), .C1(n_0_268), 
      .C2(n_0_269), .ZN(n_76));
   INV_X1 i_0_322 (.A(n_0_267), .ZN(n_0_270));
   OR3_X1 i_0_323 (.A1(n_0_254), .A2(dividend[9]), .A3(dividend[10]), .ZN(
      n_0_271));
   NAND2_X1 i_0_324 (.A1(n_0_271), .A2(dividend[12]), .ZN(n_0_272));
   XNOR2_X1 i_0_325 (.A(n_0_272), .B(dividend[11]), .ZN(n_0_273));
   INV_X1 i_0_326 (.A(n_0_257), .ZN(n_0_274));
   AOI222_X1 i_0_327 (.A1(n_0_273), .A2(n_0_182), .B1(n_0_274), .B2(n_10), 
      .C1(n_0_239), .C2(n_0_218), .ZN(n_0_275));
   AOI221_X1 i_0_328 (.A(n_0_184), .B1(n_9), .B2(n_0_270), .C1(n_0_275), 
      .C2(n_0_190), .ZN(n_0_276));
   AOI21_X1 i_0_329 (.A(n_0_276), .B1(n_0_184), .B2(n_0_273), .ZN(n_0_277));
   INV_X1 i_0_330 (.A(n_28), .ZN(n_0_278));
   OAI22_X1 i_0_331 (.A1(n_0_277), .A2(n_0_0__1), .B1(n_0_172), .B2(n_0_278), 
      .ZN(n_77));
   NAND2_X1 i_0_332 (.A1(n_0_176), .A2(n_26), .ZN(n_0_279));
   INV_X1 i_0_333 (.A(n_27), .ZN(n_0_280));
   NOR4_X1 i_0_334 (.A1(n_0_271), .A2(n_0_193), .A3(dividend[11]), .A4(n_0_33), 
      .ZN(n_0_281));
   INV_X1 i_0_335 (.A(n_0_266), .ZN(n_0_282));
   AOI22_X1 i_0_336 (.A1(n_0_282), .A2(n_10), .B1(n_0_247), .B2(n_0_218), 
      .ZN(n_0_283));
   OAI22_X1 i_0_337 (.A1(n_0_275), .A2(n_0_190), .B1(n_0_283), .B2(n_9), 
      .ZN(n_0_284));
   AOI21_X1 i_0_338 (.A(n_0_281), .B1(n_0_284), .B2(n_0_193), .ZN(n_0_285));
   OAI221_X1 i_0_339 (.A(n_0_279), .B1(n_0_280), .B2(n_0_172), .C1(n_0_285), 
      .C2(n_0_0__1), .ZN(n_78));
   INV_X1 i_0_340 (.A(n_0_181), .ZN(n_0_286));
   AOI222_X1 i_0_341 (.A1(n_0_176), .A2(n_25), .B1(n_0_286), .B2(sum3[0]), 
      .C1(n_0_173), .C2(sum2[0]), .ZN(n_0_287));
   INV_X1 i_0_342 (.A(n_0_287), .ZN(n_79));
   AOI222_X1 i_0_343 (.A1(n_0_176), .A2(n_24), .B1(n_0_286), .B2(sum3[1]), 
      .C1(n_0_173), .C2(sum2[1]), .ZN(n_0_288));
   INV_X1 i_0_344 (.A(n_0_288), .ZN(n_80));
   AOI222_X1 i_0_345 (.A1(n_0_176), .A2(n_23), .B1(n_0_286), .B2(sum3[2]), 
      .C1(n_0_173), .C2(sum2[2]), .ZN(n_0_289));
   INV_X1 i_0_346 (.A(n_0_289), .ZN(n_81));
   AOI222_X1 i_0_347 (.A1(n_0_176), .A2(n_22), .B1(n_0_286), .B2(sum3[3]), 
      .C1(n_0_173), .C2(sum2[3]), .ZN(n_0_290));
   INV_X1 i_0_348 (.A(n_0_290), .ZN(n_82));
   AOI222_X1 i_0_349 (.A1(n_0_176), .A2(n_21), .B1(n_0_286), .B2(sum3[4]), 
      .C1(n_0_173), .C2(sum2[4]), .ZN(n_0_291));
   INV_X1 i_0_350 (.A(n_0_291), .ZN(n_83));
   AOI222_X1 i_0_351 (.A1(n_0_176), .A2(n_20), .B1(n_0_286), .B2(sum3[5]), 
      .C1(n_0_173), .C2(sum2[5]), .ZN(n_0_292));
   INV_X1 i_0_352 (.A(n_0_292), .ZN(n_84));
   AOI222_X1 i_0_353 (.A1(n_0_176), .A2(n_19), .B1(n_0_286), .B2(sum3[6]), 
      .C1(n_0_173), .C2(sum2[6]), .ZN(n_0_293));
   INV_X1 i_0_354 (.A(n_0_293), .ZN(n_85));
   AOI222_X1 i_0_355 (.A1(n_0_176), .A2(n_18), .B1(n_0_286), .B2(sum3[7]), 
      .C1(n_0_173), .C2(sum2[7]), .ZN(n_0_294));
   INV_X1 i_0_356 (.A(n_0_294), .ZN(n_86));
   AOI222_X1 i_0_357 (.A1(n_0_176), .A2(n_17), .B1(n_0_286), .B2(sum3[8]), 
      .C1(n_0_173), .C2(sum2[8]), .ZN(n_0_295));
   INV_X1 i_0_358 (.A(n_0_295), .ZN(n_87));
   AOI222_X1 i_0_359 (.A1(n_0_176), .A2(n_16), .B1(n_0_286), .B2(sum3[9]), 
      .C1(n_0_173), .C2(sum2[9]), .ZN(n_0_296));
   INV_X1 i_0_360 (.A(n_0_296), .ZN(n_88));
   AOI222_X1 i_0_361 (.A1(n_0_176), .A2(n_15), .B1(n_0_286), .B2(sum3[10]), 
      .C1(n_0_173), .C2(sum2[10]), .ZN(n_0_297));
   INV_X1 i_0_362 (.A(n_0_297), .ZN(n_89));
   AOI222_X1 i_0_363 (.A1(n_0_176), .A2(n_14), .B1(n_0_286), .B2(sum3[11]), 
      .C1(n_0_173), .C2(sum2[11]), .ZN(n_0_298));
   INV_X1 i_0_364 (.A(n_0_298), .ZN(n_90));
   AOI222_X1 i_0_365 (.A1(n_0_176), .A2(n_13), .B1(n_0_286), .B2(sum3[12]), 
      .C1(n_0_173), .C2(sum2[12]), .ZN(n_0_299));
   INV_X1 i_0_366 (.A(n_0_299), .ZN(n_91));
   AOI222_X1 i_0_367 (.A1(n_0_176), .A2(n_12), .B1(n_0_286), .B2(sum3[13]), 
      .C1(n_0_173), .C2(sum2[13]), .ZN(n_0_300));
   INV_X1 i_0_368 (.A(n_0_300), .ZN(n_92));
   AOI22_X1 i_0_369 (.A1(n_0_286), .A2(sum3[14]), .B1(n_0_173), .B2(sum2[14]), 
      .ZN(n_0_301));
   INV_X1 i_0_370 (.A(n_0_301), .ZN(n_93));
   NAND2_X1 i_0_371 (.A1(n_0_170), .A2(ready), .ZN(n_94));
   INV_X1 i_0_372 (.A(n_94), .ZN(n_0_302));
   INV_X1 i_0_373 (.A(n_0_177), .ZN(n_0_303));
   AOI21_X1 i_0_374 (.A(n_0_302), .B1(n_0_170), .B2(n_0_303), .ZN(n_95));
   NAND2_X1 i_0_375 (.A1(n_0_178), .A2(n_0_0__1), .ZN(n_96));
   NOR2_X1 i_0_376 (.A1(n_0_177), .A2(reset), .ZN(n_97));
   INV_X1 i_0_377 (.A(n_0_176), .ZN(n_0_304));
   OAI21_X1 i_0_378 (.A(n_0_0__1), .B1(n_0_304), .B2(n_0_177), .ZN(n_98));
   NAND2_X1 i_0_379 (.A1(n_0_304), .A2(n_0_0__1), .ZN(n_99));
   AOI21_X1 i_0_380 (.A(n_0_137), .B1(n_118), .B2(n_117), .ZN(n_100));
   INV_X1 i_0_381 (.A(n_0_138), .ZN(n_0_305));
   INV_X1 i_0_382 (.A(n_0_136), .ZN(n_101));
   INV_X1 i_0_383 (.A(n_0_137), .ZN(n_0_306));
   AOI21_X1 i_0_384 (.A(n_0_305), .B1(n_101), .B2(n_0_306), .ZN(n_102));
   AOI21_X1 i_0_385 (.A(n_0_139), .B1(n_119), .B2(n_0_138), .ZN(n_103));
   AOI21_X1 i_0_386 (.A(n_0_143), .B1(n_0_140), .B2(n_120), .ZN(n_104));
   AOI21_X1 i_0_387 (.A(n_0_145), .B1(n_0_144), .B2(n_132), .ZN(n_105));
   INV_X1 i_0_388 (.A(n_0_149), .ZN(n_0_307));
   AOI21_X1 i_0_389 (.A(n_0_307), .B1(n_0_146), .B2(n_121), .ZN(n_106));
   AOI21_X1 i_0_390 (.A(n_0_150), .B1(n_0_149), .B2(n_131), .ZN(n_107));
   INV_X1 i_0_391 (.A(n_0_154), .ZN(n_0_308));
   AOI21_X1 i_0_392 (.A(n_0_308), .B1(n_0_151), .B2(n_130), .ZN(n_108));
   AOI21_X1 i_0_393 (.A(n_0_155), .B1(n_0_154), .B2(n_122), .ZN(n_109));
   INV_X1 i_0_394 (.A(n_0_159), .ZN(n_0_309));
   AOI21_X1 i_0_395 (.A(n_0_309), .B1(n_0_156), .B2(n_129), .ZN(n_110));
   AOI21_X1 i_0_396 (.A(n_0_160), .B1(n_0_159), .B2(n_128), .ZN(n_111));
   INV_X1 i_0_397 (.A(n_0_163), .ZN(n_0_310));
   AOI21_X1 i_0_398 (.A(n_0_310), .B1(n_0_161), .B2(n_127), .ZN(n_112));
   AOI21_X1 i_0_399 (.A(n_0_164), .B1(n_0_163), .B2(n_123), .ZN(n_113));
   AOI21_X1 i_0_401 (.A(n_0_311), .B1(n_0_165), .B2(n_124), .ZN(n_114));
   INV_X1 i_0_0 (.A(n_0_50), .ZN(n_0_311));
   NAND2_X1 i_0_69 (.A1(n_0_164), .A2(n_0_166), .ZN(n_0_50));
   INV_X1 i_0_70 (.A(n_0_161), .ZN(n_0_160));
   NAND2_X1 i_0_71 (.A1(n_0_96), .A2(n_0_318), .ZN(n_0_161));
   NAND2_X1 i_0_72 (.A1(n_0_150), .A2(n_0_323), .ZN(n_0_154));
   INV_X1 i_0_79 (.A(n_0_145), .ZN(n_0_146));
   NOR2_X1 i_0_101 (.A1(n_0_144), .A2(n_132), .ZN(n_0_145));
   NAND2_X1 i_0_102 (.A1(n_0_137), .A2(n_0_136), .ZN(n_0_138));
   NAND2_X1 i_0_106 (.A1(n_0_336), .A2(n_0_337), .ZN(n_0_100));
   INV_X1 i_0_107 (.A(n_0_98), .ZN(n_0_99));
   INV_X1 i_0_108 (.A(reset), .ZN(n_0_0__1));
   NAND2_X1 i_0_109 (.A1(n_0_92), .A2(n_0_51), .ZN(n_115));
   OAI21_X1 i_0_112 (.A(n_0_52), .B1(n_0_89), .B2(n_0_42), .ZN(n_0_51));
   AOI21_X1 i_0_113 (.A(reset), .B1(n_0_42), .B2(n_0_89), .ZN(n_0_52));
   INV_X1 i_0_114 (.A(number_of_bits_in_dividend[4]), .ZN(n_0_89));
   INV_X1 i_0_116 (.A(n_0_92), .ZN(n_116));
   NAND4_X1 i_0_117 (.A1(n_0_164), .A2(reset), .A3(n_0_166), .A4(n_0_135), 
      .ZN(n_0_92));
   NOR2_X1 i_0_118 (.A1(n_0_88), .A2(n_0_342), .ZN(n_117));
   NAND2_X1 i_0_121 (.A1(n_0_341), .A2(n_0_340), .ZN(n_118));
   NAND2_X1 i_0_122 (.A1(n_0_334), .A2(n_0_333), .ZN(n_119));
   NAND2_X1 i_0_123 (.A1(n_0_141), .A2(n_0_332), .ZN(n_120));
   INV_X1 i_0_124 (.A(n_0_327), .ZN(n_121));
   INV_X1 i_0_136 (.A(n_0_320), .ZN(n_122));
   INV_X1 i_0_142 (.A(n_0_313), .ZN(n_123));
   INV_X1 i_0_148 (.A(n_0_166), .ZN(n_124));
   NOR2_X1 i_0_154 (.A1(n_0_95), .A2(n_0_101), .ZN(n_125));
   AOI21_X1 i_0_158 (.A(n_0_135), .B1(n_0_164), .B2(n_0_166), .ZN(n_0_95));
   INV_X1 i_0_162 (.A(n_0_165), .ZN(n_0_164));
   NAND4_X1 i_0_163 (.A1(n_0_96), .A2(n_0_318), .A3(n_0_317), .A4(n_0_313), 
      .ZN(n_0_165));
   INV_X1 i_0_164 (.A(n_0_159), .ZN(n_0_96));
   NAND4_X1 i_0_165 (.A1(n_0_150), .A2(n_0_323), .A3(n_0_320), .A4(n_0_319), 
      .ZN(n_0_159));
   INV_X1 i_0_166 (.A(n_0_151), .ZN(n_0_150));
   NAND4_X1 i_0_167 (.A1(n_0_143), .A2(n_0_330), .A3(n_0_324), .A4(n_0_327), 
      .ZN(n_0_151));
   INV_X1 i_0_168 (.A(n_0_134), .ZN(n_0_101));
   NAND4_X1 i_0_169 (.A1(n_0_316), .A2(n_0_313), .A3(n_0_166), .A4(n_0_135), 
      .ZN(n_0_134));
   INV_X1 i_0_172 (.A(n_126), .ZN(n_0_135));
   AOI21_X1 i_0_173 (.A(n_0_53), .B1(n_0_133), .B2(n_0_131), .ZN(n_126));
   OAI21_X1 i_0_174 (.A(n_0_167), .B1(n_0_87), .B2(n_0_312), .ZN(n_0_166));
   INV_X1 i_0_175 (.A(n_0_130), .ZN(n_0_167));
   INV_X1 i_0_176 (.A(n_0_86), .ZN(n_0_312));
   OAI21_X1 i_0_179 (.A(n_0_314), .B1(n_0_315), .B2(n_0_87), .ZN(n_0_313));
   AOI21_X1 i_0_180 (.A(n_0_53), .B1(n_0_86), .B2(n_0_87), .ZN(n_0_314));
   INV_X1 i_0_181 (.A(n_0_74), .ZN(n_0_315));
   INV_X1 i_0_182 (.A(n_0_163), .ZN(n_0_316));
   NAND4_X1 i_0_185 (.A1(n_0_155), .A2(n_0_319), .A3(n_0_318), .A4(n_0_317), 
      .ZN(n_0_163));
   INV_X1 i_0_186 (.A(n_127), .ZN(n_0_317));
   OAI21_X1 i_0_187 (.A(n_0_162), .B1(n_0_69), .B2(n_0_88), .ZN(n_127));
   INV_X1 i_0_188 (.A(n_128), .ZN(n_0_318));
   OAI21_X1 i_0_191 (.A(n_0_126), .B1(n_0_127), .B2(n_0_88), .ZN(n_128));
   INV_X1 i_0_192 (.A(n_129), .ZN(n_0_319));
   OAI21_X1 i_0_193 (.A(n_0_157), .B1(n_0_158), .B2(n_0_88), .ZN(n_129));
   INV_X1 i_0_194 (.A(n_0_156), .ZN(n_0_155));
   NAND4_X1 i_0_196 (.A1(n_0_326), .A2(n_0_324), .A3(n_0_323), .A4(n_0_320), 
      .ZN(n_0_156));
   OAI21_X1 i_0_197 (.A(n_0_321), .B1(n_0_322), .B2(n_0_88), .ZN(n_0_320));
   INV_X1 i_0_198 (.A(n_0_122), .ZN(n_0_321));
   INV_X1 i_0_199 (.A(n_0_80), .ZN(n_0_322));
   INV_X1 i_0_200 (.A(n_130), .ZN(n_0_323));
   OAI21_X1 i_0_201 (.A(n_0_152), .B1(n_0_153), .B2(n_0_88), .ZN(n_130));
   INV_X1 i_0_202 (.A(n_131), .ZN(n_0_324));
   NAND2_X1 i_0_203 (.A1(n_0_117), .A2(n_0_325), .ZN(n_131));
   OR2_X1 i_0_400 (.A1(n_0_88), .A2(n_0_77), .ZN(n_0_325));
   INV_X1 i_0_402 (.A(n_0_149), .ZN(n_0_326));
   NAND3_X1 i_0_403 (.A1(n_0_143), .A2(n_0_330), .A3(n_0_327), .ZN(n_0_149));
   AOI21_X1 i_0_404 (.A(n_0_328), .B1(n_0_329), .B2(n_0_88), .ZN(n_0_327));
   NOR2_X1 i_0_405 (.A1(n_0_88), .A2(n_0_148), .ZN(n_0_328));
   INV_X1 i_0_406 (.A(n_0_147), .ZN(n_0_329));
   INV_X1 i_0_407 (.A(n_132), .ZN(n_0_330));
   NAND2_X1 i_0_408 (.A1(n_0_111), .A2(n_0_331), .ZN(n_132));
   OR2_X1 i_0_409 (.A1(n_0_88), .A2(n_0_112), .ZN(n_0_331));
   INV_X1 i_0_410 (.A(n_0_144), .ZN(n_0_143));
   NAND3_X1 i_0_411 (.A1(n_0_141), .A2(n_0_139), .A3(n_0_332), .ZN(n_0_144));
   OR2_X1 i_0_412 (.A1(n_0_88), .A2(n_0_142), .ZN(n_0_332));
   INV_X1 i_0_413 (.A(n_0_140), .ZN(n_0_139));
   NAND4_X1 i_0_414 (.A1(n_0_137), .A2(n_0_334), .A3(n_0_136), .A4(n_0_333), 
      .ZN(n_0_140));
   NAND2_X1 i_0_415 (.A1(n_0_53), .A2(n_0_98), .ZN(n_0_333));
   OAI21_X1 i_0_416 (.A(n_0_88), .B1(n_0_338), .B2(n_0_335), .ZN(n_0_334));
   AOI21_X1 i_0_417 (.A(n_5), .B1(n_0_336), .B2(n_0_337), .ZN(n_0_335));
   NAND2_X1 i_0_418 (.A1(n_0_83), .A2(n_0_91), .ZN(n_0_336));
   NAND2_X1 i_0_419 (.A1(n_0_349), .A2(n_0_98), .ZN(n_0_337));
   AOI21_X1 i_0_420 (.A(n_0_87), .B1(n_0_346), .B2(n_0_347), .ZN(n_0_338));
   INV_X1 i_0_421 (.A(n_0_339), .ZN(n_0_137));
   OAI211_X1 i_0_422 (.A(n_0_340), .B(n_0_341), .C1(n_0_342), .C2(n_0_88), 
      .ZN(n_0_339));
   NAND3_X1 i_0_423 (.A1(n_0_88), .A2(divisor[0]), .A3(n_0_349), .ZN(n_0_340));
   NAND2_X1 i_0_424 (.A1(n_0_53), .A2(n_0_91), .ZN(n_0_341));
   INV_X1 i_0_425 (.A(n_0_88), .ZN(n_0_53));
   INV_X1 i_0_426 (.A(divisor[0]), .ZN(n_0_342));
   OAI22_X1 i_0_427 (.A1(n_0_345), .A2(n_0_343), .B1(n_0_88), .B2(n_0_94), 
      .ZN(n_0_136));
   NAND2_X1 i_0_428 (.A1(n_0_344), .A2(n_0_88), .ZN(n_0_343));
   NAND3_X1 i_0_429 (.A1(n_0_349), .A2(n_5), .A3(n_0_91), .ZN(n_0_344));
   AOI21_X1 i_0_430 (.A(n_5), .B1(n_0_346), .B2(n_0_347), .ZN(n_0_345));
   NAND2_X1 i_0_431 (.A1(n_0_83), .A2(divisor[0]), .ZN(n_0_346));
   INV_X1 i_0_432 (.A(n_0_82), .ZN(n_0_83));
   NAND2_X1 i_0_433 (.A1(n_0_60), .A2(n_7), .ZN(n_0_82));
   INV_X1 i_0_434 (.A(n_8), .ZN(n_0_60));
   NAND2_X1 i_0_435 (.A1(n_0_349), .A2(n_0_94), .ZN(n_0_347));
   INV_X1 i_0_436 (.A(n_0_348), .ZN(n_0_94));
   XOR2_X1 i_0_437 (.A(divisor[2]), .B(n_0_93), .Z(n_0_348));
   AOI21_X1 i_0_438 (.A(n_0_49), .B1(n_0_349), .B2(n_0_87), .ZN(n_0_88));
   NOR2_X1 i_0_439 (.A1(n_8), .A2(n_7), .ZN(n_0_349));
   INV_X1 i_0_440 (.A(n_5), .ZN(n_0_87));
   MUX2_X1 overFlow_reg_enable_mux_0 (.A(overFlow), .B(n_97), .S(n_98), .Z(n_133));
   MUX2_X1 ready_reg_enable_mux_0 (.A(ready), .B(n_0_0__1), .S(n_99), .Z(n_134));
endmodule

module datapath__0_28(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_0 (.A(B[0]), .B(p_0[0]), .CO(n_0), .S(p_1[0]));
   FA_X1 i_1 (.A(B[1]), .B(p_0[1]), .CI(n_0), .CO(n_1), .S(p_1[1]));
   FA_X1 i_2 (.A(B[2]), .B(p_0[2]), .CI(n_1), .CO(n_2), .S(p_1[2]));
   FA_X1 i_3 (.A(B[3]), .B(p_0[3]), .CI(n_2), .CO(n_3), .S(p_1[3]));
   FA_X1 i_4 (.A(B[4]), .B(p_0[4]), .CI(n_3), .CO(n_4), .S(p_1[4]));
   FA_X1 i_5 (.A(B[5]), .B(p_0[5]), .CI(n_4), .CO(n_5), .S(p_1[5]));
   FA_X1 i_6 (.A(B[6]), .B(p_0[6]), .CI(n_5), .CO(n_6), .S(p_1[6]));
   FA_X1 i_7 (.A(B[7]), .B(p_0[7]), .CI(n_6), .CO(n_7), .S(p_1[7]));
   FA_X1 i_8 (.A(B[8]), .B(p_0[8]), .CI(n_7), .CO(n_8), .S(p_1[8]));
   FA_X1 i_9 (.A(B[9]), .B(p_0[9]), .CI(n_8), .CO(n_9), .S(p_1[9]));
   FA_X1 i_10 (.A(B[10]), .B(p_0[10]), .CI(n_9), .CO(n_10), .S(p_1[10]));
   FA_X1 i_11 (.A(B[11]), .B(p_0[11]), .CI(n_10), .CO(n_11), .S(p_1[11]));
   FA_X1 i_12 (.A(B[15]), .B(p_0[14]), .CI(n_11), .CO(n_12), .S(p_1[12]));
   FA_X1 i_13 (.A(B[15]), .B(p_0[14]), .CI(n_12), .CO(n_13), .S(p_1[13]));
   FA_X1 i_14 (.A(B[15]), .B(p_0[14]), .CI(n_13), .CO(n_14), .S(p_1[14]));
   XNOR2_X1 i_15 (.A(B[15]), .B(p_0[15]), .ZN(n_15));
   XNOR2_X1 i_16 (.A(n_15), .B(n_14), .ZN(p_1[15]));
endmodule

module datapath__0_33(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[14]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[14]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[14]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[14]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_34(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(p_0[13]), .B2(n_15), .ZN(p_2[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_2[15]));
   NAND2_X1 i_16 (.A1(p_0[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_1[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_1[14]), .ZN(n_16));
endmodule

module datapath__0_39(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[13]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[13]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_40(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(p_0[13]), .B2(n_15), .ZN(p_2[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_2[15]));
   NAND2_X1 i_16 (.A1(p_0[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_1[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_1[14]), .ZN(n_16));
endmodule

module datapath__0_45(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[12]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[12]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[12]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_46(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(p_0[13]), .B2(n_15), .ZN(p_2[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_2[15]));
   NAND2_X1 i_16 (.A1(p_0[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_1[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_1[14]), .ZN(n_16));
endmodule

module datapath__0_51(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[13]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[13]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_52(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(p_0[13]), .B2(n_15), .ZN(p_2[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_2[15]));
   NAND2_X1 i_16 (.A1(p_0[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_1[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_1[14]), .ZN(n_16));
endmodule

module datapath__0_57(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[12]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[12]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[12]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_58(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(p_0[13]), .B2(n_15), .ZN(p_2[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_2[15]));
   NAND2_X1 i_16 (.A1(p_0[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_1[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_1[14]), .ZN(n_16));
endmodule

module datapath__0_63(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[12]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[12]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[12]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_64(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(p_0[13]), .B2(n_15), .ZN(p_2[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_2[15]));
   NAND2_X1 i_16 (.A1(p_0[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_1[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_1[14]), .ZN(n_16));
endmodule

module datapath__0_69(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[13]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[13]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_70(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(p_0[13]), .B2(n_15), .ZN(p_2[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_2[15]));
   NAND2_X1 i_16 (.A1(p_0[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_1[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_1[14]), .ZN(n_16));
endmodule

module datapath__0_75(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[12]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[12]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[12]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_76(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(p_0[13]), .B2(n_15), .ZN(p_2[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_2[15]));
   NAND2_X1 i_16 (.A1(p_0[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_1[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_1[14]), .ZN(n_16));
endmodule

module datapath__0_81(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[12]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[12]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[12]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_82(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(p_0[13]), .B2(n_15), .ZN(p_2[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_2[15]));
   NAND2_X1 i_16 (.A1(p_0[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_1[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_1[14]), .ZN(n_16));
endmodule

module booth_16bit_multiplier(A, B, product);
   input [15:0]A;
   input [15:0]B;
   output [31:0]product;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_35;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_0;
   wire n_1_1;
   wire n_1_15;
   wire n_1_16;
   wire n_1_17;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;
   wire n_1_28;
   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;

   datapath__0_28 i_2 (.B({B[12], uc_0, uc_1, uc_2, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({n_468, n_481, uc_3, 
      uc_4, n_480, n_479, n_478, n_477, n_476, n_475, n_474, n_473, n_472, n_471, 
      n_470, n_469}), .p_1({n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, 
      n_6, n_5, n_4, n_3, n_2, n_1, n_0}));
   datapath__0_33 i_5 (.B({uc_5, B[12], uc_6, uc_7, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_8, n_467, n_466, 
      n_465, n_464, n_463, n_462, n_461, n_460, n_459, n_458, n_457, n_456, 
      n_455, n_454, n_453}), .p_1({n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
      n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16}));
   datapath__0_34 i_6 (.p_0({uc_9, uc_10, n_481, n_480, n_479, n_478, n_477, 
      n_476, n_475, n_474, n_473, n_472, n_471, n_470, n_469, B[0]}), .p_1({
      uc_11, n_467, n_466, n_465, n_464, n_463, n_462, n_461, n_460, n_459, 
      n_458, n_457, n_456, n_455, n_454, n_453}), .p_2({n_47, n_46, n_45, n_44, 
      n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32}));
   datapath__0_39 i_9 (.B({uc_12, uc_13, B[12], uc_14, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_15, n_452, 
      n_451, n_450, n_449, n_448, n_447, n_446, n_445, n_444, n_443, n_442, 
      n_441, n_440, n_439, n_438}), .p_1({n_63, n_62, n_61, n_60, n_59, n_58, 
      n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48}));
   datapath__0_40 i_10 (.p_0({uc_16, uc_17, n_481, n_480, n_479, n_478, n_477, 
      n_476, n_475, n_474, n_473, n_472, n_471, n_470, n_469, B[0]}), .p_1({
      uc_18, n_452, n_451, n_450, n_449, n_448, n_447, n_446, n_445, n_444, 
      n_443, n_442, n_441, n_440, n_439, n_438}), .p_2({n_79, n_78, n_77, n_76, 
      n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64}));
   datapath__0_45 i_13 (.B({uc_19, uc_20, uc_21, B[12], B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_22, n_437, 
      n_436, n_435, n_434, n_433, n_432, n_431, n_430, n_429, n_428, n_427, 
      n_426, n_425, n_424, n_423}), .p_1({n_95, n_94, n_93, n_92, n_91, n_90, 
      n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80}));
   datapath__0_46 i_14 (.p_0({uc_23, uc_24, n_481, n_480, n_479, n_478, n_477, 
      n_476, n_475, n_474, n_473, n_472, n_471, n_470, n_469, B[0]}), .p_1({
      uc_25, n_437, n_436, n_435, n_434, n_433, n_432, n_431, n_430, n_429, 
      n_428, n_427, n_426, n_425, n_424, n_423}), .p_2({n_111, n_110, n_109, 
      n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
      n_97, n_96}));
   datapath__0_51 i_17 (.B({uc_26, uc_27, B[12], uc_28, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_29, n_422, 
      n_421, n_420, n_419, n_418, n_417, n_416, n_415, n_414, n_413, n_412, 
      n_411, n_410, n_409, n_408}), .p_1({n_127, n_126, n_125, n_124, n_123, 
      n_122, n_121, n_120, n_119, n_118, n_117, n_116, n_115, n_114, n_113, 
      n_112}));
   datapath__0_52 i_18 (.p_0({uc_30, uc_31, n_481, n_480, n_479, n_478, n_477, 
      n_476, n_475, n_474, n_473, n_472, n_471, n_470, n_469, B[0]}), .p_1({
      uc_32, n_422, n_421, n_420, n_419, n_418, n_417, n_416, n_415, n_414, 
      n_413, n_412, n_411, n_410, n_409, n_408}), .p_2({n_143, n_142, n_141, 
      n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, n_132, n_131, 
      n_130, n_129, n_128}));
   datapath__0_57 i_21 (.B({uc_33, uc_34, uc_35, B[12], B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_36, n_407, 
      n_406, n_405, n_404, n_403, n_402, n_401, n_400, n_399, n_398, n_397, 
      n_396, n_395, n_394, n_393}), .p_1({n_159, n_158, n_157, n_156, n_155, 
      n_154, n_153, n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, 
      n_144}));
   datapath__0_58 i_22 (.p_0({uc_37, uc_38, n_481, n_480, n_479, n_478, n_477, 
      n_476, n_475, n_474, n_473, n_472, n_471, n_470, n_469, B[0]}), .p_1({
      uc_39, n_407, n_406, n_405, n_404, n_403, n_402, n_401, n_400, n_399, 
      n_398, n_397, n_396, n_395, n_394, n_393}), .p_2({n_175, n_174, n_173, 
      n_172, n_171, n_170, n_169, n_168, n_167, n_166, n_165, n_164, n_163, 
      n_162, n_161, n_160}));
   datapath__0_63 i_25 (.B({uc_40, uc_41, uc_42, B[12], B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_43, n_392, 
      n_391, n_390, n_389, n_388, n_387, n_386, n_385, n_384, n_383, n_382, 
      n_381, n_380, n_379, n_378}), .p_1({n_191, n_190, n_189, n_188, n_187, 
      n_186, n_185, n_184, n_183, n_182, n_181, n_180, n_179, n_178, n_177, 
      n_176}));
   datapath__0_64 i_26 (.p_0({uc_44, uc_45, n_481, n_480, n_479, n_478, n_477, 
      n_476, n_475, n_474, n_473, n_472, n_471, n_470, n_469, B[0]}), .p_1({
      uc_46, n_392, n_391, n_390, n_389, n_388, n_387, n_386, n_385, n_384, 
      n_383, n_382, n_381, n_380, n_379, n_378}), .p_2({n_207, n_206, n_205, 
      n_204, n_203, n_202, n_201, n_200, n_199, n_198, n_197, n_196, n_195, 
      n_194, n_193, n_192}));
   datapath__0_69 i_29 (.B({uc_47, uc_48, B[12], uc_49, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_50, n_377, 
      n_376, n_375, n_374, n_373, n_372, n_371, n_370, n_369, n_368, n_367, 
      n_366, n_365, n_364, n_363}), .p_1({n_223, n_222, n_221, n_220, n_219, 
      n_218, n_217, n_216, n_215, n_214, n_213, n_212, n_211, n_210, n_209, 
      n_208}));
   datapath__0_70 i_30 (.p_0({uc_51, uc_52, n_481, n_480, n_479, n_478, n_477, 
      n_476, n_475, n_474, n_473, n_472, n_471, n_470, n_469, B[0]}), .p_1({
      uc_53, n_377, n_376, n_375, n_374, n_373, n_372, n_371, n_370, n_369, 
      n_368, n_367, n_366, n_365, n_364, n_363}), .p_2({n_239, n_238, n_237, 
      n_236, n_235, n_234, n_233, n_232, n_231, n_230, n_229, n_228, n_227, 
      n_226, n_225, n_224}));
   datapath__0_75 i_33 (.B({uc_54, uc_55, uc_56, B[12], B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_57, n_362, 
      n_361, n_360, n_359, n_358, n_357, n_356, n_355, n_354, n_353, n_352, 
      n_351, n_350, n_349, n_348}), .p_1({n_255, n_254, n_253, n_252, n_251, 
      n_250, n_249, n_248, n_247, n_246, n_245, n_244, n_243, n_242, n_241, 
      n_240}));
   datapath__0_76 i_34 (.p_0({uc_58, uc_59, n_481, n_480, n_479, n_478, n_477, 
      n_476, n_475, n_474, n_473, n_472, n_471, n_470, n_469, B[0]}), .p_1({
      uc_60, n_362, n_361, n_360, n_359, n_358, n_357, n_356, n_355, n_354, 
      n_353, n_352, n_351, n_350, n_349, n_348}), .p_2({n_271, n_270, n_269, 
      n_268, n_267, n_266, n_265, n_264, n_263, n_262, n_261, n_260, n_259, 
      n_258, n_257, n_256}));
   datapath__0_81 i_37 (.B({uc_61, uc_62, uc_63, B[12], B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_64, n_347, 
      n_346, n_345, n_344, n_343, n_342, n_341, n_340, n_339, n_338, n_337, 
      n_336, n_335, n_334, n_333}), .p_1({n_287, n_286, n_285, n_284, n_283, 
      n_282, n_281, n_280, n_279, n_278, n_277, n_276, n_275, n_274, n_273, 
      n_272}));
   datapath__0_82 i_38 (.p_0({uc_65, uc_66, n_481, n_480, n_479, n_478, n_477, 
      n_476, n_475, n_474, n_473, n_472, n_471, n_470, n_469, B[0]}), .p_1({
      uc_67, n_347, n_346, n_345, n_344, n_343, n_342, n_341, n_340, n_339, 
      n_338, n_337, n_336, n_335, n_334, n_333}), .p_2({n_303, n_302, n_301, 
      n_300, n_299, n_298, n_297, n_296, n_295, n_294, n_293, n_292, n_291, 
      n_290, n_289, n_288}));
   INV_X1 i_0_0 (.A(n_0_0), .ZN(product[12]));
   AOI222_X1 i_0_1 (.A1(n_535), .A2(n_0_19), .B1(n_535), .B2(n_0_18), .C1(n_304), 
      .C2(n_0_17), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_1), .ZN(product[13]));
   AOI222_X1 i_0_3 (.A1(n_521), .A2(n_0_19), .B1(n_508), .B2(n_0_18), .C1(n_305), 
      .C2(n_0_17), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(n_0_2), .ZN(product[14]));
   AOI222_X1 i_0_5 (.A1(n_522), .A2(n_0_19), .B1(n_509), .B2(n_0_18), .C1(n_306), 
      .C2(n_0_17), .ZN(n_0_2));
   INV_X1 i_0_6 (.A(n_0_3), .ZN(product[15]));
   AOI222_X1 i_0_7 (.A1(n_523), .A2(n_0_19), .B1(n_510), .B2(n_0_18), .C1(n_307), 
      .C2(n_0_17), .ZN(n_0_3));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(product[16]));
   AOI222_X1 i_0_9 (.A1(n_524), .A2(n_0_19), .B1(n_511), .B2(n_0_18), .C1(n_308), 
      .C2(n_0_17), .ZN(n_0_4));
   INV_X1 i_0_10 (.A(n_0_5), .ZN(product[17]));
   AOI222_X1 i_0_11 (.A1(n_525), .A2(n_0_19), .B1(n_512), .B2(n_0_18), .C1(n_309), 
      .C2(n_0_17), .ZN(n_0_5));
   INV_X1 i_0_12 (.A(n_0_6), .ZN(product[18]));
   AOI222_X1 i_0_13 (.A1(n_526), .A2(n_0_19), .B1(n_513), .B2(n_0_18), .C1(n_310), 
      .C2(n_0_17), .ZN(n_0_6));
   INV_X1 i_0_14 (.A(n_0_7), .ZN(product[19]));
   AOI222_X1 i_0_15 (.A1(n_527), .A2(n_0_19), .B1(n_514), .B2(n_0_18), .C1(n_311), 
      .C2(n_0_17), .ZN(n_0_7));
   INV_X1 i_0_16 (.A(n_0_8), .ZN(product[20]));
   AOI222_X1 i_0_17 (.A1(n_528), .A2(n_0_19), .B1(n_515), .B2(n_0_18), .C1(n_312), 
      .C2(n_0_17), .ZN(n_0_8));
   INV_X1 i_0_18 (.A(n_0_9), .ZN(product[21]));
   AOI222_X1 i_0_19 (.A1(n_529), .A2(n_0_19), .B1(n_516), .B2(n_0_18), .C1(n_313), 
      .C2(n_0_17), .ZN(n_0_9));
   INV_X1 i_0_20 (.A(n_0_10), .ZN(product[22]));
   AOI222_X1 i_0_21 (.A1(n_530), .A2(n_0_19), .B1(n_517), .B2(n_0_18), .C1(n_314), 
      .C2(n_0_17), .ZN(n_0_10));
   INV_X1 i_0_22 (.A(n_0_11), .ZN(product[23]));
   AOI222_X1 i_0_23 (.A1(n_531), .A2(n_0_19), .B1(n_518), .B2(n_0_18), .C1(n_315), 
      .C2(n_0_17), .ZN(n_0_11));
   INV_X1 i_0_24 (.A(n_0_12), .ZN(product[24]));
   AOI222_X1 i_0_25 (.A1(n_532), .A2(n_0_19), .B1(n_519), .B2(n_0_18), .C1(n_316), 
      .C2(n_0_17), .ZN(n_0_12));
   INV_X1 i_0_26 (.A(n_0_13), .ZN(product[27]));
   AOI222_X1 i_0_27 (.A1(n_533), .A2(n_0_19), .B1(n_520), .B2(n_0_18), .C1(n_317), 
      .C2(n_0_17), .ZN(n_0_13));
   NOR2_X1 i_0_33 (.A1(n_0_19), .A2(n_0_18), .ZN(n_0_17));
   NOR2_X1 i_0_34 (.A1(A[12]), .A2(n_0_35), .ZN(n_0_18));
   AND2_X1 i_0_35 (.A1(A[12]), .A2(n_0_35), .ZN(n_0_19));
   INV_X1 i_0_36 (.A(n_0_20), .ZN(product[11]));
   AOI222_X1 i_0_37 (.A1(n_534), .A2(n_0_39), .B1(n_534), .B2(n_0_38), .C1(n_318), 
      .C2(n_0_37), .ZN(n_0_20));
   INV_X1 i_0_38 (.A(n_0_21), .ZN(n_304));
   AOI222_X1 i_0_39 (.A1(n_495), .A2(n_0_39), .B1(n_482), .B2(n_0_38), .C1(n_319), 
      .C2(n_0_37), .ZN(n_0_21));
   INV_X1 i_0_40 (.A(n_0_22), .ZN(n_305));
   AOI222_X1 i_0_41 (.A1(n_496), .A2(n_0_39), .B1(n_483), .B2(n_0_38), .C1(n_320), 
      .C2(n_0_37), .ZN(n_0_22));
   INV_X1 i_0_42 (.A(n_0_23), .ZN(n_306));
   AOI222_X1 i_0_43 (.A1(n_497), .A2(n_0_39), .B1(n_484), .B2(n_0_38), .C1(n_321), 
      .C2(n_0_37), .ZN(n_0_23));
   INV_X1 i_0_44 (.A(n_0_24), .ZN(n_307));
   AOI222_X1 i_0_45 (.A1(n_498), .A2(n_0_39), .B1(n_485), .B2(n_0_38), .C1(n_322), 
      .C2(n_0_37), .ZN(n_0_24));
   INV_X1 i_0_46 (.A(n_0_25), .ZN(n_308));
   AOI222_X1 i_0_47 (.A1(n_499), .A2(n_0_39), .B1(n_486), .B2(n_0_38), .C1(n_323), 
      .C2(n_0_37), .ZN(n_0_25));
   INV_X1 i_0_48 (.A(n_0_26), .ZN(n_309));
   AOI222_X1 i_0_49 (.A1(n_500), .A2(n_0_39), .B1(n_487), .B2(n_0_38), .C1(n_324), 
      .C2(n_0_37), .ZN(n_0_26));
   INV_X1 i_0_50 (.A(n_0_27), .ZN(n_310));
   AOI222_X1 i_0_51 (.A1(n_501), .A2(n_0_39), .B1(n_488), .B2(n_0_38), .C1(n_325), 
      .C2(n_0_37), .ZN(n_0_27));
   INV_X1 i_0_52 (.A(n_0_28), .ZN(n_311));
   AOI222_X1 i_0_53 (.A1(n_502), .A2(n_0_39), .B1(n_489), .B2(n_0_38), .C1(n_326), 
      .C2(n_0_37), .ZN(n_0_28));
   INV_X1 i_0_54 (.A(n_0_29), .ZN(n_312));
   AOI222_X1 i_0_55 (.A1(n_503), .A2(n_0_39), .B1(n_490), .B2(n_0_38), .C1(n_327), 
      .C2(n_0_37), .ZN(n_0_29));
   INV_X1 i_0_56 (.A(n_0_30), .ZN(n_313));
   AOI222_X1 i_0_57 (.A1(n_504), .A2(n_0_39), .B1(n_491), .B2(n_0_38), .C1(n_328), 
      .C2(n_0_37), .ZN(n_0_30));
   INV_X1 i_0_58 (.A(n_0_31), .ZN(n_314));
   AOI222_X1 i_0_59 (.A1(n_505), .A2(n_0_39), .B1(n_492), .B2(n_0_38), .C1(n_329), 
      .C2(n_0_37), .ZN(n_0_31));
   INV_X1 i_0_60 (.A(n_0_32), .ZN(n_315));
   AOI222_X1 i_0_61 (.A1(n_506), .A2(n_0_39), .B1(n_493), .B2(n_0_38), .C1(n_330), 
      .C2(n_0_37), .ZN(n_0_32));
   INV_X1 i_0_62 (.A(n_0_33), .ZN(n_316));
   AOI222_X1 i_0_63 (.A1(n_507), .A2(n_0_39), .B1(n_494), .B2(n_0_38), .C1(n_331), 
      .C2(n_0_37), .ZN(n_0_33));
   INV_X1 i_0_64 (.A(n_0_34), .ZN(n_317));
   AOI221_X1 i_0_65 (.A(n_0_36), .B1(n_537), .B2(n_0_38), .C1(n_536), .C2(n_0_39), 
      .ZN(n_0_34));
   AND2_X1 i_0_68 (.A1(n_332), .A2(n_0_37), .ZN(n_0_36));
   NOR2_X1 i_0_69 (.A1(n_0_39), .A2(n_0_38), .ZN(n_0_37));
   NOR2_X1 i_0_70 (.A1(A[11]), .A2(n_0_16), .ZN(n_0_38));
   NOR2_X1 i_0_71 (.A1(n_0_35), .A2(A[10]), .ZN(n_0_39));
   INV_X1 i_0_72 (.A(n_0_40), .ZN(product[10]));
   AOI222_X1 i_0_73 (.A1(n_288), .A2(n_0_59), .B1(n_272), .B2(n_0_58), .C1(n_333), 
      .C2(n_0_57), .ZN(n_0_40));
   INV_X1 i_0_74 (.A(n_0_41), .ZN(n_318));
   AOI222_X1 i_0_75 (.A1(n_289), .A2(n_0_59), .B1(n_273), .B2(n_0_58), .C1(n_334), 
      .C2(n_0_57), .ZN(n_0_41));
   INV_X1 i_0_76 (.A(n_0_42), .ZN(n_319));
   AOI222_X1 i_0_77 (.A1(n_290), .A2(n_0_59), .B1(n_274), .B2(n_0_58), .C1(n_335), 
      .C2(n_0_57), .ZN(n_0_42));
   INV_X1 i_0_78 (.A(n_0_43), .ZN(n_320));
   AOI222_X1 i_0_79 (.A1(n_291), .A2(n_0_59), .B1(n_275), .B2(n_0_58), .C1(n_336), 
      .C2(n_0_57), .ZN(n_0_43));
   INV_X1 i_0_80 (.A(n_0_44), .ZN(n_321));
   AOI222_X1 i_0_81 (.A1(n_292), .A2(n_0_59), .B1(n_276), .B2(n_0_58), .C1(n_337), 
      .C2(n_0_57), .ZN(n_0_44));
   INV_X1 i_0_82 (.A(n_0_45), .ZN(n_322));
   AOI222_X1 i_0_83 (.A1(n_293), .A2(n_0_59), .B1(n_277), .B2(n_0_58), .C1(n_338), 
      .C2(n_0_57), .ZN(n_0_45));
   INV_X1 i_0_84 (.A(n_0_46), .ZN(n_323));
   AOI222_X1 i_0_85 (.A1(n_294), .A2(n_0_59), .B1(n_278), .B2(n_0_58), .C1(n_339), 
      .C2(n_0_57), .ZN(n_0_46));
   INV_X1 i_0_86 (.A(n_0_47), .ZN(n_324));
   AOI222_X1 i_0_87 (.A1(n_295), .A2(n_0_59), .B1(n_279), .B2(n_0_58), .C1(n_340), 
      .C2(n_0_57), .ZN(n_0_47));
   INV_X1 i_0_88 (.A(n_0_48), .ZN(n_325));
   AOI222_X1 i_0_89 (.A1(n_296), .A2(n_0_59), .B1(n_280), .B2(n_0_58), .C1(n_341), 
      .C2(n_0_57), .ZN(n_0_48));
   INV_X1 i_0_90 (.A(n_0_49), .ZN(n_326));
   AOI222_X1 i_0_91 (.A1(n_297), .A2(n_0_59), .B1(n_281), .B2(n_0_58), .C1(n_342), 
      .C2(n_0_57), .ZN(n_0_49));
   INV_X1 i_0_92 (.A(n_0_50), .ZN(n_327));
   AOI222_X1 i_0_93 (.A1(n_298), .A2(n_0_59), .B1(n_282), .B2(n_0_58), .C1(n_343), 
      .C2(n_0_57), .ZN(n_0_50));
   INV_X1 i_0_94 (.A(n_0_51), .ZN(n_328));
   AOI222_X1 i_0_95 (.A1(n_299), .A2(n_0_59), .B1(n_283), .B2(n_0_58), .C1(n_344), 
      .C2(n_0_57), .ZN(n_0_51));
   INV_X1 i_0_96 (.A(n_0_52), .ZN(n_329));
   AOI222_X1 i_0_97 (.A1(n_300), .A2(n_0_59), .B1(n_284), .B2(n_0_58), .C1(n_345), 
      .C2(n_0_57), .ZN(n_0_52));
   INV_X1 i_0_98 (.A(n_0_53), .ZN(n_330));
   AOI222_X1 i_0_99 (.A1(n_301), .A2(n_0_59), .B1(n_285), .B2(n_0_58), .C1(n_346), 
      .C2(n_0_57), .ZN(n_0_53));
   INV_X1 i_0_100 (.A(n_0_54), .ZN(n_331));
   AOI221_X1 i_0_101 (.A(n_0_56), .B1(n_286), .B2(n_0_58), .C1(n_302), .C2(
      n_0_59), .ZN(n_0_54));
   INV_X1 i_0_102 (.A(n_0_55), .ZN(n_332));
   AOI221_X1 i_0_103 (.A(n_0_56), .B1(n_287), .B2(n_0_58), .C1(n_303), .C2(
      n_0_59), .ZN(n_0_55));
   AND2_X1 i_0_104 (.A1(n_347), .A2(n_0_57), .ZN(n_0_56));
   NOR2_X1 i_0_105 (.A1(n_0_59), .A2(n_0_58), .ZN(n_0_57));
   NOR2_X1 i_0_106 (.A1(A[10]), .A2(n_0_15), .ZN(n_0_58));
   NOR2_X1 i_0_107 (.A1(n_0_16), .A2(A[9]), .ZN(n_0_59));
   INV_X1 i_0_108 (.A(n_0_60), .ZN(product[9]));
   AOI222_X1 i_0_109 (.A1(n_240), .A2(n_0_78), .B1(n_256), .B2(n_0_79), .C1(
      n_348), .C2(n_0_77), .ZN(n_0_60));
   INV_X1 i_0_110 (.A(n_0_61), .ZN(n_333));
   AOI222_X1 i_0_111 (.A1(n_257), .A2(n_0_79), .B1(n_241), .B2(n_0_78), .C1(
      n_349), .C2(n_0_77), .ZN(n_0_61));
   INV_X1 i_0_112 (.A(n_0_62), .ZN(n_334));
   AOI222_X1 i_0_113 (.A1(n_258), .A2(n_0_79), .B1(n_242), .B2(n_0_78), .C1(
      n_350), .C2(n_0_77), .ZN(n_0_62));
   INV_X1 i_0_114 (.A(n_0_63), .ZN(n_335));
   AOI222_X1 i_0_115 (.A1(n_259), .A2(n_0_79), .B1(n_243), .B2(n_0_78), .C1(
      n_351), .C2(n_0_77), .ZN(n_0_63));
   INV_X1 i_0_116 (.A(n_0_64), .ZN(n_336));
   AOI222_X1 i_0_117 (.A1(n_260), .A2(n_0_79), .B1(n_244), .B2(n_0_78), .C1(
      n_352), .C2(n_0_77), .ZN(n_0_64));
   INV_X1 i_0_118 (.A(n_0_65), .ZN(n_337));
   AOI222_X1 i_0_119 (.A1(n_261), .A2(n_0_79), .B1(n_245), .B2(n_0_78), .C1(
      n_353), .C2(n_0_77), .ZN(n_0_65));
   INV_X1 i_0_120 (.A(n_0_66), .ZN(n_338));
   AOI222_X1 i_0_121 (.A1(n_262), .A2(n_0_79), .B1(n_246), .B2(n_0_78), .C1(
      n_354), .C2(n_0_77), .ZN(n_0_66));
   INV_X1 i_0_122 (.A(n_0_67), .ZN(n_339));
   AOI222_X1 i_0_123 (.A1(n_263), .A2(n_0_79), .B1(n_247), .B2(n_0_78), .C1(
      n_355), .C2(n_0_77), .ZN(n_0_67));
   INV_X1 i_0_124 (.A(n_0_68), .ZN(n_340));
   AOI222_X1 i_0_125 (.A1(n_264), .A2(n_0_79), .B1(n_248), .B2(n_0_78), .C1(
      n_356), .C2(n_0_77), .ZN(n_0_68));
   INV_X1 i_0_126 (.A(n_0_69), .ZN(n_341));
   AOI222_X1 i_0_127 (.A1(n_265), .A2(n_0_79), .B1(n_249), .B2(n_0_78), .C1(
      n_357), .C2(n_0_77), .ZN(n_0_69));
   INV_X1 i_0_128 (.A(n_0_70), .ZN(n_342));
   AOI222_X1 i_0_129 (.A1(n_266), .A2(n_0_79), .B1(n_250), .B2(n_0_78), .C1(
      n_358), .C2(n_0_77), .ZN(n_0_70));
   INV_X1 i_0_130 (.A(n_0_71), .ZN(n_343));
   AOI222_X1 i_0_131 (.A1(n_267), .A2(n_0_79), .B1(n_251), .B2(n_0_78), .C1(
      n_359), .C2(n_0_77), .ZN(n_0_71));
   INV_X1 i_0_132 (.A(n_0_72), .ZN(n_344));
   AOI222_X1 i_0_133 (.A1(n_268), .A2(n_0_79), .B1(n_252), .B2(n_0_78), .C1(
      n_360), .C2(n_0_77), .ZN(n_0_72));
   INV_X1 i_0_134 (.A(n_0_73), .ZN(n_345));
   AOI222_X1 i_0_135 (.A1(n_269), .A2(n_0_79), .B1(n_253), .B2(n_0_78), .C1(
      n_361), .C2(n_0_77), .ZN(n_0_73));
   INV_X1 i_0_136 (.A(n_0_74), .ZN(n_346));
   AOI221_X1 i_0_137 (.A(n_0_76), .B1(n_254), .B2(n_0_78), .C1(n_270), .C2(
      n_0_79), .ZN(n_0_74));
   INV_X1 i_0_138 (.A(n_0_75), .ZN(n_347));
   AOI221_X1 i_0_139 (.A(n_0_76), .B1(n_255), .B2(n_0_78), .C1(n_271), .C2(
      n_0_79), .ZN(n_0_75));
   AND2_X1 i_0_140 (.A1(n_362), .A2(n_0_77), .ZN(n_0_76));
   NOR2_X1 i_0_141 (.A1(n_0_79), .A2(n_0_78), .ZN(n_0_77));
   NOR2_X1 i_0_142 (.A1(A[9]), .A2(n_0_14), .ZN(n_0_78));
   NOR2_X1 i_0_143 (.A1(n_0_15), .A2(A[8]), .ZN(n_0_79));
   INV_X1 i_0_144 (.A(n_0_80), .ZN(product[8]));
   AOI222_X1 i_0_145 (.A1(n_208), .A2(n_0_98), .B1(n_224), .B2(n_0_99), .C1(
      n_363), .C2(n_0_97), .ZN(n_0_80));
   INV_X1 i_0_146 (.A(n_0_81), .ZN(n_348));
   AOI222_X1 i_0_147 (.A1(n_209), .A2(n_0_98), .B1(n_225), .B2(n_0_99), .C1(
      n_364), .C2(n_0_97), .ZN(n_0_81));
   INV_X1 i_0_148 (.A(n_0_82), .ZN(n_349));
   AOI222_X1 i_0_149 (.A1(n_226), .A2(n_0_99), .B1(n_210), .B2(n_0_98), .C1(
      n_365), .C2(n_0_97), .ZN(n_0_82));
   INV_X1 i_0_150 (.A(n_0_83), .ZN(n_350));
   AOI222_X1 i_0_151 (.A1(n_227), .A2(n_0_99), .B1(n_211), .B2(n_0_98), .C1(
      n_366), .C2(n_0_97), .ZN(n_0_83));
   INV_X1 i_0_152 (.A(n_0_84), .ZN(n_351));
   AOI222_X1 i_0_153 (.A1(n_228), .A2(n_0_99), .B1(n_212), .B2(n_0_98), .C1(
      n_367), .C2(n_0_97), .ZN(n_0_84));
   INV_X1 i_0_154 (.A(n_0_85), .ZN(n_352));
   AOI222_X1 i_0_155 (.A1(n_229), .A2(n_0_99), .B1(n_213), .B2(n_0_98), .C1(
      n_368), .C2(n_0_97), .ZN(n_0_85));
   INV_X1 i_0_156 (.A(n_0_86), .ZN(n_353));
   AOI222_X1 i_0_157 (.A1(n_230), .A2(n_0_99), .B1(n_214), .B2(n_0_98), .C1(
      n_369), .C2(n_0_97), .ZN(n_0_86));
   INV_X1 i_0_158 (.A(n_0_87), .ZN(n_354));
   AOI222_X1 i_0_159 (.A1(n_231), .A2(n_0_99), .B1(n_215), .B2(n_0_98), .C1(
      n_370), .C2(n_0_97), .ZN(n_0_87));
   INV_X1 i_0_160 (.A(n_0_88), .ZN(n_355));
   AOI222_X1 i_0_161 (.A1(n_232), .A2(n_0_99), .B1(n_216), .B2(n_0_98), .C1(
      n_371), .C2(n_0_97), .ZN(n_0_88));
   INV_X1 i_0_162 (.A(n_0_89), .ZN(n_356));
   AOI222_X1 i_0_163 (.A1(n_233), .A2(n_0_99), .B1(n_217), .B2(n_0_98), .C1(
      n_372), .C2(n_0_97), .ZN(n_0_89));
   INV_X1 i_0_164 (.A(n_0_90), .ZN(n_357));
   AOI222_X1 i_0_165 (.A1(n_234), .A2(n_0_99), .B1(n_218), .B2(n_0_98), .C1(
      n_373), .C2(n_0_97), .ZN(n_0_90));
   INV_X1 i_0_166 (.A(n_0_91), .ZN(n_358));
   AOI222_X1 i_0_167 (.A1(n_235), .A2(n_0_99), .B1(n_219), .B2(n_0_98), .C1(
      n_374), .C2(n_0_97), .ZN(n_0_91));
   INV_X1 i_0_168 (.A(n_0_92), .ZN(n_359));
   AOI222_X1 i_0_169 (.A1(n_236), .A2(n_0_99), .B1(n_220), .B2(n_0_98), .C1(
      n_375), .C2(n_0_97), .ZN(n_0_92));
   INV_X1 i_0_170 (.A(n_0_93), .ZN(n_360));
   AOI222_X1 i_0_171 (.A1(n_237), .A2(n_0_99), .B1(n_221), .B2(n_0_98), .C1(
      n_376), .C2(n_0_97), .ZN(n_0_93));
   INV_X1 i_0_172 (.A(n_0_94), .ZN(n_361));
   AOI221_X1 i_0_173 (.A(n_0_96), .B1(n_222), .B2(n_0_98), .C1(n_238), .C2(
      n_0_99), .ZN(n_0_94));
   INV_X1 i_0_174 (.A(n_0_95), .ZN(n_362));
   AOI221_X1 i_0_175 (.A(n_0_96), .B1(n_223), .B2(n_0_98), .C1(n_239), .C2(
      n_0_99), .ZN(n_0_95));
   AND2_X1 i_0_176 (.A1(n_377), .A2(n_0_97), .ZN(n_0_96));
   NOR2_X1 i_0_177 (.A1(n_0_99), .A2(n_0_98), .ZN(n_0_97));
   NOR2_X1 i_0_178 (.A1(A[8]), .A2(n_0_269), .ZN(n_0_98));
   NOR2_X1 i_0_179 (.A1(n_0_14), .A2(A[7]), .ZN(n_0_99));
   INV_X1 i_0_180 (.A(n_0_100), .ZN(product[7]));
   AOI222_X1 i_0_181 (.A1(n_176), .A2(n_0_118), .B1(n_192), .B2(n_0_119), 
      .C1(n_378), .C2(n_0_117), .ZN(n_0_100));
   INV_X1 i_0_182 (.A(n_0_101), .ZN(n_363));
   AOI222_X1 i_0_183 (.A1(n_177), .A2(n_0_118), .B1(n_193), .B2(n_0_119), 
      .C1(n_379), .C2(n_0_117), .ZN(n_0_101));
   INV_X1 i_0_184 (.A(n_0_102), .ZN(n_364));
   AOI222_X1 i_0_185 (.A1(n_178), .A2(n_0_118), .B1(n_194), .B2(n_0_119), 
      .C1(n_380), .C2(n_0_117), .ZN(n_0_102));
   INV_X1 i_0_186 (.A(n_0_103), .ZN(n_365));
   AOI222_X1 i_0_187 (.A1(n_179), .A2(n_0_118), .B1(n_195), .B2(n_0_119), 
      .C1(n_381), .C2(n_0_117), .ZN(n_0_103));
   INV_X1 i_0_188 (.A(n_0_104), .ZN(n_366));
   AOI222_X1 i_0_189 (.A1(n_196), .A2(n_0_119), .B1(n_180), .B2(n_0_118), 
      .C1(n_382), .C2(n_0_117), .ZN(n_0_104));
   INV_X1 i_0_190 (.A(n_0_105), .ZN(n_367));
   AOI222_X1 i_0_191 (.A1(n_197), .A2(n_0_119), .B1(n_181), .B2(n_0_118), 
      .C1(n_383), .C2(n_0_117), .ZN(n_0_105));
   INV_X1 i_0_192 (.A(n_0_106), .ZN(n_368));
   AOI222_X1 i_0_193 (.A1(n_198), .A2(n_0_119), .B1(n_182), .B2(n_0_118), 
      .C1(n_384), .C2(n_0_117), .ZN(n_0_106));
   INV_X1 i_0_194 (.A(n_0_107), .ZN(n_369));
   AOI222_X1 i_0_195 (.A1(n_199), .A2(n_0_119), .B1(n_183), .B2(n_0_118), 
      .C1(n_385), .C2(n_0_117), .ZN(n_0_107));
   INV_X1 i_0_196 (.A(n_0_108), .ZN(n_370));
   AOI222_X1 i_0_197 (.A1(n_200), .A2(n_0_119), .B1(n_184), .B2(n_0_118), 
      .C1(n_386), .C2(n_0_117), .ZN(n_0_108));
   INV_X1 i_0_198 (.A(n_0_109), .ZN(n_371));
   AOI222_X1 i_0_199 (.A1(n_201), .A2(n_0_119), .B1(n_185), .B2(n_0_118), 
      .C1(n_387), .C2(n_0_117), .ZN(n_0_109));
   INV_X1 i_0_200 (.A(n_0_110), .ZN(n_372));
   AOI222_X1 i_0_201 (.A1(n_202), .A2(n_0_119), .B1(n_186), .B2(n_0_118), 
      .C1(n_388), .C2(n_0_117), .ZN(n_0_110));
   INV_X1 i_0_202 (.A(n_0_111), .ZN(n_373));
   AOI222_X1 i_0_203 (.A1(n_203), .A2(n_0_119), .B1(n_187), .B2(n_0_118), 
      .C1(n_389), .C2(n_0_117), .ZN(n_0_111));
   INV_X1 i_0_204 (.A(n_0_112), .ZN(n_374));
   AOI222_X1 i_0_205 (.A1(n_204), .A2(n_0_119), .B1(n_188), .B2(n_0_118), 
      .C1(n_390), .C2(n_0_117), .ZN(n_0_112));
   INV_X1 i_0_206 (.A(n_0_113), .ZN(n_375));
   AOI222_X1 i_0_207 (.A1(n_205), .A2(n_0_119), .B1(n_189), .B2(n_0_118), 
      .C1(n_391), .C2(n_0_117), .ZN(n_0_113));
   INV_X1 i_0_208 (.A(n_0_114), .ZN(n_376));
   AOI221_X1 i_0_209 (.A(n_0_116), .B1(n_190), .B2(n_0_118), .C1(n_206), 
      .C2(n_0_119), .ZN(n_0_114));
   INV_X1 i_0_210 (.A(n_0_115), .ZN(n_377));
   AOI221_X1 i_0_211 (.A(n_0_116), .B1(n_191), .B2(n_0_118), .C1(n_207), 
      .C2(n_0_119), .ZN(n_0_115));
   AND2_X1 i_0_212 (.A1(n_392), .A2(n_0_117), .ZN(n_0_116));
   NOR2_X1 i_0_213 (.A1(n_0_119), .A2(n_0_118), .ZN(n_0_117));
   NOR2_X1 i_0_214 (.A1(A[7]), .A2(n_0_268), .ZN(n_0_118));
   NOR2_X1 i_0_215 (.A1(n_0_269), .A2(A[6]), .ZN(n_0_119));
   INV_X1 i_0_216 (.A(n_0_120), .ZN(product[6]));
   AOI222_X1 i_0_217 (.A1(n_144), .A2(n_0_138), .B1(n_160), .B2(n_0_139), 
      .C1(n_393), .C2(n_0_137), .ZN(n_0_120));
   INV_X1 i_0_218 (.A(n_0_121), .ZN(n_378));
   AOI222_X1 i_0_219 (.A1(n_145), .A2(n_0_138), .B1(n_161), .B2(n_0_139), 
      .C1(n_394), .C2(n_0_137), .ZN(n_0_121));
   INV_X1 i_0_220 (.A(n_0_122), .ZN(n_379));
   AOI222_X1 i_0_221 (.A1(n_146), .A2(n_0_138), .B1(n_162), .B2(n_0_139), 
      .C1(n_395), .C2(n_0_137), .ZN(n_0_122));
   INV_X1 i_0_222 (.A(n_0_123), .ZN(n_380));
   AOI222_X1 i_0_223 (.A1(n_147), .A2(n_0_138), .B1(n_163), .B2(n_0_139), 
      .C1(n_396), .C2(n_0_137), .ZN(n_0_123));
   INV_X1 i_0_224 (.A(n_0_124), .ZN(n_381));
   AOI222_X1 i_0_225 (.A1(n_148), .A2(n_0_138), .B1(n_164), .B2(n_0_139), 
      .C1(n_397), .C2(n_0_137), .ZN(n_0_124));
   INV_X1 i_0_226 (.A(n_0_125), .ZN(n_382));
   AOI222_X1 i_0_227 (.A1(n_165), .A2(n_0_139), .B1(n_149), .B2(n_0_138), 
      .C1(n_398), .C2(n_0_137), .ZN(n_0_125));
   INV_X1 i_0_228 (.A(n_0_126), .ZN(n_383));
   AOI222_X1 i_0_229 (.A1(n_166), .A2(n_0_139), .B1(n_150), .B2(n_0_138), 
      .C1(n_399), .C2(n_0_137), .ZN(n_0_126));
   INV_X1 i_0_230 (.A(n_0_127), .ZN(n_384));
   AOI222_X1 i_0_231 (.A1(n_167), .A2(n_0_139), .B1(n_151), .B2(n_0_138), 
      .C1(n_400), .C2(n_0_137), .ZN(n_0_127));
   INV_X1 i_0_232 (.A(n_0_128), .ZN(n_385));
   AOI222_X1 i_0_233 (.A1(n_168), .A2(n_0_139), .B1(n_152), .B2(n_0_138), 
      .C1(n_401), .C2(n_0_137), .ZN(n_0_128));
   INV_X1 i_0_234 (.A(n_0_129), .ZN(n_386));
   AOI222_X1 i_0_235 (.A1(n_169), .A2(n_0_139), .B1(n_153), .B2(n_0_138), 
      .C1(n_402), .C2(n_0_137), .ZN(n_0_129));
   INV_X1 i_0_236 (.A(n_0_130), .ZN(n_387));
   AOI222_X1 i_0_237 (.A1(n_170), .A2(n_0_139), .B1(n_154), .B2(n_0_138), 
      .C1(n_403), .C2(n_0_137), .ZN(n_0_130));
   INV_X1 i_0_238 (.A(n_0_131), .ZN(n_388));
   AOI222_X1 i_0_239 (.A1(n_171), .A2(n_0_139), .B1(n_155), .B2(n_0_138), 
      .C1(n_404), .C2(n_0_137), .ZN(n_0_131));
   INV_X1 i_0_240 (.A(n_0_132), .ZN(n_389));
   AOI222_X1 i_0_241 (.A1(n_172), .A2(n_0_139), .B1(n_156), .B2(n_0_138), 
      .C1(n_405), .C2(n_0_137), .ZN(n_0_132));
   INV_X1 i_0_242 (.A(n_0_133), .ZN(n_390));
   AOI222_X1 i_0_243 (.A1(n_173), .A2(n_0_139), .B1(n_157), .B2(n_0_138), 
      .C1(n_406), .C2(n_0_137), .ZN(n_0_133));
   INV_X1 i_0_244 (.A(n_0_134), .ZN(n_391));
   AOI221_X1 i_0_245 (.A(n_0_136), .B1(n_158), .B2(n_0_138), .C1(n_174), 
      .C2(n_0_139), .ZN(n_0_134));
   INV_X1 i_0_246 (.A(n_0_135), .ZN(n_392));
   AOI221_X1 i_0_247 (.A(n_0_136), .B1(n_159), .B2(n_0_138), .C1(n_175), 
      .C2(n_0_139), .ZN(n_0_135));
   AND2_X1 i_0_248 (.A1(n_407), .A2(n_0_137), .ZN(n_0_136));
   NOR2_X1 i_0_249 (.A1(n_0_139), .A2(n_0_138), .ZN(n_0_137));
   NOR2_X1 i_0_250 (.A1(A[6]), .A2(n_0_267), .ZN(n_0_138));
   NOR2_X1 i_0_251 (.A1(n_0_268), .A2(A[5]), .ZN(n_0_139));
   INV_X1 i_0_252 (.A(n_0_140), .ZN(product[5]));
   AOI222_X1 i_0_253 (.A1(n_112), .A2(n_0_158), .B1(n_128), .B2(n_0_159), 
      .C1(n_408), .C2(n_0_157), .ZN(n_0_140));
   INV_X1 i_0_254 (.A(n_0_141), .ZN(n_393));
   AOI222_X1 i_0_255 (.A1(n_113), .A2(n_0_158), .B1(n_129), .B2(n_0_159), 
      .C1(n_409), .C2(n_0_157), .ZN(n_0_141));
   INV_X1 i_0_256 (.A(n_0_142), .ZN(n_394));
   AOI222_X1 i_0_257 (.A1(n_114), .A2(n_0_158), .B1(n_130), .B2(n_0_159), 
      .C1(n_410), .C2(n_0_157), .ZN(n_0_142));
   INV_X1 i_0_258 (.A(n_0_143), .ZN(n_395));
   AOI222_X1 i_0_259 (.A1(n_115), .A2(n_0_158), .B1(n_131), .B2(n_0_159), 
      .C1(n_411), .C2(n_0_157), .ZN(n_0_143));
   INV_X1 i_0_260 (.A(n_0_144), .ZN(n_396));
   AOI222_X1 i_0_261 (.A1(n_116), .A2(n_0_158), .B1(n_132), .B2(n_0_159), 
      .C1(n_412), .C2(n_0_157), .ZN(n_0_144));
   INV_X1 i_0_262 (.A(n_0_145), .ZN(n_397));
   AOI222_X1 i_0_263 (.A1(n_117), .A2(n_0_158), .B1(n_133), .B2(n_0_159), 
      .C1(n_413), .C2(n_0_157), .ZN(n_0_145));
   INV_X1 i_0_264 (.A(n_0_146), .ZN(n_398));
   AOI222_X1 i_0_265 (.A1(n_134), .A2(n_0_159), .B1(n_118), .B2(n_0_158), 
      .C1(n_414), .C2(n_0_157), .ZN(n_0_146));
   INV_X1 i_0_266 (.A(n_0_147), .ZN(n_399));
   AOI222_X1 i_0_267 (.A1(n_135), .A2(n_0_159), .B1(n_119), .B2(n_0_158), 
      .C1(n_415), .C2(n_0_157), .ZN(n_0_147));
   INV_X1 i_0_268 (.A(n_0_148), .ZN(n_400));
   AOI222_X1 i_0_269 (.A1(n_136), .A2(n_0_159), .B1(n_120), .B2(n_0_158), 
      .C1(n_416), .C2(n_0_157), .ZN(n_0_148));
   INV_X1 i_0_270 (.A(n_0_149), .ZN(n_401));
   AOI222_X1 i_0_271 (.A1(n_137), .A2(n_0_159), .B1(n_121), .B2(n_0_158), 
      .C1(n_417), .C2(n_0_157), .ZN(n_0_149));
   INV_X1 i_0_272 (.A(n_0_150), .ZN(n_402));
   AOI222_X1 i_0_273 (.A1(n_138), .A2(n_0_159), .B1(n_122), .B2(n_0_158), 
      .C1(n_418), .C2(n_0_157), .ZN(n_0_150));
   INV_X1 i_0_274 (.A(n_0_151), .ZN(n_403));
   AOI222_X1 i_0_275 (.A1(n_139), .A2(n_0_159), .B1(n_123), .B2(n_0_158), 
      .C1(n_419), .C2(n_0_157), .ZN(n_0_151));
   INV_X1 i_0_276 (.A(n_0_152), .ZN(n_404));
   AOI222_X1 i_0_277 (.A1(n_140), .A2(n_0_159), .B1(n_124), .B2(n_0_158), 
      .C1(n_420), .C2(n_0_157), .ZN(n_0_152));
   INV_X1 i_0_278 (.A(n_0_153), .ZN(n_405));
   AOI222_X1 i_0_279 (.A1(n_141), .A2(n_0_159), .B1(n_125), .B2(n_0_158), 
      .C1(n_421), .C2(n_0_157), .ZN(n_0_153));
   INV_X1 i_0_280 (.A(n_0_154), .ZN(n_406));
   AOI221_X1 i_0_281 (.A(n_0_156), .B1(n_126), .B2(n_0_158), .C1(n_142), 
      .C2(n_0_159), .ZN(n_0_154));
   INV_X1 i_0_282 (.A(n_0_155), .ZN(n_407));
   AOI221_X1 i_0_283 (.A(n_0_156), .B1(n_127), .B2(n_0_158), .C1(n_143), 
      .C2(n_0_159), .ZN(n_0_155));
   AND2_X1 i_0_284 (.A1(n_422), .A2(n_0_157), .ZN(n_0_156));
   NOR2_X1 i_0_285 (.A1(n_0_159), .A2(n_0_158), .ZN(n_0_157));
   NOR2_X1 i_0_286 (.A1(A[5]), .A2(n_0_266), .ZN(n_0_158));
   NOR2_X1 i_0_287 (.A1(n_0_267), .A2(A[4]), .ZN(n_0_159));
   INV_X1 i_0_288 (.A(n_0_160), .ZN(product[4]));
   AOI222_X1 i_0_289 (.A1(n_80), .A2(n_0_178), .B1(n_96), .B2(n_0_179), .C1(
      n_423), .C2(n_0_177), .ZN(n_0_160));
   INV_X1 i_0_290 (.A(n_0_161), .ZN(n_408));
   AOI222_X1 i_0_291 (.A1(n_81), .A2(n_0_178), .B1(n_97), .B2(n_0_179), .C1(
      n_424), .C2(n_0_177), .ZN(n_0_161));
   INV_X1 i_0_292 (.A(n_0_162), .ZN(n_409));
   AOI222_X1 i_0_293 (.A1(n_82), .A2(n_0_178), .B1(n_98), .B2(n_0_179), .C1(
      n_425), .C2(n_0_177), .ZN(n_0_162));
   INV_X1 i_0_294 (.A(n_0_163), .ZN(n_410));
   AOI222_X1 i_0_295 (.A1(n_83), .A2(n_0_178), .B1(n_99), .B2(n_0_179), .C1(
      n_426), .C2(n_0_177), .ZN(n_0_163));
   INV_X1 i_0_296 (.A(n_0_164), .ZN(n_411));
   AOI222_X1 i_0_297 (.A1(n_84), .A2(n_0_178), .B1(n_100), .B2(n_0_179), 
      .C1(n_427), .C2(n_0_177), .ZN(n_0_164));
   INV_X1 i_0_298 (.A(n_0_165), .ZN(n_412));
   AOI222_X1 i_0_299 (.A1(n_85), .A2(n_0_178), .B1(n_101), .B2(n_0_179), 
      .C1(n_428), .C2(n_0_177), .ZN(n_0_165));
   INV_X1 i_0_300 (.A(n_0_166), .ZN(n_413));
   AOI222_X1 i_0_301 (.A1(n_86), .A2(n_0_178), .B1(n_102), .B2(n_0_179), 
      .C1(n_429), .C2(n_0_177), .ZN(n_0_166));
   INV_X1 i_0_302 (.A(n_0_167), .ZN(n_414));
   AOI222_X1 i_0_303 (.A1(n_87), .A2(n_0_178), .B1(n_103), .B2(n_0_179), 
      .C1(n_430), .C2(n_0_177), .ZN(n_0_167));
   INV_X1 i_0_304 (.A(n_0_168), .ZN(n_415));
   AOI222_X1 i_0_305 (.A1(n_104), .A2(n_0_179), .B1(n_88), .B2(n_0_178), 
      .C1(n_431), .C2(n_0_177), .ZN(n_0_168));
   INV_X1 i_0_306 (.A(n_0_169), .ZN(n_416));
   AOI222_X1 i_0_307 (.A1(n_105), .A2(n_0_179), .B1(n_89), .B2(n_0_178), 
      .C1(n_432), .C2(n_0_177), .ZN(n_0_169));
   INV_X1 i_0_308 (.A(n_0_170), .ZN(n_417));
   AOI222_X1 i_0_309 (.A1(n_106), .A2(n_0_179), .B1(n_90), .B2(n_0_178), 
      .C1(n_433), .C2(n_0_177), .ZN(n_0_170));
   INV_X1 i_0_310 (.A(n_0_171), .ZN(n_418));
   AOI222_X1 i_0_311 (.A1(n_107), .A2(n_0_179), .B1(n_91), .B2(n_0_178), 
      .C1(n_434), .C2(n_0_177), .ZN(n_0_171));
   INV_X1 i_0_312 (.A(n_0_172), .ZN(n_419));
   AOI222_X1 i_0_313 (.A1(n_108), .A2(n_0_179), .B1(n_92), .B2(n_0_178), 
      .C1(n_435), .C2(n_0_177), .ZN(n_0_172));
   INV_X1 i_0_314 (.A(n_0_173), .ZN(n_420));
   AOI222_X1 i_0_315 (.A1(n_109), .A2(n_0_179), .B1(n_93), .B2(n_0_178), 
      .C1(n_436), .C2(n_0_177), .ZN(n_0_173));
   INV_X1 i_0_316 (.A(n_0_174), .ZN(n_421));
   AOI221_X1 i_0_317 (.A(n_0_176), .B1(n_94), .B2(n_0_178), .C1(n_110), .C2(
      n_0_179), .ZN(n_0_174));
   INV_X1 i_0_318 (.A(n_0_175), .ZN(n_422));
   AOI221_X1 i_0_319 (.A(n_0_176), .B1(n_95), .B2(n_0_178), .C1(n_111), .C2(
      n_0_179), .ZN(n_0_175));
   AND2_X1 i_0_320 (.A1(n_437), .A2(n_0_177), .ZN(n_0_176));
   NOR2_X1 i_0_321 (.A1(n_0_179), .A2(n_0_178), .ZN(n_0_177));
   NOR2_X1 i_0_322 (.A1(A[4]), .A2(n_0_265), .ZN(n_0_178));
   NOR2_X1 i_0_323 (.A1(n_0_266), .A2(A[3]), .ZN(n_0_179));
   INV_X1 i_0_324 (.A(n_0_180), .ZN(product[3]));
   AOI222_X1 i_0_325 (.A1(n_48), .A2(n_0_198), .B1(n_64), .B2(n_0_199), .C1(
      n_438), .C2(n_0_197), .ZN(n_0_180));
   INV_X1 i_0_326 (.A(n_0_181), .ZN(n_423));
   AOI222_X1 i_0_327 (.A1(n_49), .A2(n_0_198), .B1(n_65), .B2(n_0_199), .C1(
      n_439), .C2(n_0_197), .ZN(n_0_181));
   INV_X1 i_0_328 (.A(n_0_182), .ZN(n_424));
   AOI222_X1 i_0_329 (.A1(n_50), .A2(n_0_198), .B1(n_66), .B2(n_0_199), .C1(
      n_440), .C2(n_0_197), .ZN(n_0_182));
   INV_X1 i_0_330 (.A(n_0_183), .ZN(n_425));
   AOI222_X1 i_0_331 (.A1(n_51), .A2(n_0_198), .B1(n_67), .B2(n_0_199), .C1(
      n_441), .C2(n_0_197), .ZN(n_0_183));
   INV_X1 i_0_332 (.A(n_0_184), .ZN(n_426));
   AOI222_X1 i_0_333 (.A1(n_52), .A2(n_0_198), .B1(n_68), .B2(n_0_199), .C1(
      n_442), .C2(n_0_197), .ZN(n_0_184));
   INV_X1 i_0_334 (.A(n_0_185), .ZN(n_427));
   AOI222_X1 i_0_335 (.A1(n_53), .A2(n_0_198), .B1(n_69), .B2(n_0_199), .C1(
      n_443), .C2(n_0_197), .ZN(n_0_185));
   INV_X1 i_0_336 (.A(n_0_186), .ZN(n_428));
   AOI222_X1 i_0_337 (.A1(n_54), .A2(n_0_198), .B1(n_70), .B2(n_0_199), .C1(
      n_444), .C2(n_0_197), .ZN(n_0_186));
   INV_X1 i_0_338 (.A(n_0_187), .ZN(n_429));
   AOI222_X1 i_0_339 (.A1(n_55), .A2(n_0_198), .B1(n_71), .B2(n_0_199), .C1(
      n_445), .C2(n_0_197), .ZN(n_0_187));
   INV_X1 i_0_340 (.A(n_0_188), .ZN(n_430));
   AOI222_X1 i_0_341 (.A1(n_56), .A2(n_0_198), .B1(n_72), .B2(n_0_199), .C1(
      n_446), .C2(n_0_197), .ZN(n_0_188));
   INV_X1 i_0_342 (.A(n_0_189), .ZN(n_431));
   AOI222_X1 i_0_343 (.A1(n_73), .A2(n_0_199), .B1(n_57), .B2(n_0_198), .C1(
      n_447), .C2(n_0_197), .ZN(n_0_189));
   INV_X1 i_0_344 (.A(n_0_190), .ZN(n_432));
   AOI222_X1 i_0_345 (.A1(n_74), .A2(n_0_199), .B1(n_58), .B2(n_0_198), .C1(
      n_448), .C2(n_0_197), .ZN(n_0_190));
   INV_X1 i_0_346 (.A(n_0_191), .ZN(n_433));
   AOI222_X1 i_0_347 (.A1(n_75), .A2(n_0_199), .B1(n_59), .B2(n_0_198), .C1(
      n_449), .C2(n_0_197), .ZN(n_0_191));
   INV_X1 i_0_348 (.A(n_0_192), .ZN(n_434));
   AOI222_X1 i_0_349 (.A1(n_76), .A2(n_0_199), .B1(n_60), .B2(n_0_198), .C1(
      n_450), .C2(n_0_197), .ZN(n_0_192));
   INV_X1 i_0_350 (.A(n_0_193), .ZN(n_435));
   AOI222_X1 i_0_351 (.A1(n_77), .A2(n_0_199), .B1(n_61), .B2(n_0_198), .C1(
      n_451), .C2(n_0_197), .ZN(n_0_193));
   INV_X1 i_0_352 (.A(n_0_194), .ZN(n_436));
   AOI221_X1 i_0_353 (.A(n_0_196), .B1(n_62), .B2(n_0_198), .C1(n_78), .C2(
      n_0_199), .ZN(n_0_194));
   INV_X1 i_0_354 (.A(n_0_195), .ZN(n_437));
   AOI221_X1 i_0_355 (.A(n_0_196), .B1(n_63), .B2(n_0_198), .C1(n_79), .C2(
      n_0_199), .ZN(n_0_195));
   AND2_X1 i_0_356 (.A1(n_452), .A2(n_0_197), .ZN(n_0_196));
   NOR2_X1 i_0_357 (.A1(n_0_199), .A2(n_0_198), .ZN(n_0_197));
   NOR2_X1 i_0_358 (.A1(A[3]), .A2(n_0_264), .ZN(n_0_198));
   NOR2_X1 i_0_359 (.A1(n_0_265), .A2(A[2]), .ZN(n_0_199));
   INV_X1 i_0_360 (.A(n_0_200), .ZN(product[2]));
   AOI222_X1 i_0_361 (.A1(n_16), .A2(n_0_218), .B1(n_32), .B2(n_0_219), .C1(
      n_453), .C2(n_0_217), .ZN(n_0_200));
   INV_X1 i_0_362 (.A(n_0_201), .ZN(n_438));
   AOI222_X1 i_0_363 (.A1(n_17), .A2(n_0_218), .B1(n_33), .B2(n_0_219), .C1(
      n_454), .C2(n_0_217), .ZN(n_0_201));
   INV_X1 i_0_364 (.A(n_0_202), .ZN(n_439));
   AOI222_X1 i_0_365 (.A1(n_18), .A2(n_0_218), .B1(n_34), .B2(n_0_219), .C1(
      n_455), .C2(n_0_217), .ZN(n_0_202));
   INV_X1 i_0_366 (.A(n_0_203), .ZN(n_440));
   AOI222_X1 i_0_367 (.A1(n_19), .A2(n_0_218), .B1(n_35), .B2(n_0_219), .C1(
      n_456), .C2(n_0_217), .ZN(n_0_203));
   INV_X1 i_0_368 (.A(n_0_204), .ZN(n_441));
   AOI222_X1 i_0_369 (.A1(n_20), .A2(n_0_218), .B1(n_36), .B2(n_0_219), .C1(
      n_457), .C2(n_0_217), .ZN(n_0_204));
   INV_X1 i_0_370 (.A(n_0_205), .ZN(n_442));
   AOI222_X1 i_0_371 (.A1(n_21), .A2(n_0_218), .B1(n_37), .B2(n_0_219), .C1(
      n_458), .C2(n_0_217), .ZN(n_0_205));
   INV_X1 i_0_372 (.A(n_0_206), .ZN(n_443));
   AOI222_X1 i_0_373 (.A1(n_22), .A2(n_0_218), .B1(n_38), .B2(n_0_219), .C1(
      n_459), .C2(n_0_217), .ZN(n_0_206));
   INV_X1 i_0_374 (.A(n_0_207), .ZN(n_444));
   AOI222_X1 i_0_375 (.A1(n_23), .A2(n_0_218), .B1(n_39), .B2(n_0_219), .C1(
      n_460), .C2(n_0_217), .ZN(n_0_207));
   INV_X1 i_0_376 (.A(n_0_208), .ZN(n_445));
   AOI222_X1 i_0_377 (.A1(n_24), .A2(n_0_218), .B1(n_40), .B2(n_0_219), .C1(
      n_461), .C2(n_0_217), .ZN(n_0_208));
   INV_X1 i_0_378 (.A(n_0_209), .ZN(n_446));
   AOI222_X1 i_0_379 (.A1(n_25), .A2(n_0_218), .B1(n_41), .B2(n_0_219), .C1(
      n_462), .C2(n_0_217), .ZN(n_0_209));
   INV_X1 i_0_380 (.A(n_0_210), .ZN(n_447));
   AOI222_X1 i_0_381 (.A1(n_42), .A2(n_0_219), .B1(n_26), .B2(n_0_218), .C1(
      n_463), .C2(n_0_217), .ZN(n_0_210));
   INV_X1 i_0_382 (.A(n_0_211), .ZN(n_448));
   AOI222_X1 i_0_383 (.A1(n_43), .A2(n_0_219), .B1(n_27), .B2(n_0_218), .C1(
      n_464), .C2(n_0_217), .ZN(n_0_211));
   INV_X1 i_0_384 (.A(n_0_212), .ZN(n_449));
   AOI222_X1 i_0_385 (.A1(n_28), .A2(n_0_218), .B1(n_44), .B2(n_0_219), .C1(
      n_465), .C2(n_0_217), .ZN(n_0_212));
   INV_X1 i_0_386 (.A(n_0_213), .ZN(n_450));
   AOI222_X1 i_0_387 (.A1(n_29), .A2(n_0_218), .B1(n_45), .B2(n_0_219), .C1(
      n_466), .C2(n_0_217), .ZN(n_0_213));
   INV_X1 i_0_388 (.A(n_0_214), .ZN(n_451));
   AOI221_X1 i_0_389 (.A(n_0_216), .B1(n_30), .B2(n_0_218), .C1(n_46), .C2(
      n_0_219), .ZN(n_0_214));
   INV_X1 i_0_390 (.A(n_0_215), .ZN(n_452));
   AOI221_X1 i_0_391 (.A(n_0_216), .B1(n_31), .B2(n_0_218), .C1(n_47), .C2(
      n_0_219), .ZN(n_0_215));
   AND2_X1 i_0_392 (.A1(n_467), .A2(n_0_217), .ZN(n_0_216));
   NOR2_X1 i_0_393 (.A1(n_0_219), .A2(n_0_218), .ZN(n_0_217));
   NOR2_X1 i_0_394 (.A1(A[2]), .A2(n_0_263), .ZN(n_0_218));
   NOR2_X1 i_0_395 (.A1(n_0_264), .A2(A[1]), .ZN(n_0_219));
   INV_X1 i_0_396 (.A(n_0_220), .ZN(product[1]));
   AOI222_X1 i_0_397 (.A1(n_0), .A2(n_0_239), .B1(B[0]), .B2(n_0_237), .C1(n_469), 
      .C2(n_0_236), .ZN(n_0_220));
   INV_X1 i_0_398 (.A(n_0_221), .ZN(n_453));
   AOI222_X1 i_0_399 (.A1(n_1), .A2(n_0_239), .B1(n_469), .B2(n_0_237), .C1(
      n_470), .C2(n_0_236), .ZN(n_0_221));
   INV_X1 i_0_400 (.A(n_0_222), .ZN(n_454));
   AOI222_X1 i_0_401 (.A1(n_2), .A2(n_0_239), .B1(n_470), .B2(n_0_237), .C1(
      n_471), .C2(n_0_236), .ZN(n_0_222));
   INV_X1 i_0_402 (.A(n_0_223), .ZN(n_455));
   AOI222_X1 i_0_403 (.A1(n_3), .A2(n_0_239), .B1(n_471), .B2(n_0_237), .C1(
      n_472), .C2(n_0_236), .ZN(n_0_223));
   INV_X1 i_0_404 (.A(n_0_224), .ZN(n_456));
   AOI222_X1 i_0_405 (.A1(n_4), .A2(n_0_239), .B1(n_472), .B2(n_0_237), .C1(
      n_473), .C2(n_0_236), .ZN(n_0_224));
   INV_X1 i_0_406 (.A(n_0_225), .ZN(n_457));
   AOI222_X1 i_0_407 (.A1(n_473), .A2(n_0_237), .B1(n_5), .B2(n_0_239), .C1(
      n_474), .C2(n_0_236), .ZN(n_0_225));
   INV_X1 i_0_408 (.A(n_0_226), .ZN(n_458));
   AOI222_X1 i_0_409 (.A1(n_6), .A2(n_0_239), .B1(n_474), .B2(n_0_237), .C1(
      n_475), .C2(n_0_236), .ZN(n_0_226));
   INV_X1 i_0_410 (.A(n_0_227), .ZN(n_459));
   AOI222_X1 i_0_411 (.A1(n_7), .A2(n_0_239), .B1(n_475), .B2(n_0_237), .C1(
      n_476), .C2(n_0_236), .ZN(n_0_227));
   INV_X1 i_0_412 (.A(n_0_228), .ZN(n_460));
   AOI222_X1 i_0_413 (.A1(n_8), .A2(n_0_239), .B1(n_476), .B2(n_0_237), .C1(
      n_477), .C2(n_0_236), .ZN(n_0_228));
   INV_X1 i_0_414 (.A(n_0_229), .ZN(n_461));
   AOI222_X1 i_0_415 (.A1(n_9), .A2(n_0_239), .B1(n_477), .B2(n_0_237), .C1(
      n_478), .C2(n_0_236), .ZN(n_0_229));
   INV_X1 i_0_416 (.A(n_0_230), .ZN(n_462));
   AOI222_X1 i_0_417 (.A1(n_10), .A2(n_0_239), .B1(n_478), .B2(n_0_237), 
      .C1(n_479), .C2(n_0_236), .ZN(n_0_230));
   INV_X1 i_0_418 (.A(n_0_231), .ZN(n_463));
   AOI222_X1 i_0_419 (.A1(n_11), .A2(n_0_239), .B1(n_479), .B2(n_0_237), 
      .C1(n_480), .C2(n_0_236), .ZN(n_0_231));
   INV_X1 i_0_420 (.A(n_0_232), .ZN(n_464));
   AOI222_X1 i_0_421 (.A1(n_481), .A2(n_0_236), .B1(n_12), .B2(n_0_239), 
      .C1(n_480), .C2(n_0_237), .ZN(n_0_232));
   INV_X1 i_0_422 (.A(n_0_233), .ZN(n_465));
   AOI21_X1 i_0_423 (.A(n_0_238), .B1(n_13), .B2(n_0_239), .ZN(n_0_233));
   INV_X1 i_0_424 (.A(n_0_234), .ZN(n_466));
   AOI21_X1 i_0_425 (.A(n_0_238), .B1(n_14), .B2(n_0_239), .ZN(n_0_234));
   INV_X1 i_0_426 (.A(n_0_235), .ZN(n_467));
   AOI21_X1 i_0_427 (.A(n_0_238), .B1(n_15), .B2(n_0_239), .ZN(n_0_235));
   NOR2_X1 i_0_428 (.A1(n_0_262), .A2(n_0_239), .ZN(n_0_236));
   NOR2_X1 i_0_429 (.A1(n_0_263), .A2(A[0]), .ZN(n_0_237));
   NOR3_X1 i_0_430 (.A1(B[12]), .A2(n_0_241), .A3(n_0_263), .ZN(n_0_238));
   NOR2_X1 i_0_431 (.A1(A[1]), .A2(n_0_262), .ZN(n_0_239));
   AND2_X1 i_0_432 (.A1(B[0]), .A2(A[0]), .ZN(product[0]));
   NOR3_X1 i_0_433 (.A1(B[12]), .A2(n_0_241), .A3(n_0_262), .ZN(n_468));
   AOI21_X1 i_0_434 (.A(n_0_261), .B1(B[1]), .B2(B[0]), .ZN(n_469));
   AOI21_X1 i_0_435 (.A(n_0_259), .B1(B[2]), .B2(n_0_260), .ZN(n_470));
   AOI21_X1 i_0_436 (.A(n_0_257), .B1(B[3]), .B2(n_0_258), .ZN(n_471));
   AOI21_X1 i_0_437 (.A(n_0_255), .B1(B[4]), .B2(n_0_256), .ZN(n_472));
   AOI21_X1 i_0_438 (.A(n_0_253), .B1(B[5]), .B2(n_0_254), .ZN(n_473));
   AOI21_X1 i_0_439 (.A(n_0_251), .B1(B[6]), .B2(n_0_252), .ZN(n_474));
   AOI21_X1 i_0_440 (.A(n_0_249), .B1(B[7]), .B2(n_0_250), .ZN(n_475));
   AOI21_X1 i_0_441 (.A(n_0_247), .B1(B[8]), .B2(n_0_248), .ZN(n_476));
   AOI21_X1 i_0_442 (.A(n_0_245), .B1(B[9]), .B2(n_0_246), .ZN(n_477));
   AOI21_X1 i_0_443 (.A(n_0_243), .B1(B[10]), .B2(n_0_244), .ZN(n_478));
   AOI21_X1 i_0_444 (.A(n_0_241), .B1(B[11]), .B2(n_0_242), .ZN(n_479));
   INV_X1 i_0_445 (.A(n_0_240), .ZN(n_480));
   AOI21_X1 i_0_446 (.A(n_481), .B1(B[12]), .B2(n_0_241), .ZN(n_0_240));
   NOR2_X1 i_0_447 (.A1(B[12]), .A2(n_0_241), .ZN(n_481));
   NOR2_X1 i_0_448 (.A1(B[11]), .A2(n_0_242), .ZN(n_0_241));
   INV_X1 i_0_449 (.A(n_0_243), .ZN(n_0_242));
   NOR2_X1 i_0_450 (.A1(B[10]), .A2(n_0_244), .ZN(n_0_243));
   INV_X1 i_0_451 (.A(n_0_245), .ZN(n_0_244));
   NOR2_X1 i_0_452 (.A1(B[9]), .A2(n_0_246), .ZN(n_0_245));
   INV_X1 i_0_453 (.A(n_0_247), .ZN(n_0_246));
   NOR2_X1 i_0_454 (.A1(B[8]), .A2(n_0_248), .ZN(n_0_247));
   INV_X1 i_0_455 (.A(n_0_249), .ZN(n_0_248));
   NOR2_X1 i_0_456 (.A1(B[7]), .A2(n_0_250), .ZN(n_0_249));
   INV_X1 i_0_457 (.A(n_0_251), .ZN(n_0_250));
   NOR2_X1 i_0_458 (.A1(B[6]), .A2(n_0_252), .ZN(n_0_251));
   INV_X1 i_0_459 (.A(n_0_253), .ZN(n_0_252));
   NOR2_X1 i_0_460 (.A1(B[5]), .A2(n_0_254), .ZN(n_0_253));
   INV_X1 i_0_461 (.A(n_0_255), .ZN(n_0_254));
   NOR2_X1 i_0_462 (.A1(B[4]), .A2(n_0_256), .ZN(n_0_255));
   INV_X1 i_0_463 (.A(n_0_257), .ZN(n_0_256));
   NOR2_X1 i_0_464 (.A1(B[3]), .A2(n_0_258), .ZN(n_0_257));
   INV_X1 i_0_465 (.A(n_0_259), .ZN(n_0_258));
   NOR2_X1 i_0_466 (.A1(B[2]), .A2(n_0_260), .ZN(n_0_259));
   INV_X1 i_0_467 (.A(n_0_261), .ZN(n_0_260));
   NOR2_X1 i_0_468 (.A1(B[1]), .A2(B[0]), .ZN(n_0_261));
   INV_X1 i_0_469 (.A(A[0]), .ZN(n_0_262));
   INV_X1 i_0_470 (.A(A[1]), .ZN(n_0_263));
   INV_X1 i_0_471 (.A(A[2]), .ZN(n_0_264));
   INV_X1 i_0_472 (.A(A[3]), .ZN(n_0_265));
   INV_X1 i_0_473 (.A(A[4]), .ZN(n_0_266));
   INV_X1 i_0_474 (.A(A[5]), .ZN(n_0_267));
   INV_X1 i_0_475 (.A(A[6]), .ZN(n_0_268));
   INV_X1 i_0_476 (.A(A[7]), .ZN(n_0_269));
   INV_X1 i_0_477 (.A(A[8]), .ZN(n_0_14));
   INV_X1 i_0_478 (.A(A[9]), .ZN(n_0_15));
   INV_X1 i_0_479 (.A(A[10]), .ZN(n_0_16));
   INV_X1 i_0_480 (.A(A[11]), .ZN(n_0_35));
   FA_X1 i_1_0 (.A(B[1]), .B(n_319), .CI(n_1_52), .CO(n_1_2), .S(n_482));
   FA_X1 i_1_1 (.A(B[2]), .B(n_320), .CI(n_1_2), .CO(n_1_3), .S(n_483));
   FA_X1 i_1_2 (.A(B[3]), .B(n_321), .CI(n_1_3), .CO(n_1_4), .S(n_484));
   FA_X1 i_1_3 (.A(B[4]), .B(n_322), .CI(n_1_4), .CO(n_1_5), .S(n_485));
   FA_X1 i_1_4 (.A(B[5]), .B(n_323), .CI(n_1_5), .CO(n_1_6), .S(n_486));
   FA_X1 i_1_5 (.A(B[6]), .B(n_324), .CI(n_1_6), .CO(n_1_7), .S(n_487));
   FA_X1 i_1_6 (.A(B[7]), .B(n_325), .CI(n_1_7), .CO(n_1_8), .S(n_488));
   FA_X1 i_1_7 (.A(B[8]), .B(n_326), .CI(n_1_8), .CO(n_1_9), .S(n_489));
   FA_X1 i_1_8 (.A(B[9]), .B(n_327), .CI(n_1_9), .CO(n_1_10), .S(n_490));
   FA_X1 i_1_9 (.A(B[10]), .B(n_328), .CI(n_1_10), .CO(n_1_11), .S(n_491));
   FA_X1 i_1_10 (.A(B[11]), .B(n_329), .CI(n_1_11), .CO(n_1_12), .S(n_492));
   FA_X1 i_1_11 (.A(B[12]), .B(n_330), .CI(n_1_12), .CO(n_1_13), .S(n_493));
   FA_X1 i_1_12 (.A(B[12]), .B(n_331), .CI(n_1_13), .CO(n_1_14), .S(n_494));
   FA_X1 i_1_13 (.A(n_469), .B(n_319), .CI(n_1_52), .CO(n_1_0), .S(n_495));
   FA_X1 i_1_14 (.A(n_470), .B(n_320), .CI(n_1_0), .CO(n_1_1), .S(n_496));
   FA_X1 i_1_15 (.A(n_471), .B(n_321), .CI(n_1_1), .CO(n_1_15), .S(n_497));
   FA_X1 i_1_16 (.A(n_472), .B(n_322), .CI(n_1_15), .CO(n_1_16), .S(n_498));
   FA_X1 i_1_17 (.A(n_473), .B(n_323), .CI(n_1_16), .CO(n_1_17), .S(n_499));
   FA_X1 i_1_18 (.A(n_474), .B(n_324), .CI(n_1_17), .CO(n_1_18), .S(n_500));
   FA_X1 i_1_19 (.A(n_475), .B(n_325), .CI(n_1_18), .CO(n_1_19), .S(n_501));
   FA_X1 i_1_20 (.A(n_476), .B(n_326), .CI(n_1_19), .CO(n_1_20), .S(n_502));
   FA_X1 i_1_21 (.A(n_477), .B(n_327), .CI(n_1_20), .CO(n_1_21), .S(n_503));
   FA_X1 i_1_22 (.A(n_478), .B(n_328), .CI(n_1_21), .CO(n_1_22), .S(n_504));
   FA_X1 i_1_23 (.A(n_479), .B(n_329), .CI(n_1_22), .CO(n_1_23), .S(n_505));
   FA_X1 i_1_24 (.A(n_480), .B(n_330), .CI(n_1_23), .CO(n_1_24), .S(n_506));
   FA_X1 i_1_25 (.A(n_481), .B(n_331), .CI(n_1_24), .CO(n_1_25), .S(n_507));
   FA_X1 i_1_26 (.A(B[1]), .B(n_305), .CI(n_1_53), .CO(n_1_26), .S(n_508));
   FA_X1 i_1_27 (.A(B[2]), .B(n_306), .CI(n_1_26), .CO(n_1_27), .S(n_509));
   FA_X1 i_1_28 (.A(B[3]), .B(n_307), .CI(n_1_27), .CO(n_1_28), .S(n_510));
   FA_X1 i_1_29 (.A(B[4]), .B(n_308), .CI(n_1_28), .CO(n_1_29), .S(n_511));
   FA_X1 i_1_30 (.A(B[5]), .B(n_309), .CI(n_1_29), .CO(n_1_30), .S(n_512));
   FA_X1 i_1_31 (.A(B[6]), .B(n_310), .CI(n_1_30), .CO(n_1_31), .S(n_513));
   FA_X1 i_1_32 (.A(B[7]), .B(n_311), .CI(n_1_31), .CO(n_1_32), .S(n_514));
   FA_X1 i_1_33 (.A(B[8]), .B(n_312), .CI(n_1_32), .CO(n_1_33), .S(n_515));
   FA_X1 i_1_34 (.A(B[9]), .B(n_313), .CI(n_1_33), .CO(n_1_34), .S(n_516));
   FA_X1 i_1_35 (.A(B[10]), .B(n_314), .CI(n_1_34), .CO(n_1_35), .S(n_517));
   FA_X1 i_1_36 (.A(B[11]), .B(n_315), .CI(n_1_35), .CO(n_1_36), .S(n_518));
   FA_X1 i_1_37 (.A(B[12]), .B(n_316), .CI(n_1_36), .CO(n_1_37), .S(n_519));
   FA_X1 i_1_38 (.A(B[12]), .B(n_317), .CI(n_1_37), .CO(n_1_38), .S(n_520));
   FA_X1 i_1_39 (.A(n_469), .B(n_305), .CI(n_1_53), .CO(n_1_39), .S(n_521));
   FA_X1 i_1_40 (.A(n_470), .B(n_306), .CI(n_1_39), .CO(n_1_40), .S(n_522));
   FA_X1 i_1_41 (.A(n_471), .B(n_307), .CI(n_1_40), .CO(n_1_41), .S(n_523));
   FA_X1 i_1_42 (.A(n_472), .B(n_308), .CI(n_1_41), .CO(n_1_42), .S(n_524));
   FA_X1 i_1_43 (.A(n_473), .B(n_309), .CI(n_1_42), .CO(n_1_43), .S(n_525));
   FA_X1 i_1_44 (.A(n_474), .B(n_310), .CI(n_1_43), .CO(n_1_44), .S(n_526));
   FA_X1 i_1_45 (.A(n_475), .B(n_311), .CI(n_1_44), .CO(n_1_45), .S(n_527));
   FA_X1 i_1_46 (.A(n_476), .B(n_312), .CI(n_1_45), .CO(n_1_46), .S(n_528));
   FA_X1 i_1_47 (.A(n_477), .B(n_313), .CI(n_1_46), .CO(n_1_47), .S(n_529));
   FA_X1 i_1_48 (.A(n_478), .B(n_314), .CI(n_1_47), .CO(n_1_48), .S(n_530));
   FA_X1 i_1_49 (.A(n_479), .B(n_315), .CI(n_1_48), .CO(n_1_49), .S(n_531));
   FA_X1 i_1_50 (.A(n_480), .B(n_316), .CI(n_1_49), .CO(n_1_50), .S(n_532));
   FA_X1 i_1_51 (.A(n_481), .B(n_317), .CI(n_1_50), .CO(n_1_51), .S(n_533));
   HA_X1 i_1_52 (.A(B[0]), .B(n_318), .CO(n_1_52), .S(n_534));
   HA_X1 i_1_53 (.A(B[0]), .B(n_304), .CO(n_1_53), .S(n_535));
   XNOR2_X1 i_1_54 (.A(n_332), .B(n_1_54), .ZN(n_536));
   XNOR2_X1 i_1_55 (.A(n_481), .B(n_1_25), .ZN(n_1_54));
   XNOR2_X1 i_1_56 (.A(B[12]), .B(n_1_55), .ZN(n_537));
   XNOR2_X1 i_1_57 (.A(n_332), .B(n_1_14), .ZN(n_1_55));
endmodule

module multiplier_16bit(first_operand, second_operand, out, enable, overflow);
   input [15:0]first_operand;
   input [15:0]second_operand;
   output [15:0]out;
   input enable;
   output overflow;

   wire [31:0]temp_result_wire;
   wire [15:0]second_operand_number;
   wire [15:0]first_operand_number;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_25;
   wire n_0_26;
   wire n_0_56;
   wire n_0_57;
   wire n_0_74;
   wire n_0_75;
   wire n_0_83;

   booth_16bit_multiplier mult (.A({uc_0, uc_1, uc_2, first_operand_number[12], 
      first_operand_number[11], first_operand_number[10], 
      first_operand_number[9], first_operand_number[8], first_operand_number[7], 
      first_operand_number[6], first_operand_number[5], first_operand_number[4], 
      first_operand_number[3], first_operand_number[2], first_operand_number[1], 
      first_operand_number[0]}), .B({uc_3, uc_4, uc_5, second_operand_number[12], 
      second_operand_number[11], second_operand_number[10], 
      second_operand_number[9], second_operand_number[8], 
      second_operand_number[7], second_operand_number[6], 
      second_operand_number[5], second_operand_number[4], 
      second_operand_number[3], second_operand_number[2], 
      second_operand_number[1], second_operand_number[0]}), .product({uc_6, uc_7, 
      uc_8, uc_9, temp_result_wire[25], uc_10, uc_11, temp_result_wire[24], 
      temp_result_wire[23], temp_result_wire[22], temp_result_wire[21], 
      temp_result_wire[20], temp_result_wire[19], temp_result_wire[18], 
      temp_result_wire[17], temp_result_wire[16], temp_result_wire[15], 
      temp_result_wire[14], temp_result_wire[13], temp_result_wire[12], 
      temp_result_wire[11], temp_result_wire[10], temp_result_wire[9], 
      temp_result_wire[8], temp_result_wire[7], temp_result_wire[6], 
      temp_result_wire[5], temp_result_wire[4], temp_result_wire[3], 
      temp_result_wire[2], temp_result_wire[1], temp_result_wire[0]}));
   DLH_X1 overflow_reg (.D(n_13), .G(enable), .Q(overflow));
   DLH_X1 \out_reg[15]  (.D(n_16), .G(enable), .Q(out[15]));
   DLH_X1 \out_reg[14]  (.D(n_15), .G(enable), .Q(out[14]));
   DLH_X1 \out_reg[13]  (.D(n_14), .G(enable), .Q(out[13]));
   DLH_X1 \out_reg[12]  (.D(n_12), .G(enable), .Q(out[12]));
   DLH_X1 \out_reg[11]  (.D(n_11), .G(enable), .Q(out[11]));
   DLH_X1 \out_reg[10]  (.D(n_10), .G(enable), .Q(out[10]));
   DLH_X1 \out_reg[9]  (.D(n_9), .G(enable), .Q(out[9]));
   DLH_X1 \out_reg[8]  (.D(n_8), .G(enable), .Q(out[8]));
   DLH_X1 \out_reg[7]  (.D(n_7), .G(enable), .Q(out[7]));
   DLH_X1 \out_reg[6]  (.D(n_6), .G(enable), .Q(out[6]));
   DLH_X1 \out_reg[5]  (.D(n_5), .G(enable), .Q(out[5]));
   DLH_X1 \out_reg[4]  (.D(n_4), .G(enable), .Q(out[4]));
   DLH_X1 \out_reg[3]  (.D(n_3), .G(enable), .Q(out[3]));
   DLH_X1 \out_reg[2]  (.D(n_2), .G(enable), .Q(out[2]));
   DLH_X1 \out_reg[1]  (.D(n_1), .G(enable), .Q(out[1]));
   DLH_X1 \out_reg[0]  (.D(n_0), .G(enable), .Q(out[0]));
   DLH_X1 \second_operand_number_reg[12]  (.D(second_operand[12]), .G(enable), 
      .Q(second_operand_number[12]));
   DLH_X1 \second_operand_number_reg[11]  (.D(second_operand[11]), .G(enable), 
      .Q(second_operand_number[11]));
   DLH_X1 \second_operand_number_reg[10]  (.D(second_operand[10]), .G(enable), 
      .Q(second_operand_number[10]));
   DLH_X1 \second_operand_number_reg[9]  (.D(second_operand[9]), .G(enable), 
      .Q(second_operand_number[9]));
   DLH_X1 \second_operand_number_reg[8]  (.D(second_operand[8]), .G(enable), 
      .Q(second_operand_number[8]));
   DLH_X1 \second_operand_number_reg[7]  (.D(second_operand[7]), .G(enable), 
      .Q(second_operand_number[7]));
   DLH_X1 \second_operand_number_reg[6]  (.D(second_operand[6]), .G(enable), 
      .Q(second_operand_number[6]));
   DLH_X1 \second_operand_number_reg[5]  (.D(second_operand[5]), .G(enable), 
      .Q(second_operand_number[5]));
   DLH_X1 \second_operand_number_reg[4]  (.D(second_operand[4]), .G(enable), 
      .Q(second_operand_number[4]));
   DLH_X1 \second_operand_number_reg[3]  (.D(second_operand[3]), .G(enable), 
      .Q(second_operand_number[3]));
   DLH_X1 \second_operand_number_reg[2]  (.D(second_operand[2]), .G(enable), 
      .Q(second_operand_number[2]));
   DLH_X1 \second_operand_number_reg[1]  (.D(second_operand[1]), .G(enable), 
      .Q(second_operand_number[1]));
   DLH_X1 \second_operand_number_reg[0]  (.D(second_operand[0]), .G(enable), 
      .Q(second_operand_number[0]));
   DLH_X1 \first_operand_number_reg[12]  (.D(first_operand[12]), .G(enable), 
      .Q(first_operand_number[12]));
   DLH_X1 \first_operand_number_reg[11]  (.D(first_operand[11]), .G(enable), 
      .Q(first_operand_number[11]));
   DLH_X1 \first_operand_number_reg[10]  (.D(first_operand[10]), .G(enable), 
      .Q(first_operand_number[10]));
   DLH_X1 \first_operand_number_reg[9]  (.D(first_operand[9]), .G(enable), 
      .Q(first_operand_number[9]));
   DLH_X1 \first_operand_number_reg[8]  (.D(first_operand[8]), .G(enable), 
      .Q(first_operand_number[8]));
   DLH_X1 \first_operand_number_reg[7]  (.D(first_operand[7]), .G(enable), 
      .Q(first_operand_number[7]));
   DLH_X1 \first_operand_number_reg[6]  (.D(first_operand[6]), .G(enable), 
      .Q(first_operand_number[6]));
   DLH_X1 \first_operand_number_reg[5]  (.D(first_operand[5]), .G(enable), 
      .Q(first_operand_number[5]));
   DLH_X1 \first_operand_number_reg[4]  (.D(first_operand[4]), .G(enable), 
      .Q(first_operand_number[4]));
   DLH_X1 \first_operand_number_reg[3]  (.D(first_operand[3]), .G(enable), 
      .Q(first_operand_number[3]));
   DLH_X1 \first_operand_number_reg[2]  (.D(first_operand[2]), .G(enable), 
      .Q(first_operand_number[2]));
   DLH_X1 \first_operand_number_reg[1]  (.D(first_operand[1]), .G(enable), 
      .Q(first_operand_number[1]));
   DLH_X1 \first_operand_number_reg[0]  (.D(first_operand[0]), .G(enable), 
      .Q(first_operand_number[0]));
   MUX2_X1 i_0_0 (.A(temp_result_wire[0]), .B(temp_result_wire[4]), .S(n_0_79), 
      .Z(n_0_0));
   MUX2_X1 i_0_1 (.A(temp_result_wire[1]), .B(temp_result_wire[5]), .S(n_0_79), 
      .Z(n_0_1));
   MUX2_X1 i_0_2 (.A(temp_result_wire[2]), .B(temp_result_wire[6]), .S(n_0_79), 
      .Z(n_0_2));
   MUX2_X1 i_0_3 (.A(temp_result_wire[3]), .B(temp_result_wire[7]), .S(n_0_79), 
      .Z(n_0_3));
   MUX2_X1 i_0_4 (.A(temp_result_wire[4]), .B(temp_result_wire[8]), .S(n_0_79), 
      .Z(n_0_4));
   MUX2_X1 i_0_5 (.A(temp_result_wire[5]), .B(temp_result_wire[9]), .S(n_0_79), 
      .Z(n_0_5));
   MUX2_X1 i_0_6 (.A(temp_result_wire[6]), .B(temp_result_wire[10]), .S(n_0_79), 
      .Z(n_0_6));
   MUX2_X1 i_0_7 (.A(temp_result_wire[7]), .B(temp_result_wire[11]), .S(n_0_79), 
      .Z(n_0_7));
   MUX2_X1 i_0_8 (.A(temp_result_wire[8]), .B(temp_result_wire[12]), .S(n_0_79), 
      .Z(n_0_8));
   MUX2_X1 i_0_9 (.A(temp_result_wire[9]), .B(temp_result_wire[13]), .S(n_0_79), 
      .Z(n_0_9));
   MUX2_X1 i_0_10 (.A(temp_result_wire[10]), .B(temp_result_wire[14]), .S(n_0_79), 
      .Z(n_0_10));
   MUX2_X1 i_0_11 (.A(temp_result_wire[11]), .B(temp_result_wire[15]), .S(n_0_79), 
      .Z(n_0_11));
   MUX2_X1 i_0_12 (.A(temp_result_wire[12]), .B(temp_result_wire[16]), .S(n_0_79), 
      .Z(n_0_12));
   MUX2_X1 i_0_13 (.A(temp_result_wire[13]), .B(temp_result_wire[17]), .S(n_0_79), 
      .Z(n_0_13));
   MUX2_X1 i_0_14 (.A(temp_result_wire[14]), .B(temp_result_wire[18]), .S(n_0_79), 
      .Z(n_0_14));
   MUX2_X1 i_0_15 (.A(temp_result_wire[15]), .B(temp_result_wire[19]), .S(n_0_79), 
      .Z(n_0_15));
   MUX2_X1 i_0_16 (.A(temp_result_wire[16]), .B(temp_result_wire[20]), .S(n_0_79), 
      .Z(n_0_16));
   MUX2_X1 i_0_17 (.A(temp_result_wire[17]), .B(temp_result_wire[21]), .S(n_0_79), 
      .Z(n_0_17));
   MUX2_X1 i_0_18 (.A(temp_result_wire[18]), .B(temp_result_wire[22]), .S(n_0_79), 
      .Z(n_0_18));
   MUX2_X1 i_0_19 (.A(temp_result_wire[19]), .B(temp_result_wire[23]), .S(n_0_79), 
      .Z(n_0_19));
   MUX2_X1 i_0_20 (.A(temp_result_wire[20]), .B(temp_result_wire[24]), .S(n_0_79), 
      .Z(n_0_20));
   MUX2_X1 i_0_21 (.A(temp_result_wire[21]), .B(temp_result_wire[25]), .S(n_0_79), 
      .Z(n_0_21));
   MUX2_X1 i_0_22 (.A(temp_result_wire[22]), .B(temp_result_wire[25]), .S(n_0_79), 
      .Z(n_0_22));
   MUX2_X1 i_0_23 (.A(temp_result_wire[23]), .B(temp_result_wire[25]), .S(n_0_79), 
      .Z(n_0_23));
   MUX2_X1 i_0_24 (.A(temp_result_wire[24]), .B(temp_result_wire[25]), .S(n_0_79), 
      .Z(n_0_24));
   MUX2_X1 i_0_27 (.A(n_0_0), .B(n_0_2), .S(n_0_78), .Z(n_0_31));
   MUX2_X1 i_0_28 (.A(n_0_1), .B(n_0_3), .S(n_0_78), .Z(n_0_32));
   MUX2_X1 i_0_29 (.A(n_0_2), .B(n_0_4), .S(n_0_78), .Z(n_0_33));
   MUX2_X1 i_0_30 (.A(n_0_3), .B(n_0_5), .S(n_0_78), .Z(n_0_34));
   MUX2_X1 i_0_31 (.A(n_0_4), .B(n_0_6), .S(n_0_78), .Z(n_0_35));
   MUX2_X1 i_0_32 (.A(n_0_5), .B(n_0_7), .S(n_0_78), .Z(n_0_36));
   MUX2_X1 i_0_33 (.A(n_0_6), .B(n_0_8), .S(n_0_78), .Z(n_0_37));
   MUX2_X1 i_0_34 (.A(n_0_7), .B(n_0_9), .S(n_0_78), .Z(n_0_38));
   MUX2_X1 i_0_35 (.A(n_0_8), .B(n_0_10), .S(n_0_78), .Z(n_0_39));
   MUX2_X1 i_0_36 (.A(n_0_9), .B(n_0_11), .S(n_0_78), .Z(n_0_40));
   MUX2_X1 i_0_37 (.A(n_0_10), .B(n_0_12), .S(n_0_78), .Z(n_0_41));
   MUX2_X1 i_0_38 (.A(n_0_11), .B(n_0_13), .S(n_0_78), .Z(n_0_42));
   MUX2_X1 i_0_39 (.A(n_0_12), .B(n_0_14), .S(n_0_78), .Z(n_0_43));
   MUX2_X1 i_0_40 (.A(n_0_13), .B(n_0_15), .S(n_0_78), .Z(n_0_44));
   MUX2_X1 i_0_41 (.A(n_0_14), .B(n_0_16), .S(n_0_78), .Z(n_0_45));
   MUX2_X1 i_0_42 (.A(n_0_15), .B(n_0_17), .S(n_0_78), .Z(n_0_46));
   MUX2_X1 i_0_43 (.A(n_0_16), .B(n_0_18), .S(n_0_78), .Z(n_0_47));
   MUX2_X1 i_0_44 (.A(n_0_17), .B(n_0_19), .S(n_0_78), .Z(n_0_48));
   MUX2_X1 i_0_45 (.A(n_0_18), .B(n_0_20), .S(n_0_78), .Z(n_0_49));
   MUX2_X1 i_0_46 (.A(n_0_19), .B(n_0_21), .S(n_0_78), .Z(n_0_50));
   MUX2_X1 i_0_47 (.A(n_0_20), .B(n_0_22), .S(n_0_78), .Z(n_0_51));
   MUX2_X1 i_0_48 (.A(n_0_21), .B(n_0_23), .S(n_0_78), .Z(n_0_52));
   MUX2_X1 i_0_49 (.A(n_0_22), .B(n_0_24), .S(n_0_78), .Z(n_0_53));
   MUX2_X1 i_0_50 (.A(n_0_23), .B(temp_result_wire[25]), .S(n_0_78), .Z(n_0_54));
   MUX2_X1 i_0_51 (.A(n_0_24), .B(temp_result_wire[25]), .S(n_0_78), .Z(n_0_55));
   MUX2_X1 i_0_54 (.A(n_0_31), .B(n_0_32), .S(n_0_77), .Z(n_0));
   MUX2_X1 i_0_55 (.A(n_0_32), .B(n_0_33), .S(n_0_77), .Z(n_1));
   MUX2_X1 i_0_56 (.A(n_0_33), .B(n_0_34), .S(n_0_77), .Z(n_2));
   MUX2_X1 i_0_57 (.A(n_0_34), .B(n_0_35), .S(n_0_77), .Z(n_3));
   MUX2_X1 i_0_58 (.A(n_0_35), .B(n_0_36), .S(n_0_77), .Z(n_4));
   MUX2_X1 i_0_59 (.A(n_0_36), .B(n_0_37), .S(n_0_77), .Z(n_5));
   MUX2_X1 i_0_60 (.A(n_0_37), .B(n_0_38), .S(n_0_77), .Z(n_6));
   MUX2_X1 i_0_61 (.A(n_0_38), .B(n_0_39), .S(n_0_77), .Z(n_7));
   MUX2_X1 i_0_62 (.A(n_0_39), .B(n_0_40), .S(n_0_77), .Z(n_8));
   MUX2_X1 i_0_63 (.A(n_0_40), .B(n_0_41), .S(n_0_77), .Z(n_9));
   MUX2_X1 i_0_64 (.A(n_0_41), .B(n_0_42), .S(n_0_77), .Z(n_10));
   MUX2_X1 i_0_65 (.A(n_0_42), .B(n_0_43), .S(n_0_77), .Z(n_11));
   MUX2_X1 i_0_66 (.A(n_0_43), .B(n_0_44), .S(n_0_77), .Z(n_12));
   MUX2_X1 i_0_67 (.A(n_0_44), .B(n_0_45), .S(n_0_77), .Z(n_0_62));
   MUX2_X1 i_0_68 (.A(n_0_45), .B(n_0_46), .S(n_0_77), .Z(n_0_63));
   MUX2_X1 i_0_69 (.A(n_0_46), .B(n_0_47), .S(n_0_77), .Z(n_0_64));
   MUX2_X1 i_0_70 (.A(n_0_47), .B(n_0_48), .S(n_0_77), .Z(n_0_65));
   MUX2_X1 i_0_71 (.A(n_0_48), .B(n_0_49), .S(n_0_77), .Z(n_0_66));
   MUX2_X1 i_0_72 (.A(n_0_49), .B(n_0_50), .S(n_0_77), .Z(n_0_67));
   MUX2_X1 i_0_73 (.A(n_0_50), .B(n_0_51), .S(n_0_77), .Z(n_0_68));
   MUX2_X1 i_0_74 (.A(n_0_51), .B(n_0_52), .S(n_0_77), .Z(n_0_69));
   MUX2_X1 i_0_75 (.A(n_0_52), .B(n_0_53), .S(n_0_77), .Z(n_0_70));
   MUX2_X1 i_0_76 (.A(n_0_53), .B(n_0_54), .S(n_0_77), .Z(n_0_71));
   MUX2_X1 i_0_77 (.A(n_0_54), .B(n_0_55), .S(n_0_77), .Z(n_0_72));
   MUX2_X1 i_0_78 (.A(n_0_55), .B(temp_result_wire[25]), .S(n_0_77), .Z(n_0_73));
   INV_X1 i_0_81 (.A(second_operand[13]), .ZN(n_0_27));
   INV_X1 i_0_82 (.A(second_operand[14]), .ZN(n_0_28));
   OAI211_X1 i_0_83 (.A(n_0_27), .B(first_operand[13]), .C1(n_0_28), .C2(
      first_operand[14]), .ZN(n_0_29));
   INV_X1 i_0_84 (.A(first_operand[14]), .ZN(n_0_30));
   OAI21_X1 i_0_85 (.A(n_0_29), .B1(second_operand[14]), .B2(n_0_30), .ZN(n_0_58));
   INV_X1 i_0_86 (.A(second_operand[15]), .ZN(n_0_59));
   OAI21_X1 i_0_87 (.A(n_0_58), .B1(first_operand[15]), .B2(n_0_59), .ZN(n_0_60));
   INV_X1 i_0_88 (.A(first_operand[15]), .ZN(n_0_61));
   OAI21_X1 i_0_89 (.A(n_0_60), .B1(second_operand[15]), .B2(n_0_61), .ZN(n_0_76));
   MUX2_X1 i_0_90 (.A(first_operand[13]), .B(second_operand[13]), .S(n_0_76), 
      .Z(n_0_77));
   MUX2_X1 i_0_91 (.A(first_operand[14]), .B(second_operand[14]), .S(n_0_76), 
      .Z(n_0_78));
   MUX2_X1 i_0_92 (.A(first_operand[15]), .B(second_operand[15]), .S(n_0_76), 
      .Z(n_0_79));
   NAND4_X1 i_0_93 (.A1(n_12), .A2(n_0_64), .A3(n_0_63), .A4(n_0_62), .ZN(n_0_80));
   NAND4_X1 i_0_94 (.A1(n_0_67), .A2(n_0_66), .A3(n_0_65), .A4(n_0_70), .ZN(
      n_0_81));
   NAND4_X1 i_0_95 (.A1(n_0_69), .A2(n_0_68), .A3(n_0_73), .A4(n_0_72), .ZN(
      n_0_82));
   NOR3_X1 i_0_97 (.A1(n_0_80), .A2(n_0_81), .A3(n_0_82), .ZN(n_0_84));
   NOR2_X1 i_0_98 (.A1(n_0_83), .A2(n_0_74), .ZN(n_0_85));
   NAND2_X1 i_0_99 (.A1(n_0_85), .A2(n_0_84), .ZN(n_0_86));
   NOR4_X1 i_0_100 (.A1(n_12), .A2(n_0_64), .A3(n_0_63), .A4(n_0_62), .ZN(n_0_87));
   NOR4_X1 i_0_101 (.A1(n_0_67), .A2(n_0_66), .A3(n_0_65), .A4(n_0_70), .ZN(
      n_0_88));
   NOR4_X1 i_0_102 (.A1(n_0_69), .A2(n_0_68), .A3(n_0_73), .A4(n_0_72), .ZN(
      n_0_25));
   AND3_X1 i_0_104 (.A1(n_0_87), .A2(n_0_88), .A3(n_0_25), .ZN(n_0_26));
   NAND3_X1 i_0_105 (.A1(n_0_26), .A2(n_0_75), .A3(n_0_74), .ZN(n_0_56));
   NAND2_X1 i_0_106 (.A1(n_0_56), .A2(n_0_86), .ZN(n_0_57));
   INV_X1 i_0_107 (.A(temp_result_wire[25]), .ZN(n_0_74));
   NOR2_X1 i_0_25 (.A1(n_0_71), .A2(temp_result_wire[25]), .ZN(n_0_75));
   NAND2_X1 i_0_26 (.A1(n_0_71), .A2(temp_result_wire[25]), .ZN(n_0_83));
   NAND2_X1 i_0_108 (.A1(n_0_57), .A2(enable), .ZN(n_13));
   MUX2_X1 i_0_109 (.A(second_operand[13]), .B(first_operand[13]), .S(n_0_76), 
      .Z(n_14));
   MUX2_X1 i_0_110 (.A(second_operand[14]), .B(first_operand[14]), .S(n_0_76), 
      .Z(n_15));
   MUX2_X1 i_0_111 (.A(second_operand[15]), .B(first_operand[15]), .S(n_0_76), 
      .Z(n_16));
endmodule

module Step_Module(RST, CLK, Step_Memory_WR_Enable, RAM_Data_RD_A, RAM_Data_RD_B, 
      RAM_Address_RD_A, RAM_Address_RD_B, RAM_Data_WR, RAM_Address_WR, 
      Euler_Enable, Euler_End, Error_Flag);
   input RST;
   input CLK;
   output Step_Memory_WR_Enable;
   input [63:0]RAM_Data_RD_A;
   input [63:0]RAM_Data_RD_B;
   output [12:0]RAM_Address_RD_A;
   output [12:0]RAM_Address_RD_B;
   output [63:0]RAM_Data_WR;
   output [12:0]RAM_Address_WR;
   output Euler_Enable;
   input Euler_End;
   output Error_Flag;

   wire n_1_0;
   wire [3:0]State;
   wire [15:0]second_operand;
   wire [2:0]hstate;
   wire n_1_1;
   wire [15:0]dividend;
   wire [15:0]first_operand;
   wire n_1_2;
   wire [63:0]N;
   wire division_operation;
   wire n_1_3;
   wire [15:0]in11;
   wire n_1_4;
   wire n_1_1_0;
   wire n_1_1_1;
   wire n_1_1_2;
   wire n_1_1_3;
   wire n_1_1_4;
   wire n_1_1_5;
   wire n_1_1_6;
   wire n_1_1_7;
   wire n_1_1_8;
   wire n_1_1_9;
   wire n_1_1_10;
   wire n_1_1_11;
   wire n_1_1_12;
   wire n_1_1_13;
   wire n_1_1_21;
   wire n_1_1_22;
   wire n_1_1_24;
   wire n_1_1_25;
   wire n_1_1_27;
   wire n_1_1_28;
   wire n_1_1_30;
   wire n_1_1_31;
   wire n_1_1_32;
   wire n_1_6;
   wire n_1_7;
   wire n_1_1_33;
   wire n_1_11;
   wire n_1_15;
   wire n_1_1_34;
   wire n_1_1_35;
   wire n_1_1_36;
   wire n_1_1_37;
   wire n_1_1_38;
   wire n_1_1_39;
   wire n_1_1_40;
   wire n_1_1_41;
   wire n_1_1_42;
   wire n_1_1_43;
   wire n_1_1_44;
   wire n_1_1_45;
   wire n_1_1_46;
   wire n_1_1_47;
   wire n_1_1_48;
   wire n_1_1_49;
   wire n_1_1_50;
   wire n_1_1_51;
   wire n_1_1_52;
   wire n_1_1_53;
   wire n_1_1_54;
   wire n_1_16;
   wire n_1_18;
   wire n_1_20;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;
   wire n_1_28;
   wire n_1_80;
   wire n_1_1_57;
   wire n_1_8;
   wire n_1_9;
   wire n_1_1_58;
   wire n_1_1_59;
   wire n_1_83;
   wire n_1_1_60;
   wire n_1_84;
   wire n_1_1_61;
   wire n_1_85;
   wire n_1_1_62;
   wire n_1_86;
   wire n_1_1_63;
   wire n_1_87;
   wire n_1_1_64;
   wire n_1_88;
   wire n_1_1_65;
   wire n_1_89;
   wire n_1_1_66;
   wire n_1_90;
   wire n_1_1_67;
   wire n_1_91;
   wire n_1_1_68;
   wire n_1_92;
   wire n_1_1_69;
   wire n_1_93;
   wire n_1_1_70;
   wire n_1_94;
   wire n_1_1_71;
   wire n_1_95;
   wire n_1_1_72;
   wire n_1_96;
   wire n_1_1_73;
   wire n_1_97;
   wire n_1_1_74;
   wire n_1_98;
   wire n_1_1_75;
   wire n_1_1_76;
   wire n_1_1_77;
   wire n_1_17;
   wire n_1_1_78;
   wire n_1_1_79;
   wire n_1_19;
   wire n_1_1_80;
   wire n_1_1_81;
   wire n_1_21;
   wire n_1_1_82;
   wire n_1_22;
   wire n_1_1_83;
   wire n_1_1_84;
   wire n_1_1_85;
   wire n_1_1_86;
   wire n_1_1_87;
   wire n_1_1_88;
   wire n_1_1_89;
   wire n_1_1_90;
   wire n_1_1_91;
   wire n_1_1_92;
   wire n_1_1_93;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire n_1_60;
   wire n_1_61;
   wire n_1_62;
   wire n_1_63;
   wire n_1_64;
   wire n_1_65;
   wire n_1_66;
   wire n_1_67;
   wire n_1_68;
   wire n_1_69;
   wire n_1_70;
   wire n_1_71;
   wire n_1_72;
   wire n_1_73;
   wire n_1_74;
   wire n_1_75;
   wire n_1_76;
   wire n_1_77;
   wire n_1_78;
   wire n_1_79;
   wire n_1_1_98;
   wire n_1_1_99;
   wire n_1_1_100;
   wire n_1_1_101;
   wire n_1_1_102;
   wire n_1_1_103;
   wire n_1_99;
   wire n_1_1_104;
   wire n_1_100;
   wire n_1_1_105;
   wire n_1_101;
   wire n_1_102;
   wire n_1_103;
   wire n_1_1_106;
   wire n_1_104;
   wire n_1_1_107;
   wire n_1_105;
   wire n_1_1_108;
   wire n_1_106;
   wire n_1_107;
   wire n_1_108;
   wire n_1_109;
   wire n_1_110;
   wire n_1_111;
   wire n_1_112;
   wire n_1_1_109;
   wire n_1_113;
   wire n_1_1_110;
   wire n_1_114;
   wire n_1_1_111;
   wire n_1_116;
   wire n_1_1_112;
   wire n_1_117;
   wire n_1_1_113;
   wire n_1_118;
   wire n_1_1_114;
   wire n_1_119;
   wire n_1_1_115;
   wire n_1_120;
   wire n_1_1_116;
   wire n_1_121;
   wire n_1_1_117;
   wire n_1_122;
   wire n_1_1_118;
   wire n_1_123;
   wire n_1_1_119;
   wire n_1_124;
   wire n_1_1_120;
   wire n_1_125;
   wire n_1_1_121;
   wire n_1_126;
   wire n_1_1_122;
   wire n_1_127;
   wire n_1_1_123;
   wire n_1_128;
   wire n_1_1_124;
   wire n_1_129;
   wire n_1_1_125;
   wire n_1_130;
   wire n_1_1_126;
   wire n_1_131;
   wire n_1_1_127;
   wire n_1_1_132;
   wire n_1_1_133;
   wire n_1_1_134;
   wire n_1_1_135;
   wire n_1_1_136;
   wire n_1_1_137;
   wire n_1_1_138;
   wire n_1_1_139;
   wire n_1_1_140;
   wire n_1_1_141;
   wire n_1_1_142;
   wire n_1_1_143;
   wire n_1_1_144;
   wire n_1_1_145;
   wire n_1_1_146;
   wire n_1_1_147;
   wire n_1_1_148;
   wire n_1_1_149;
   wire n_1_1_150;
   wire n_1_1_151;
   wire n_1_1_152;
   wire n_1_1_153;
   wire n_1_1_154;
   wire n_1_1_155;
   wire n_1_1_156;
   wire n_1_1_157;
   wire n_1_1_158;
   wire n_1_132;
   wire n_1_1_165;
   wire n_1_1_166;
   wire n_1_133;
   wire n_1_1_167;
   wire n_1_134;
   wire n_1_1_168;
   wire n_1_1_169;
   wire n_1_1_170;
   wire n_1_135;
   wire n_1_1_171;
   wire n_1_136;
   wire n_1_1_172;
   wire n_1_137;
   wire n_1_1_173;
   wire n_1_138;
   wire n_1_1_174;
   wire n_1_139;
   wire n_1_1_175;
   wire n_1_140;
   wire n_1_1_176;
   wire n_1_141;
   wire n_1_1_177;
   wire n_1_142;
   wire n_1_1_178;
   wire n_1_143;
   wire n_1_1_179;
   wire n_1_1_180;
   wire n_1_1_181;
   wire n_1_1_182;
   wire n_1_144;
   wire n_1_1_183;
   wire n_1_145;
   wire n_1_1_184;
   wire n_1_146;
   wire n_1_1_185;
   wire n_1_147;
   wire n_1_1_186;
   wire n_1_1_187;
   wire n_1_1_189;
   wire n_1_1_190;
   wire n_1_1_191;
   wire n_1_1_192;
   wire n_1_1_193;
   wire n_1_1_194;
   wire n_1_1_195;
   wire n_1_1_196;
   wire n_1_1_197;
   wire n_1_1_198;
   wire n_1_1_199;
   wire n_1_1_200;
   wire n_1_1_201;
   wire n_1_1_202;
   wire n_1_1_203;
   wire n_1_1_204;
   wire n_1_1_205;
   wire n_1_1_206;
   wire n_1_1_207;
   wire n_1_1_208;
   wire n_1_1_209;
   wire n_1_1_210;
   wire n_1_1_211;
   wire n_1_1_212;
   wire n_1_1_213;
   wire n_1_1_214;
   wire n_1_1_215;
   wire n_1_1_216;
   wire n_1_1_217;
   wire n_1_1_219;
   wire n_1_1_221;
   wire n_1_1_222;
   wire n_1_1_223;
   wire n_1_1_224;
   wire n_1_1_225;
   wire n_1_1_226;
   wire n_1_1_227;
   wire n_1_1_228;
   wire n_1_1_229;
   wire n_1_1_230;
   wire n_1_1_231;
   wire n_1_1_232;
   wire n_1_1_233;
   wire n_1_1_234;
   wire n_1_29;
   wire n_1_1_235;
   wire n_1_1_236;
   wire n_1_30;
   wire n_1_1_237;
   wire n_1_1_238;
   wire n_1_1_239;
   wire n_1_31;
   wire n_1_1_240;
   wire n_1_1_242;
   wire n_1_1_243;
   wire n_1_1_244;
   wire n_1_1_245;
   wire n_1_1_246;
   wire n_1_1_247;
   wire n_1_1_249;
   wire n_1_1_250;
   wire n_1_1_251;
   wire n_1_1_252;
   wire n_1_1_254;
   wire n_1_1_259;
   wire n_1_1_260;
   wire n_1_1_265;
   wire n_1_1_266;
   wire n_1_1_267;
   wire n_1_1_268;
   wire n_1_12;
   wire n_1_1_269;
   wire n_1_1_270;
   wire n_1_1_273;
   wire n_1_1_274;
   wire n_1_1_275;
   wire n_1_1_276;
   wire n_1_1_277;
   wire n_1_1_278;
   wire n_1_1_280;
   wire n_1_1_281;
   wire n_1_1_282;
   wire n_1_1_283;
   wire n_1_1_284;
   wire n_1_1_285;
   wire n_1_1_286;
   wire n_1_1_287;
   wire n_1_1_288;
   wire n_1_1_289;
   wire n_1_1_290;
   wire n_1_1_291;
   wire n_1_1_292;
   wire n_1_1_293;
   wire n_1_1_294;
   wire n_1_1_295;
   wire n_1_1_296;
   wire n_1_1_297;
   wire n_1_1_298;
   wire n_1_1_299;
   wire n_1_1_300;
   wire n_1_1_304;
   wire n_1_1_325;
   wire n_1_1_331;
   wire n_1_1_344;
   wire n_1_1_349;
   wire n_1_1_350;
   wire n_1_1_351;
   wire n_1_1_352;
   wire n_1_1_353;
   wire n_1_1_354;
   wire n_1_5;
   wire n_1_1_450;
   wire n_1_1_457;
   wire n_1_1_458;
   wire n_1_1_459;
   wire n_1_1_461;
   wire n_1_1_462;
   wire n_1_1_463;
   wire n_1_1_464;
   wire n_1_1_465;
   wire n_1_1_466;
   wire n_1_1_467;
   wire n_1_1_468;
   wire n_1_1_469;
   wire n_1_1_470;
   wire n_1_1_471;
   wire n_1_1_472;
   wire n_1_1_473;
   wire n_1_1_474;
   wire n_1_1_475;
   wire n_1_1_476;
   wire n_1_1_477;
   wire n_1_1_478;
   wire n_1_1_479;
   wire n_1_1_480;
   wire n_1_13;
   wire n_1_1_481;
   wire n_1_1_483;
   wire n_1_1_485;
   wire n_1_1_487;
   wire n_1_1_488;
   wire n_1_1_489;
   wire n_1_1_490;
   wire n_1_1_491;
   wire n_1_1_492;
   wire n_1_1_493;
   wire n_1_1_494;
   wire n_1_1_495;
   wire n_1_1_496;
   wire n_1_1_497;
   wire n_1_1_498;
   wire n_1_1_499;
   wire n_1_1_500;
   wire n_1_1_501;
   wire n_1_1_502;
   wire n_1_1_503;
   wire n_1_1_504;
   wire n_1_1_505;
   wire n_1_1_506;
   wire n_1_1_507;
   wire n_1_1_508;
   wire n_1_1_509;
   wire n_1_1_510;
   wire n_1_1_511;
   wire n_1_1_512;
   wire n_1_1_513;
   wire n_1_1_514;
   wire n_1_1_515;
   wire n_1_1_516;
   wire n_1_1_517;
   wire n_1_1_518;
   wire n_1_1_519;
   wire n_1_1_520;
   wire n_1_1_521;
   wire n_1_1_522;
   wire n_1_1_523;
   wire n_1_1_524;
   wire n_1_1_525;
   wire n_1_1_526;
   wire n_1_1_527;
   wire n_1_1_528;
   wire n_1_1_529;
   wire n_1_1_530;
   wire n_1_1_531;
   wire n_1_1_532;
   wire n_1_1_533;
   wire n_1_1_534;
   wire n_1_1_536;
   wire n_1_14;
   wire n_1_1_547;
   wire n_1_1_548;
   wire n_1_1_549;
   wire n_1_1_550;
   wire n_1_1_551;
   wire n_1_1_552;
   wire n_1_1_553;
   wire n_1_1_554;
   wire n_1_1_555;
   wire n_1_1_556;
   wire n_1_1_557;
   wire n_1_1_558;
   wire n_1_1_559;
   wire n_1_1_560;
   wire n_1_1_561;
   wire n_1_1_562;
   wire n_1_1_584;
   wire n_1_1_585;
   wire n_1_1_586;
   wire n_1_1_587;
   wire n_1_1_588;
   wire n_1_1_589;
   wire n_1_1_590;
   wire n_1_1_592;
   wire n_1_1_595;
   wire n_1_1_596;
   wire n_1_1_599;
   wire n_1_1_600;
   wire n_1_1_601;
   wire n_1_1_603;
   wire n_1_1_606;
   wire n_1_1_607;
   wire n_1_1_608;
   wire n_1_1_609;
   wire n_1_1_611;
   wire n_1_1_612;
   wire n_1_1_642;
   wire n_1_1_643;
   wire n_1_1_644;
   wire n_1_1_645;
   wire n_1_1_646;
   wire n_1_1_647;
   wire n_1_1_648;
   wire n_1_1_649;
   wire n_1_1_650;
   wire n_1_1_651;
   wire n_1_1_652;
   wire n_1_1_653;
   wire n_1_1_654;
   wire n_1_1_655;
   wire n_1_1_656;
   wire n_1_1_657;
   wire n_1_1_658;
   wire n_1_1_597;
   wire n_1_1_19;
   wire n_1_1_159;
   wire n_1_1_23;
   wire n_1_1_20;
   wire n_1_1_95;
   wire n_1_1_55;
   wire n_1_1_56;
   wire n_1_1_97;
   wire n_1_1_272;
   wire n_1_1_164;
   wire n_1_1_188;
   wire n_1_1_220;
   wire n_1_1_255;
   wire n_1_1_256;
   wire n_1_1_94;
   wire n_1_1_257;
   wire n_1_1_258;
   wire n_1_1_241;
   wire n_1_1_660;
   wire n_1_1_271;
   wire n_1_1_661;
   wire n_1_1_662;
   wire n_1_1_663;
   wire n_1_1_664;
   wire n_1_1_665;
   wire n_1_1_666;
   wire n_1_1_668;
   wire n_1_1_669;
   wire n_1_1_670;
   wire n_1_1_598;
   wire n_1_1_671;
   wire n_1_1_672;
   wire n_1_1_591;
   wire n_1_1_673;
   wire n_1_1_674;
   wire n_1_1_675;
   wire n_1_1_621;
   wire n_1_1_620;
   wire n_1_1_617;
   wire n_1_1_616;
   wire n_1_1_613;
   wire n_1_1_631;
   wire n_1_1_486;
   wire n_1_1_635;
   wire n_1_1_624;
   wire n_1_1_623;
   wire n_1_1_160;
   wire n_1_1_610;
   wire n_1_1_14;
   wire n_1_1_29;
   wire n_1_1_26;
   wire n_1_1_15;
   wire n_1_1_16;
   wire n_1_1_17;
   wire n_1_1_18;
   wire n_1_1_128;
   wire n_1_1_129;
   wire n_1_1_130;
   wire n_1_1_131;
   wire n_1_1_161;
   wire n_1_1_163;
   wire n_1_1_262;
   wire n_1_1_604;
   wire n_1_1_263;
   wire n_1_1_218;
   wire n_1_1_96;
   wire n_1_1_301;
   wire n_1_115;
   wire n_1_1_253;
   wire n_1_1_593;
   wire n_1_1_248;
   wire n_1_1_302;
   wire n_1_1_303;
   wire n_1_1_305;
   wire n_1_1_306;
   wire n_1_1_261;
   wire n_1_1_162;
   wire n_1_1_279;
   wire n_1_1_307;
   wire n_1_1_308;
   wire n_1_1_667;
   wire n_1_1_309;
   wire n_1_1_310;
   wire n_1_1_311;
   wire n_1_1_312;
   wire n_1_1_264;
   wire n_1_1_313;
   wire n_1_1_314;
   wire n_1_1_315;
   wire n_1_1_316;
   wire n_1_1_317;
   wire n_1_1_318;
   wire n_1_1_319;
   wire n_1_1_320;
   wire n_1_1_321;
   wire n_1_1_322;
   wire n_1_1_323;
   wire n_1_1_324;
   wire n_1_1_326;
   wire n_1_1_327;
   wire n_1_1_328;
   wire n_1_1_329;
   wire n_1_1_330;
   wire n_1_1_332;
   wire n_1_1_333;
   wire n_1_1_334;
   wire n_1_1_335;
   wire n_1_1_336;
   wire n_1_1_337;
   wire n_1_1_338;
   wire n_1_1_339;
   wire n_1_1_340;
   wire n_1_1_341;
   wire n_1_1_342;
   wire n_1_1_343;
   wire n_1_1_345;
   wire n_1_1_346;
   wire n_1_1_347;
   wire n_1_1_348;
   wire n_1_1_355;
   wire n_1_1_356;
   wire n_1_1_357;
   wire n_1_1_358;
   wire n_1_1_359;
   wire n_1_1_360;
   wire n_1_1_361;
   wire n_1_1_362;
   wire n_1_1_363;
   wire n_1_1_364;
   wire n_1_1_365;
   wire n_1_1_366;
   wire n_1_1_367;
   wire n_1_1_368;
   wire n_1_1_369;
   wire n_1_1_370;
   wire n_1_1_371;
   wire n_1_1_372;
   wire n_1_1_373;
   wire n_1_1_374;
   wire n_1_1_375;
   wire n_1_1_376;
   wire n_1_1_377;
   wire n_1_1_378;
   wire n_1_1_379;
   wire n_1_1_380;
   wire n_1_1_381;
   wire n_1_1_382;
   wire n_1_1_383;
   wire n_1_1_384;
   wire n_1_1_385;
   wire n_1_1_386;
   wire n_1_1_387;
   wire n_1_1_388;
   wire n_1_1_389;
   wire n_1_1_390;
   wire n_1_1_391;
   wire n_1_1_392;
   wire n_1_1_393;
   wire n_1_1_394;
   wire n_1_1_455;
   wire n_1_1_395;
   wire n_1_1_396;
   wire n_1_1_397;
   wire n_1_1_398;
   wire n_1_1_399;
   wire n_1_1_400;
   wire n_1_1_401;
   wire n_1_1_402;
   wire n_1_1_403;
   wire n_1_1_404;
   wire n_1_1_405;
   wire n_1_1_406;
   wire n_1_1_407;
   wire n_1_1_408;
   wire n_1_1_409;
   wire n_1_1_410;
   wire n_1_1_411;
   wire n_1_1_412;
   wire n_1_1_413;
   wire n_1_1_414;
   wire n_1_1_415;
   wire n_1_1_416;
   wire n_1_1_417;
   wire n_1_1_418;
   wire n_1_1_419;
   wire n_1_1_420;
   wire n_1_1_421;
   wire n_1_1_422;
   wire n_1_1_423;
   wire n_1_1_424;
   wire n_1_1_425;
   wire n_1_1_426;
   wire n_1_1_427;
   wire n_1_1_428;
   wire n_1_1_429;
   wire n_1_1_430;
   wire n_1_1_431;
   wire n_1_1_432;
   wire n_1_1_433;
   wire n_1_1_434;
   wire n_1_1_435;
   wire n_1_1_436;
   wire n_1_1_437;
   wire n_1_1_438;
   wire n_1_1_439;
   wire n_1_1_440;
   wire n_1_1_441;
   wire n_1_1_442;
   wire n_1_1_443;
   wire n_1_1_444;
   wire n_1_1_445;
   wire n_1_1_446;
   wire n_1_1_447;
   wire n_1_1_448;
   wire n_1_1_449;
   wire n_1_1_453;
   wire n_1_1_454;
   wire n_1_1_456;
   wire n_1_1_484;
   wire n_1_1_537;
   wire n_1_1_538;
   wire n_1_1_539;
   wire n_1_1_542;
   wire n_1_1_543;
   wire n_1_1_564;
   wire n_1_1_565;
   wire n_1_1_566;
   wire n_1_1_567;
   wire n_1_1_568;
   wire n_1_1_569;
   wire n_1_1_570;
   wire n_1_1_571;
   wire n_1_1_572;
   wire n_1_1_573;
   wire n_1_1_574;
   wire n_1_1_575;
   wire n_1_1_576;
   wire n_1_1_577;
   wire n_1_1_578;
   wire n_1_1_579;
   wire n_1_1_580;
   wire n_1_1_602;
   wire n_1_1_659;
   wire n_1_1_676;
   wire n_1_1_677;
   wire n_1_1_678;
   wire n_1_1_679;
   wire n_1_1_680;
   wire n_1_1_681;
   wire n_1_1_682;
   wire n_1_1_683;
   wire n_1_1_684;
   wire n_1_1_685;
   wire n_1_1_686;
   wire n_1_1_687;
   wire n_1_1_688;
   wire n_1_1_689;
   wire n_1_1_690;
   wire n_1_1_691;
   wire n_1_1_692;
   wire n_1_1_693;
   wire n_1_1_694;
   wire n_1_1_695;
   wire n_1_1_696;
   wire n_1_1_697;
   wire n_1_1_698;
   wire n_1_1_699;
   wire n_1_1_700;
   wire n_1_1_701;
   wire n_1_1_702;
   wire n_1_1_703;
   wire n_1_1_704;
   wire n_1_1_705;
   wire n_1_1_706;
   wire n_1_1_707;
   wire n_1_1_708;
   wire n_1_1_709;
   wire n_1_1_710;
   wire n_1_1_711;
   wire n_1_1_712;
   wire n_1_1_713;
   wire n_1_1_714;
   wire n_1_1_715;
   wire n_1_1_716;
   wire n_1_1_717;
   wire n_1_1_718;
   wire n_1_1_719;
   wire n_1_1_720;
   wire n_1_1_721;
   wire n_1_1_722;
   wire n_1_1_723;
   wire n_1_1_724;
   wire n_1_1_725;
   wire n_1_1_726;
   wire n_1_1_727;
   wire n_1_1_728;
   wire n_1_1_729;
   wire n_1_1_730;
   wire n_1_1_731;
   wire n_1_1_732;
   wire n_1_1_733;
   wire n_1_1_734;
   wire n_1_1_735;
   wire n_1_1_736;
   wire n_1_1_737;
   wire n_1_1_738;
   wire n_1_1_739;
   wire n_1_1_740;
   wire n_1_1_741;
   wire n_1_1_742;
   wire n_1_1_743;
   wire n_1_1_744;
   wire n_1_1_745;
   wire n_1_1_746;
   wire n_1_1_747;
   wire n_1_1_748;
   wire n_1_1_749;
   wire n_1_1_750;
   wire n_1_1_751;
   wire n_1_1_752;
   wire n_1_1_753;
   wire n_1_1_754;
   wire n_1_1_755;
   wire n_1_1_756;
   wire n_1_1_757;
   wire n_1_1_758;
   wire n_1_1_759;
   wire n_1_1_760;
   wire n_1_1_761;
   wire n_1_1_762;
   wire n_1_1_763;
   wire n_1_1_764;
   wire n_1_1_765;
   wire n_1_1_766;
   wire n_1_1_767;
   wire n_1_1_768;
   wire n_1_1_769;
   wire n_1_1_770;
   wire n_1_1_771;
   wire n_1_1_772;
   wire n_1_1_773;
   wire n_1_1_774;
   wire n_1_1_775;
   wire n_1_1_776;
   wire n_1_1_777;
   wire n_1_1_778;
   wire n_1_1_779;
   wire n_1_1_780;
   wire n_1_1_781;
   wire n_1_1_782;
   wire n_1_1_783;
   wire n_1_1_784;
   wire n_1_1_785;
   wire n_1_1_786;
   wire n_1_1_787;
   wire n_1_1_788;
   wire n_1_1_789;
   wire n_1_1_790;
   wire n_1_1_791;
   wire n_1_1_792;
   wire n_1_1_793;
   wire n_1_1_794;
   wire n_1_1_795;
   wire n_1_1_796;
   wire n_1_1_797;
   wire n_1_1_798;
   wire n_1_1_799;
   wire n_1_1_800;
   wire n_1_1_801;
   wire n_1_1_802;
   wire n_1_1_803;
   wire n_1_1_804;
   wire n_1_1_805;
   wire n_1_1_806;
   wire n_1_1_807;
   wire n_1_1_808;
   wire n_1_1_809;
   wire n_1_1_810;
   wire n_1_1_811;
   wire n_1_1_812;
   wire n_1_1_813;
   wire n_1_1_814;
   wire n_1_1_815;
   wire n_1_1_816;
   wire n_1_1_817;
   wire n_1_1_818;
   wire n_1_1_819;
   wire n_1_1_820;
   wire n_1_1_821;
   wire n_1_1_822;
   wire n_1_1_823;
   wire n_1_1_824;
   wire n_1_1_825;
   wire n_1_1_452;
   wire n_1_1_826;
   wire n_1_1_827;
   wire n_1_1_828;
   wire n_1_1_829;
   wire n_1_1_460;
   wire n_1_1_830;
   wire n_1_1_451;
   wire n_1_1_535;
   wire n_1_1_545;
   wire n_1_1_831;
   wire n_1_1_832;
   wire n_1_1_833;
   wire n_1_1_834;
   wire n_1_1_544;
   wire n_1_1_482;
   wire n_1_1_835;
   wire n_1_1_836;
   wire n_1_1_605;
   wire n_1_1_837;
   wire n_1_1_838;
   wire n_1_1_839;
   wire n_1_1_540;
   wire n_1_1_541;
   wire n_1_1_581;
   wire n_1_1_840;
   wire n_1_1_582;
   wire n_1_1_841;
   wire n_1_1_594;
   wire n_1_1_842;
   wire n_1_1_583;
   wire n_1_1_843;
   wire n_1_1_844;
   wire n_1_1_845;
   wire n_1_1_846;
   wire n_1_1_847;
   wire n_1_1_546;
   wire n_1_1_848;
   wire n_1_1_563;
   wire n_1_1_849;
   wire n_1_1_625;
   wire n_1_1_850;
   wire n_1_1_851;
   wire n_1_1_641;
   wire n_1_1_852;
   wire n_1_1_640;
   wire n_1_1_853;
   wire n_1_1_854;
   wire n_1_1_622;
   wire n_1_1_855;
   wire n_1_1_856;
   wire n_1_1_638;
   wire n_1_1_857;
   wire n_1_1_637;
   wire n_1_1_858;
   wire n_1_1_859;
   wire n_1_1_860;
   wire n_1_1_618;
   wire n_1_1_619;
   wire n_1_1_861;
   wire n_1_1_862;
   wire n_1_1_634;
   wire n_1_1_863;
   wire n_1_1_633;
   wire n_1_1_864;
   wire n_1_1_865;
   wire n_1_1_866;
   wire n_1_1_614;
   wire n_1_1_615;
   wire n_1_1_867;
   wire n_1_1_868;
   wire n_1_1_630;
   wire n_1_1_869;
   wire n_1_1_629;
   wire n_1_1_870;
   wire n_1_1_871;
   wire n_1_1_628;
   wire n_1_1_872;
   wire n_1_1_626;
   wire n_1_1_627;
   wire n_1_1_632;
   wire n_1_1_636;
   wire n_1_1_639;
   wire n_1_81;
   wire n_1_10;
   wire n_1_82;
   wire n_2_0;
   wire [63:0]htemp;
   wire n_2_1;
   wire n_2_2;
   wire [63:0]Temp;
   wire n_2_3;
   wire [15:0]in22;
   wire [15:0]in12;
   wire n_2_4;
   wire [15:0]divisor;
   wire n_2_5;
   wire n_2_6;
   wire n_2_7;
   wire mult_enable;
   wire reset;
   wire sub2;
   wire n_3_0;
   wire [3:0]NextState;
   wire sub1;
   wire n_3_1;
   wire [15:0]in21;
   wire n_3_2;
   wire [12:0]count;
   wire n_3_6;
   wire n_3_3;
   wire n_3_4;
   wire [63:0]Errortemp;
   wire n_3_5;
   wire n_3_7;
   wire reset_reg_enable_mux_n_0;
   wire reset_reg_enable_mux_n_1;
   wire reset_reg_enable_mux_n_2;
   wire n_3_8;
   wire n_3_10;
   wire n_3_9;
   wire n_3_11;
   wire n_3_12;
   wire n_3_13;
   wire n_3_14;
   wire invalid1;
   wire [15:0]adder_out1;
   wire invalid2;
   wire [15:0]adder_out2;
   wire divideByZero;
   wire div_overflow;
   wire ready;
   wire [15:0]Q;
   wire mult_overflow;
   wire [15:0]out;
   wire n_0_0_0;

   CLKGATETST_X1 clk_gate_State_reg (.CK(CLK), .E(n_1_15), .SE(1'b0), .GCK(n_1_0));
   DFF_X1 \State_reg[3]  (.D(n_1_14), .CK(n_1_0), .Q(State[3]), .QN());
   DFF_X1 \State_reg[2]  (.D(n_1_13), .CK(n_1_0), .Q(State[2]), .QN());
   DFF_X1 \State_reg[1]  (.D(n_1_12), .CK(n_1_0), .Q(State[1]), .QN());
   DFF_X1 \State_reg[0]  (.D(n_1_11), .CK(n_1_0), .Q(State[0]), .QN());
   DFF_X1 \second_operand_reg[15]  (.D(n_1_131), .CK(n_1_4), .Q(
      second_operand[15]), .QN());
   DFF_X1 \second_operand_reg[14]  (.D(n_1_130), .CK(n_1_4), .Q(
      second_operand[14]), .QN());
   DFF_X1 \second_operand_reg[13]  (.D(n_1_129), .CK(n_1_4), .Q(
      second_operand[13]), .QN());
   DFF_X1 \second_operand_reg[12]  (.D(n_1_128), .CK(n_1_4), .Q(
      second_operand[12]), .QN());
   DFF_X1 \second_operand_reg[11]  (.D(n_1_127), .CK(n_1_4), .Q(
      second_operand[11]), .QN());
   DFF_X1 \second_operand_reg[10]  (.D(n_1_126), .CK(n_1_4), .Q(
      second_operand[10]), .QN());
   DFF_X1 \second_operand_reg[9]  (.D(n_1_125), .CK(n_1_4), .Q(second_operand[9]), 
      .QN());
   DFF_X1 \second_operand_reg[8]  (.D(n_1_124), .CK(n_1_4), .Q(second_operand[8]), 
      .QN());
   DFF_X1 \second_operand_reg[7]  (.D(n_1_123), .CK(n_1_4), .Q(second_operand[7]), 
      .QN());
   DFF_X1 \second_operand_reg[6]  (.D(n_1_122), .CK(n_1_4), .Q(second_operand[6]), 
      .QN());
   DFF_X1 \second_operand_reg[5]  (.D(n_1_121), .CK(n_1_4), .Q(second_operand[5]), 
      .QN());
   DFF_X1 \second_operand_reg[4]  (.D(n_1_120), .CK(n_1_4), .Q(second_operand[4]), 
      .QN());
   DFF_X1 \second_operand_reg[3]  (.D(n_1_119), .CK(n_1_4), .Q(second_operand[3]), 
      .QN());
   DFF_X1 \second_operand_reg[2]  (.D(n_1_118), .CK(n_1_4), .Q(second_operand[2]), 
      .QN());
   DFF_X1 \second_operand_reg[1]  (.D(n_1_117), .CK(n_1_4), .Q(second_operand[1]), 
      .QN());
   DFF_X1 \second_operand_reg[0]  (.D(n_1_116), .CK(n_1_4), .Q(second_operand[0]), 
      .QN());
   DFF_X1 \hstate_reg[0]  (.D(n_1_81), .CK(CLK), .Q(hstate[0]), .QN());
   DFF_X1 \hstate_reg[1]  (.D(n_1_10), .CK(CLK), .Q(hstate[1]), .QN());
   CLKGATETST_X1 clk_gate_dividend_reg (.CK(CLK), .E(n_242), .SE(1'b0), .GCK(
      n_1_1));
   DFF_X1 \dividend_reg[15]  (.D(n_1_98), .CK(n_1_1), .Q(dividend[15]), .QN());
   DFF_X1 \dividend_reg[14]  (.D(n_1_97), .CK(n_1_1), .Q(dividend[14]), .QN());
   DFF_X1 \dividend_reg[13]  (.D(n_1_96), .CK(n_1_1), .Q(dividend[13]), .QN());
   DFF_X1 \dividend_reg[12]  (.D(n_1_95), .CK(n_1_1), .Q(dividend[12]), .QN());
   DFF_X1 \dividend_reg[11]  (.D(n_1_94), .CK(n_1_1), .Q(dividend[11]), .QN());
   DFF_X1 \dividend_reg[10]  (.D(n_1_93), .CK(n_1_1), .Q(dividend[10]), .QN());
   DFF_X1 \dividend_reg[9]  (.D(n_1_92), .CK(n_1_1), .Q(dividend[9]), .QN());
   DFF_X1 \dividend_reg[8]  (.D(n_1_91), .CK(n_1_1), .Q(dividend[8]), .QN());
   DFF_X1 \dividend_reg[7]  (.D(n_1_90), .CK(n_1_1), .Q(dividend[7]), .QN());
   DFF_X1 \dividend_reg[6]  (.D(n_1_89), .CK(n_1_1), .Q(dividend[6]), .QN());
   DFF_X1 \dividend_reg[5]  (.D(n_1_88), .CK(n_1_1), .Q(dividend[5]), .QN());
   DFF_X1 \dividend_reg[4]  (.D(n_1_87), .CK(n_1_1), .Q(dividend[4]), .QN());
   DFF_X1 \dividend_reg[3]  (.D(n_1_86), .CK(n_1_1), .Q(dividend[3]), .QN());
   DFF_X1 \dividend_reg[2]  (.D(n_1_85), .CK(n_1_1), .Q(dividend[2]), .QN());
   DFF_X1 \dividend_reg[1]  (.D(n_1_84), .CK(n_1_1), .Q(dividend[1]), .QN());
   DFF_X1 \dividend_reg[0]  (.D(n_1_83), .CK(n_1_1), .Q(dividend[0]), .QN());
   DFF_X1 \first_operand_reg[15]  (.D(n_1_114), .CK(n_1_4), .Q(first_operand[15]), 
      .QN());
   DFF_X1 \first_operand_reg[14]  (.D(n_1_113), .CK(n_1_4), .Q(first_operand[14]), 
      .QN());
   DFF_X1 \first_operand_reg[13]  (.D(n_1_112), .CK(n_1_4), .Q(first_operand[13]), 
      .QN());
   DFF_X1 \first_operand_reg[12]  (.D(n_1_111), .CK(n_1_4), .Q(first_operand[12]), 
      .QN());
   DFF_X1 \first_operand_reg[11]  (.D(n_1_110), .CK(n_1_4), .Q(first_operand[11]), 
      .QN());
   DFF_X1 \first_operand_reg[10]  (.D(n_1_109), .CK(n_1_4), .Q(first_operand[10]), 
      .QN());
   DFF_X1 \first_operand_reg[9]  (.D(n_1_108), .CK(n_1_4), .Q(first_operand[9]), 
      .QN());
   DFF_X1 \first_operand_reg[8]  (.D(n_1_107), .CK(n_1_4), .Q(first_operand[8]), 
      .QN());
   DFF_X1 \first_operand_reg[7]  (.D(n_1_106), .CK(n_1_4), .Q(first_operand[7]), 
      .QN());
   DFF_X1 \first_operand_reg[6]  (.D(n_1_105), .CK(n_1_4), .Q(first_operand[6]), 
      .QN());
   DFF_X1 \first_operand_reg[5]  (.D(n_1_104), .CK(n_1_4), .Q(first_operand[5]), 
      .QN());
   DFF_X1 \first_operand_reg[4]  (.D(n_1_103), .CK(n_1_4), .Q(first_operand[4]), 
      .QN());
   DFF_X1 \first_operand_reg[3]  (.D(n_1_102), .CK(n_1_4), .Q(first_operand[3]), 
      .QN());
   DFF_X1 \first_operand_reg[2]  (.D(n_1_101), .CK(n_1_4), .Q(first_operand[2]), 
      .QN());
   DFF_X1 \first_operand_reg[1]  (.D(n_1_100), .CK(n_1_4), .Q(first_operand[1]), 
      .QN());
   DFF_X1 \first_operand_reg[0]  (.D(n_1_99), .CK(n_1_4), .Q(first_operand[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_N_reg (.CK(CLK), .E(n_1_80), .SE(1'b0), .GCK(n_1_2));
   DFF_X1 \N_reg[63]  (.D(n_1_79), .CK(n_1_2), .Q(N[63]), .QN());
   DFF_X1 \N_reg[62]  (.D(n_1_78), .CK(n_1_2), .Q(N[62]), .QN());
   DFF_X1 \N_reg[61]  (.D(n_1_77), .CK(n_1_2), .Q(N[61]), .QN());
   DFF_X1 \N_reg[60]  (.D(n_1_76), .CK(n_1_2), .Q(N[60]), .QN());
   DFF_X1 \N_reg[59]  (.D(n_1_75), .CK(n_1_2), .Q(N[59]), .QN());
   DFF_X1 \N_reg[58]  (.D(n_1_74), .CK(n_1_2), .Q(N[58]), .QN());
   DFF_X1 \N_reg[57]  (.D(n_1_73), .CK(n_1_2), .Q(N[57]), .QN());
   DFF_X1 \N_reg[56]  (.D(n_1_72), .CK(n_1_2), .Q(N[56]), .QN());
   DFF_X1 \N_reg[55]  (.D(n_1_71), .CK(n_1_2), .Q(N[55]), .QN());
   DFF_X1 \N_reg[54]  (.D(n_1_70), .CK(n_1_2), .Q(N[54]), .QN());
   DFF_X1 \N_reg[53]  (.D(n_1_69), .CK(n_1_2), .Q(N[53]), .QN());
   DFF_X1 \N_reg[52]  (.D(n_1_68), .CK(n_1_2), .Q(N[52]), .QN());
   DFF_X1 \N_reg[51]  (.D(n_1_67), .CK(n_1_2), .Q(N[51]), .QN());
   DFF_X1 \N_reg[50]  (.D(n_1_66), .CK(n_1_2), .Q(N[50]), .QN());
   DFF_X1 \N_reg[49]  (.D(n_1_65), .CK(n_1_2), .Q(N[49]), .QN());
   DFF_X1 \N_reg[48]  (.D(n_1_64), .CK(n_1_2), .Q(N[48]), .QN());
   DFF_X1 \N_reg[47]  (.D(n_1_63), .CK(n_1_2), .Q(N[47]), .QN());
   DFF_X1 \N_reg[46]  (.D(n_1_62), .CK(n_1_2), .Q(N[46]), .QN());
   DFF_X1 \N_reg[45]  (.D(n_1_61), .CK(n_1_2), .Q(N[45]), .QN());
   DFF_X1 \N_reg[44]  (.D(n_1_60), .CK(n_1_2), .Q(N[44]), .QN());
   DFF_X1 \N_reg[43]  (.D(n_1_59), .CK(n_1_2), .Q(N[43]), .QN());
   DFF_X1 \N_reg[42]  (.D(n_1_58), .CK(n_1_2), .Q(N[42]), .QN());
   DFF_X1 \N_reg[41]  (.D(n_1_57), .CK(n_1_2), .Q(N[41]), .QN());
   DFF_X1 \N_reg[40]  (.D(n_1_56), .CK(n_1_2), .Q(N[40]), .QN());
   DFF_X1 \N_reg[39]  (.D(n_1_55), .CK(n_1_2), .Q(N[39]), .QN());
   DFF_X1 \N_reg[38]  (.D(n_1_54), .CK(n_1_2), .Q(N[38]), .QN());
   DFF_X1 \N_reg[37]  (.D(n_1_53), .CK(n_1_2), .Q(N[37]), .QN());
   DFF_X1 \N_reg[36]  (.D(n_1_52), .CK(n_1_2), .Q(N[36]), .QN());
   DFF_X1 \N_reg[35]  (.D(n_1_51), .CK(n_1_2), .Q(N[35]), .QN());
   DFF_X1 \N_reg[34]  (.D(n_1_50), .CK(n_1_2), .Q(N[34]), .QN());
   DFF_X1 \N_reg[33]  (.D(n_1_49), .CK(n_1_2), .Q(N[33]), .QN());
   DFF_X1 \N_reg[32]  (.D(n_1_48), .CK(n_1_2), .Q(N[32]), .QN());
   DFF_X1 \N_reg[31]  (.D(n_1_47), .CK(n_1_2), .Q(N[31]), .QN());
   DFF_X1 \N_reg[30]  (.D(n_1_46), .CK(n_1_2), .Q(N[30]), .QN());
   DFF_X1 \N_reg[29]  (.D(n_1_45), .CK(n_1_2), .Q(N[29]), .QN());
   DFF_X1 \N_reg[28]  (.D(n_1_44), .CK(n_1_2), .Q(N[28]), .QN());
   DFF_X1 \N_reg[27]  (.D(n_1_43), .CK(n_1_2), .Q(N[27]), .QN());
   DFF_X1 \N_reg[26]  (.D(n_1_42), .CK(n_1_2), .Q(N[26]), .QN());
   DFF_X1 \N_reg[25]  (.D(n_1_41), .CK(n_1_2), .Q(N[25]), .QN());
   DFF_X1 \N_reg[24]  (.D(n_1_40), .CK(n_1_2), .Q(N[24]), .QN());
   DFF_X1 \N_reg[23]  (.D(n_1_39), .CK(n_1_2), .Q(N[23]), .QN());
   DFF_X1 \N_reg[22]  (.D(n_1_38), .CK(n_1_2), .Q(N[22]), .QN());
   DFF_X1 \N_reg[21]  (.D(n_1_37), .CK(n_1_2), .Q(N[21]), .QN());
   DFF_X1 \N_reg[20]  (.D(n_1_36), .CK(n_1_2), .Q(N[20]), .QN());
   DFF_X1 \N_reg[19]  (.D(n_1_35), .CK(n_1_2), .Q(N[19]), .QN());
   DFF_X1 \N_reg[18]  (.D(n_1_34), .CK(n_1_2), .Q(N[18]), .QN());
   DFF_X1 \N_reg[17]  (.D(n_1_33), .CK(n_1_2), .Q(N[17]), .QN());
   DFF_X1 \N_reg[16]  (.D(n_1_32), .CK(n_1_2), .Q(N[16]), .QN());
   DFF_X1 \N_reg[15]  (.D(n_1_31), .CK(n_1_2), .Q(N[15]), .QN());
   DFF_X1 \N_reg[14]  (.D(n_1_30), .CK(n_1_2), .Q(N[14]), .QN());
   DFF_X1 \N_reg[13]  (.D(n_1_29), .CK(n_1_2), .Q(N[13]), .QN());
   DFF_X1 \N_reg[12]  (.D(n_1_28), .CK(n_1_2), .Q(N[12]), .QN());
   DFF_X1 \N_reg[11]  (.D(n_1_27), .CK(n_1_2), .Q(N[11]), .QN());
   DFF_X1 \N_reg[10]  (.D(n_1_26), .CK(n_1_2), .Q(N[10]), .QN());
   DFF_X1 \N_reg[9]  (.D(n_1_25), .CK(n_1_2), .Q(N[9]), .QN());
   DFF_X1 \N_reg[8]  (.D(n_1_24), .CK(n_1_2), .Q(N[8]), .QN());
   DFF_X1 \N_reg[7]  (.D(n_1_23), .CK(n_1_2), .Q(N[7]), .QN());
   DFF_X1 \N_reg[6]  (.D(n_1_22), .CK(n_1_2), .Q(N[6]), .QN());
   DFF_X1 \N_reg[5]  (.D(n_1_21), .CK(n_1_2), .Q(N[5]), .QN());
   DFF_X1 \N_reg[4]  (.D(n_1_20), .CK(n_1_2), .Q(N[4]), .QN());
   DFF_X1 \N_reg[3]  (.D(n_1_19), .CK(n_1_2), .Q(N[3]), .QN());
   DFF_X1 \N_reg[2]  (.D(n_1_18), .CK(n_1_2), .Q(N[2]), .QN());
   DFF_X1 \N_reg[1]  (.D(n_1_17), .CK(n_1_2), .Q(N[1]), .QN());
   DFF_X1 \N_reg[0]  (.D(n_1_16), .CK(n_1_2), .Q(N[0]), .QN());
   DFF_X1 division_operation_reg (.D(n_1_82), .CK(CLK), .Q(division_operation), 
      .QN());
   CLKGATETST_X1 clk_gate_in11_reg (.CK(CLK), .E(n_236), .SE(1'b0), .GCK(n_1_3));
   DFF_X1 \in11_reg[15]  (.D(n_1_147), .CK(n_1_3), .Q(in11[15]), .QN());
   DFF_X1 \in11_reg[14]  (.D(n_1_146), .CK(n_1_3), .Q(in11[14]), .QN());
   DFF_X1 \in11_reg[13]  (.D(n_1_145), .CK(n_1_3), .Q(in11[13]), .QN());
   DFF_X1 \in11_reg[12]  (.D(n_1_144), .CK(n_1_3), .Q(in11[12]), .QN());
   DFF_X1 \in11_reg[11]  (.D(n_1_143), .CK(n_1_3), .Q(in11[11]), .QN());
   DFF_X1 \in11_reg[10]  (.D(n_1_142), .CK(n_1_3), .Q(in11[10]), .QN());
   DFF_X1 \in11_reg[9]  (.D(n_1_141), .CK(n_1_3), .Q(in11[9]), .QN());
   DFF_X1 \in11_reg[8]  (.D(n_1_140), .CK(n_1_3), .Q(in11[8]), .QN());
   DFF_X1 \in11_reg[7]  (.D(n_1_139), .CK(n_1_3), .Q(in11[7]), .QN());
   DFF_X1 \in11_reg[6]  (.D(n_1_138), .CK(n_1_3), .Q(in11[6]), .QN());
   DFF_X1 \in11_reg[5]  (.D(n_1_137), .CK(n_1_3), .Q(in11[5]), .QN());
   DFF_X1 \in11_reg[4]  (.D(n_1_136), .CK(n_1_3), .Q(in11[4]), .QN());
   DFF_X1 \in11_reg[3]  (.D(n_1_135), .CK(n_1_3), .Q(in11[3]), .QN());
   DFF_X1 \in11_reg[2]  (.D(n_1_134), .CK(n_1_3), .Q(in11[2]), .QN());
   DFF_X1 \in11_reg[1]  (.D(n_1_133), .CK(n_1_3), .Q(in11[1]), .QN());
   DFF_X1 \in11_reg[0]  (.D(n_1_132), .CK(n_1_3), .Q(in11[0]), .QN());
   CLKGATETST_X1 clk_gate_second_operand_reg (.CK(CLK), .E(n_1_115), .SE(1'b0), 
      .GCK(n_1_4));
   OAI22_X1 i_1_1_0 (.A1(n_1_1_0), .A2(n_1_1_460), .B1(n_1_1_480), .B2(n_1_1_595), 
      .ZN(n_0));
   NOR3_X1 i_1_1_1 (.A1(n_312), .A2(n_311), .A3(n_1_1_545), .ZN(n_1_1_0));
   OAI21_X1 i_1_1_2 (.A(n_1_1_7), .B1(n_1_1_5), .B2(n_1_1_1), .ZN(n_1));
   NAND3_X1 i_1_1_3 (.A1(n_1_1_2), .A2(n_1_1_3), .A3(n_1_1_94), .ZN(n_1_1_1));
   AOI21_X1 i_1_1_4 (.A(n_1_1_23), .B1(n_1_1_4), .B2(n_1_1_254), .ZN(n_1_1_2));
   OAI21_X1 i_1_1_5 (.A(n_1_1_609), .B1(n_1_1_608), .B2(NextState[0]), .ZN(
      n_1_1_3));
   OAI21_X1 i_1_1_6 (.A(n_1_1_610), .B1(n_1_1_251), .B2(n_1_1_244), .ZN(n_1_1_4));
   AOI211_X1 i_1_1_7 (.A(NextState[2]), .B(n_1_1_533), .C1(n_1_1_6), .C2(n_312), 
      .ZN(n_1_1_5));
   NOR2_X1 i_1_1_8 (.A1(n_1_1_261), .A2(division_operation), .ZN(n_1_1_6));
   OAI21_X1 i_1_1_9 (.A(n_1_1_605), .B1(n_1_1_30), .B2(n_1_1_8), .ZN(n_1_1_7));
   NOR4_X1 i_1_1_10 (.A1(n_1_1_588), .A2(n_1_1_586), .A3(n_1_1_546), .A4(n_1_1_9), 
      .ZN(n_1_1_8));
   NAND4_X1 i_1_1_11 (.A1(n_1_1_13), .A2(n_1_1_12), .A3(n_1_1_11), .A4(n_1_1_10), 
      .ZN(n_1_1_9));
   NOR4_X1 i_1_1_12 (.A1(RAM_Data_RD_A[2]), .A2(n_1_1_626), .A3(RAM_Data_RD_A[1]), 
      .A4(RAM_Data_RD_A[3]), .ZN(n_1_1_10));
   NOR4_X1 i_1_1_13 (.A1(RAM_Data_RD_A[7]), .A2(RAM_Data_RD_A[6]), .A3(
      RAM_Data_RD_A[5]), .A4(RAM_Data_RD_A[4]), .ZN(n_1_1_11));
   NOR4_X1 i_1_1_14 (.A1(RAM_Data_RD_A[11]), .A2(RAM_Data_RD_A[10]), .A3(
      RAM_Data_RD_A[9]), .A4(RAM_Data_RD_A[8]), .ZN(n_1_1_12));
   NOR4_X1 i_1_1_15 (.A1(RAM_Data_RD_A[15]), .A2(RAM_Data_RD_A[14]), .A3(
      RAM_Data_RD_A[13]), .A4(RAM_Data_RD_A[12]), .ZN(n_1_1_13));
   OAI21_X1 i_1_1_25 (.A(n_1_1_610), .B1(n_1_1_249), .B2(n_1_1_243), .ZN(
      n_1_1_21));
   AOI21_X1 i_1_1_26 (.A(NextState[2]), .B1(n_1_1_584), .B2(NextState[3]), 
      .ZN(n_1_1_22));
   NAND2_X1 i_1_1_28 (.A1(n_1_1_598), .A2(n_1_1_96), .ZN(n_1_1_24));
   OAI22_X1 i_1_1_29 (.A1(n_1_1_26), .A2(n_1_1_25), .B1(n_1_1_159), .B2(n_1_1_29), 
      .ZN(n_2));
   AOI21_X1 i_1_1_30 (.A(NextState[3]), .B1(NextState[2]), .B2(n_1_1_533), 
      .ZN(n_1_1_25));
   NOR2_X1 i_1_1_32 (.A1(n_1_1_29), .A2(n_1_1_28), .ZN(n_1_1_27));
   NOR2_X1 i_1_1_33 (.A1(n_1_1_586), .A2(n_1_1_533), .ZN(n_1_1_28));
   AOI22_X1 i_1_1_35 (.A1(n_1_1_485), .A2(n_1_1_31), .B1(Euler_End), .B2(
      n_1_1_585), .ZN(n_1_1_30));
   AOI22_X1 i_1_1_36 (.A1(n_1_1_32), .A2(n_1_1_587), .B1(n_1_1_544), .B2(
      n_1_1_482), .ZN(n_1_1_31));
   OAI21_X1 i_1_1_37 (.A(NextState[1]), .B1(n_1_1_606), .B2(n_1_1_54), .ZN(
      n_1_1_32));
   NOR3_X1 i_1_1_38 (.A1(n_1_1_272), .A2(n_1_1_54), .A3(RST), .ZN(n_1_6));
   AOI22_X1 i_1_1_39 (.A1(n_1_1_268), .A2(n_1_1_485), .B1(n_1_1_605), .B2(
      n_1_1_271), .ZN(n_1_7));
   AND2_X1 i_1_1_40 (.A1(n_1_1_33), .A2(adder_out1[0]), .ZN(n_3));
   AND2_X1 i_1_1_41 (.A1(n_1_1_33), .A2(adder_out1[1]), .ZN(n_4));
   AND2_X1 i_1_1_42 (.A1(n_1_1_33), .A2(adder_out1[2]), .ZN(n_5));
   AND2_X1 i_1_1_43 (.A1(n_1_1_33), .A2(adder_out1[3]), .ZN(n_6));
   AND2_X1 i_1_1_44 (.A1(n_1_1_33), .A2(adder_out1[4]), .ZN(n_7));
   AND2_X1 i_1_1_45 (.A1(n_1_1_33), .A2(adder_out1[5]), .ZN(n_8));
   AND2_X1 i_1_1_46 (.A1(n_1_1_33), .A2(adder_out1[6]), .ZN(n_9));
   AND2_X1 i_1_1_47 (.A1(n_1_1_33), .A2(adder_out1[7]), .ZN(n_10));
   AND2_X1 i_1_1_48 (.A1(n_1_1_33), .A2(adder_out1[8]), .ZN(n_11));
   AND2_X1 i_1_1_49 (.A1(n_1_1_33), .A2(adder_out1[9]), .ZN(n_12));
   AND2_X1 i_1_1_50 (.A1(n_1_1_33), .A2(adder_out1[10]), .ZN(n_13));
   AND2_X1 i_1_1_51 (.A1(n_1_1_33), .A2(adder_out1[11]), .ZN(n_14));
   AND2_X1 i_1_1_52 (.A1(n_1_1_33), .A2(adder_out1[12]), .ZN(n_15));
   AND2_X1 i_1_1_53 (.A1(n_1_1_33), .A2(adder_out1[13]), .ZN(n_16));
   AND2_X1 i_1_1_54 (.A1(n_1_1_33), .A2(adder_out1[14]), .ZN(n_17));
   AND2_X1 i_1_1_55 (.A1(n_1_1_33), .A2(adder_out1[15]), .ZN(n_18));
   AOI21_X1 i_1_1_56 (.A(RST), .B1(n_1_1_590), .B2(n_1_1_530), .ZN(n_1_1_33));
   AOI21_X1 i_1_1_57 (.A(RST), .B1(n_1_1_241), .B2(n_1_1_224), .ZN(n_19));
   NOR2_X1 i_1_1_58 (.A1(n_1_1_606), .A2(RST), .ZN(n_1_11));
   NAND3_X1 i_1_1_59 (.A1(n_1_1_251), .A2(n_1_1_605), .A3(n_1_1_254), .ZN(n_1_15));
   OAI22_X1 i_1_1_60 (.A1(n_1_1_460), .A2(n_1_1_34), .B1(n_1_1_239), .B2(
      n_1_1_249), .ZN(n_20));
   AOI21_X1 i_1_1_61 (.A(n_1_1_603), .B1(n_311), .B2(n_1_1_604), .ZN(n_1_1_34));
   OAI21_X1 i_1_1_62 (.A(n_1_1_35), .B1(n_1_1_248), .B2(n_1_1_239), .ZN(n_21));
   NAND2_X1 i_1_1_63 (.A1(n_1_1_461), .A2(n_1_1_36), .ZN(n_1_1_35));
   AOI21_X1 i_1_1_64 (.A(n_1_1_603), .B1(n_311), .B2(division_operation), 
      .ZN(n_1_1_36));
   AND2_X1 i_1_1_65 (.A1(adder_out2[0]), .A2(n_183), .ZN(n_22));
   AND2_X1 i_1_1_66 (.A1(adder_out2[1]), .A2(n_183), .ZN(n_23));
   AND2_X1 i_1_1_67 (.A1(adder_out2[2]), .A2(n_183), .ZN(n_24));
   AND2_X1 i_1_1_68 (.A1(adder_out2[3]), .A2(n_183), .ZN(n_25));
   AND2_X1 i_1_1_69 (.A1(adder_out2[4]), .A2(n_183), .ZN(n_26));
   AND2_X1 i_1_1_70 (.A1(adder_out2[5]), .A2(n_183), .ZN(n_27));
   AND2_X1 i_1_1_71 (.A1(adder_out2[6]), .A2(n_183), .ZN(n_28));
   AND2_X1 i_1_1_72 (.A1(adder_out2[7]), .A2(n_183), .ZN(n_29));
   AND2_X1 i_1_1_73 (.A1(adder_out2[8]), .A2(n_183), .ZN(n_30));
   AND2_X1 i_1_1_74 (.A1(adder_out2[9]), .A2(n_183), .ZN(n_31));
   AND2_X1 i_1_1_75 (.A1(adder_out2[10]), .A2(n_183), .ZN(n_32));
   AND2_X1 i_1_1_76 (.A1(adder_out2[11]), .A2(n_183), .ZN(n_33));
   AND2_X1 i_1_1_77 (.A1(adder_out2[12]), .A2(n_183), .ZN(n_34));
   AND2_X1 i_1_1_78 (.A1(adder_out2[13]), .A2(n_183), .ZN(n_35));
   AND2_X1 i_1_1_79 (.A1(adder_out2[14]), .A2(n_183), .ZN(n_36));
   AND2_X1 i_1_1_80 (.A1(adder_out2[15]), .A2(n_183), .ZN(n_37));
   OAI21_X1 i_1_1_82 (.A(n_1_1_38), .B1(n_1_1_37), .B2(n_1_1_480), .ZN(n_38));
   AOI21_X1 i_1_1_83 (.A(n_1_1_596), .B1(n_1_1_589), .B2(count[0]), .ZN(n_1_1_37));
   OAI211_X1 i_1_1_84 (.A(n_1_1_594), .B(n_1_1_479), .C1(Errortemp[0]), .C2(
      n_1_1_607), .ZN(n_1_1_38));
   INV_X1 i_1_1_85 (.A(n_1_1_39), .ZN(n_39));
   AOI221_X1 i_1_1_86 (.A(n_183), .B1(n_1_1_187), .B2(Errortemp[1]), .C1(
      n_1_1_145), .C2(count[1]), .ZN(n_1_1_39));
   INV_X1 i_1_1_87 (.A(n_1_1_40), .ZN(n_40));
   AOI22_X1 i_1_1_88 (.A1(Errortemp[2]), .A2(n_1_1_187), .B1(n_1_1_145), 
      .B2(count[2]), .ZN(n_1_1_40));
   NAND2_X1 i_1_1_89 (.A1(n_1_1_43), .A2(n_1_1_41), .ZN(n_41));
   AOI22_X1 i_1_1_90 (.A1(Errortemp[3]), .A2(n_1_1_187), .B1(n_1_1_145), 
      .B2(count[3]), .ZN(n_1_1_41));
   INV_X1 i_1_1_91 (.A(n_1_1_42), .ZN(n_42));
   AOI221_X1 i_1_1_92 (.A(n_1_5), .B1(n_1_1_187), .B2(Errortemp[4]), .C1(
      n_1_1_145), .C2(count[4]), .ZN(n_1_1_42));
   NAND2_X1 i_1_1_93 (.A1(n_1_1_44), .A2(n_1_1_43), .ZN(n_43));
   AOI21_X1 i_1_1_94 (.A(n_1_5), .B1(n_1_1_268), .B2(n_1_1_222), .ZN(n_1_1_43));
   AOI22_X1 i_1_1_95 (.A1(Errortemp[5]), .A2(n_1_1_187), .B1(n_1_1_145), 
      .B2(count[5]), .ZN(n_1_1_44));
   INV_X1 i_1_1_96 (.A(n_1_1_45), .ZN(n_44));
   AOI222_X1 i_1_1_97 (.A1(Errortemp[6]), .A2(n_1_1_187), .B1(n_1_1_145), 
      .B2(count[6]), .C1(n_1_1_268), .C2(n_1_1_222), .ZN(n_1_1_45));
   INV_X1 i_1_1_98 (.A(n_1_1_46), .ZN(n_45));
   AOI22_X1 i_1_1_99 (.A1(Errortemp[7]), .A2(n_1_1_187), .B1(n_1_1_145), 
      .B2(count[7]), .ZN(n_1_1_46));
   INV_X1 i_1_1_100 (.A(n_1_1_47), .ZN(n_46));
   AOI22_X1 i_1_1_101 (.A1(Errortemp[8]), .A2(n_1_1_187), .B1(n_1_1_145), 
      .B2(count[8]), .ZN(n_1_1_47));
   INV_X1 i_1_1_102 (.A(n_1_1_48), .ZN(n_47));
   AOI22_X1 i_1_1_103 (.A1(Errortemp[9]), .A2(n_1_1_187), .B1(n_1_1_145), 
      .B2(count[9]), .ZN(n_1_1_48));
   INV_X1 i_1_1_104 (.A(n_1_1_49), .ZN(n_48));
   AOI22_X1 i_1_1_105 (.A1(Errortemp[10]), .A2(n_1_1_187), .B1(n_1_1_145), 
      .B2(count[10]), .ZN(n_1_1_49));
   INV_X1 i_1_1_106 (.A(n_1_1_50), .ZN(n_49));
   AOI22_X1 i_1_1_107 (.A1(Errortemp[11]), .A2(n_1_1_187), .B1(n_1_1_145), 
      .B2(count[11]), .ZN(n_1_1_50));
   INV_X1 i_1_1_108 (.A(n_1_1_51), .ZN(n_50));
   AOI22_X1 i_1_1_109 (.A1(Errortemp[12]), .A2(n_1_1_187), .B1(n_1_1_145), 
      .B2(count[12]), .ZN(n_1_1_51));
   NOR3_X1 i_1_1_110 (.A1(n_1_1_623), .A2(n_1_1_590), .A3(RST), .ZN(n_51));
   NOR3_X1 i_1_1_111 (.A1(n_1_1_624), .A2(n_1_1_590), .A3(RST), .ZN(n_52));
   NOR3_X1 i_1_1_112 (.A1(n_1_1_625), .A2(n_1_1_590), .A3(RST), .ZN(n_53));
   AND2_X1 i_1_1_113 (.A1(adder_out2[0]), .A2(n_1_1_52), .ZN(n_54));
   AND2_X1 i_1_1_114 (.A1(adder_out2[1]), .A2(n_1_1_52), .ZN(n_55));
   AND2_X1 i_1_1_115 (.A1(adder_out2[2]), .A2(n_1_1_52), .ZN(n_56));
   AND2_X1 i_1_1_116 (.A1(adder_out2[3]), .A2(n_1_1_52), .ZN(n_57));
   AND2_X1 i_1_1_117 (.A1(adder_out2[4]), .A2(n_1_1_52), .ZN(n_58));
   AND2_X1 i_1_1_118 (.A1(adder_out2[5]), .A2(n_1_1_52), .ZN(n_59));
   AND2_X1 i_1_1_119 (.A1(adder_out2[6]), .A2(n_1_1_52), .ZN(n_60));
   AND2_X1 i_1_1_120 (.A1(adder_out2[7]), .A2(n_1_1_52), .ZN(n_61));
   AND2_X1 i_1_1_121 (.A1(adder_out2[8]), .A2(n_1_1_52), .ZN(n_62));
   AND2_X1 i_1_1_122 (.A1(adder_out2[9]), .A2(n_1_1_52), .ZN(n_63));
   AND2_X1 i_1_1_123 (.A1(adder_out2[10]), .A2(n_1_1_52), .ZN(n_64));
   AND2_X1 i_1_1_124 (.A1(adder_out2[11]), .A2(n_1_1_52), .ZN(n_65));
   AND2_X1 i_1_1_125 (.A1(adder_out2[12]), .A2(n_1_1_52), .ZN(n_66));
   AOI21_X1 i_1_1_126 (.A(n_1_1_267), .B1(n_1_1_241), .B2(n_1_1_475), .ZN(
      n_1_1_52));
   INV_X1 i_1_1_127 (.A(n_1_1_53), .ZN(n_67));
   AOI211_X1 i_1_1_128 (.A(RST), .B(n_1_1_189), .C1(n_1_1_54), .C2(n_1_1_476), 
      .ZN(n_1_1_53));
   NAND2_X1 i_1_1_129 (.A1(n_1_1_599), .A2(hstate[0]), .ZN(n_1_1_54));
   NOR2_X1 i_1_1_133 (.A1(n_1_1_626), .A2(RST), .ZN(n_1_16));
   NOR2_X1 i_1_1_134 (.A1(n_1_1_628), .A2(RST), .ZN(n_1_18));
   NOR2_X1 i_1_1_135 (.A1(n_1_1_630), .A2(RST), .ZN(n_1_20));
   NOR2_X1 i_1_1_136 (.A1(n_1_1_633), .A2(RST), .ZN(n_1_23));
   NOR2_X1 i_1_1_137 (.A1(n_1_1_634), .A2(RST), .ZN(n_1_24));
   NOR2_X1 i_1_1_138 (.A1(n_1_1_635), .A2(RST), .ZN(n_1_25));
   NOR2_X1 i_1_1_139 (.A1(n_1_1_636), .A2(RST), .ZN(n_1_26));
   NOR2_X1 i_1_1_140 (.A1(n_1_1_637), .A2(RST), .ZN(n_1_27));
   NOR2_X1 i_1_1_141 (.A1(n_1_1_638), .A2(RST), .ZN(n_1_28));
   INV_X1 i_1_1_142 (.A(n_1_1_57), .ZN(n_1_80));
   AOI21_X1 i_1_1_143 (.A(RST), .B1(n_1_1_587), .B2(n_1_1_533), .ZN(n_1_1_57));
   NAND3_X1 i_1_1_144 (.A1(n_1_1_486), .A2(n_1_1_261), .A3(n_1_1_58), .ZN(n_68));
   NOR2_X1 i_1_1_146 (.A1(n_1_1_95), .A2(RST), .ZN(n_1_8));
   NAND3_X1 i_1_1_147 (.A1(n_1_1_485), .A2(n_1_1_59), .A3(n_1_1_58), .ZN(n_1_9));
   AOI21_X1 i_1_1_148 (.A(RST), .B1(ready), .B2(n_1_1_96), .ZN(n_1_1_58));
   NAND2_X1 i_1_1_149 (.A1(n_1_1_254), .A2(n_1_1_251), .ZN(n_1_1_59));
   INV_X1 i_1_1_150 (.A(n_1_1_60), .ZN(n_1_83));
   AOI221_X1 i_1_1_151 (.A(RST), .B1(out[0]), .B2(n_1_1_582), .C1(n_1_1_531), 
      .C2(htemp[0]), .ZN(n_1_1_60));
   INV_X1 i_1_1_152 (.A(n_1_1_61), .ZN(n_1_84));
   AOI22_X1 i_1_1_153 (.A1(out[1]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[1]), 
      .ZN(n_1_1_61));
   INV_X1 i_1_1_154 (.A(n_1_1_62), .ZN(n_1_85));
   AOI22_X1 i_1_1_155 (.A1(out[2]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[2]), 
      .ZN(n_1_1_62));
   INV_X1 i_1_1_156 (.A(n_1_1_63), .ZN(n_1_86));
   AOI22_X1 i_1_1_157 (.A1(out[3]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[3]), 
      .ZN(n_1_1_63));
   INV_X1 i_1_1_158 (.A(n_1_1_64), .ZN(n_1_87));
   AOI22_X1 i_1_1_159 (.A1(out[4]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[4]), 
      .ZN(n_1_1_64));
   INV_X1 i_1_1_160 (.A(n_1_1_65), .ZN(n_1_88));
   AOI22_X1 i_1_1_161 (.A1(out[5]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[5]), 
      .ZN(n_1_1_65));
   INV_X1 i_1_1_162 (.A(n_1_1_66), .ZN(n_1_89));
   AOI22_X1 i_1_1_163 (.A1(out[6]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[6]), 
      .ZN(n_1_1_66));
   INV_X1 i_1_1_164 (.A(n_1_1_67), .ZN(n_1_90));
   AOI22_X1 i_1_1_165 (.A1(out[7]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[7]), 
      .ZN(n_1_1_67));
   INV_X1 i_1_1_166 (.A(n_1_1_68), .ZN(n_1_91));
   AOI22_X1 i_1_1_167 (.A1(out[8]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[8]), 
      .ZN(n_1_1_68));
   INV_X1 i_1_1_168 (.A(n_1_1_69), .ZN(n_1_92));
   AOI22_X1 i_1_1_169 (.A1(out[9]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[9]), 
      .ZN(n_1_1_69));
   INV_X1 i_1_1_170 (.A(n_1_1_70), .ZN(n_1_93));
   AOI22_X1 i_1_1_171 (.A1(out[10]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[10]), 
      .ZN(n_1_1_70));
   INV_X1 i_1_1_172 (.A(n_1_1_71), .ZN(n_1_94));
   AOI22_X1 i_1_1_173 (.A1(out[11]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[11]), 
      .ZN(n_1_1_71));
   INV_X1 i_1_1_174 (.A(n_1_1_72), .ZN(n_1_95));
   AOI22_X1 i_1_1_175 (.A1(out[12]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[12]), 
      .ZN(n_1_1_72));
   INV_X1 i_1_1_176 (.A(n_1_1_73), .ZN(n_1_96));
   AOI22_X1 i_1_1_177 (.A1(out[13]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[13]), 
      .ZN(n_1_1_73));
   INV_X1 i_1_1_178 (.A(n_1_1_74), .ZN(n_1_97));
   AOI22_X1 i_1_1_179 (.A1(out[14]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[14]), 
      .ZN(n_1_1_74));
   INV_X1 i_1_1_180 (.A(n_1_1_75), .ZN(n_1_98));
   AOI22_X1 i_1_1_181 (.A1(out[15]), .A2(n_1_1_461), .B1(n_1_5), .B2(htemp[15]), 
      .ZN(n_1_1_75));
   INV_X1 i_1_1_182 (.A(n_1_1_76), .ZN(n_69));
   AOI222_X1 i_1_1_183 (.A1(RAM_Data_RD_A[0]), .A2(n_1_5), .B1(n_1_1_187), 
      .B2(adder_out1[0]), .C1(n_1_1_92), .C2(Q[0]), .ZN(n_1_1_76));
   INV_X1 i_1_1_184 (.A(n_1_1_77), .ZN(n_70));
   AOI222_X1 i_1_1_185 (.A1(adder_out1[1]), .A2(n_1_1_187), .B1(n_1_1_92), 
      .B2(Q[1]), .C1(n_1_17), .C2(n_1_1_531), .ZN(n_1_1_77));
   NOR2_X1 i_1_1_186 (.A1(n_1_1_627), .A2(RST), .ZN(n_1_17));
   INV_X1 i_1_1_187 (.A(n_1_1_78), .ZN(n_71));
   AOI222_X1 i_1_1_188 (.A1(RAM_Data_RD_A[2]), .A2(n_1_5), .B1(n_1_1_187), 
      .B2(adder_out1[2]), .C1(n_1_1_92), .C2(Q[2]), .ZN(n_1_1_78));
   INV_X1 i_1_1_189 (.A(n_1_1_79), .ZN(n_72));
   AOI222_X1 i_1_1_190 (.A1(adder_out1[3]), .A2(n_1_1_187), .B1(n_1_1_92), 
      .B2(Q[3]), .C1(n_1_19), .C2(n_1_1_531), .ZN(n_1_1_79));
   NOR2_X1 i_1_1_191 (.A1(n_1_1_629), .A2(RST), .ZN(n_1_19));
   INV_X1 i_1_1_192 (.A(n_1_1_80), .ZN(n_73));
   AOI222_X1 i_1_1_193 (.A1(RAM_Data_RD_A[4]), .A2(n_1_5), .B1(n_1_1_187), 
      .B2(adder_out1[4]), .C1(n_1_1_92), .C2(Q[4]), .ZN(n_1_1_80));
   INV_X1 i_1_1_194 (.A(n_1_1_81), .ZN(n_74));
   AOI222_X1 i_1_1_195 (.A1(adder_out1[5]), .A2(n_1_1_187), .B1(n_1_1_92), 
      .B2(Q[5]), .C1(n_1_21), .C2(n_1_1_531), .ZN(n_1_1_81));
   NOR2_X1 i_1_1_196 (.A1(n_1_1_631), .A2(RST), .ZN(n_1_21));
   INV_X1 i_1_1_197 (.A(n_1_1_82), .ZN(n_75));
   AOI222_X1 i_1_1_198 (.A1(adder_out1[6]), .A2(n_1_1_187), .B1(n_1_1_92), 
      .B2(Q[6]), .C1(n_1_22), .C2(n_1_1_531), .ZN(n_1_1_82));
   NOR2_X1 i_1_1_199 (.A1(n_1_1_632), .A2(RST), .ZN(n_1_22));
   INV_X1 i_1_1_200 (.A(n_1_1_83), .ZN(n_76));
   AOI222_X1 i_1_1_201 (.A1(RAM_Data_RD_A[7]), .A2(n_1_5), .B1(n_1_1_187), 
      .B2(adder_out1[7]), .C1(n_1_1_92), .C2(Q[7]), .ZN(n_1_1_83));
   INV_X1 i_1_1_202 (.A(n_1_1_84), .ZN(n_77));
   AOI222_X1 i_1_1_203 (.A1(RAM_Data_RD_A[8]), .A2(n_1_5), .B1(n_1_1_187), 
      .B2(adder_out1[8]), .C1(n_1_1_92), .C2(Q[8]), .ZN(n_1_1_84));
   INV_X1 i_1_1_204 (.A(n_1_1_85), .ZN(n_78));
   AOI222_X1 i_1_1_205 (.A1(RAM_Data_RD_A[9]), .A2(n_1_5), .B1(n_1_1_187), 
      .B2(adder_out1[9]), .C1(n_1_1_92), .C2(Q[9]), .ZN(n_1_1_85));
   INV_X1 i_1_1_206 (.A(n_1_1_86), .ZN(n_79));
   AOI222_X1 i_1_1_207 (.A1(RAM_Data_RD_A[10]), .A2(n_1_5), .B1(n_1_1_187), 
      .B2(adder_out1[10]), .C1(n_1_1_92), .C2(Q[10]), .ZN(n_1_1_86));
   INV_X1 i_1_1_208 (.A(n_1_1_87), .ZN(n_80));
   AOI222_X1 i_1_1_209 (.A1(RAM_Data_RD_A[11]), .A2(n_1_5), .B1(n_1_1_187), 
      .B2(adder_out1[11]), .C1(n_1_1_92), .C2(Q[11]), .ZN(n_1_1_87));
   INV_X1 i_1_1_210 (.A(n_1_1_88), .ZN(n_81));
   AOI222_X1 i_1_1_211 (.A1(RAM_Data_RD_A[12]), .A2(n_1_5), .B1(n_1_1_187), 
      .B2(adder_out1[12]), .C1(n_1_1_92), .C2(Q[12]), .ZN(n_1_1_88));
   NAND2_X1 i_1_1_212 (.A1(n_1_1_89), .A2(n_1_1_91), .ZN(n_82));
   AOI21_X1 i_1_1_213 (.A(n_163), .B1(n_1_5), .B2(RAM_Data_RD_A[13]), .ZN(
      n_1_1_89));
   NAND2_X1 i_1_1_214 (.A1(n_1_1_90), .A2(n_1_1_91), .ZN(n_83));
   AOI21_X1 i_1_1_215 (.A(n_164), .B1(n_1_5), .B2(RAM_Data_RD_A[14]), .ZN(
      n_1_1_90));
   NAND2_X1 i_1_1_216 (.A1(Q[14]), .A2(n_1_1_92), .ZN(n_1_1_91));
   NOR3_X1 i_1_1_217 (.A1(n_1_1_583), .A2(n_1_1_483), .A3(RST), .ZN(n_1_1_92));
   INV_X1 i_1_1_218 (.A(n_1_1_93), .ZN(n_84));
   AOI21_X1 i_1_1_219 (.A(n_165), .B1(n_1_5), .B2(RAM_Data_RD_A[15]), .ZN(
      n_1_1_93));
   AND2_X1 i_1_1_220 (.A1(n_1_1_531), .A2(n_1_32), .ZN(n_85));
   NOR2_X1 i_1_1_221 (.A1(n_1_1_642), .A2(RST), .ZN(n_1_32));
   AND2_X1 i_1_1_222 (.A1(n_1_1_531), .A2(n_1_33), .ZN(n_86));
   NOR2_X1 i_1_1_223 (.A1(n_1_1_643), .A2(RST), .ZN(n_1_33));
   AND2_X1 i_1_1_224 (.A1(n_1_1_531), .A2(n_1_34), .ZN(n_87));
   NOR2_X1 i_1_1_225 (.A1(n_1_1_644), .A2(RST), .ZN(n_1_34));
   AND2_X1 i_1_1_226 (.A1(n_1_1_531), .A2(n_1_35), .ZN(n_88));
   NOR2_X1 i_1_1_227 (.A1(n_1_1_645), .A2(RST), .ZN(n_1_35));
   AND2_X1 i_1_1_228 (.A1(n_1_1_531), .A2(n_1_36), .ZN(n_89));
   NOR2_X1 i_1_1_229 (.A1(n_1_1_646), .A2(RST), .ZN(n_1_36));
   AND2_X1 i_1_1_230 (.A1(n_1_1_531), .A2(n_1_37), .ZN(n_90));
   NOR2_X1 i_1_1_231 (.A1(n_1_1_647), .A2(RST), .ZN(n_1_37));
   AND2_X1 i_1_1_232 (.A1(n_1_1_531), .A2(n_1_38), .ZN(n_91));
   NOR2_X1 i_1_1_233 (.A1(n_1_1_648), .A2(RST), .ZN(n_1_38));
   AND2_X1 i_1_1_234 (.A1(n_1_1_531), .A2(n_1_39), .ZN(n_92));
   NOR2_X1 i_1_1_235 (.A1(n_1_1_649), .A2(RST), .ZN(n_1_39));
   AND2_X1 i_1_1_236 (.A1(n_1_1_531), .A2(n_1_40), .ZN(n_93));
   NOR2_X1 i_1_1_237 (.A1(n_1_1_650), .A2(RST), .ZN(n_1_40));
   AND2_X1 i_1_1_238 (.A1(n_1_1_531), .A2(n_1_41), .ZN(n_94));
   NOR2_X1 i_1_1_239 (.A1(n_1_1_651), .A2(RST), .ZN(n_1_41));
   AND2_X1 i_1_1_240 (.A1(n_1_1_531), .A2(n_1_42), .ZN(n_95));
   NOR2_X1 i_1_1_241 (.A1(n_1_1_652), .A2(RST), .ZN(n_1_42));
   AND2_X1 i_1_1_242 (.A1(n_1_1_531), .A2(n_1_43), .ZN(n_96));
   NOR2_X1 i_1_1_243 (.A1(n_1_1_653), .A2(RST), .ZN(n_1_43));
   AND2_X1 i_1_1_244 (.A1(n_1_1_531), .A2(n_1_44), .ZN(n_97));
   AND2_X1 i_1_1_245 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[28]), .ZN(n_1_44));
   AND2_X1 i_1_1_246 (.A1(n_1_1_531), .A2(n_1_45), .ZN(n_98));
   AND2_X1 i_1_1_247 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[29]), .ZN(n_1_45));
   AND2_X1 i_1_1_248 (.A1(n_1_1_531), .A2(n_1_46), .ZN(n_99));
   AND2_X1 i_1_1_249 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[30]), .ZN(n_1_46));
   AND2_X1 i_1_1_250 (.A1(n_1_1_531), .A2(n_1_47), .ZN(n_100));
   AND2_X1 i_1_1_251 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[31]), .ZN(n_1_47));
   AND2_X1 i_1_1_252 (.A1(n_1_1_531), .A2(n_1_48), .ZN(n_101));
   AND2_X1 i_1_1_253 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[32]), .ZN(n_1_48));
   AND2_X1 i_1_1_254 (.A1(n_1_1_531), .A2(n_1_49), .ZN(n_102));
   AND2_X1 i_1_1_255 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[33]), .ZN(n_1_49));
   AND2_X1 i_1_1_256 (.A1(n_1_1_531), .A2(n_1_50), .ZN(n_103));
   AND2_X1 i_1_1_257 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[34]), .ZN(n_1_50));
   AND2_X1 i_1_1_258 (.A1(n_1_1_531), .A2(n_1_51), .ZN(n_104));
   AND2_X1 i_1_1_259 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[35]), .ZN(n_1_51));
   AND2_X1 i_1_1_260 (.A1(n_1_1_531), .A2(n_1_52), .ZN(n_105));
   NOR2_X1 i_1_1_261 (.A1(n_1_1_654), .A2(RST), .ZN(n_1_52));
   AND2_X1 i_1_1_262 (.A1(n_1_1_531), .A2(n_1_53), .ZN(n_106));
   NOR2_X1 i_1_1_263 (.A1(n_1_1_655), .A2(RST), .ZN(n_1_53));
   AND2_X1 i_1_1_264 (.A1(n_1_1_531), .A2(n_1_54), .ZN(n_107));
   NOR2_X1 i_1_1_265 (.A1(n_1_1_656), .A2(RST), .ZN(n_1_54));
   AND2_X1 i_1_1_266 (.A1(n_1_1_531), .A2(n_1_55), .ZN(n_108));
   NOR2_X1 i_1_1_267 (.A1(n_1_1_657), .A2(RST), .ZN(n_1_55));
   AND2_X1 i_1_1_268 (.A1(n_1_1_531), .A2(n_1_56), .ZN(n_109));
   AND2_X1 i_1_1_269 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[40]), .ZN(n_1_56));
   AND2_X1 i_1_1_270 (.A1(n_1_1_531), .A2(n_1_57), .ZN(n_110));
   AND2_X1 i_1_1_271 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[41]), .ZN(n_1_57));
   AND2_X1 i_1_1_272 (.A1(n_1_1_531), .A2(n_1_58), .ZN(n_111));
   AND2_X1 i_1_1_273 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[42]), .ZN(n_1_58));
   AND2_X1 i_1_1_274 (.A1(n_1_1_531), .A2(n_1_59), .ZN(n_112));
   AND2_X1 i_1_1_275 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[43]), .ZN(n_1_59));
   AND2_X1 i_1_1_276 (.A1(n_1_1_531), .A2(n_1_60), .ZN(n_113));
   AND2_X1 i_1_1_277 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[44]), .ZN(n_1_60));
   AND2_X1 i_1_1_278 (.A1(n_1_1_531), .A2(n_1_61), .ZN(n_114));
   AND2_X1 i_1_1_279 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[45]), .ZN(n_1_61));
   AND2_X1 i_1_1_280 (.A1(n_1_1_531), .A2(n_1_62), .ZN(n_115));
   AND2_X1 i_1_1_281 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[46]), .ZN(n_1_62));
   AND2_X1 i_1_1_282 (.A1(n_1_1_531), .A2(n_1_63), .ZN(n_116));
   AND2_X1 i_1_1_283 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[47]), .ZN(n_1_63));
   AND2_X1 i_1_1_284 (.A1(n_1_1_531), .A2(n_1_64), .ZN(n_117));
   AND2_X1 i_1_1_285 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[48]), .ZN(n_1_64));
   AND2_X1 i_1_1_286 (.A1(n_1_1_531), .A2(n_1_65), .ZN(n_118));
   AND2_X1 i_1_1_287 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[49]), .ZN(n_1_65));
   AND2_X1 i_1_1_288 (.A1(n_1_1_531), .A2(n_1_66), .ZN(n_119));
   AND2_X1 i_1_1_289 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[50]), .ZN(n_1_66));
   AND2_X1 i_1_1_290 (.A1(n_1_1_531), .A2(n_1_67), .ZN(n_120));
   AND2_X1 i_1_1_291 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[51]), .ZN(n_1_67));
   AND2_X1 i_1_1_292 (.A1(n_1_1_531), .A2(n_1_68), .ZN(n_121));
   AND2_X1 i_1_1_293 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[52]), .ZN(n_1_68));
   AND2_X1 i_1_1_294 (.A1(n_1_1_531), .A2(n_1_69), .ZN(n_122));
   AND2_X1 i_1_1_295 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[53]), .ZN(n_1_69));
   AND2_X1 i_1_1_296 (.A1(n_1_1_531), .A2(n_1_70), .ZN(n_123));
   AND2_X1 i_1_1_297 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[54]), .ZN(n_1_70));
   AND2_X1 i_1_1_298 (.A1(n_1_1_531), .A2(n_1_71), .ZN(n_124));
   AND2_X1 i_1_1_299 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[55]), .ZN(n_1_71));
   AND2_X1 i_1_1_300 (.A1(n_1_1_531), .A2(n_1_72), .ZN(n_125));
   AND2_X1 i_1_1_301 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[56]), .ZN(n_1_72));
   AND2_X1 i_1_1_302 (.A1(n_1_1_531), .A2(n_1_73), .ZN(n_126));
   AND2_X1 i_1_1_303 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[57]), .ZN(n_1_73));
   AND2_X1 i_1_1_304 (.A1(n_1_1_531), .A2(n_1_74), .ZN(n_127));
   AND2_X1 i_1_1_305 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[58]), .ZN(n_1_74));
   AND2_X1 i_1_1_306 (.A1(n_1_1_531), .A2(n_1_75), .ZN(n_128));
   AND2_X1 i_1_1_307 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[59]), .ZN(n_1_75));
   AND2_X1 i_1_1_308 (.A1(n_1_1_531), .A2(n_1_76), .ZN(n_129));
   AND2_X1 i_1_1_309 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[60]), .ZN(n_1_76));
   AND2_X1 i_1_1_310 (.A1(n_1_1_531), .A2(n_1_77), .ZN(n_130));
   AND2_X1 i_1_1_311 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[61]), .ZN(n_1_77));
   AND2_X1 i_1_1_312 (.A1(n_1_1_531), .A2(n_1_78), .ZN(n_131));
   AND2_X1 i_1_1_313 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[62]), .ZN(n_1_78));
   AND2_X1 i_1_1_314 (.A1(n_1_1_531), .A2(n_1_79), .ZN(n_132));
   AND2_X1 i_1_1_315 (.A1(n_1_1_605), .A2(RAM_Data_RD_A[63]), .ZN(n_1_79));
   NOR2_X1 i_1_1_322 (.A1(Temp[5]), .A2(Temp[4]), .ZN(n_1_1_98));
   NOR2_X1 i_1_1_323 (.A1(Temp[7]), .A2(Temp[6]), .ZN(n_1_1_99));
   NOR4_X1 i_1_1_324 (.A1(Temp[3]), .A2(Temp[2]), .A3(Temp[1]), .A4(Temp[0]), 
      .ZN(n_1_1_100));
   NOR4_X1 i_1_1_325 (.A1(n_1_1_103), .A2(n_1_1_102), .A3(Temp[13]), .A4(
      Temp[12]), .ZN(n_1_1_101));
   OR2_X1 i_1_1_326 (.A1(Temp[15]), .A2(Temp[14]), .ZN(n_1_1_102));
   OR4_X1 i_1_1_327 (.A1(Temp[11]), .A2(Temp[10]), .A3(Temp[9]), .A4(Temp[8]), 
      .ZN(n_1_1_103));
   INV_X1 i_1_1_328 (.A(n_1_1_104), .ZN(n_1_99));
   AOI21_X1 i_1_1_329 (.A(n_1_1_461), .B1(n_183), .B2(out[0]), .ZN(n_1_1_104));
   INV_X1 i_1_1_330 (.A(n_1_1_105), .ZN(n_1_100));
   AOI21_X1 i_1_1_331 (.A(n_1_1_461), .B1(n_183), .B2(out[1]), .ZN(n_1_1_105));
   AND2_X1 i_1_1_332 (.A1(out[2]), .A2(n_183), .ZN(n_1_101));
   AND2_X1 i_1_1_333 (.A1(out[3]), .A2(n_183), .ZN(n_1_102));
   INV_X1 i_1_1_334 (.A(n_1_1_106), .ZN(n_1_103));
   AOI21_X1 i_1_1_335 (.A(n_1_1_461), .B1(n_183), .B2(out[4]), .ZN(n_1_1_106));
   INV_X1 i_1_1_336 (.A(n_1_1_107), .ZN(n_1_104));
   AOI21_X1 i_1_1_337 (.A(n_1_1_461), .B1(n_183), .B2(out[5]), .ZN(n_1_1_107));
   INV_X1 i_1_1_338 (.A(n_1_1_108), .ZN(n_1_105));
   AOI21_X1 i_1_1_339 (.A(n_1_1_461), .B1(n_183), .B2(out[6]), .ZN(n_1_1_108));
   AND2_X1 i_1_1_340 (.A1(out[7]), .A2(n_183), .ZN(n_1_106));
   AND2_X1 i_1_1_341 (.A1(out[8]), .A2(n_183), .ZN(n_1_107));
   AND2_X1 i_1_1_342 (.A1(out[9]), .A2(n_183), .ZN(n_1_108));
   AND2_X1 i_1_1_343 (.A1(out[10]), .A2(n_183), .ZN(n_1_109));
   AND2_X1 i_1_1_344 (.A1(out[11]), .A2(n_183), .ZN(n_1_110));
   AND2_X1 i_1_1_345 (.A1(out[12]), .A2(n_183), .ZN(n_1_111));
   INV_X1 i_1_1_346 (.A(n_1_1_109), .ZN(n_1_112));
   AOI21_X1 i_1_1_347 (.A(n_1_1_461), .B1(n_183), .B2(out[13]), .ZN(n_1_1_109));
   INV_X1 i_1_1_348 (.A(n_1_1_110), .ZN(n_1_113));
   AOI21_X1 i_1_1_349 (.A(n_1_1_461), .B1(n_183), .B2(out[14]), .ZN(n_1_1_110));
   INV_X1 i_1_1_350 (.A(n_1_1_111), .ZN(n_1_114));
   AOI21_X1 i_1_1_351 (.A(n_1_1_461), .B1(n_183), .B2(out[15]), .ZN(n_1_1_111));
   INV_X1 i_1_1_353 (.A(n_1_1_112), .ZN(n_1_116));
   AOI22_X1 i_1_1_354 (.A1(RAM_Data_RD_A[0]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[0]), .ZN(n_1_1_112));
   INV_X1 i_1_1_355 (.A(n_1_1_113), .ZN(n_1_117));
   AOI22_X1 i_1_1_356 (.A1(RAM_Data_RD_A[1]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[1]), .ZN(n_1_1_113));
   INV_X1 i_1_1_357 (.A(n_1_1_114), .ZN(n_1_118));
   AOI22_X1 i_1_1_358 (.A1(RAM_Data_RD_A[2]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[2]), .ZN(n_1_1_114));
   INV_X1 i_1_1_359 (.A(n_1_1_115), .ZN(n_1_119));
   AOI22_X1 i_1_1_360 (.A1(RAM_Data_RD_A[3]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[3]), .ZN(n_1_1_115));
   INV_X1 i_1_1_361 (.A(n_1_1_116), .ZN(n_1_120));
   AOI22_X1 i_1_1_362 (.A1(RAM_Data_RD_A[4]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[4]), .ZN(n_1_1_116));
   INV_X1 i_1_1_363 (.A(n_1_1_117), .ZN(n_1_121));
   AOI22_X1 i_1_1_364 (.A1(RAM_Data_RD_A[5]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[5]), .ZN(n_1_1_117));
   INV_X1 i_1_1_365 (.A(n_1_1_118), .ZN(n_1_122));
   AOI22_X1 i_1_1_366 (.A1(RAM_Data_RD_A[6]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[6]), .ZN(n_1_1_118));
   INV_X1 i_1_1_367 (.A(n_1_1_119), .ZN(n_1_123));
   AOI22_X1 i_1_1_368 (.A1(RAM_Data_RD_A[7]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[7]), .ZN(n_1_1_119));
   INV_X1 i_1_1_369 (.A(n_1_1_120), .ZN(n_1_124));
   AOI22_X1 i_1_1_370 (.A1(RAM_Data_RD_A[8]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[8]), .ZN(n_1_1_120));
   INV_X1 i_1_1_371 (.A(n_1_1_121), .ZN(n_1_125));
   AOI22_X1 i_1_1_372 (.A1(RAM_Data_RD_A[9]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[9]), .ZN(n_1_1_121));
   INV_X1 i_1_1_373 (.A(n_1_1_122), .ZN(n_1_126));
   AOI22_X1 i_1_1_374 (.A1(RAM_Data_RD_A[10]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[10]), .ZN(n_1_1_122));
   INV_X1 i_1_1_375 (.A(n_1_1_123), .ZN(n_1_127));
   AOI22_X1 i_1_1_376 (.A1(RAM_Data_RD_A[11]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[11]), .ZN(n_1_1_123));
   INV_X1 i_1_1_377 (.A(n_1_1_124), .ZN(n_1_128));
   AOI22_X1 i_1_1_378 (.A1(RAM_Data_RD_A[12]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[12]), .ZN(n_1_1_124));
   INV_X1 i_1_1_379 (.A(n_1_1_125), .ZN(n_1_129));
   AOI22_X1 i_1_1_380 (.A1(RAM_Data_RD_A[13]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[13]), .ZN(n_1_1_125));
   INV_X1 i_1_1_381 (.A(n_1_1_126), .ZN(n_1_130));
   AOI22_X1 i_1_1_382 (.A1(RAM_Data_RD_A[14]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[14]), .ZN(n_1_1_126));
   INV_X1 i_1_1_383 (.A(n_1_1_127), .ZN(n_1_131));
   AOI22_X1 i_1_1_384 (.A1(RAM_Data_RD_A[15]), .A2(n_1_1_461), .B1(n_183), 
      .B2(RAM_Data_RD_B[15]), .ZN(n_1_1_127));
   OAI21_X1 i_1_1_385 (.A(n_1_1_605), .B1(n_1_1_563), .B2(n_1_1_546), .ZN(n_133));
   INV_X1 i_1_1_392 (.A(n_1_1_132), .ZN(n_134));
   AOI21_X1 i_1_1_393 (.A(RST), .B1(n_1_1_582), .B2(Errortemp[0]), .ZN(n_1_1_132));
   INV_X1 i_1_1_394 (.A(n_1_1_133), .ZN(n_135));
   AOI21_X1 i_1_1_395 (.A(n_1_5), .B1(n_1_1_461), .B2(Errortemp[1]), .ZN(
      n_1_1_133));
   NOR2_X1 i_1_1_396 (.A1(n_1_1_612), .A2(n_1_1_460), .ZN(n_136));
   NOR2_X1 i_1_1_397 (.A1(n_1_1_613), .A2(n_1_1_460), .ZN(n_137));
   NOR2_X1 i_1_1_398 (.A1(n_1_1_614), .A2(n_1_1_460), .ZN(n_138));
   NOR2_X1 i_1_1_399 (.A1(n_1_1_615), .A2(n_1_1_460), .ZN(n_139));
   NOR2_X1 i_1_1_400 (.A1(n_1_1_616), .A2(n_1_1_460), .ZN(n_140));
   NOR2_X1 i_1_1_401 (.A1(n_1_1_617), .A2(n_1_1_460), .ZN(n_141));
   NOR2_X1 i_1_1_402 (.A1(n_1_1_618), .A2(n_1_1_460), .ZN(n_142));
   NOR2_X1 i_1_1_403 (.A1(n_1_1_619), .A2(n_1_1_460), .ZN(n_143));
   NOR2_X1 i_1_1_404 (.A1(n_1_1_620), .A2(n_1_1_460), .ZN(n_144));
   NOR2_X1 i_1_1_405 (.A1(n_1_1_621), .A2(n_1_1_460), .ZN(n_145));
   NOR2_X1 i_1_1_406 (.A1(n_1_1_622), .A2(n_1_1_460), .ZN(n_146));
   NOR2_X1 i_1_1_407 (.A1(n_1_1_623), .A2(n_1_1_460), .ZN(n_147));
   NOR2_X1 i_1_1_408 (.A1(n_1_1_624), .A2(n_1_1_460), .ZN(n_148));
   NOR2_X1 i_1_1_409 (.A1(n_1_1_625), .A2(n_1_1_460), .ZN(n_149));
   AOI211_X1 i_1_1_410 (.A(n_1_1_478), .B(n_1_1_135), .C1(n_1_1_134), .C2(
      n_1_1_536), .ZN(n_150));
   OAI22_X1 i_1_1_411 (.A1(n_1_1_594), .A2(n_1_1_535), .B1(n_1_1_607), .B2(
      adder_out1[0]), .ZN(n_1_1_134));
   AOI211_X1 i_1_1_412 (.A(count[0]), .B(n_1_1_219), .C1(n_1_1_591), .C2(
      adder_out1[0]), .ZN(n_1_1_135));
   NAND2_X1 i_1_1_413 (.A1(n_1_1_137), .A2(n_1_1_136), .ZN(n_151));
   OAI21_X1 i_1_1_414 (.A(n_1_1_146), .B1(n_1_1_145), .B2(count[1]), .ZN(
      n_1_1_136));
   NAND2_X1 i_1_1_415 (.A1(adder_out1[1]), .A2(n_1_1_187), .ZN(n_1_1_137));
   INV_X1 i_1_1_416 (.A(n_1_1_138), .ZN(n_152));
   AOI22_X1 i_1_1_417 (.A1(n_1_1_154), .A2(count[2]), .B1(adder_out1[2]), 
      .B2(n_1_1_187), .ZN(n_1_1_138));
   NAND2_X1 i_1_1_418 (.A1(n_1_1_140), .A2(n_1_1_139), .ZN(n_153));
   OAI21_X1 i_1_1_419 (.A(n_1_1_146), .B1(n_1_1_145), .B2(count[3]), .ZN(
      n_1_1_139));
   NAND2_X1 i_1_1_420 (.A1(adder_out1[3]), .A2(n_1_1_187), .ZN(n_1_1_140));
   INV_X1 i_1_1_421 (.A(n_1_1_141), .ZN(n_154));
   AOI22_X1 i_1_1_422 (.A1(n_1_1_154), .A2(count[4]), .B1(adder_out1[4]), 
      .B2(n_1_1_187), .ZN(n_1_1_141));
   NAND2_X1 i_1_1_423 (.A1(n_1_1_143), .A2(n_1_1_142), .ZN(n_155));
   OAI21_X1 i_1_1_424 (.A(n_1_1_146), .B1(n_1_1_145), .B2(count[5]), .ZN(
      n_1_1_142));
   NAND2_X1 i_1_1_425 (.A1(adder_out1[5]), .A2(n_1_1_187), .ZN(n_1_1_143));
   NAND2_X1 i_1_1_426 (.A1(n_1_1_147), .A2(n_1_1_144), .ZN(n_156));
   OAI21_X1 i_1_1_427 (.A(n_1_1_146), .B1(n_1_1_145), .B2(count[6]), .ZN(
      n_1_1_144));
   NOR2_X1 i_1_1_428 (.A1(n_1_1_298), .A2(n_1_1_267), .ZN(n_1_1_145));
   OAI21_X1 i_1_1_429 (.A(n_1_1_155), .B1(n_1_1_480), .B2(n_1_1_584), .ZN(
      n_1_1_146));
   NAND2_X1 i_1_1_430 (.A1(adder_out1[6]), .A2(n_1_1_187), .ZN(n_1_1_147));
   INV_X1 i_1_1_431 (.A(n_1_1_148), .ZN(n_157));
   AOI22_X1 i_1_1_432 (.A1(n_1_1_154), .A2(count[7]), .B1(adder_out1[7]), 
      .B2(n_1_1_187), .ZN(n_1_1_148));
   INV_X1 i_1_1_433 (.A(n_1_1_149), .ZN(n_158));
   AOI22_X1 i_1_1_434 (.A1(n_1_1_154), .A2(count[8]), .B1(adder_out1[8]), 
      .B2(n_1_1_187), .ZN(n_1_1_149));
   INV_X1 i_1_1_435 (.A(n_1_1_150), .ZN(n_159));
   AOI22_X1 i_1_1_436 (.A1(n_1_1_154), .A2(count[9]), .B1(adder_out1[9]), 
      .B2(n_1_1_187), .ZN(n_1_1_150));
   INV_X1 i_1_1_437 (.A(n_1_1_151), .ZN(n_160));
   AOI22_X1 i_1_1_438 (.A1(n_1_1_154), .A2(count[10]), .B1(adder_out1[10]), 
      .B2(n_1_1_187), .ZN(n_1_1_151));
   INV_X1 i_1_1_439 (.A(n_1_1_152), .ZN(n_161));
   AOI22_X1 i_1_1_440 (.A1(n_1_1_154), .A2(count[11]), .B1(adder_out1[11]), 
      .B2(n_1_1_187), .ZN(n_1_1_152));
   INV_X1 i_1_1_441 (.A(n_1_1_153), .ZN(n_162));
   AOI22_X1 i_1_1_442 (.A1(n_1_1_154), .A2(count[12]), .B1(adder_out1[12]), 
      .B2(n_1_1_187), .ZN(n_1_1_153));
   OAI21_X1 i_1_1_443 (.A(n_1_1_155), .B1(n_1_1_480), .B2(NextState[0]), 
      .ZN(n_1_1_154));
   AOI21_X1 i_1_1_444 (.A(n_1_1_156), .B1(n_1_1_157), .B2(n_1_1_596), .ZN(
      n_1_1_155));
   NOR2_X1 i_1_1_445 (.A1(n_1_1_299), .A2(RST), .ZN(n_1_1_156));
   NOR2_X1 i_1_1_446 (.A1(n_1_1_243), .A2(n_1_1_481), .ZN(n_1_1_157));
   AND2_X1 i_1_1_447 (.A1(adder_out1[13]), .A2(n_1_1_187), .ZN(n_163));
   AND2_X1 i_1_1_448 (.A1(adder_out1[14]), .A2(n_1_1_187), .ZN(n_164));
   AND2_X1 i_1_1_449 (.A1(adder_out1[15]), .A2(n_1_1_187), .ZN(n_165));
   NAND2_X1 i_1_1_450 (.A1(n_1_1_158), .A2(n_1_1_159), .ZN(n_166));
   NOR2_X1 i_1_1_451 (.A1(RST), .A2(n_1_1_160), .ZN(n_1_1_158));
   NOR4_X1 i_1_1_460 (.A1(n_1_1_182), .A2(n_1_1_165), .A3(n_1_1_166), .A4(
      n_1_1_222), .ZN(n_1_132));
   OAI221_X1 i_1_1_461 (.A(n_1_1_530), .B1(n_1_1_475), .B2(Temp[0]), .C1(
      n_1_1_241), .C2(RAM_Data_RD_A[0]), .ZN(n_1_1_165));
   NOR2_X1 i_1_1_462 (.A1(n_1_1_180), .A2(RAM_Data_RD_B[0]), .ZN(n_1_1_166));
   NOR2_X1 i_1_1_463 (.A1(n_1_1_170), .A2(n_1_1_167), .ZN(n_1_133));
   OAI222_X1 i_1_1_464 (.A1(n_1_1_180), .A2(RAM_Data_RD_B[1]), .B1(n_1_1_241), 
      .B2(RAM_Data_RD_A[1]), .C1(Temp[1]), .C2(n_1_1_475), .ZN(n_1_1_167));
   NOR3_X1 i_1_1_465 (.A1(n_1_1_170), .A2(n_1_1_169), .A3(n_1_1_168), .ZN(
      n_1_134));
   OAI21_X1 i_1_1_466 (.A(n_1_1_224), .B1(n_1_1_180), .B2(RAM_Data_RD_B[2]), 
      .ZN(n_1_1_168));
   OAI22_X1 i_1_1_467 (.A1(Temp[2]), .A2(n_1_1_475), .B1(n_1_1_241), .B2(
      RAM_Data_RD_A[2]), .ZN(n_1_1_169));
   OAI21_X1 i_1_1_468 (.A(n_1_1_218), .B1(n_1_1_225), .B2(n_1_1_473), .ZN(
      n_1_1_170));
   NOR2_X1 i_1_1_469 (.A1(n_1_1_181), .A2(n_1_1_171), .ZN(n_1_135));
   OAI222_X1 i_1_1_470 (.A1(n_1_1_180), .A2(RAM_Data_RD_B[3]), .B1(n_1_1_241), 
      .B2(RAM_Data_RD_A[3]), .C1(Temp[3]), .C2(n_1_1_475), .ZN(n_1_1_171));
   NOR2_X1 i_1_1_471 (.A1(n_1_1_181), .A2(n_1_1_172), .ZN(n_1_136));
   OAI222_X1 i_1_1_472 (.A1(n_1_1_180), .A2(RAM_Data_RD_B[4]), .B1(n_1_1_241), 
      .B2(RAM_Data_RD_A[4]), .C1(Temp[4]), .C2(n_1_1_475), .ZN(n_1_1_172));
   NOR2_X1 i_1_1_473 (.A1(n_1_1_181), .A2(n_1_1_173), .ZN(n_1_137));
   OAI222_X1 i_1_1_474 (.A1(n_1_1_180), .A2(RAM_Data_RD_B[5]), .B1(n_1_1_241), 
      .B2(RAM_Data_RD_A[5]), .C1(Temp[5]), .C2(n_1_1_475), .ZN(n_1_1_173));
   NOR2_X1 i_1_1_475 (.A1(n_1_1_181), .A2(n_1_1_174), .ZN(n_1_138));
   OAI222_X1 i_1_1_476 (.A1(n_1_1_180), .A2(RAM_Data_RD_B[6]), .B1(n_1_1_241), 
      .B2(RAM_Data_RD_A[6]), .C1(Temp[6]), .C2(n_1_1_475), .ZN(n_1_1_174));
   NOR2_X1 i_1_1_477 (.A1(n_1_1_181), .A2(n_1_1_175), .ZN(n_1_139));
   OAI222_X1 i_1_1_478 (.A1(n_1_1_180), .A2(RAM_Data_RD_B[7]), .B1(n_1_1_241), 
      .B2(RAM_Data_RD_A[7]), .C1(Temp[7]), .C2(n_1_1_475), .ZN(n_1_1_175));
   NOR2_X1 i_1_1_479 (.A1(n_1_1_181), .A2(n_1_1_176), .ZN(n_1_140));
   OAI222_X1 i_1_1_480 (.A1(n_1_1_180), .A2(RAM_Data_RD_B[8]), .B1(n_1_1_241), 
      .B2(RAM_Data_RD_A[8]), .C1(Temp[8]), .C2(n_1_1_475), .ZN(n_1_1_176));
   AOI211_X1 i_1_1_481 (.A(n_1_1_181), .B(n_1_1_177), .C1(n_1_1_635), .C2(
      n_1_1_658), .ZN(n_1_141));
   OAI22_X1 i_1_1_482 (.A1(n_1_1_180), .A2(RAM_Data_RD_B[9]), .B1(Temp[9]), 
      .B2(n_1_1_475), .ZN(n_1_1_177));
   NOR2_X1 i_1_1_483 (.A1(n_1_1_181), .A2(n_1_1_178), .ZN(n_1_142));
   OAI222_X1 i_1_1_484 (.A1(n_1_1_180), .A2(RAM_Data_RD_B[10]), .B1(n_1_1_241), 
      .B2(RAM_Data_RD_A[10]), .C1(Temp[10]), .C2(n_1_1_475), .ZN(n_1_1_178));
   AOI211_X1 i_1_1_485 (.A(n_1_1_181), .B(n_1_1_179), .C1(n_1_1_637), .C2(
      n_1_1_658), .ZN(n_1_143));
   OAI22_X1 i_1_1_486 (.A1(n_1_1_180), .A2(RAM_Data_RD_B[11]), .B1(Temp[11]), 
      .B2(n_1_1_475), .ZN(n_1_1_179));
   NAND2_X1 i_1_1_487 (.A1(n_1_1_226), .A2(n_1_1_475), .ZN(n_1_1_180));
   OR2_X1 i_1_1_488 (.A1(n_1_1_182), .A2(n_1_1_229), .ZN(n_1_1_181));
   NOR2_X1 i_1_1_489 (.A1(n_1_1_473), .A2(n_1_1_225), .ZN(n_1_1_182));
   NOR2_X1 i_1_1_490 (.A1(n_1_1_183), .A2(n_1_1_267), .ZN(n_1_144));
   AOI222_X1 i_1_1_491 (.A1(Temp[12]), .A2(n_1_1_474), .B1(n_1_1_658), .B2(
      RAM_Data_RD_A[12]), .C1(RAM_Data_RD_B[12]), .C2(n_1_1_591), .ZN(n_1_1_183));
   INV_X1 i_1_1_492 (.A(n_1_1_184), .ZN(n_1_145));
   AOI222_X1 i_1_1_493 (.A1(Temp[13]), .A2(n_1_1_473), .B1(n_1_1_658), .B2(
      n_1_29), .C1(n_1_1_187), .C2(RAM_Data_RD_B[13]), .ZN(n_1_1_184));
   INV_X1 i_1_1_494 (.A(n_1_1_185), .ZN(n_1_146));
   AOI222_X1 i_1_1_495 (.A1(Temp[14]), .A2(n_1_1_473), .B1(n_1_1_658), .B2(
      n_1_30), .C1(n_1_1_187), .C2(RAM_Data_RD_B[14]), .ZN(n_1_1_185));
   INV_X1 i_1_1_496 (.A(n_1_1_186), .ZN(n_1_147));
   AOI222_X1 i_1_1_497 (.A1(Temp[15]), .A2(n_1_1_473), .B1(n_1_1_240), .B2(
      RAM_Data_RD_A[15]), .C1(n_1_1_187), .C2(RAM_Data_RD_B[15]), .ZN(n_1_1_186));
   NOR2_X1 i_1_1_498 (.A1(n_1_1_590), .A2(RST), .ZN(n_1_1_187));
   NAND2_X1 i_1_1_501 (.A1(n_1_1_475), .A2(n_1_1_241), .ZN(n_1_1_189));
   NOR2_X1 i_1_1_502 (.A1(RST), .A2(n_1_1_190), .ZN(n_167));
   NOR2_X1 i_1_1_503 (.A1(n_1_1_273), .A2(n_1_1_191), .ZN(n_1_1_190));
   AOI22_X1 i_1_1_504 (.A1(n_1_1_195), .A2(n_1_1_194), .B1(n_1_1_193), .B2(
      n_1_1_192), .ZN(n_1_1_191));
   OAI22_X1 i_1_1_505 (.A1(RAM_Data_RD_A[0]), .A2(NextState[2]), .B1(n_1_1_593), 
      .B2(n_1_1_474), .ZN(n_1_1_192));
   AOI22_X1 i_1_1_506 (.A1(count[0]), .A2(n_1_1_531), .B1(n_1_1_658), .B2(
      RAM_Data_RD_B[0]), .ZN(n_1_1_193));
   AOI22_X1 i_1_1_507 (.A1(RAM_Data_RD_B[0]), .A2(n_1_1_243), .B1(n_1_1_233), 
      .B2(count[0]), .ZN(n_1_1_194));
   AOI21_X1 i_1_1_508 (.A(n_1_1_253), .B1(n_1_1_244), .B2(adder_out1[0]), 
      .ZN(n_1_1_195));
   NOR2_X1 i_1_1_509 (.A1(n_1_1_197), .A2(n_1_1_196), .ZN(n_168));
   OAI22_X1 i_1_1_510 (.A1(count[1]), .A2(n_1_1_221), .B1(n_1_1_217), .B2(
      RAM_Data_RD_B[1]), .ZN(n_1_1_196));
   OAI221_X1 i_1_1_511 (.A(n_1_1_225), .B1(n_1_1_224), .B2(adder_out1[1]), 
      .C1(n_1_1_227), .C2(RAM_Data_RD_A[1]), .ZN(n_1_1_197));
   NOR2_X1 i_1_1_512 (.A1(n_1_1_199), .A2(n_1_1_198), .ZN(n_169));
   OAI22_X1 i_1_1_513 (.A1(count[2]), .A2(n_1_1_221), .B1(n_1_1_217), .B2(
      RAM_Data_RD_B[2]), .ZN(n_1_1_198));
   OAI221_X1 i_1_1_514 (.A(n_1_1_225), .B1(n_1_1_224), .B2(adder_out1[2]), 
      .C1(n_1_1_227), .C2(RAM_Data_RD_A[2]), .ZN(n_1_1_199));
   NOR2_X1 i_1_1_515 (.A1(n_1_1_201), .A2(n_1_1_200), .ZN(n_170));
   OAI22_X1 i_1_1_516 (.A1(count[3]), .A2(n_1_1_221), .B1(n_1_1_217), .B2(
      RAM_Data_RD_B[3]), .ZN(n_1_1_200));
   OAI221_X1 i_1_1_517 (.A(n_1_1_225), .B1(n_1_1_224), .B2(adder_out1[3]), 
      .C1(n_1_1_227), .C2(RAM_Data_RD_A[3]), .ZN(n_1_1_201));
   NOR2_X1 i_1_1_518 (.A1(n_1_1_203), .A2(n_1_1_202), .ZN(n_171));
   OAI22_X1 i_1_1_519 (.A1(count[4]), .A2(n_1_1_221), .B1(n_1_1_217), .B2(
      RAM_Data_RD_B[4]), .ZN(n_1_1_202));
   OAI221_X1 i_1_1_520 (.A(n_1_1_225), .B1(n_1_1_224), .B2(adder_out1[4]), 
      .C1(n_1_1_227), .C2(RAM_Data_RD_A[4]), .ZN(n_1_1_203));
   NOR2_X1 i_1_1_521 (.A1(n_1_1_205), .A2(n_1_1_204), .ZN(n_172));
   OAI22_X1 i_1_1_522 (.A1(count[5]), .A2(n_1_1_221), .B1(n_1_1_217), .B2(
      RAM_Data_RD_B[5]), .ZN(n_1_1_204));
   OAI221_X1 i_1_1_523 (.A(n_1_1_225), .B1(n_1_1_224), .B2(adder_out1[5]), 
      .C1(n_1_1_227), .C2(RAM_Data_RD_A[5]), .ZN(n_1_1_205));
   NOR2_X1 i_1_1_524 (.A1(n_1_1_207), .A2(n_1_1_206), .ZN(n_173));
   OAI22_X1 i_1_1_525 (.A1(count[6]), .A2(n_1_1_221), .B1(n_1_1_217), .B2(
      RAM_Data_RD_B[6]), .ZN(n_1_1_206));
   OAI221_X1 i_1_1_526 (.A(n_1_1_225), .B1(n_1_1_224), .B2(adder_out1[6]), 
      .C1(n_1_1_227), .C2(RAM_Data_RD_A[6]), .ZN(n_1_1_207));
   NOR2_X1 i_1_1_527 (.A1(n_1_1_209), .A2(n_1_1_208), .ZN(n_174));
   OAI22_X1 i_1_1_528 (.A1(count[7]), .A2(n_1_1_221), .B1(n_1_1_217), .B2(
      RAM_Data_RD_B[7]), .ZN(n_1_1_208));
   OAI221_X1 i_1_1_529 (.A(n_1_1_225), .B1(n_1_1_224), .B2(adder_out1[7]), 
      .C1(n_1_1_227), .C2(RAM_Data_RD_A[7]), .ZN(n_1_1_209));
   NOR2_X1 i_1_1_530 (.A1(n_1_1_211), .A2(n_1_1_210), .ZN(n_175));
   OAI22_X1 i_1_1_531 (.A1(count[8]), .A2(n_1_1_221), .B1(n_1_1_217), .B2(
      RAM_Data_RD_B[8]), .ZN(n_1_1_210));
   OAI221_X1 i_1_1_532 (.A(n_1_1_225), .B1(n_1_1_224), .B2(adder_out1[8]), 
      .C1(n_1_1_227), .C2(RAM_Data_RD_A[8]), .ZN(n_1_1_211));
   NOR2_X1 i_1_1_533 (.A1(n_1_1_213), .A2(n_1_1_212), .ZN(n_176));
   OAI22_X1 i_1_1_534 (.A1(count[9]), .A2(n_1_1_221), .B1(n_1_1_217), .B2(
      RAM_Data_RD_B[9]), .ZN(n_1_1_212));
   OAI221_X1 i_1_1_535 (.A(n_1_1_225), .B1(n_1_1_224), .B2(adder_out1[9]), 
      .C1(n_1_1_227), .C2(RAM_Data_RD_A[9]), .ZN(n_1_1_213));
   NOR2_X1 i_1_1_536 (.A1(n_1_1_215), .A2(n_1_1_214), .ZN(n_177));
   OAI22_X1 i_1_1_537 (.A1(count[10]), .A2(n_1_1_221), .B1(n_1_1_217), .B2(
      RAM_Data_RD_B[10]), .ZN(n_1_1_214));
   OAI221_X1 i_1_1_538 (.A(n_1_1_225), .B1(n_1_1_224), .B2(adder_out1[10]), 
      .C1(n_1_1_227), .C2(RAM_Data_RD_A[10]), .ZN(n_1_1_215));
   NOR2_X1 i_1_1_539 (.A1(n_1_1_223), .A2(n_1_1_216), .ZN(n_178));
   OAI22_X1 i_1_1_540 (.A1(count[11]), .A2(n_1_1_221), .B1(n_1_1_217), .B2(
      RAM_Data_RD_B[11]), .ZN(n_1_1_216));
   NOR2_X1 i_1_1_541 (.A1(n_1_1_658), .A2(n_1_1_219), .ZN(n_1_1_217));
   AND2_X1 i_1_1_543 (.A1(n_1_1_254), .A2(n_1_1_243), .ZN(n_1_1_219));
   AOI22_X1 i_1_1_545 (.A1(n_1_1_254), .A2(n_1_1_233), .B1(n_1_1_595), .B2(
      n_1_1_452), .ZN(n_1_1_221));
   NOR2_X1 i_1_1_546 (.A1(n_1_1_253), .A2(n_1_1_243), .ZN(n_1_1_222));
   OAI221_X1 i_1_1_547 (.A(n_1_1_225), .B1(n_1_1_224), .B2(adder_out1[11]), 
      .C1(n_1_1_227), .C2(RAM_Data_RD_A[11]), .ZN(n_1_1_223));
   NAND2_X1 i_1_1_548 (.A1(n_1_1_254), .A2(n_1_1_244), .ZN(n_1_1_224));
   AOI21_X1 i_1_1_549 (.A(n_1_1_267), .B1(n_1_1_226), .B2(n_1_1_590), .ZN(
      n_1_1_225));
   INV_X1 i_1_1_550 (.A(n_1_1_227), .ZN(n_1_1_226));
   NAND3_X1 i_1_1_551 (.A1(n_1_1_530), .A2(n_1_1_253), .A3(n_1_1_241), .ZN(
      n_1_1_227));
   AOI211_X1 i_1_1_552 (.A(n_1_1_230), .B(n_1_1_228), .C1(n_1_1_232), .C2(
      n_1_1_231), .ZN(n_179));
   AOI221_X1 i_1_1_553 (.A(n_1_1_229), .B1(n_1_1_658), .B2(RAM_Data_RD_B[12]), 
      .C1(RAM_Data_RD_A[12]), .C2(n_1_1_591), .ZN(n_1_1_228));
   NAND2_X1 i_1_1_554 (.A1(n_1_1_530), .A2(n_1_1_253), .ZN(n_1_1_229));
   OAI221_X1 i_1_1_555 (.A(n_1_1_605), .B1(n_1_1_583), .B2(NextState[3]), 
      .C1(n_1_1_530), .C2(count[12]), .ZN(n_1_1_230));
   AOI221_X1 i_1_1_556 (.A(n_1_1_253), .B1(n_1_1_244), .B2(adder_out1[12]), 
      .C1(n_1_1_243), .C2(RAM_Data_RD_B[12]), .ZN(n_1_1_231));
   NAND2_X1 i_1_1_557 (.A1(count[12]), .A2(n_1_1_233), .ZN(n_1_1_232));
   NOR2_X1 i_1_1_558 (.A1(n_1_1_244), .A2(n_1_1_243), .ZN(n_1_1_233));
   AOI22_X1 i_1_1_559 (.A1(n_1_1_246), .A2(n_1_1_235), .B1(n_1_1_234), .B2(
      n_1_1_239), .ZN(n_180));
   AOI22_X1 i_1_1_560 (.A1(RAM_Data_RD_B[13]), .A2(n_1_1_240), .B1(n_1_29), 
      .B2(n_1_1_593), .ZN(n_1_1_234));
   NOR2_X1 i_1_1_561 (.A1(n_1_1_639), .A2(RST), .ZN(n_1_29));
   AOI22_X1 i_1_1_562 (.A1(adder_out1[13]), .A2(n_1_1_244), .B1(n_1_1_243), 
      .B2(RAM_Data_RD_B[13]), .ZN(n_1_1_235));
   AOI22_X1 i_1_1_563 (.A1(n_1_1_246), .A2(n_1_1_237), .B1(n_1_1_236), .B2(
      n_1_1_239), .ZN(n_181));
   AOI22_X1 i_1_1_564 (.A1(RAM_Data_RD_B[14]), .A2(n_1_1_240), .B1(n_1_30), 
      .B2(n_1_1_593), .ZN(n_1_1_236));
   NOR2_X1 i_1_1_565 (.A1(n_1_1_640), .A2(RST), .ZN(n_1_30));
   AOI22_X1 i_1_1_566 (.A1(adder_out1[14]), .A2(n_1_1_244), .B1(n_1_1_243), 
      .B2(RAM_Data_RD_B[14]), .ZN(n_1_1_237));
   AOI22_X1 i_1_1_567 (.A1(n_1_1_246), .A2(n_1_1_242), .B1(n_1_1_239), .B2(
      n_1_1_238), .ZN(n_182));
   AOI22_X1 i_1_1_568 (.A1(RAM_Data_RD_B[15]), .A2(n_1_1_240), .B1(n_1_31), 
      .B2(n_1_1_593), .ZN(n_1_1_238));
   INV_X1 i_1_1_569 (.A(n_1_1_239), .ZN(n_183));
   NAND2_X1 i_1_1_570 (.A1(n_1_1_593), .A2(n_1_13), .ZN(n_1_1_239));
   NOR2_X1 i_1_1_571 (.A1(n_1_1_641), .A2(RST), .ZN(n_1_31));
   NOR2_X1 i_1_1_572 (.A1(n_1_1_241), .A2(RST), .ZN(n_1_1_240));
   AOI22_X1 i_1_1_574 (.A1(adder_out1[15]), .A2(n_1_1_244), .B1(n_1_1_243), 
      .B2(RAM_Data_RD_B[15]), .ZN(n_1_1_242));
   NOR3_X1 i_1_1_575 (.A1(n_1_1_245), .A2(State[2]), .A3(n_1_1_611), .ZN(
      n_1_1_243));
   AND2_X1 i_1_1_576 (.A1(n_313), .A2(n_1_1_252), .ZN(n_1_1_244));
   NAND3_X1 i_1_1_577 (.A1(State[3]), .A2(State[1]), .A3(n_313), .ZN(n_1_1_245));
   INV_X1 i_1_1_578 (.A(n_1_1_247), .ZN(n_1_1_246));
   NAND2_X1 i_1_1_579 (.A1(n_1_1_254), .A2(n_1_1_248), .ZN(n_1_1_247));
   NOR3_X1 i_1_1_581 (.A1(n_1_1_250), .A2(State[2]), .A3(n_1_1_611), .ZN(
      n_1_1_249));
   NAND3_X1 i_1_1_582 (.A1(State[3]), .A2(State[1]), .A3(n_315), .ZN(n_1_1_250));
   AND2_X1 i_1_1_583 (.A1(n_314), .A2(n_1_1_252), .ZN(n_1_1_251));
   AND4_X1 i_1_1_584 (.A1(n_1_1_611), .A2(State[1]), .A3(State[2]), .A4(State[3]), 
      .ZN(n_1_1_252));
   NOR2_X1 i_1_1_586 (.A1(n_1_1_608), .A2(n_1_1_592), .ZN(n_1_1_254));
   NAND3_X1 i_1_1_592 (.A1(n_1_1_582), .A2(n_1_1_545), .A3(n_1_1_259), .ZN(n_184));
   NOR4_X1 i_1_1_593 (.A1(n_1_1_260), .A2(n_1_1_540), .A3(n_1_1_544), .A4(RST), 
      .ZN(n_1_1_259));
   NAND2_X1 i_1_1_594 (.A1(n_1_1_536), .A2(n_1_1_300), .ZN(n_1_1_260));
   AOI21_X1 i_1_1_600 (.A(RST), .B1(n_1_1_277), .B2(n_1_1_265), .ZN(n_185));
   NAND2_X1 i_1_1_601 (.A1(n_1_1_297), .A2(adder_out1[0]), .ZN(n_1_1_265));
   AOI21_X1 i_1_1_602 (.A(n_1_1_267), .B1(n_1_1_277), .B2(n_1_1_266), .ZN(n_186));
   AOI22_X1 i_1_1_603 (.A1(n_1_1_297), .A2(adder_out1[1]), .B1(NextState[0]), 
      .B2(n_1_1_587), .ZN(n_1_1_266));
   NAND2_X1 i_1_1_604 (.A1(n_1_1_605), .A2(n_1_1_272), .ZN(n_1_1_267));
   NOR2_X1 i_1_1_605 (.A1(RST), .A2(n_1_1_273), .ZN(n_1_1_268));
   OAI21_X1 i_1_1_606 (.A(n_1_1_269), .B1(n_1_1_272), .B2(RST), .ZN(n_187));
   NOR2_X1 i_1_1_607 (.A1(n_1_1_607), .A2(RST), .ZN(n_1_12));
   NAND2_X1 i_1_1_608 (.A1(adder_out1[2]), .A2(n_1_1_278), .ZN(n_1_1_269));
   AND2_X1 i_1_1_609 (.A1(adder_out1[3]), .A2(n_1_1_278), .ZN(n_188));
   AND2_X1 i_1_1_610 (.A1(adder_out1[4]), .A2(n_1_1_278), .ZN(n_189));
   AND2_X1 i_1_1_611 (.A1(adder_out1[5]), .A2(n_1_1_278), .ZN(n_190));
   AND2_X1 i_1_1_612 (.A1(adder_out1[6]), .A2(n_1_1_278), .ZN(n_191));
   AND2_X1 i_1_1_613 (.A1(adder_out1[7]), .A2(n_1_1_278), .ZN(n_192));
   AND2_X1 i_1_1_614 (.A1(adder_out1[8]), .A2(n_1_1_278), .ZN(n_193));
   AND2_X1 i_1_1_615 (.A1(adder_out1[9]), .A2(n_1_1_278), .ZN(n_194));
   AND2_X1 i_1_1_616 (.A1(adder_out1[10]), .A2(n_1_1_278), .ZN(n_195));
   AND2_X1 i_1_1_617 (.A1(adder_out1[11]), .A2(n_1_1_278), .ZN(n_196));
   AND2_X1 i_1_1_618 (.A1(adder_out1[12]), .A2(n_1_1_278), .ZN(n_197));
   OR3_X1 i_1_1_619 (.A1(n_1_1_275), .A2(n_1_1_271), .A3(n_1_1_270), .ZN(n_198));
   OAI33_X1 i_1_1_620 (.A1(n_1_1_299), .A2(invalid2), .A3(invalid1), .B1(
      n_1_1_606), .B2(NextState[3]), .B3(NextState[1]), .ZN(n_1_1_270));
   NOR2_X1 i_1_1_623 (.A1(n_1_1_586), .A2(n_1_1_583), .ZN(n_1_1_273));
   INV_X1 i_1_1_624 (.A(n_1_1_274), .ZN(n_199));
   AOI21_X1 i_1_1_625 (.A(n_1_1_275), .B1(n_1_1_297), .B2(adder_out2[0]), 
      .ZN(n_1_1_274));
   NAND2_X1 i_1_1_626 (.A1(n_1_1_605), .A2(n_1_1_277), .ZN(n_1_1_275));
   AND2_X1 i_1_1_627 (.A1(adder_out2[1]), .A2(n_1_1_278), .ZN(n_200));
   AOI21_X1 i_1_1_628 (.A(RST), .B1(n_1_1_277), .B2(n_1_1_276), .ZN(n_201));
   NAND2_X1 i_1_1_629 (.A1(n_1_1_297), .A2(adder_out2[2]), .ZN(n_1_1_276));
   OR2_X1 i_1_1_630 (.A1(n_1_1_299), .A2(n_1_1_280), .ZN(n_1_1_277));
   AND2_X1 i_1_1_631 (.A1(adder_out2[3]), .A2(n_1_1_278), .ZN(n_202));
   AND2_X1 i_1_1_632 (.A1(adder_out2[4]), .A2(n_1_1_278), .ZN(n_203));
   AND2_X1 i_1_1_633 (.A1(adder_out2[5]), .A2(n_1_1_278), .ZN(n_204));
   AND2_X1 i_1_1_634 (.A1(adder_out2[6]), .A2(n_1_1_278), .ZN(n_205));
   AND2_X1 i_1_1_635 (.A1(adder_out2[7]), .A2(n_1_1_278), .ZN(n_206));
   AND2_X1 i_1_1_636 (.A1(adder_out2[8]), .A2(n_1_1_278), .ZN(n_207));
   AND2_X1 i_1_1_637 (.A1(adder_out2[9]), .A2(n_1_1_278), .ZN(n_208));
   AND2_X1 i_1_1_638 (.A1(adder_out2[10]), .A2(n_1_1_278), .ZN(n_209));
   AND2_X1 i_1_1_639 (.A1(adder_out2[11]), .A2(n_1_1_278), .ZN(n_210));
   AND2_X1 i_1_1_640 (.A1(adder_out2[12]), .A2(n_1_1_278), .ZN(n_211));
   AOI21_X1 i_1_1_641 (.A(RST), .B1(n_1_1_298), .B2(n_1_1_279), .ZN(n_1_1_278));
   NAND4_X1 i_1_1_643 (.A1(n_1_1_296), .A2(n_1_1_294), .A3(n_1_1_282), .A4(
      n_1_1_281), .ZN(n_1_1_280));
   NOR4_X1 i_1_1_644 (.A1(n_1_1_295), .A2(n_1_1_291), .A3(n_1_1_290), .A4(
      n_1_1_286), .ZN(n_1_1_281));
   NOR4_X1 i_1_1_645 (.A1(n_1_1_284), .A2(n_1_1_283), .A3(n_1_1_293), .A4(
      n_1_1_289), .ZN(n_1_1_282));
   NAND4_X1 i_1_1_646 (.A1(n_1_1_292), .A2(n_1_1_288), .A3(n_1_1_287), .A4(
      n_1_1_285), .ZN(n_1_1_283));
   XOR2_X1 i_1_1_647 (.A(N[6]), .B(count[6]), .Z(n_1_1_284));
   XNOR2_X1 i_1_1_648 (.A(N[4]), .B(count[4]), .ZN(n_1_1_285));
   XOR2_X1 i_1_1_649 (.A(N[2]), .B(count[2]), .Z(n_1_1_286));
   XNOR2_X1 i_1_1_650 (.A(N[10]), .B(count[10]), .ZN(n_1_1_287));
   XNOR2_X1 i_1_1_651 (.A(N[9]), .B(count[9]), .ZN(n_1_1_288));
   XOR2_X1 i_1_1_652 (.A(N[12]), .B(count[12]), .Z(n_1_1_289));
   XOR2_X1 i_1_1_653 (.A(N[1]), .B(count[1]), .Z(n_1_1_290));
   XOR2_X1 i_1_1_654 (.A(N[8]), .B(count[8]), .Z(n_1_1_291));
   XNOR2_X1 i_1_1_655 (.A(N[0]), .B(count[0]), .ZN(n_1_1_292));
   XOR2_X1 i_1_1_656 (.A(N[5]), .B(count[5]), .Z(n_1_1_293));
   XNOR2_X1 i_1_1_657 (.A(N[11]), .B(count[11]), .ZN(n_1_1_294));
   XOR2_X1 i_1_1_658 (.A(N[7]), .B(count[7]), .Z(n_1_1_295));
   XNOR2_X1 i_1_1_659 (.A(N[3]), .B(count[3]), .ZN(n_1_1_296));
   NAND3_X1 i_1_1_660 (.A1(n_1_1_605), .A2(n_1_1_299), .A3(n_1_1_298), .ZN(n_212));
   NAND2_X1 i_1_1_661 (.A1(n_1_1_299), .A2(n_1_1_298), .ZN(n_1_1_297));
   NAND2_X1 i_1_1_662 (.A1(n_1_1_589), .A2(n_1_1_535), .ZN(n_1_1_298));
   NAND2_X1 i_1_1_663 (.A1(n_1_1_594), .A2(n_1_1_533), .ZN(n_1_1_299));
   NAND2_X1 i_1_1_664 (.A1(n_1_1_608), .A2(n_1_1_607), .ZN(n_1_1_300));
   AOI222_X1 i_1_1_669 (.A1(RAM_Data_RD_A[0]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(RAM_Data_RD_B[0]), .C1(n_1_5), .C2(htemp[0]), .ZN(n_1_1_304));
   AOI222_X1 i_1_1_697 (.A1(RAM_Data_RD_A[7]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(RAM_Data_RD_B[7]), .C1(n_1_5), .C2(htemp[7]), .ZN(n_1_1_325));
   AOI222_X1 i_1_1_705 (.A1(RAM_Data_RD_A[9]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(RAM_Data_RD_B[9]), .C1(n_1_5), .C2(htemp[9]), .ZN(n_1_1_331));
   AOI222_X1 i_1_1_722 (.A1(RAM_Data_RD_A[13]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(RAM_Data_RD_B[13]), .C1(n_1_5), .C2(htemp[13]), .ZN(n_1_1_344));
   AOI21_X1 i_1_1_728 (.A(n_1_1_350), .B1(n_1_1_349), .B2(n_1_1_460), .ZN(n_213));
   AOI222_X1 i_1_1_729 (.A1(RAM_Data_RD_A[15]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(RAM_Data_RD_B[15]), .C1(n_1_5), .C2(htemp[15]), .ZN(n_1_1_349));
   AOI21_X1 i_1_1_730 (.A(n_1_1_351), .B1(n_1_1_455), .B2(RAM_Data_RD_B[15]), 
      .ZN(n_1_1_350));
   OAI21_X1 i_1_1_731 (.A(n_1_1_451), .B1(n_1_1_545), .B2(n_1_1_352), .ZN(
      n_1_1_351));
   NAND2_X1 i_1_1_732 (.A1(adder_out1[12]), .A2(adder_out2[15]), .ZN(n_1_1_352));
   AOI21_X1 i_1_1_733 (.A(n_1_1_354), .B1(n_1_1_353), .B2(n_1_1_460), .ZN(n_214));
   AOI222_X1 i_1_1_734 (.A1(RAM_Data_RD_A[16]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(RAM_Data_RD_B[16]), .C1(n_1_5), .C2(htemp[16]), .ZN(n_1_1_353));
   AOI21_X1 i_1_1_735 (.A(n_1_1_452), .B1(n_1_1_455), .B2(RAM_Data_RD_B[16]), 
      .ZN(n_1_1_354));
   NOR2_X1 i_1_1_877 (.A1(n_1_1_530), .A2(RST), .ZN(n_1_5));
   NOR3_X1 i_1_1_879 (.A1(n_1_1_563), .A2(n_1_1_546), .A3(n_1_1_452), .ZN(
      n_1_1_450));
   AOI211_X1 i_1_1_887 (.A(n_1_1_481), .B(n_1_1_457), .C1(NextState[3]), 
      .C2(n_1_1_532), .ZN(n_215));
   AOI221_X1 i_1_1_888 (.A(NextState[3]), .B1(adder_out2[0]), .B2(n_1_1_596), 
      .C1(n_1_1_584), .C2(adder_out1[0]), .ZN(n_1_1_457));
   INV_X1 i_1_1_889 (.A(n_1_1_458), .ZN(n_216));
   AOI22_X1 i_1_1_890 (.A1(adder_out2[1]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(adder_out1[1]), .ZN(n_1_1_458));
   OAI211_X1 i_1_1_891 (.A(n_1_1_462), .B(n_1_1_460), .C1(n_1_1_459), .C2(
      n_1_1_481), .ZN(n_217));
   AOI21_X1 i_1_1_892 (.A(n_1_1_533), .B1(n_1_1_476), .B2(adder_out1[2]), 
      .ZN(n_1_1_459));
   NOR2_X1 i_1_1_894 (.A1(n_1_1_581), .A2(RST), .ZN(n_1_1_461));
   NAND3_X1 i_1_1_895 (.A1(adder_out2[2]), .A2(n_1_1_535), .A3(n_1_1_479), 
      .ZN(n_1_1_462));
   INV_X1 i_1_1_896 (.A(n_1_1_463), .ZN(n_218));
   AOI22_X1 i_1_1_897 (.A1(adder_out2[3]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(adder_out1[3]), .ZN(n_1_1_463));
   INV_X1 i_1_1_898 (.A(n_1_1_464), .ZN(n_219));
   AOI22_X1 i_1_1_899 (.A1(adder_out2[4]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(adder_out1[4]), .ZN(n_1_1_464));
   INV_X1 i_1_1_900 (.A(n_1_1_465), .ZN(n_220));
   AOI22_X1 i_1_1_901 (.A1(adder_out2[5]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(adder_out1[5]), .ZN(n_1_1_465));
   INV_X1 i_1_1_902 (.A(n_1_1_466), .ZN(n_221));
   AOI22_X1 i_1_1_903 (.A1(adder_out2[6]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(adder_out1[6]), .ZN(n_1_1_466));
   INV_X1 i_1_1_904 (.A(n_1_1_467), .ZN(n_222));
   AOI22_X1 i_1_1_905 (.A1(adder_out2[7]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(adder_out1[7]), .ZN(n_1_1_467));
   INV_X1 i_1_1_906 (.A(n_1_1_468), .ZN(n_223));
   AOI22_X1 i_1_1_907 (.A1(adder_out2[8]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(adder_out1[8]), .ZN(n_1_1_468));
   INV_X1 i_1_1_908 (.A(n_1_1_469), .ZN(n_224));
   AOI22_X1 i_1_1_909 (.A1(adder_out2[9]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(adder_out1[9]), .ZN(n_1_1_469));
   INV_X1 i_1_1_910 (.A(n_1_1_470), .ZN(n_225));
   AOI22_X1 i_1_1_911 (.A1(adder_out2[10]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(adder_out1[10]), .ZN(n_1_1_470));
   INV_X1 i_1_1_912 (.A(n_1_1_471), .ZN(n_226));
   AOI22_X1 i_1_1_913 (.A1(adder_out2[11]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(adder_out1[11]), .ZN(n_1_1_471));
   INV_X1 i_1_1_914 (.A(n_1_1_472), .ZN(n_227));
   AOI22_X1 i_1_1_915 (.A1(adder_out2[12]), .A2(n_1_1_477), .B1(n_1_1_473), 
      .B2(adder_out1[12]), .ZN(n_1_1_472));
   NOR2_X1 i_1_1_916 (.A1(n_1_1_475), .A2(RST), .ZN(n_1_1_473));
   INV_X1 i_1_1_917 (.A(n_1_1_475), .ZN(n_1_1_474));
   NAND2_X1 i_1_1_918 (.A1(n_1_1_584), .A2(n_1_1_535), .ZN(n_1_1_475));
   NOR2_X1 i_1_1_919 (.A1(n_1_1_583), .A2(NextState[3]), .ZN(n_1_1_476));
   NOR2_X1 i_1_1_920 (.A1(n_1_1_595), .A2(n_1_1_480), .ZN(n_1_1_477));
   INV_X1 i_1_1_921 (.A(n_1_1_479), .ZN(n_1_1_478));
   NOR2_X1 i_1_1_922 (.A1(NextState[0]), .A2(RST), .ZN(n_1_1_479));
   NAND2_X1 i_1_1_923 (.A1(n_1_13), .A2(n_1_1_609), .ZN(n_1_1_480));
   INV_X1 i_1_1_924 (.A(n_1_1_481), .ZN(n_1_13));
   NAND2_X1 i_1_1_925 (.A1(n_1_1_605), .A2(NextState[2]), .ZN(n_1_1_481));
   NAND2_X1 i_1_1_928 (.A1(NextState[3]), .A2(NextState[2]), .ZN(n_1_1_483));
   NAND3_X1 i_1_1_931 (.A1(division_operation), .A2(n_1_1_531), .A3(n_1_1_487), 
      .ZN(n_1_1_485));
   AND3_X1 i_1_1_933 (.A1(n_1_1_508), .A2(n_1_1_501), .A3(n_1_1_488), .ZN(
      n_1_1_487));
   NOR4_X1 i_1_1_934 (.A1(n_1_1_496), .A2(n_1_1_493), .A3(n_1_1_489), .A4(
      n_1_1_529), .ZN(n_1_1_488));
   NAND4_X1 i_1_1_935 (.A1(n_1_1_492), .A2(n_1_1_491), .A3(n_1_1_490), .A4(
      n_1_1_524), .ZN(n_1_1_489));
   NOR4_X1 i_1_1_936 (.A1(N[54]), .A2(N[53]), .A3(N[51]), .A4(N[48]), .ZN(
      n_1_1_490));
   NOR4_X1 i_1_1_937 (.A1(N[63]), .A2(N[60]), .A3(N[58]), .A4(N[57]), .ZN(
      n_1_1_491));
   XNOR2_X1 i_1_1_938 (.A(N[10]), .B(Temp[10]), .ZN(n_1_1_492));
   NAND4_X1 i_1_1_939 (.A1(n_1_1_528), .A2(n_1_1_527), .A3(n_1_1_495), .A4(
      n_1_1_494), .ZN(n_1_1_493));
   XNOR2_X1 i_1_1_940 (.A(N[7]), .B(Temp[7]), .ZN(n_1_1_494));
   XNOR2_X1 i_1_1_941 (.A(N[13]), .B(Temp[13]), .ZN(n_1_1_495));
   NAND4_X1 i_1_1_942 (.A1(n_1_1_500), .A2(n_1_1_499), .A3(n_1_1_498), .A4(
      n_1_1_497), .ZN(n_1_1_496));
   NOR4_X1 i_1_1_943 (.A1(N[38]), .A2(N[37]), .A3(N[35]), .A4(N[32]), .ZN(
      n_1_1_497));
   NOR4_X1 i_1_1_944 (.A1(N[47]), .A2(N[44]), .A3(N[42]), .A4(N[41]), .ZN(
      n_1_1_498));
   NOR4_X1 i_1_1_945 (.A1(N[23]), .A2(N[20]), .A3(N[18]), .A4(N[17]), .ZN(
      n_1_1_499));
   NOR4_X1 i_1_1_946 (.A1(N[30]), .A2(N[29]), .A3(N[27]), .A4(N[24]), .ZN(
      n_1_1_500));
   NOR2_X1 i_1_1_947 (.A1(n_1_1_506), .A2(n_1_1_502), .ZN(n_1_1_501));
   NAND4_X1 i_1_1_948 (.A1(n_1_1_505), .A2(n_1_1_504), .A3(n_1_1_503), .A4(
      n_1_1_525), .ZN(n_1_1_502));
   XNOR2_X1 i_1_1_949 (.A(N[3]), .B(Temp[3]), .ZN(n_1_1_503));
   NOR4_X1 i_1_1_950 (.A1(N[55]), .A2(N[52]), .A3(N[50]), .A4(N[49]), .ZN(
      n_1_1_504));
   NOR4_X1 i_1_1_951 (.A1(N[62]), .A2(N[61]), .A3(N[59]), .A4(N[56]), .ZN(
      n_1_1_505));
   NAND4_X1 i_1_1_952 (.A1(n_1_1_526), .A2(n_1_1_523), .A3(n_1_1_522), .A4(
      n_1_1_507), .ZN(n_1_1_506));
   XNOR2_X1 i_1_1_953 (.A(N[14]), .B(Temp[14]), .ZN(n_1_1_507));
   NOR3_X1 i_1_1_954 (.A1(n_1_1_518), .A2(n_1_1_513), .A3(n_1_1_509), .ZN(
      n_1_1_508));
   NAND3_X1 i_1_1_955 (.A1(n_1_1_512), .A2(n_1_1_511), .A3(n_1_1_510), .ZN(
      n_1_1_509));
   NOR2_X1 i_1_1_956 (.A1(N[39]), .A2(N[36]), .ZN(n_1_1_510));
   NOR2_X1 i_1_1_957 (.A1(N[34]), .A2(N[33]), .ZN(n_1_1_511));
   NOR4_X1 i_1_1_958 (.A1(N[46]), .A2(N[45]), .A3(N[43]), .A4(N[40]), .ZN(
      n_1_1_512));
   NAND4_X1 i_1_1_959 (.A1(n_1_1_517), .A2(n_1_1_516), .A3(n_1_1_515), .A4(
      n_1_1_514), .ZN(n_1_1_513));
   NOR2_X1 i_1_1_960 (.A1(N[19]), .A2(N[16]), .ZN(n_1_1_514));
   NOR2_X1 i_1_1_961 (.A1(N[22]), .A2(N[21]), .ZN(n_1_1_515));
   NOR2_X1 i_1_1_962 (.A1(N[31]), .A2(N[28]), .ZN(n_1_1_516));
   NOR2_X1 i_1_1_963 (.A1(N[26]), .A2(N[25]), .ZN(n_1_1_517));
   NAND3_X1 i_1_1_964 (.A1(n_1_1_521), .A2(n_1_1_520), .A3(n_1_1_519), .ZN(
      n_1_1_518));
   XNOR2_X1 i_1_1_965 (.A(N[8]), .B(Temp[8]), .ZN(n_1_1_519));
   XNOR2_X1 i_1_1_966 (.A(N[6]), .B(Temp[6]), .ZN(n_1_1_520));
   XNOR2_X1 i_1_1_967 (.A(N[4]), .B(Temp[4]), .ZN(n_1_1_521));
   XNOR2_X1 i_1_1_968 (.A(N[1]), .B(Temp[1]), .ZN(n_1_1_522));
   XNOR2_X1 i_1_1_969 (.A(N[0]), .B(Temp[0]), .ZN(n_1_1_523));
   XNOR2_X1 i_1_1_970 (.A(N[5]), .B(Temp[5]), .ZN(n_1_1_524));
   XNOR2_X1 i_1_1_971 (.A(N[12]), .B(Temp[12]), .ZN(n_1_1_525));
   XNOR2_X1 i_1_1_972 (.A(N[11]), .B(Temp[11]), .ZN(n_1_1_526));
   XNOR2_X1 i_1_1_973 (.A(N[2]), .B(Temp[2]), .ZN(n_1_1_527));
   XNOR2_X1 i_1_1_974 (.A(N[9]), .B(Temp[9]), .ZN(n_1_1_528));
   XOR2_X1 i_1_1_975 (.A(N[15]), .B(Temp[15]), .Z(n_1_1_529));
   NAND2_X1 i_1_1_976 (.A1(n_1_1_535), .A2(n_1_1_533), .ZN(n_1_1_530));
   NOR2_X1 i_1_1_977 (.A1(n_1_1_534), .A2(n_1_1_532), .ZN(n_1_1_531));
   NAND2_X1 i_1_1_978 (.A1(n_1_1_607), .A2(n_1_1_606), .ZN(n_1_1_532));
   NOR2_X1 i_1_1_979 (.A1(NextState[1]), .A2(NextState[0]), .ZN(n_1_1_533));
   NAND2_X1 i_1_1_980 (.A1(n_1_1_609), .A2(NextState[2]), .ZN(n_1_1_534));
   NAND2_X1 i_1_1_982 (.A1(NextState[2]), .A2(NextState[1]), .ZN(n_1_1_536));
   NOR2_X1 i_1_1_983 (.A1(n_1_1_609), .A2(RST), .ZN(n_1_14));
   NOR3_X1 i_1_1_994 (.A1(n_1_1_555), .A2(n_1_1_553), .A3(n_1_1_548), .ZN(
      n_1_1_547));
   NAND4_X1 i_1_1_995 (.A1(n_1_1_552), .A2(n_1_1_551), .A3(n_1_1_550), .A4(
      n_1_1_549), .ZN(n_1_1_548));
   NOR4_X1 i_1_1_996 (.A1(RAM_Data_RD_A[51]), .A2(RAM_Data_RD_A[50]), .A3(
      RAM_Data_RD_A[49]), .A4(RAM_Data_RD_A[48]), .ZN(n_1_1_549));
   NOR4_X1 i_1_1_997 (.A1(RAM_Data_RD_A[55]), .A2(RAM_Data_RD_A[54]), .A3(
      RAM_Data_RD_A[53]), .A4(RAM_Data_RD_A[52]), .ZN(n_1_1_550));
   NOR4_X1 i_1_1_998 (.A1(RAM_Data_RD_A[63]), .A2(RAM_Data_RD_A[62]), .A3(
      RAM_Data_RD_A[61]), .A4(RAM_Data_RD_A[60]), .ZN(n_1_1_551));
   NOR4_X1 i_1_1_999 (.A1(RAM_Data_RD_A[59]), .A2(RAM_Data_RD_A[58]), .A3(
      RAM_Data_RD_A[57]), .A4(RAM_Data_RD_A[56]), .ZN(n_1_1_552));
   NAND3_X1 i_1_1_1000 (.A1(n_1_1_557), .A2(n_1_1_556), .A3(n_1_1_554), .ZN(
      n_1_1_553));
   NOR4_X1 i_1_1_1001 (.A1(RAM_Data_RD_A[35]), .A2(RAM_Data_RD_A[34]), .A3(
      RAM_Data_RD_A[33]), .A4(RAM_Data_RD_A[32]), .ZN(n_1_1_554));
   NAND4_X1 i_1_1_1002 (.A1(n_1_1_657), .A2(n_1_1_656), .A3(n_1_1_655), .A4(
      n_1_1_654), .ZN(n_1_1_555));
   NOR4_X1 i_1_1_1003 (.A1(RAM_Data_RD_A[47]), .A2(RAM_Data_RD_A[46]), .A3(
      RAM_Data_RD_A[45]), .A4(RAM_Data_RD_A[44]), .ZN(n_1_1_556));
   NOR4_X1 i_1_1_1004 (.A1(RAM_Data_RD_A[43]), .A2(RAM_Data_RD_A[42]), .A3(
      RAM_Data_RD_A[41]), .A4(RAM_Data_RD_A[40]), .ZN(n_1_1_557));
   NOR3_X1 i_1_1_1005 (.A1(n_1_1_562), .A2(n_1_1_561), .A3(n_1_1_559), .ZN(
      n_1_1_558));
   NAND4_X1 i_1_1_1006 (.A1(n_1_1_653), .A2(n_1_1_652), .A3(n_1_1_651), .A4(
      n_1_1_650), .ZN(n_1_1_559));
   NOR4_X1 i_1_1_1007 (.A1(RAM_Data_RD_A[31]), .A2(RAM_Data_RD_A[30]), .A3(
      RAM_Data_RD_A[29]), .A4(RAM_Data_RD_A[28]), .ZN(n_1_1_560));
   NAND4_X1 i_1_1_1008 (.A1(n_1_1_649), .A2(n_1_1_648), .A3(n_1_1_647), .A4(
      n_1_1_646), .ZN(n_1_1_561));
   NAND4_X1 i_1_1_1009 (.A1(n_1_1_645), .A2(n_1_1_644), .A3(n_1_1_643), .A4(
      n_1_1_642), .ZN(n_1_1_562));
   NOR2_X1 i_1_1_1031 (.A1(n_1_1_607), .A2(n_1_1_606), .ZN(n_1_1_584));
   NOR2_X1 i_1_1_1032 (.A1(Euler_End), .A2(RST), .ZN(n_228));
   OAI21_X1 i_1_1_1033 (.A(n_1_1_605), .B1(n_1_1_588), .B2(n_1_1_586), .ZN(n_229));
   NOR2_X1 i_1_1_1034 (.A1(n_1_1_588), .A2(n_1_1_586), .ZN(n_1_1_585));
   NAND2_X1 i_1_1_1035 (.A1(n_1_1_609), .A2(n_1_1_608), .ZN(n_1_1_586));
   NOR2_X1 i_1_1_1036 (.A1(NextState[3]), .A2(NextState[2]), .ZN(n_1_1_587));
   NAND2_X1 i_1_1_1037 (.A1(n_1_1_607), .A2(NextState[0]), .ZN(n_1_1_588));
   NOR2_X1 i_1_1_1038 (.A1(n_1_1_606), .A2(NextState[1]), .ZN(n_1_1_589));
   NOR2_X1 i_1_1_1039 (.A1(RST), .A2(n_1_1_597), .ZN(n_230));
   OAI21_X1 i_1_1_1040 (.A(n_1_1_605), .B1(n_1_1_597), .B2(n_1_1_590), .ZN(n_231));
   NAND2_X1 i_1_1_1041 (.A1(n_1_1_596), .A2(n_1_1_594), .ZN(n_1_1_590));
   NAND2_X1 i_1_1_1043 (.A1(NextState[3]), .A2(n_1_1_596), .ZN(n_1_1_592));
   NAND2_X1 i_1_1_1046 (.A1(n_1_1_606), .A2(NextState[1]), .ZN(n_1_1_595));
   NOR2_X1 i_1_1_1047 (.A1(n_1_1_607), .A2(NextState[0]), .ZN(n_1_1_596));
   INV_X1 i_1_1_1050 (.A(hstate[1]), .ZN(n_1_1_599));
   INV_X1 i_1_1_1051 (.A(Q[7]), .ZN(n_1_1_600));
   INV_X1 i_1_1_1052 (.A(Q[9]), .ZN(n_1_1_601));
   INV_X1 i_1_1_1054 (.A(n_312), .ZN(n_1_1_603));
   INV_X1 i_1_1_1057 (.A(NextState[0]), .ZN(n_1_1_606));
   INV_X1 i_1_1_1058 (.A(NextState[1]), .ZN(n_1_1_607));
   INV_X1 i_1_1_1059 (.A(NextState[2]), .ZN(n_1_1_608));
   INV_X1 i_1_1_1060 (.A(NextState[3]), .ZN(n_1_1_609));
   INV_X1 i_1_1_1062 (.A(State[0]), .ZN(n_1_1_611));
   INV_X1 i_1_1_1063 (.A(Errortemp[2]), .ZN(n_1_1_612));
   INV_X1 i_1_1_1093 (.A(RAM_Data_RD_A[16]), .ZN(n_1_1_642));
   INV_X1 i_1_1_1094 (.A(RAM_Data_RD_A[17]), .ZN(n_1_1_643));
   INV_X1 i_1_1_1095 (.A(RAM_Data_RD_A[18]), .ZN(n_1_1_644));
   INV_X1 i_1_1_1096 (.A(RAM_Data_RD_A[19]), .ZN(n_1_1_645));
   INV_X1 i_1_1_1097 (.A(RAM_Data_RD_A[20]), .ZN(n_1_1_646));
   INV_X1 i_1_1_1098 (.A(RAM_Data_RD_A[21]), .ZN(n_1_1_647));
   INV_X1 i_1_1_1099 (.A(RAM_Data_RD_A[22]), .ZN(n_1_1_648));
   INV_X1 i_1_1_1100 (.A(RAM_Data_RD_A[23]), .ZN(n_1_1_649));
   INV_X1 i_1_1_1101 (.A(RAM_Data_RD_A[24]), .ZN(n_1_1_650));
   INV_X1 i_1_1_1102 (.A(RAM_Data_RD_A[25]), .ZN(n_1_1_651));
   INV_X1 i_1_1_1103 (.A(RAM_Data_RD_A[26]), .ZN(n_1_1_652));
   INV_X1 i_1_1_1104 (.A(RAM_Data_RD_A[27]), .ZN(n_1_1_653));
   INV_X1 i_1_1_1105 (.A(RAM_Data_RD_A[36]), .ZN(n_1_1_654));
   INV_X1 i_1_1_1106 (.A(RAM_Data_RD_A[37]), .ZN(n_1_1_655));
   INV_X1 i_1_1_1107 (.A(RAM_Data_RD_A[38]), .ZN(n_1_1_656));
   INV_X1 i_1_1_1108 (.A(RAM_Data_RD_A[39]), .ZN(n_1_1_657));
   INV_X1 i_1_1_1109 (.A(n_1_1_241), .ZN(n_1_1_658));
   INV_X1 i_1_1_22 (.A(n_1_1_19), .ZN(n_1_1_597));
   NAND3_X1 i_1_1_23 (.A1(n_1_1_673), .A2(n_1_1_674), .A3(n_1_1_670), .ZN(
      n_1_1_19));
   NAND2_X1 i_1_1_27 (.A1(n_1_1_273), .A2(hstate[1]), .ZN(n_1_1_159));
   NAND2_X1 i_1_1_34 (.A1(n_1_1_27), .A2(n_1_1_24), .ZN(n_1_1_23));
   OAI21_X1 i_1_1_130 (.A(n_1_1_97), .B1(n_1_1_55), .B2(n_1_1_20), .ZN(n_232));
   OAI211_X1 i_1_1_131 (.A(n_1_1_27), .B(n_1_1_24), .C1(n_1_1_541), .C2(n_1_1_95), 
      .ZN(n_1_1_20));
   NAND2_X1 i_1_1_132 (.A1(n_1_1_96), .A2(ready), .ZN(n_1_1_95));
   AOI21_X1 i_1_1_316 (.A(n_1_1_56), .B1(n_1_1_668), .B2(n_1_1_675), .ZN(
      n_1_1_55));
   AOI21_X1 i_1_1_317 (.A(n_1_1_22), .B1(n_1_1_21), .B2(n_1_1_593), .ZN(n_1_1_56));
   OR2_X1 i_1_1_318 (.A1(n_1_1_29), .A2(n_1_1_272), .ZN(n_1_1_97));
   NAND2_X1 i_1_1_321 (.A1(n_1_1_584), .A2(n_1_1_587), .ZN(n_1_1_272));
   NAND4_X1 i_1_1_452 (.A1(n_1_1_667), .A2(n_1_1_664), .A3(n_1_1_256), .A4(
      n_1_1_164), .ZN(n_233));
   AOI221_X1 i_1_1_456 (.A(n_1_1_188), .B1(hstate[1]), .B2(n_1_1_273), .C1(
      n_1_1_243), .C2(n_1_1_220), .ZN(n_1_1_164));
   NOR3_X1 i_1_1_458 (.A1(n_1_1_584), .A2(n_1_1_533), .A3(n_1_1_534), .ZN(
      n_1_1_188));
   INV_X1 i_1_1_459 (.A(n_1_1_255), .ZN(n_1_1_220));
   NAND2_X1 i_1_1_499 (.A1(n_1_1_596), .A2(NextState[2]), .ZN(n_1_1_255));
   INV_X1 i_1_1_500 (.A(n_1_1_162), .ZN(n_1_1_256));
   NAND4_X1 i_1_1_573 (.A1(n_1_1_667), .A2(n_1_1_605), .A3(n_1_1_257), .A4(
      n_1_1_94), .ZN(n_234));
   NAND3_X1 i_1_1_587 (.A1(n_1_1_96), .A2(ready), .A3(n_1_1_541), .ZN(n_1_1_94));
   NAND3_X1 i_1_1_589 (.A1(n_1_1_667), .A2(n_1_1_605), .A3(n_1_1_257), .ZN(n_235));
   OR2_X1 i_1_1_590 (.A1(n_1_1_264), .A2(n_1_1_258), .ZN(n_1_1_257));
   NAND4_X1 i_1_1_591 (.A1(n_1_1_101), .A2(n_1_1_100), .A3(n_1_1_99), .A4(
      n_1_1_98), .ZN(n_1_1_258));
   NAND2_X1 i_1_1_988 (.A1(n_1_1_594), .A2(n_1_1_589), .ZN(n_1_1_241));
   OAI211_X1 i_1_1_1048 (.A(n_1_1_664), .B(n_1_1_660), .C1(n_1_1_669), .C2(
      n_1_1_675), .ZN(n_236));
   NOR3_X1 i_1_1_1049 (.A1(n_1_1_246), .A2(n_1_1_189), .A3(n_1_1_271), .ZN(
      n_1_1_660));
   INV_X1 i_1_1_1053 (.A(n_1_1_661), .ZN(n_1_1_271));
   NAND3_X1 i_1_1_1056 (.A1(n_1_1_667), .A2(n_1_1_664), .A3(n_1_1_661), .ZN(
      n_237));
   NAND4_X1 i_1_1_1061 (.A1(n_1_1_584), .A2(n_1_1_663), .A3(n_1_1_662), .A4(
      n_1_1_587), .ZN(n_1_1_661));
   INV_X1 i_1_1_1110 (.A(hstate[0]), .ZN(n_1_1_662));
   INV_X1 i_1_1_1111 (.A(hstate[1]), .ZN(n_1_1_663));
   AOI21_X1 i_1_1_1112 (.A(RST), .B1(n_1_1_665), .B2(n_1_1_666), .ZN(n_1_1_664));
   INV_X1 i_1_1_1113 (.A(n_1_1_487), .ZN(n_1_1_665));
   INV_X1 i_1_1_1114 (.A(n_1_1_530), .ZN(n_1_1_666));
   INV_X1 i_1_1_1116 (.A(n_1_1_669), .ZN(n_1_1_668));
   NAND4_X1 i_1_1_1117 (.A1(n_1_1_673), .A2(n_1_1_674), .A3(n_1_1_591), .A4(
      n_1_1_670), .ZN(n_1_1_669));
   INV_X1 i_1_1_1118 (.A(n_1_1_598), .ZN(n_1_1_670));
   NAND3_X1 i_1_1_1119 (.A1(n_1_1_672), .A2(n_1_1_671), .A3(n_1_1_610), .ZN(
      n_1_1_598));
   INV_X1 i_1_1_1120 (.A(divideByZero), .ZN(n_1_1_671));
   INV_X1 i_1_1_1121 (.A(div_overflow), .ZN(n_1_1_672));
   NOR2_X1 i_1_1_1123 (.A1(n_1_1_592), .A2(NextState[2]), .ZN(n_1_1_591));
   INV_X1 i_1_1_1124 (.A(invalid2), .ZN(n_1_1_673));
   INV_X1 i_1_1_1125 (.A(invalid1), .ZN(n_1_1_674));
   INV_X1 i_1_1_1126 (.A(adder_out1[12]), .ZN(n_1_1_675));
   INV_X1 i_1_1_16 (.A(Errortemp[11]), .ZN(n_1_1_621));
   INV_X1 i_1_1_17 (.A(Errortemp[10]), .ZN(n_1_1_620));
   INV_X1 i_1_1_18 (.A(Errortemp[7]), .ZN(n_1_1_617));
   INV_X1 i_1_1_19 (.A(Errortemp[6]), .ZN(n_1_1_616));
   INV_X1 i_1_1_20 (.A(Errortemp[3]), .ZN(n_1_1_613));
   INV_X1 i_1_1_21 (.A(RAM_Data_RD_A[5]), .ZN(n_1_1_631));
   NAND2_X1 i_1_1_24 (.A1(n_1_1_487), .A2(n_1_1_531), .ZN(n_1_1_486));
   INV_X1 i_1_1_31 (.A(RAM_Data_RD_A[9]), .ZN(n_1_1_635));
   INV_X1 i_1_1_81 (.A(Errortemp[14]), .ZN(n_1_1_624));
   INV_X1 i_1_1_145 (.A(Errortemp[13]), .ZN(n_1_1_623));
   INV_X1 i_1_1_319 (.A(n_1_1_18), .ZN(n_1_1_160));
   INV_X1 i_1_1_320 (.A(mult_overflow), .ZN(n_1_1_610));
   OAI22_X1 i_1_1_352 (.A1(n_1_1_15), .A2(n_1_1_26), .B1(n_1_1_29), .B2(n_1_1_14), 
      .ZN(n_238));
   OAI21_X1 i_1_1_386 (.A(n_1_1_28), .B1(hstate[1]), .B2(n_1_1_583), .ZN(
      n_1_1_14));
   OR2_X1 i_1_1_387 (.A1(n_1_1_30), .A2(RST), .ZN(n_1_1_29));
   OAI211_X1 i_1_1_388 (.A(n_1_1_27), .B(n_1_1_264), .C1(n_1_1_94), .C2(
      n_1_1_598), .ZN(n_1_1_26));
   AOI221_X1 i_1_1_389 (.A(n_1_1_96), .B1(n_1_1_583), .B2(n_1_1_535), .C1(
      n_1_1_131), .C2(n_1_1_16), .ZN(n_1_1_15));
   INV_X1 i_1_1_390 (.A(n_1_1_17), .ZN(n_1_1_16));
   OAI21_X1 i_1_1_391 (.A(n_1_1_279), .B1(n_1_1_18), .B2(mult_overflow), 
      .ZN(n_1_1_17));
   NAND3_X1 i_1_1_453 (.A1(n_1_1_128), .A2(n_1_1_130), .A3(n_1_1_129), .ZN(
      n_1_1_18));
   INV_X1 i_1_1_454 (.A(n_1_1_247), .ZN(n_1_1_128));
   INV_X1 i_1_1_455 (.A(n_1_1_243), .ZN(n_1_1_129));
   INV_X1 i_1_1_457 (.A(n_1_1_244), .ZN(n_1_1_130));
   OAI21_X1 i_1_1_542 (.A(n_1_1_161), .B1(n_1_1_595), .B2(n_1_1_609), .ZN(
      n_1_1_131));
   OAI21_X1 i_1_1_544 (.A(n_1_1_594), .B1(n_1_1_163), .B2(n_1_1_263), .ZN(
      n_1_1_161));
   AOI21_X1 i_1_1_580 (.A(n_1_1_262), .B1(n_1_1_846), .B2(n_1_1_843), .ZN(
      n_1_1_163));
   NOR2_X1 i_1_1_585 (.A1(n_1_1_603), .A2(n_1_1_604), .ZN(n_1_1_262));
   INV_X1 i_1_1_588 (.A(division_operation), .ZN(n_1_1_604));
   INV_X1 i_1_1_595 (.A(NextState[1]), .ZN(n_1_1_263));
   NAND3_X1 i_1_1_596 (.A1(n_1_1_840), .A2(n_1_1_605), .A3(n_1_1_218), .ZN(n_239));
   INV_X1 i_1_1_597 (.A(n_1_1_219), .ZN(n_1_1_218));
   OR2_X1 i_1_1_598 (.A1(n_242), .A2(n_1_1_96), .ZN(n_240));
   INV_X1 i_1_1_599 (.A(n_1_1_301), .ZN(n_1_1_96));
   OR2_X1 i_1_1_621 (.A1(n_1_1_583), .A2(n_1_1_483), .ZN(n_1_1_301));
   OAI221_X1 i_1_1_622 (.A(n_1_1_605), .B1(n_1_1_248), .B2(n_1_1_253), .C1(
      n_1_1_261), .C2(n_1_1_843), .ZN(n_1_115));
   NAND2_X1 i_1_1_642 (.A1(n_1_1_593), .A2(NextState[2]), .ZN(n_1_1_253));
   NOR2_X1 i_1_1_665 (.A1(n_1_1_595), .A2(n_1_1_609), .ZN(n_1_1_593));
   NOR2_X1 i_1_1_666 (.A1(n_1_1_249), .A2(n_1_1_251), .ZN(n_1_1_248));
   OAI21_X1 i_1_1_667 (.A(n_1_1_605), .B1(n_1_1_261), .B2(n_1_1_843), .ZN(n_241));
   OAI21_X1 i_1_1_668 (.A(n_1_1_605), .B1(n_1_1_302), .B2(division_operation), 
      .ZN(n_242));
   AOI22_X1 i_1_1_670 (.A1(n_1_1_303), .A2(n_1_1_540), .B1(n_1_1_531), .B2(
      n_1_1_487), .ZN(n_1_1_302));
   INV_X1 i_1_1_671 (.A(n_1_1_261), .ZN(n_1_1_303));
   OR2_X1 i_1_1_672 (.A1(n_1_1_305), .A2(RST), .ZN(n_243));
   AOI21_X1 i_1_1_673 (.A(n_1_1_162), .B1(n_1_1_261), .B2(n_1_1_306), .ZN(
      n_1_1_305));
   NAND3_X1 i_1_1_674 (.A1(n_1_1_260), .A2(NextState[3]), .A3(n_1_1_606), 
      .ZN(n_1_1_306));
   NAND2_X1 i_1_1_675 (.A1(n_1_1_545), .A2(n_1_1_582), .ZN(n_1_1_261));
   OAI21_X1 i_1_1_676 (.A(n_1_1_279), .B1(n_1_1_247), .B2(n_1_1_244), .ZN(
      n_1_1_162));
   NAND3_X1 i_1_1_677 (.A1(n_1_1_280), .A2(n_1_1_533), .A3(n_1_1_594), .ZN(
      n_1_1_279));
   NAND4_X1 i_1_1_678 (.A1(n_1_1_667), .A2(n_1_1_605), .A3(n_1_1_840), .A4(
      n_1_1_307), .ZN(n_244));
   AND2_X1 i_1_1_679 (.A1(n_1_1_308), .A2(n_1_1_241), .ZN(n_1_1_307));
   OR2_X1 i_1_1_680 (.A1(n_1_1_224), .A2(n_314), .ZN(n_1_1_308));
   NAND2_X1 i_1_1_681 (.A1(n_1_1_668), .A2(n_1_1_675), .ZN(n_1_1_667));
   NAND3_X1 i_1_1_682 (.A1(n_1_1_837), .A2(n_1_1_264), .A3(n_1_1_309), .ZN(n_245));
   INV_X1 i_1_1_683 (.A(n_1_1_310), .ZN(n_1_1_309));
   OAI211_X1 i_1_1_684 (.A(n_1_1_312), .B(n_1_1_605), .C1(n_1_1_536), .C2(
      n_1_1_311), .ZN(n_1_1_310));
   OR2_X1 i_1_1_685 (.A1(NextState[3]), .A2(NextState[0]), .ZN(n_1_1_311));
   OR3_X1 i_1_1_686 (.A1(n_1_1_594), .A2(n_1_1_535), .A3(n_1_1_588), .ZN(
      n_1_1_312));
   NAND2_X1 i_1_1_687 (.A1(n_1_1_665), .A2(n_1_1_666), .ZN(n_1_1_264));
   INV_X1 i_1_1_688 (.A(n_1_1_313), .ZN(n_246));
   OAI221_X1 i_1_1_689 (.A(n_1_1_314), .B1(Q[0]), .B2(n_1_1_830), .C1(
      RAM_Data_RD_B[0]), .C2(n_1_1_394), .ZN(n_1_1_313));
   INV_X1 i_1_1_690 (.A(n_1_1_315), .ZN(n_1_1_314));
   OAI21_X1 i_1_1_691 (.A(n_1_1_316), .B1(n_1_1_393), .B2(adder_out2[0]), 
      .ZN(n_1_1_315));
   NAND2_X1 i_1_1_692 (.A1(n_1_1_304), .A2(n_1_1_460), .ZN(n_1_1_316));
   INV_X1 i_1_1_693 (.A(n_1_1_317), .ZN(n_247));
   OAI221_X1 i_1_1_694 (.A(n_1_1_318), .B1(adder_out2[1]), .B2(n_1_1_393), 
      .C1(RAM_Data_RD_B[1]), .C2(n_1_1_394), .ZN(n_1_1_317));
   AOI22_X1 i_1_1_695 (.A1(n_1_1_382), .A2(n_1_1_321), .B1(n_1_1_320), .B2(
      n_1_1_319), .ZN(n_1_1_318));
   AOI221_X1 i_1_1_696 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[1]), .C1(
      RAM_Data_RD_B[1]), .C2(n_1_1_473), .ZN(n_1_1_319));
   NAND2_X1 i_1_1_698 (.A1(RAM_Data_RD_A[1]), .A2(n_1_1_477), .ZN(n_1_1_320));
   INV_X1 i_1_1_699 (.A(Q[1]), .ZN(n_1_1_321));
   INV_X1 i_1_1_700 (.A(n_1_1_322), .ZN(n_248));
   OAI221_X1 i_1_1_701 (.A(n_1_1_323), .B1(adder_out2[2]), .B2(n_1_1_393), 
      .C1(RAM_Data_RD_B[2]), .C2(n_1_1_394), .ZN(n_1_1_322));
   AOI22_X1 i_1_1_702 (.A1(n_1_1_382), .A2(n_1_1_327), .B1(n_1_1_326), .B2(
      n_1_1_324), .ZN(n_1_1_323));
   AOI221_X1 i_1_1_703 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[2]), .C1(
      RAM_Data_RD_B[2]), .C2(n_1_1_473), .ZN(n_1_1_324));
   NAND2_X1 i_1_1_704 (.A1(RAM_Data_RD_A[2]), .A2(n_1_1_477), .ZN(n_1_1_326));
   INV_X1 i_1_1_706 (.A(Q[2]), .ZN(n_1_1_327));
   INV_X1 i_1_1_707 (.A(n_1_1_328), .ZN(n_249));
   OAI221_X1 i_1_1_708 (.A(n_1_1_329), .B1(adder_out2[3]), .B2(n_1_1_393), 
      .C1(RAM_Data_RD_B[3]), .C2(n_1_1_394), .ZN(n_1_1_328));
   AOI22_X1 i_1_1_709 (.A1(n_1_1_382), .A2(n_1_1_333), .B1(n_1_1_332), .B2(
      n_1_1_330), .ZN(n_1_1_329));
   AOI221_X1 i_1_1_710 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[3]), .C1(
      RAM_Data_RD_B[3]), .C2(n_1_1_473), .ZN(n_1_1_330));
   NAND2_X1 i_1_1_711 (.A1(RAM_Data_RD_A[3]), .A2(n_1_1_477), .ZN(n_1_1_332));
   INV_X1 i_1_1_712 (.A(Q[3]), .ZN(n_1_1_333));
   INV_X1 i_1_1_713 (.A(n_1_1_334), .ZN(n_250));
   OAI221_X1 i_1_1_714 (.A(n_1_1_335), .B1(adder_out2[4]), .B2(n_1_1_393), 
      .C1(RAM_Data_RD_B[4]), .C2(n_1_1_394), .ZN(n_1_1_334));
   AOI22_X1 i_1_1_715 (.A1(n_1_1_382), .A2(n_1_1_338), .B1(n_1_1_337), .B2(
      n_1_1_336), .ZN(n_1_1_335));
   AOI221_X1 i_1_1_716 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[4]), .C1(
      RAM_Data_RD_B[4]), .C2(n_1_1_473), .ZN(n_1_1_336));
   NAND2_X1 i_1_1_717 (.A1(RAM_Data_RD_A[4]), .A2(n_1_1_477), .ZN(n_1_1_337));
   INV_X1 i_1_1_718 (.A(Q[4]), .ZN(n_1_1_338));
   INV_X1 i_1_1_719 (.A(n_1_1_339), .ZN(n_251));
   OAI221_X1 i_1_1_720 (.A(n_1_1_340), .B1(adder_out2[5]), .B2(n_1_1_393), 
      .C1(RAM_Data_RD_B[5]), .C2(n_1_1_394), .ZN(n_1_1_339));
   AOI22_X1 i_1_1_721 (.A1(n_1_1_382), .A2(n_1_1_343), .B1(n_1_1_342), .B2(
      n_1_1_341), .ZN(n_1_1_340));
   AOI221_X1 i_1_1_723 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[5]), .C1(
      RAM_Data_RD_B[5]), .C2(n_1_1_473), .ZN(n_1_1_341));
   NAND2_X1 i_1_1_724 (.A1(RAM_Data_RD_A[5]), .A2(n_1_1_477), .ZN(n_1_1_342));
   INV_X1 i_1_1_725 (.A(Q[5]), .ZN(n_1_1_343));
   INV_X1 i_1_1_726 (.A(n_1_1_345), .ZN(n_252));
   OAI221_X1 i_1_1_727 (.A(n_1_1_346), .B1(adder_out2[6]), .B2(n_1_1_393), 
      .C1(RAM_Data_RD_B[6]), .C2(n_1_1_394), .ZN(n_1_1_345));
   AOI22_X1 i_1_1_736 (.A1(n_1_1_382), .A2(n_1_1_355), .B1(n_1_1_348), .B2(
      n_1_1_347), .ZN(n_1_1_346));
   AOI221_X1 i_1_1_737 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[6]), .C1(
      RAM_Data_RD_B[6]), .C2(n_1_1_473), .ZN(n_1_1_347));
   NAND2_X1 i_1_1_738 (.A1(RAM_Data_RD_A[6]), .A2(n_1_1_477), .ZN(n_1_1_348));
   INV_X1 i_1_1_739 (.A(Q[6]), .ZN(n_1_1_355));
   AOI21_X1 i_1_1_740 (.A(n_1_1_356), .B1(n_1_1_450), .B2(n_1_1_600), .ZN(n_253));
   OAI221_X1 i_1_1_741 (.A(n_1_1_357), .B1(n_1_1_393), .B2(adder_out2[7]), 
      .C1(n_1_1_394), .C2(RAM_Data_RD_B[7]), .ZN(n_1_1_356));
   NAND2_X1 i_1_1_742 (.A1(n_1_1_325), .A2(n_1_1_460), .ZN(n_1_1_357));
   INV_X1 i_1_1_743 (.A(n_1_1_358), .ZN(n_254));
   OAI221_X1 i_1_1_744 (.A(n_1_1_359), .B1(adder_out2[8]), .B2(n_1_1_393), 
      .C1(RAM_Data_RD_B[8]), .C2(n_1_1_394), .ZN(n_1_1_358));
   AOI22_X1 i_1_1_745 (.A1(n_1_1_382), .A2(n_1_1_362), .B1(n_1_1_361), .B2(
      n_1_1_360), .ZN(n_1_1_359));
   AOI221_X1 i_1_1_746 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[8]), .C1(
      RAM_Data_RD_B[8]), .C2(n_1_1_473), .ZN(n_1_1_360));
   NAND2_X1 i_1_1_747 (.A1(RAM_Data_RD_A[8]), .A2(n_1_1_477), .ZN(n_1_1_361));
   INV_X1 i_1_1_748 (.A(Q[8]), .ZN(n_1_1_362));
   AOI21_X1 i_1_1_749 (.A(n_1_1_363), .B1(n_1_1_450), .B2(n_1_1_601), .ZN(n_255));
   OAI221_X1 i_1_1_750 (.A(n_1_1_364), .B1(n_1_1_393), .B2(adder_out2[9]), 
      .C1(n_1_1_394), .C2(RAM_Data_RD_B[9]), .ZN(n_1_1_363));
   NAND2_X1 i_1_1_751 (.A1(n_1_1_331), .A2(n_1_1_460), .ZN(n_1_1_364));
   INV_X1 i_1_1_752 (.A(n_1_1_365), .ZN(n_256));
   OAI221_X1 i_1_1_753 (.A(n_1_1_366), .B1(adder_out2[10]), .B2(n_1_1_393), 
      .C1(RAM_Data_RD_B[10]), .C2(n_1_1_394), .ZN(n_1_1_365));
   AOI22_X1 i_1_1_754 (.A1(n_1_1_382), .A2(n_1_1_369), .B1(n_1_1_368), .B2(
      n_1_1_367), .ZN(n_1_1_366));
   AOI221_X1 i_1_1_755 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[10]), .C1(
      RAM_Data_RD_B[10]), .C2(n_1_1_473), .ZN(n_1_1_367));
   NAND2_X1 i_1_1_756 (.A1(RAM_Data_RD_A[10]), .A2(n_1_1_477), .ZN(n_1_1_368));
   INV_X1 i_1_1_757 (.A(Q[10]), .ZN(n_1_1_369));
   INV_X1 i_1_1_758 (.A(n_1_1_370), .ZN(n_257));
   OAI221_X1 i_1_1_759 (.A(n_1_1_371), .B1(adder_out2[11]), .B2(n_1_1_393), 
      .C1(RAM_Data_RD_B[11]), .C2(n_1_1_394), .ZN(n_1_1_370));
   AOI22_X1 i_1_1_760 (.A1(n_1_1_382), .A2(n_1_1_374), .B1(n_1_1_373), .B2(
      n_1_1_372), .ZN(n_1_1_371));
   AOI221_X1 i_1_1_761 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[11]), .C1(
      RAM_Data_RD_B[11]), .C2(n_1_1_473), .ZN(n_1_1_372));
   NAND2_X1 i_1_1_762 (.A1(RAM_Data_RD_A[11]), .A2(n_1_1_477), .ZN(n_1_1_373));
   INV_X1 i_1_1_763 (.A(Q[11]), .ZN(n_1_1_374));
   INV_X1 i_1_1_764 (.A(n_1_1_375), .ZN(n_258));
   OAI221_X1 i_1_1_765 (.A(n_1_1_376), .B1(adder_out2[12]), .B2(n_1_1_393), 
      .C1(RAM_Data_RD_B[12]), .C2(n_1_1_394), .ZN(n_1_1_375));
   AOI22_X1 i_1_1_766 (.A1(n_1_1_382), .A2(n_1_1_379), .B1(n_1_1_378), .B2(
      n_1_1_377), .ZN(n_1_1_376));
   AOI221_X1 i_1_1_767 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[12]), .C1(
      RAM_Data_RD_B[12]), .C2(n_1_1_473), .ZN(n_1_1_377));
   NAND2_X1 i_1_1_768 (.A1(RAM_Data_RD_A[12]), .A2(n_1_1_477), .ZN(n_1_1_378));
   INV_X1 i_1_1_769 (.A(Q[12]), .ZN(n_1_1_379));
   INV_X1 i_1_1_770 (.A(n_1_1_380), .ZN(n_259));
   OAI221_X1 i_1_1_771 (.A(n_1_1_381), .B1(adder_out2[13]), .B2(n_1_1_393), 
      .C1(RAM_Data_RD_B[13]), .C2(n_1_1_394), .ZN(n_1_1_380));
   AOI22_X1 i_1_1_772 (.A1(n_1_1_382), .A2(n_1_1_383), .B1(n_1_1_344), .B2(
      n_1_1_460), .ZN(n_1_1_381));
   INV_X1 i_1_1_773 (.A(n_1_1_830), .ZN(n_1_1_382));
   INV_X1 i_1_1_774 (.A(Q[14]), .ZN(n_1_1_383));
   INV_X1 i_1_1_775 (.A(n_1_1_384), .ZN(n_260));
   OAI221_X1 i_1_1_776 (.A(n_1_1_385), .B1(RAM_Data_RD_B[14]), .B2(n_1_1_394), 
      .C1(Q[14]), .C2(n_1_1_830), .ZN(n_1_1_384));
   INV_X1 i_1_1_777 (.A(n_1_1_386), .ZN(n_1_1_385));
   NAND2_X1 i_1_1_778 (.A1(n_1_1_392), .A2(n_1_1_387), .ZN(n_1_1_386));
   OAI221_X1 i_1_1_779 (.A(n_1_1_388), .B1(n_1_1_640), .B2(n_1_1_389), .C1(
      n_1_1_391), .C2(n_1_1_390), .ZN(n_1_1_387));
   AOI21_X1 i_1_1_780 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[14]), .ZN(n_1_1_388));
   INV_X1 i_1_1_781 (.A(n_1_1_477), .ZN(n_1_1_389));
   INV_X1 i_1_1_782 (.A(n_1_1_473), .ZN(n_1_1_390));
   INV_X1 i_1_1_783 (.A(RAM_Data_RD_B[14]), .ZN(n_1_1_391));
   OR2_X1 i_1_1_784 (.A1(n_1_1_393), .A2(adder_out2[14]), .ZN(n_1_1_392));
   NAND3_X1 i_1_1_785 (.A1(n_1_1_846), .A2(adder_out1[12]), .A3(n_1_1_451), 
      .ZN(n_1_1_393));
   NAND2_X1 i_1_1_786 (.A1(n_1_1_455), .A2(n_1_1_451), .ZN(n_1_1_394));
   INV_X1 i_1_1_787 (.A(n_1_1_833), .ZN(n_1_1_455));
   INV_X1 i_1_1_788 (.A(n_1_1_395), .ZN(n_261));
   NAND2_X1 i_1_1_789 (.A1(n_1_1_830), .A2(n_1_1_396), .ZN(n_1_1_395));
   OAI21_X1 i_1_1_790 (.A(n_1_1_397), .B1(n_1_1_825), .B2(n_1_1_399), .ZN(
      n_1_1_396));
   OAI21_X1 i_1_1_791 (.A(RAM_Data_RD_B[17]), .B1(n_1_1_398), .B2(n_1_1_473), 
      .ZN(n_1_1_397));
   INV_X1 i_1_1_792 (.A(n_1_1_399), .ZN(n_1_1_398));
   AOI221_X1 i_1_1_793 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[17]), .C1(
      RAM_Data_RD_A[17]), .C2(n_1_1_477), .ZN(n_1_1_399));
   INV_X1 i_1_1_794 (.A(n_1_1_400), .ZN(n_262));
   NAND2_X1 i_1_1_795 (.A1(n_1_1_830), .A2(n_1_1_401), .ZN(n_1_1_400));
   OAI21_X1 i_1_1_796 (.A(n_1_1_402), .B1(n_1_1_825), .B2(n_1_1_404), .ZN(
      n_1_1_401));
   OAI21_X1 i_1_1_797 (.A(RAM_Data_RD_B[18]), .B1(n_1_1_403), .B2(n_1_1_473), 
      .ZN(n_1_1_402));
   INV_X1 i_1_1_798 (.A(n_1_1_404), .ZN(n_1_1_403));
   AOI221_X1 i_1_1_799 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[18]), .C1(
      RAM_Data_RD_A[18]), .C2(n_1_1_477), .ZN(n_1_1_404));
   INV_X1 i_1_1_800 (.A(n_1_1_405), .ZN(n_263));
   NAND2_X1 i_1_1_801 (.A1(n_1_1_830), .A2(n_1_1_406), .ZN(n_1_1_405));
   OAI21_X1 i_1_1_802 (.A(n_1_1_407), .B1(n_1_1_825), .B2(n_1_1_409), .ZN(
      n_1_1_406));
   OAI21_X1 i_1_1_803 (.A(RAM_Data_RD_B[19]), .B1(n_1_1_408), .B2(n_1_1_473), 
      .ZN(n_1_1_407));
   INV_X1 i_1_1_804 (.A(n_1_1_409), .ZN(n_1_1_408));
   AOI221_X1 i_1_1_805 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[19]), .C1(
      RAM_Data_RD_A[19]), .C2(n_1_1_477), .ZN(n_1_1_409));
   INV_X1 i_1_1_806 (.A(n_1_1_410), .ZN(n_264));
   NAND2_X1 i_1_1_807 (.A1(n_1_1_830), .A2(n_1_1_411), .ZN(n_1_1_410));
   OAI21_X1 i_1_1_808 (.A(n_1_1_412), .B1(n_1_1_825), .B2(n_1_1_414), .ZN(
      n_1_1_411));
   OAI21_X1 i_1_1_809 (.A(RAM_Data_RD_B[20]), .B1(n_1_1_413), .B2(n_1_1_473), 
      .ZN(n_1_1_412));
   INV_X1 i_1_1_810 (.A(n_1_1_414), .ZN(n_1_1_413));
   AOI221_X1 i_1_1_811 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[20]), .C1(
      RAM_Data_RD_A[20]), .C2(n_1_1_477), .ZN(n_1_1_414));
   INV_X1 i_1_1_812 (.A(n_1_1_415), .ZN(n_265));
   NAND2_X1 i_1_1_813 (.A1(n_1_1_830), .A2(n_1_1_416), .ZN(n_1_1_415));
   OAI21_X1 i_1_1_814 (.A(n_1_1_417), .B1(n_1_1_825), .B2(n_1_1_419), .ZN(
      n_1_1_416));
   OAI21_X1 i_1_1_815 (.A(RAM_Data_RD_B[21]), .B1(n_1_1_418), .B2(n_1_1_473), 
      .ZN(n_1_1_417));
   INV_X1 i_1_1_816 (.A(n_1_1_419), .ZN(n_1_1_418));
   AOI221_X1 i_1_1_817 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[21]), .C1(
      RAM_Data_RD_A[21]), .C2(n_1_1_477), .ZN(n_1_1_419));
   INV_X1 i_1_1_818 (.A(n_1_1_420), .ZN(n_266));
   NAND2_X1 i_1_1_819 (.A1(n_1_1_830), .A2(n_1_1_421), .ZN(n_1_1_420));
   OAI21_X1 i_1_1_820 (.A(n_1_1_422), .B1(n_1_1_825), .B2(n_1_1_424), .ZN(
      n_1_1_421));
   OAI21_X1 i_1_1_821 (.A(RAM_Data_RD_B[22]), .B1(n_1_1_423), .B2(n_1_1_473), 
      .ZN(n_1_1_422));
   INV_X1 i_1_1_822 (.A(n_1_1_424), .ZN(n_1_1_423));
   AOI221_X1 i_1_1_823 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[22]), .C1(
      RAM_Data_RD_A[22]), .C2(n_1_1_477), .ZN(n_1_1_424));
   INV_X1 i_1_1_824 (.A(n_1_1_425), .ZN(n_267));
   NAND2_X1 i_1_1_825 (.A1(n_1_1_830), .A2(n_1_1_426), .ZN(n_1_1_425));
   OAI21_X1 i_1_1_826 (.A(n_1_1_427), .B1(n_1_1_825), .B2(n_1_1_429), .ZN(
      n_1_1_426));
   OAI21_X1 i_1_1_827 (.A(RAM_Data_RD_B[23]), .B1(n_1_1_428), .B2(n_1_1_473), 
      .ZN(n_1_1_427));
   INV_X1 i_1_1_828 (.A(n_1_1_429), .ZN(n_1_1_428));
   AOI221_X1 i_1_1_829 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[23]), .C1(
      RAM_Data_RD_A[23]), .C2(n_1_1_477), .ZN(n_1_1_429));
   INV_X1 i_1_1_830 (.A(n_1_1_430), .ZN(n_268));
   NAND2_X1 i_1_1_831 (.A1(n_1_1_830), .A2(n_1_1_431), .ZN(n_1_1_430));
   OAI21_X1 i_1_1_832 (.A(n_1_1_432), .B1(n_1_1_825), .B2(n_1_1_434), .ZN(
      n_1_1_431));
   OAI21_X1 i_1_1_833 (.A(RAM_Data_RD_B[24]), .B1(n_1_1_433), .B2(n_1_1_473), 
      .ZN(n_1_1_432));
   INV_X1 i_1_1_834 (.A(n_1_1_434), .ZN(n_1_1_433));
   AOI221_X1 i_1_1_835 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[24]), .C1(
      RAM_Data_RD_A[24]), .C2(n_1_1_477), .ZN(n_1_1_434));
   INV_X1 i_1_1_836 (.A(n_1_1_435), .ZN(n_269));
   NAND2_X1 i_1_1_837 (.A1(n_1_1_830), .A2(n_1_1_436), .ZN(n_1_1_435));
   OAI21_X1 i_1_1_838 (.A(n_1_1_437), .B1(n_1_1_825), .B2(n_1_1_439), .ZN(
      n_1_1_436));
   OAI21_X1 i_1_1_839 (.A(RAM_Data_RD_B[25]), .B1(n_1_1_438), .B2(n_1_1_473), 
      .ZN(n_1_1_437));
   INV_X1 i_1_1_840 (.A(n_1_1_439), .ZN(n_1_1_438));
   AOI221_X1 i_1_1_841 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[25]), .C1(
      RAM_Data_RD_A[25]), .C2(n_1_1_477), .ZN(n_1_1_439));
   INV_X1 i_1_1_842 (.A(n_1_1_440), .ZN(n_270));
   NAND2_X1 i_1_1_843 (.A1(n_1_1_830), .A2(n_1_1_441), .ZN(n_1_1_440));
   OAI21_X1 i_1_1_844 (.A(n_1_1_442), .B1(n_1_1_825), .B2(n_1_1_444), .ZN(
      n_1_1_441));
   OAI21_X1 i_1_1_845 (.A(RAM_Data_RD_B[26]), .B1(n_1_1_443), .B2(n_1_1_473), 
      .ZN(n_1_1_442));
   INV_X1 i_1_1_846 (.A(n_1_1_444), .ZN(n_1_1_443));
   AOI221_X1 i_1_1_847 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[26]), .C1(
      RAM_Data_RD_A[26]), .C2(n_1_1_477), .ZN(n_1_1_444));
   INV_X1 i_1_1_848 (.A(n_1_1_445), .ZN(n_271));
   NAND2_X1 i_1_1_849 (.A1(n_1_1_830), .A2(n_1_1_446), .ZN(n_1_1_445));
   OAI21_X1 i_1_1_850 (.A(n_1_1_447), .B1(n_1_1_825), .B2(n_1_1_449), .ZN(
      n_1_1_446));
   OAI21_X1 i_1_1_851 (.A(RAM_Data_RD_B[27]), .B1(n_1_1_448), .B2(n_1_1_473), 
      .ZN(n_1_1_447));
   INV_X1 i_1_1_852 (.A(n_1_1_449), .ZN(n_1_1_448));
   AOI221_X1 i_1_1_853 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[27]), .C1(
      RAM_Data_RD_A[27]), .C2(n_1_1_477), .ZN(n_1_1_449));
   INV_X1 i_1_1_854 (.A(n_1_1_453), .ZN(n_272));
   NAND2_X1 i_1_1_855 (.A1(n_1_1_830), .A2(n_1_1_454), .ZN(n_1_1_453));
   OAI21_X1 i_1_1_856 (.A(n_1_1_456), .B1(n_1_1_825), .B2(n_1_1_537), .ZN(
      n_1_1_454));
   OAI21_X1 i_1_1_857 (.A(RAM_Data_RD_B[28]), .B1(n_1_1_484), .B2(n_1_1_473), 
      .ZN(n_1_1_456));
   INV_X1 i_1_1_858 (.A(n_1_1_537), .ZN(n_1_1_484));
   AOI221_X1 i_1_1_859 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[28]), .C1(
      RAM_Data_RD_A[28]), .C2(n_1_1_477), .ZN(n_1_1_537));
   INV_X1 i_1_1_860 (.A(n_1_1_538), .ZN(n_273));
   NAND2_X1 i_1_1_861 (.A1(n_1_1_830), .A2(n_1_1_539), .ZN(n_1_1_538));
   OAI21_X1 i_1_1_862 (.A(n_1_1_542), .B1(n_1_1_825), .B2(n_1_1_564), .ZN(
      n_1_1_539));
   OAI21_X1 i_1_1_863 (.A(RAM_Data_RD_B[29]), .B1(n_1_1_543), .B2(n_1_1_473), 
      .ZN(n_1_1_542));
   INV_X1 i_1_1_864 (.A(n_1_1_564), .ZN(n_1_1_543));
   AOI221_X1 i_1_1_865 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[29]), .C1(
      RAM_Data_RD_A[29]), .C2(n_1_1_477), .ZN(n_1_1_564));
   INV_X1 i_1_1_866 (.A(n_1_1_565), .ZN(n_274));
   NAND2_X1 i_1_1_867 (.A1(n_1_1_830), .A2(n_1_1_566), .ZN(n_1_1_565));
   OAI21_X1 i_1_1_868 (.A(n_1_1_567), .B1(n_1_1_825), .B2(n_1_1_569), .ZN(
      n_1_1_566));
   OAI21_X1 i_1_1_869 (.A(RAM_Data_RD_B[30]), .B1(n_1_1_568), .B2(n_1_1_473), 
      .ZN(n_1_1_567));
   INV_X1 i_1_1_870 (.A(n_1_1_569), .ZN(n_1_1_568));
   AOI221_X1 i_1_1_871 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[30]), .C1(
      RAM_Data_RD_A[30]), .C2(n_1_1_477), .ZN(n_1_1_569));
   INV_X1 i_1_1_872 (.A(n_1_1_570), .ZN(n_275));
   NAND2_X1 i_1_1_873 (.A1(n_1_1_830), .A2(n_1_1_571), .ZN(n_1_1_570));
   OAI21_X1 i_1_1_874 (.A(n_1_1_572), .B1(n_1_1_825), .B2(n_1_1_574), .ZN(
      n_1_1_571));
   OAI21_X1 i_1_1_875 (.A(RAM_Data_RD_B[31]), .B1(n_1_1_573), .B2(n_1_1_473), 
      .ZN(n_1_1_572));
   INV_X1 i_1_1_876 (.A(n_1_1_574), .ZN(n_1_1_573));
   AOI221_X1 i_1_1_878 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[31]), .C1(
      RAM_Data_RD_A[31]), .C2(n_1_1_477), .ZN(n_1_1_574));
   INV_X1 i_1_1_880 (.A(n_1_1_575), .ZN(n_276));
   NAND2_X1 i_1_1_881 (.A1(n_1_1_830), .A2(n_1_1_576), .ZN(n_1_1_575));
   OAI21_X1 i_1_1_882 (.A(n_1_1_577), .B1(n_1_1_825), .B2(n_1_1_579), .ZN(
      n_1_1_576));
   OAI21_X1 i_1_1_883 (.A(RAM_Data_RD_B[32]), .B1(n_1_1_578), .B2(n_1_1_473), 
      .ZN(n_1_1_577));
   INV_X1 i_1_1_884 (.A(n_1_1_579), .ZN(n_1_1_578));
   AOI221_X1 i_1_1_885 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[32]), .C1(
      RAM_Data_RD_A[32]), .C2(n_1_1_477), .ZN(n_1_1_579));
   INV_X1 i_1_1_886 (.A(n_1_1_580), .ZN(n_277));
   NAND2_X1 i_1_1_893 (.A1(n_1_1_830), .A2(n_1_1_602), .ZN(n_1_1_580));
   OAI21_X1 i_1_1_926 (.A(n_1_1_659), .B1(n_1_1_825), .B2(n_1_1_677), .ZN(
      n_1_1_602));
   OAI21_X1 i_1_1_927 (.A(RAM_Data_RD_B[33]), .B1(n_1_1_676), .B2(n_1_1_473), 
      .ZN(n_1_1_659));
   INV_X1 i_1_1_929 (.A(n_1_1_677), .ZN(n_1_1_676));
   AOI221_X1 i_1_1_930 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[33]), .C1(
      RAM_Data_RD_A[33]), .C2(n_1_1_477), .ZN(n_1_1_677));
   INV_X1 i_1_1_932 (.A(n_1_1_678), .ZN(n_278));
   NAND2_X1 i_1_1_981 (.A1(n_1_1_830), .A2(n_1_1_679), .ZN(n_1_1_678));
   OAI21_X1 i_1_1_984 (.A(n_1_1_680), .B1(n_1_1_825), .B2(n_1_1_682), .ZN(
      n_1_1_679));
   OAI21_X1 i_1_1_985 (.A(RAM_Data_RD_B[34]), .B1(n_1_1_681), .B2(n_1_1_473), 
      .ZN(n_1_1_680));
   INV_X1 i_1_1_986 (.A(n_1_1_682), .ZN(n_1_1_681));
   AOI221_X1 i_1_1_987 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[34]), .C1(
      RAM_Data_RD_A[34]), .C2(n_1_1_477), .ZN(n_1_1_682));
   INV_X1 i_1_1_989 (.A(n_1_1_683), .ZN(n_279));
   NAND2_X1 i_1_1_990 (.A1(n_1_1_830), .A2(n_1_1_684), .ZN(n_1_1_683));
   OAI21_X1 i_1_1_991 (.A(n_1_1_685), .B1(n_1_1_825), .B2(n_1_1_687), .ZN(
      n_1_1_684));
   OAI21_X1 i_1_1_992 (.A(RAM_Data_RD_B[35]), .B1(n_1_1_686), .B2(n_1_1_473), 
      .ZN(n_1_1_685));
   INV_X1 i_1_1_993 (.A(n_1_1_687), .ZN(n_1_1_686));
   AOI221_X1 i_1_1_1010 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[35]), .C1(
      RAM_Data_RD_A[35]), .C2(n_1_1_477), .ZN(n_1_1_687));
   INV_X1 i_1_1_1011 (.A(n_1_1_688), .ZN(n_280));
   NAND2_X1 i_1_1_1012 (.A1(n_1_1_830), .A2(n_1_1_689), .ZN(n_1_1_688));
   OAI21_X1 i_1_1_1013 (.A(n_1_1_690), .B1(n_1_1_825), .B2(n_1_1_692), .ZN(
      n_1_1_689));
   OAI21_X1 i_1_1_1014 (.A(RAM_Data_RD_B[36]), .B1(n_1_1_691), .B2(n_1_1_473), 
      .ZN(n_1_1_690));
   INV_X1 i_1_1_1015 (.A(n_1_1_692), .ZN(n_1_1_691));
   AOI221_X1 i_1_1_1016 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[36]), .C1(
      RAM_Data_RD_A[36]), .C2(n_1_1_477), .ZN(n_1_1_692));
   INV_X1 i_1_1_1017 (.A(n_1_1_693), .ZN(n_281));
   NAND2_X1 i_1_1_1018 (.A1(n_1_1_830), .A2(n_1_1_694), .ZN(n_1_1_693));
   OAI21_X1 i_1_1_1019 (.A(n_1_1_695), .B1(n_1_1_825), .B2(n_1_1_697), .ZN(
      n_1_1_694));
   OAI21_X1 i_1_1_1020 (.A(RAM_Data_RD_B[37]), .B1(n_1_1_696), .B2(n_1_1_473), 
      .ZN(n_1_1_695));
   INV_X1 i_1_1_1021 (.A(n_1_1_697), .ZN(n_1_1_696));
   AOI221_X1 i_1_1_1022 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[37]), .C1(
      RAM_Data_RD_A[37]), .C2(n_1_1_477), .ZN(n_1_1_697));
   INV_X1 i_1_1_1023 (.A(n_1_1_698), .ZN(n_282));
   NAND2_X1 i_1_1_1024 (.A1(n_1_1_830), .A2(n_1_1_699), .ZN(n_1_1_698));
   OAI21_X1 i_1_1_1025 (.A(n_1_1_700), .B1(n_1_1_825), .B2(n_1_1_702), .ZN(
      n_1_1_699));
   OAI21_X1 i_1_1_1026 (.A(RAM_Data_RD_B[38]), .B1(n_1_1_701), .B2(n_1_1_473), 
      .ZN(n_1_1_700));
   INV_X1 i_1_1_1027 (.A(n_1_1_702), .ZN(n_1_1_701));
   AOI221_X1 i_1_1_1028 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[38]), .C1(
      RAM_Data_RD_A[38]), .C2(n_1_1_477), .ZN(n_1_1_702));
   INV_X1 i_1_1_1029 (.A(n_1_1_703), .ZN(n_283));
   NAND2_X1 i_1_1_1030 (.A1(n_1_1_830), .A2(n_1_1_704), .ZN(n_1_1_703));
   OAI21_X1 i_1_1_1042 (.A(n_1_1_705), .B1(n_1_1_825), .B2(n_1_1_707), .ZN(
      n_1_1_704));
   OAI21_X1 i_1_1_1044 (.A(RAM_Data_RD_B[39]), .B1(n_1_1_706), .B2(n_1_1_473), 
      .ZN(n_1_1_705));
   INV_X1 i_1_1_1045 (.A(n_1_1_707), .ZN(n_1_1_706));
   AOI221_X1 i_1_1_1055 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[39]), .C1(
      RAM_Data_RD_A[39]), .C2(n_1_1_477), .ZN(n_1_1_707));
   INV_X1 i_1_1_1064 (.A(n_1_1_708), .ZN(n_284));
   NAND2_X1 i_1_1_1065 (.A1(n_1_1_830), .A2(n_1_1_709), .ZN(n_1_1_708));
   OAI21_X1 i_1_1_1066 (.A(n_1_1_710), .B1(n_1_1_825), .B2(n_1_1_712), .ZN(
      n_1_1_709));
   OAI21_X1 i_1_1_1067 (.A(RAM_Data_RD_B[40]), .B1(n_1_1_711), .B2(n_1_1_473), 
      .ZN(n_1_1_710));
   INV_X1 i_1_1_1068 (.A(n_1_1_712), .ZN(n_1_1_711));
   AOI221_X1 i_1_1_1069 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[40]), .C1(
      RAM_Data_RD_A[40]), .C2(n_1_1_477), .ZN(n_1_1_712));
   INV_X1 i_1_1_1070 (.A(n_1_1_713), .ZN(n_285));
   NAND2_X1 i_1_1_1071 (.A1(n_1_1_830), .A2(n_1_1_714), .ZN(n_1_1_713));
   OAI21_X1 i_1_1_1072 (.A(n_1_1_715), .B1(n_1_1_825), .B2(n_1_1_717), .ZN(
      n_1_1_714));
   OAI21_X1 i_1_1_1073 (.A(RAM_Data_RD_B[41]), .B1(n_1_1_716), .B2(n_1_1_473), 
      .ZN(n_1_1_715));
   INV_X1 i_1_1_1074 (.A(n_1_1_717), .ZN(n_1_1_716));
   AOI221_X1 i_1_1_1075 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[41]), .C1(
      RAM_Data_RD_A[41]), .C2(n_1_1_477), .ZN(n_1_1_717));
   INV_X1 i_1_1_1076 (.A(n_1_1_718), .ZN(n_286));
   NAND2_X1 i_1_1_1077 (.A1(n_1_1_830), .A2(n_1_1_719), .ZN(n_1_1_718));
   OAI21_X1 i_1_1_1078 (.A(n_1_1_720), .B1(n_1_1_825), .B2(n_1_1_722), .ZN(
      n_1_1_719));
   OAI21_X1 i_1_1_1079 (.A(RAM_Data_RD_B[42]), .B1(n_1_1_721), .B2(n_1_1_473), 
      .ZN(n_1_1_720));
   INV_X1 i_1_1_1080 (.A(n_1_1_722), .ZN(n_1_1_721));
   AOI221_X1 i_1_1_1081 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[42]), .C1(
      RAM_Data_RD_A[42]), .C2(n_1_1_477), .ZN(n_1_1_722));
   INV_X1 i_1_1_1082 (.A(n_1_1_723), .ZN(n_287));
   NAND2_X1 i_1_1_1083 (.A1(n_1_1_830), .A2(n_1_1_724), .ZN(n_1_1_723));
   OAI21_X1 i_1_1_1084 (.A(n_1_1_725), .B1(n_1_1_825), .B2(n_1_1_727), .ZN(
      n_1_1_724));
   OAI21_X1 i_1_1_1085 (.A(RAM_Data_RD_B[43]), .B1(n_1_1_726), .B2(n_1_1_473), 
      .ZN(n_1_1_725));
   INV_X1 i_1_1_1086 (.A(n_1_1_727), .ZN(n_1_1_726));
   AOI221_X1 i_1_1_1087 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[43]), .C1(
      RAM_Data_RD_A[43]), .C2(n_1_1_477), .ZN(n_1_1_727));
   INV_X1 i_1_1_1088 (.A(n_1_1_728), .ZN(n_288));
   NAND2_X1 i_1_1_1089 (.A1(n_1_1_830), .A2(n_1_1_729), .ZN(n_1_1_728));
   OAI21_X1 i_1_1_1090 (.A(n_1_1_730), .B1(n_1_1_825), .B2(n_1_1_732), .ZN(
      n_1_1_729));
   OAI21_X1 i_1_1_1091 (.A(RAM_Data_RD_B[44]), .B1(n_1_1_731), .B2(n_1_1_473), 
      .ZN(n_1_1_730));
   INV_X1 i_1_1_1092 (.A(n_1_1_732), .ZN(n_1_1_731));
   AOI221_X1 i_1_1_1115 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[44]), .C1(
      RAM_Data_RD_A[44]), .C2(n_1_1_477), .ZN(n_1_1_732));
   INV_X1 i_1_1_1122 (.A(n_1_1_733), .ZN(n_289));
   NAND2_X1 i_1_1_1127 (.A1(n_1_1_830), .A2(n_1_1_734), .ZN(n_1_1_733));
   OAI21_X1 i_1_1_1128 (.A(n_1_1_735), .B1(n_1_1_825), .B2(n_1_1_737), .ZN(
      n_1_1_734));
   OAI21_X1 i_1_1_1129 (.A(RAM_Data_RD_B[45]), .B1(n_1_1_736), .B2(n_1_1_473), 
      .ZN(n_1_1_735));
   INV_X1 i_1_1_1130 (.A(n_1_1_737), .ZN(n_1_1_736));
   AOI221_X1 i_1_1_1131 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[45]), .C1(
      RAM_Data_RD_A[45]), .C2(n_1_1_477), .ZN(n_1_1_737));
   INV_X1 i_1_1_1132 (.A(n_1_1_738), .ZN(n_290));
   NAND2_X1 i_1_1_1133 (.A1(n_1_1_830), .A2(n_1_1_739), .ZN(n_1_1_738));
   OAI21_X1 i_1_1_1134 (.A(n_1_1_740), .B1(n_1_1_825), .B2(n_1_1_742), .ZN(
      n_1_1_739));
   OAI21_X1 i_1_1_1135 (.A(RAM_Data_RD_B[46]), .B1(n_1_1_741), .B2(n_1_1_473), 
      .ZN(n_1_1_740));
   INV_X1 i_1_1_1136 (.A(n_1_1_742), .ZN(n_1_1_741));
   AOI221_X1 i_1_1_1137 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[46]), .C1(
      RAM_Data_RD_A[46]), .C2(n_1_1_477), .ZN(n_1_1_742));
   INV_X1 i_1_1_1138 (.A(n_1_1_743), .ZN(n_291));
   NAND2_X1 i_1_1_1139 (.A1(n_1_1_830), .A2(n_1_1_744), .ZN(n_1_1_743));
   OAI21_X1 i_1_1_1140 (.A(n_1_1_745), .B1(n_1_1_825), .B2(n_1_1_747), .ZN(
      n_1_1_744));
   OAI21_X1 i_1_1_1141 (.A(RAM_Data_RD_B[47]), .B1(n_1_1_746), .B2(n_1_1_473), 
      .ZN(n_1_1_745));
   INV_X1 i_1_1_1142 (.A(n_1_1_747), .ZN(n_1_1_746));
   AOI221_X1 i_1_1_1143 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[47]), .C1(
      RAM_Data_RD_A[47]), .C2(n_1_1_477), .ZN(n_1_1_747));
   INV_X1 i_1_1_1144 (.A(n_1_1_748), .ZN(n_292));
   NAND2_X1 i_1_1_1145 (.A1(n_1_1_830), .A2(n_1_1_749), .ZN(n_1_1_748));
   OAI21_X1 i_1_1_1146 (.A(n_1_1_750), .B1(n_1_1_825), .B2(n_1_1_752), .ZN(
      n_1_1_749));
   OAI21_X1 i_1_1_1147 (.A(RAM_Data_RD_B[48]), .B1(n_1_1_751), .B2(n_1_1_473), 
      .ZN(n_1_1_750));
   INV_X1 i_1_1_1148 (.A(n_1_1_752), .ZN(n_1_1_751));
   AOI221_X1 i_1_1_1149 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[48]), .C1(
      RAM_Data_RD_A[48]), .C2(n_1_1_477), .ZN(n_1_1_752));
   INV_X1 i_1_1_1150 (.A(n_1_1_753), .ZN(n_293));
   NAND2_X1 i_1_1_1151 (.A1(n_1_1_830), .A2(n_1_1_754), .ZN(n_1_1_753));
   OAI21_X1 i_1_1_1152 (.A(n_1_1_755), .B1(n_1_1_825), .B2(n_1_1_757), .ZN(
      n_1_1_754));
   OAI21_X1 i_1_1_1153 (.A(RAM_Data_RD_B[49]), .B1(n_1_1_756), .B2(n_1_1_473), 
      .ZN(n_1_1_755));
   INV_X1 i_1_1_1154 (.A(n_1_1_757), .ZN(n_1_1_756));
   AOI221_X1 i_1_1_1155 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[49]), .C1(
      RAM_Data_RD_A[49]), .C2(n_1_1_477), .ZN(n_1_1_757));
   INV_X1 i_1_1_1156 (.A(n_1_1_758), .ZN(n_294));
   NAND2_X1 i_1_1_1157 (.A1(n_1_1_830), .A2(n_1_1_759), .ZN(n_1_1_758));
   OAI21_X1 i_1_1_1158 (.A(n_1_1_760), .B1(n_1_1_825), .B2(n_1_1_762), .ZN(
      n_1_1_759));
   OAI21_X1 i_1_1_1159 (.A(RAM_Data_RD_B[50]), .B1(n_1_1_761), .B2(n_1_1_473), 
      .ZN(n_1_1_760));
   INV_X1 i_1_1_1160 (.A(n_1_1_762), .ZN(n_1_1_761));
   AOI221_X1 i_1_1_1161 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[50]), .C1(
      RAM_Data_RD_A[50]), .C2(n_1_1_477), .ZN(n_1_1_762));
   INV_X1 i_1_1_1162 (.A(n_1_1_763), .ZN(n_295));
   NAND2_X1 i_1_1_1163 (.A1(n_1_1_830), .A2(n_1_1_764), .ZN(n_1_1_763));
   OAI21_X1 i_1_1_1164 (.A(n_1_1_765), .B1(n_1_1_825), .B2(n_1_1_767), .ZN(
      n_1_1_764));
   OAI21_X1 i_1_1_1165 (.A(RAM_Data_RD_B[51]), .B1(n_1_1_766), .B2(n_1_1_473), 
      .ZN(n_1_1_765));
   INV_X1 i_1_1_1166 (.A(n_1_1_767), .ZN(n_1_1_766));
   AOI221_X1 i_1_1_1167 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[51]), .C1(
      RAM_Data_RD_A[51]), .C2(n_1_1_477), .ZN(n_1_1_767));
   INV_X1 i_1_1_1168 (.A(n_1_1_768), .ZN(n_296));
   NAND2_X1 i_1_1_1169 (.A1(n_1_1_830), .A2(n_1_1_769), .ZN(n_1_1_768));
   OAI21_X1 i_1_1_1170 (.A(n_1_1_770), .B1(n_1_1_825), .B2(n_1_1_772), .ZN(
      n_1_1_769));
   OAI21_X1 i_1_1_1171 (.A(RAM_Data_RD_B[52]), .B1(n_1_1_771), .B2(n_1_1_473), 
      .ZN(n_1_1_770));
   INV_X1 i_1_1_1172 (.A(n_1_1_772), .ZN(n_1_1_771));
   AOI221_X1 i_1_1_1173 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[52]), .C1(
      RAM_Data_RD_A[52]), .C2(n_1_1_477), .ZN(n_1_1_772));
   INV_X1 i_1_1_1174 (.A(n_1_1_773), .ZN(n_297));
   NAND2_X1 i_1_1_1175 (.A1(n_1_1_830), .A2(n_1_1_774), .ZN(n_1_1_773));
   OAI21_X1 i_1_1_1176 (.A(n_1_1_775), .B1(n_1_1_825), .B2(n_1_1_777), .ZN(
      n_1_1_774));
   OAI21_X1 i_1_1_1177 (.A(RAM_Data_RD_B[53]), .B1(n_1_1_776), .B2(n_1_1_473), 
      .ZN(n_1_1_775));
   INV_X1 i_1_1_1178 (.A(n_1_1_777), .ZN(n_1_1_776));
   AOI221_X1 i_1_1_1179 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[53]), .C1(
      RAM_Data_RD_A[53]), .C2(n_1_1_477), .ZN(n_1_1_777));
   INV_X1 i_1_1_1180 (.A(n_1_1_778), .ZN(n_298));
   NAND2_X1 i_1_1_1181 (.A1(n_1_1_830), .A2(n_1_1_779), .ZN(n_1_1_778));
   OAI21_X1 i_1_1_1182 (.A(n_1_1_780), .B1(n_1_1_825), .B2(n_1_1_782), .ZN(
      n_1_1_779));
   OAI21_X1 i_1_1_1183 (.A(RAM_Data_RD_B[54]), .B1(n_1_1_781), .B2(n_1_1_473), 
      .ZN(n_1_1_780));
   INV_X1 i_1_1_1184 (.A(n_1_1_782), .ZN(n_1_1_781));
   AOI221_X1 i_1_1_1185 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[54]), .C1(
      RAM_Data_RD_A[54]), .C2(n_1_1_477), .ZN(n_1_1_782));
   INV_X1 i_1_1_1186 (.A(n_1_1_783), .ZN(n_299));
   NAND2_X1 i_1_1_1187 (.A1(n_1_1_830), .A2(n_1_1_784), .ZN(n_1_1_783));
   OAI21_X1 i_1_1_1188 (.A(n_1_1_785), .B1(n_1_1_825), .B2(n_1_1_787), .ZN(
      n_1_1_784));
   OAI21_X1 i_1_1_1189 (.A(RAM_Data_RD_B[55]), .B1(n_1_1_786), .B2(n_1_1_473), 
      .ZN(n_1_1_785));
   INV_X1 i_1_1_1190 (.A(n_1_1_787), .ZN(n_1_1_786));
   AOI221_X1 i_1_1_1191 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[55]), .C1(
      RAM_Data_RD_A[55]), .C2(n_1_1_477), .ZN(n_1_1_787));
   INV_X1 i_1_1_1192 (.A(n_1_1_788), .ZN(n_300));
   NAND2_X1 i_1_1_1193 (.A1(n_1_1_830), .A2(n_1_1_789), .ZN(n_1_1_788));
   OAI21_X1 i_1_1_1194 (.A(n_1_1_790), .B1(n_1_1_825), .B2(n_1_1_792), .ZN(
      n_1_1_789));
   OAI21_X1 i_1_1_1195 (.A(RAM_Data_RD_B[56]), .B1(n_1_1_791), .B2(n_1_1_473), 
      .ZN(n_1_1_790));
   INV_X1 i_1_1_1196 (.A(n_1_1_792), .ZN(n_1_1_791));
   AOI221_X1 i_1_1_1197 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[56]), .C1(
      RAM_Data_RD_A[56]), .C2(n_1_1_477), .ZN(n_1_1_792));
   INV_X1 i_1_1_1198 (.A(n_1_1_793), .ZN(n_301));
   NAND2_X1 i_1_1_1199 (.A1(n_1_1_830), .A2(n_1_1_794), .ZN(n_1_1_793));
   OAI21_X1 i_1_1_1200 (.A(n_1_1_795), .B1(n_1_1_825), .B2(n_1_1_797), .ZN(
      n_1_1_794));
   OAI21_X1 i_1_1_1201 (.A(RAM_Data_RD_B[57]), .B1(n_1_1_796), .B2(n_1_1_473), 
      .ZN(n_1_1_795));
   INV_X1 i_1_1_1202 (.A(n_1_1_797), .ZN(n_1_1_796));
   AOI221_X1 i_1_1_1203 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[57]), .C1(
      RAM_Data_RD_A[57]), .C2(n_1_1_477), .ZN(n_1_1_797));
   INV_X1 i_1_1_1204 (.A(n_1_1_798), .ZN(n_302));
   NAND2_X1 i_1_1_1205 (.A1(n_1_1_830), .A2(n_1_1_799), .ZN(n_1_1_798));
   OAI21_X1 i_1_1_1206 (.A(n_1_1_800), .B1(n_1_1_825), .B2(n_1_1_802), .ZN(
      n_1_1_799));
   OAI21_X1 i_1_1_1207 (.A(RAM_Data_RD_B[58]), .B1(n_1_1_801), .B2(n_1_1_473), 
      .ZN(n_1_1_800));
   INV_X1 i_1_1_1208 (.A(n_1_1_802), .ZN(n_1_1_801));
   AOI221_X1 i_1_1_1209 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[58]), .C1(
      RAM_Data_RD_A[58]), .C2(n_1_1_477), .ZN(n_1_1_802));
   INV_X1 i_1_1_1210 (.A(n_1_1_803), .ZN(n_303));
   NAND2_X1 i_1_1_1211 (.A1(n_1_1_830), .A2(n_1_1_804), .ZN(n_1_1_803));
   OAI21_X1 i_1_1_1212 (.A(n_1_1_805), .B1(n_1_1_825), .B2(n_1_1_807), .ZN(
      n_1_1_804));
   OAI21_X1 i_1_1_1213 (.A(RAM_Data_RD_B[59]), .B1(n_1_1_806), .B2(n_1_1_473), 
      .ZN(n_1_1_805));
   INV_X1 i_1_1_1214 (.A(n_1_1_807), .ZN(n_1_1_806));
   AOI221_X1 i_1_1_1215 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[59]), .C1(
      RAM_Data_RD_A[59]), .C2(n_1_1_477), .ZN(n_1_1_807));
   INV_X1 i_1_1_1216 (.A(n_1_1_808), .ZN(n_304));
   NAND2_X1 i_1_1_1217 (.A1(n_1_1_830), .A2(n_1_1_809), .ZN(n_1_1_808));
   OAI21_X1 i_1_1_1218 (.A(n_1_1_810), .B1(n_1_1_825), .B2(n_1_1_812), .ZN(
      n_1_1_809));
   OAI21_X1 i_1_1_1219 (.A(RAM_Data_RD_B[60]), .B1(n_1_1_811), .B2(n_1_1_473), 
      .ZN(n_1_1_810));
   INV_X1 i_1_1_1220 (.A(n_1_1_812), .ZN(n_1_1_811));
   AOI221_X1 i_1_1_1221 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[60]), .C1(
      RAM_Data_RD_A[60]), .C2(n_1_1_477), .ZN(n_1_1_812));
   INV_X1 i_1_1_1222 (.A(n_1_1_813), .ZN(n_305));
   NAND2_X1 i_1_1_1223 (.A1(n_1_1_830), .A2(n_1_1_814), .ZN(n_1_1_813));
   OAI21_X1 i_1_1_1224 (.A(n_1_1_815), .B1(n_1_1_825), .B2(n_1_1_817), .ZN(
      n_1_1_814));
   OAI21_X1 i_1_1_1225 (.A(RAM_Data_RD_B[61]), .B1(n_1_1_816), .B2(n_1_1_473), 
      .ZN(n_1_1_815));
   INV_X1 i_1_1_1226 (.A(n_1_1_817), .ZN(n_1_1_816));
   AOI221_X1 i_1_1_1227 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[61]), .C1(
      RAM_Data_RD_A[61]), .C2(n_1_1_477), .ZN(n_1_1_817));
   INV_X1 i_1_1_1228 (.A(n_1_1_818), .ZN(n_306));
   NAND2_X1 i_1_1_1229 (.A1(n_1_1_830), .A2(n_1_1_819), .ZN(n_1_1_818));
   OAI21_X1 i_1_1_1230 (.A(n_1_1_820), .B1(n_1_1_825), .B2(n_1_1_822), .ZN(
      n_1_1_819));
   OAI21_X1 i_1_1_1231 (.A(RAM_Data_RD_B[62]), .B1(n_1_1_821), .B2(n_1_1_473), 
      .ZN(n_1_1_820));
   INV_X1 i_1_1_1232 (.A(n_1_1_822), .ZN(n_1_1_821));
   AOI221_X1 i_1_1_1233 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[62]), .C1(
      RAM_Data_RD_A[62]), .C2(n_1_1_477), .ZN(n_1_1_822));
   INV_X1 i_1_1_1234 (.A(n_1_1_823), .ZN(n_307));
   NAND2_X1 i_1_1_1235 (.A1(n_1_1_830), .A2(n_1_1_824), .ZN(n_1_1_823));
   OAI21_X1 i_1_1_1236 (.A(n_1_1_826), .B1(n_1_1_828), .B2(n_1_1_825), .ZN(
      n_1_1_824));
   INV_X1 i_1_1_1237 (.A(n_1_1_452), .ZN(n_1_1_825));
   NOR2_X1 i_1_1_1238 (.A1(n_1_1_589), .A2(n_1_1_534), .ZN(n_1_1_452));
   OAI21_X1 i_1_1_1239 (.A(RAM_Data_RD_B[63]), .B1(n_1_1_827), .B2(n_1_1_473), 
      .ZN(n_1_1_826));
   INV_X1 i_1_1_1240 (.A(n_1_1_828), .ZN(n_1_1_827));
   AOI221_X1 i_1_1_1241 (.A(n_1_1_829), .B1(n_1_5), .B2(htemp[63]), .C1(
      RAM_Data_RD_A[63]), .C2(n_1_1_477), .ZN(n_1_1_828));
   INV_X1 i_1_1_1242 (.A(n_1_1_460), .ZN(n_1_1_829));
   NAND2_X1 i_1_1_1243 (.A1(n_1_1_582), .A2(n_1_1_605), .ZN(n_1_1_460));
   NAND2_X1 i_1_1_1244 (.A1(n_1_1_545), .A2(n_1_1_451), .ZN(n_1_1_830));
   NAND2_X1 i_1_1_1245 (.A1(n_1_1_535), .A2(n_1_1_588), .ZN(n_1_1_451));
   NOR2_X1 i_1_1_1246 (.A1(n_1_1_608), .A2(NextState[3]), .ZN(n_1_1_535));
   INV_X1 i_1_1_1247 (.A(n_1_1_846), .ZN(n_1_1_545));
   OAI21_X1 i_1_1_1248 (.A(n_1_1_835), .B1(n_1_1_831), .B2(n_1_1_581), .ZN(n_308));
   INV_X1 i_1_1_1249 (.A(n_1_1_832), .ZN(n_1_1_831));
   OAI22_X1 i_1_1_1250 (.A1(n_1_1_833), .A2(n_1_1_544), .B1(n_1_1_846), .B2(
      n_1_1_839), .ZN(n_1_1_832));
   NAND2_X1 i_1_1_1251 (.A1(n_1_1_846), .A2(n_1_1_834), .ZN(n_1_1_833));
   INV_X1 i_1_1_1252 (.A(adder_out1[12]), .ZN(n_1_1_834));
   INV_X1 i_1_1_1253 (.A(n_1_1_843), .ZN(n_1_1_544));
   OR2_X1 i_1_1_1254 (.A1(n_310), .A2(n_1_1_482), .ZN(n_309));
   NOR2_X1 i_1_1_1255 (.A1(n_1_1_532), .A2(n_1_1_483), .ZN(n_1_1_482));
   NAND2_X1 i_1_1_1256 (.A1(n_1_1_837), .A2(n_1_1_835), .ZN(n_310));
   INV_X1 i_1_1_1257 (.A(n_1_1_836), .ZN(n_1_1_835));
   OAI211_X1 i_1_1_1258 (.A(n_1_1_485), .B(n_1_1_605), .C1(n_1_1_607), .C2(
      n_1_1_534), .ZN(n_1_1_836));
   INV_X1 i_1_1_1259 (.A(RST), .ZN(n_1_1_605));
   INV_X1 i_1_1_1260 (.A(n_1_1_838), .ZN(n_1_1_837));
   OAI21_X1 i_1_1_1261 (.A(n_1_1_840), .B1(n_1_1_581), .B2(n_1_1_839), .ZN(
      n_1_1_838));
   NAND2_X1 i_1_1_1262 (.A1(n_1_1_540), .A2(division_operation), .ZN(n_1_1_839));
   INV_X1 i_1_1_1263 (.A(n_1_1_541), .ZN(n_1_1_540));
   NAND2_X1 i_1_1_1264 (.A1(n_312), .A2(n_311), .ZN(n_1_1_541));
   NAND2_X1 i_1_1_1265 (.A1(n_1_1_584), .A2(n_1_1_594), .ZN(n_1_1_581));
   NAND3_X1 i_1_1_1266 (.A1(n_1_1_846), .A2(n_1_1_843), .A3(n_1_1_582), .ZN(
      n_1_1_840));
   INV_X1 i_1_1_1267 (.A(n_1_1_841), .ZN(n_1_1_582));
   NAND2_X1 i_1_1_1268 (.A1(n_1_1_594), .A2(n_1_1_842), .ZN(n_1_1_841));
   NOR2_X1 i_1_1_1269 (.A1(n_1_1_609), .A2(NextState[2]), .ZN(n_1_1_594));
   INV_X1 i_1_1_1270 (.A(n_1_1_583), .ZN(n_1_1_842));
   NAND2_X1 i_1_1_1271 (.A1(NextState[0]), .A2(NextState[1]), .ZN(n_1_1_583));
   NAND2_X1 i_1_1_1272 (.A1(n_1_1_845), .A2(n_1_1_844), .ZN(n_1_1_843));
   INV_X1 i_1_1_1273 (.A(n_311), .ZN(n_1_1_844));
   INV_X1 i_1_1_1274 (.A(n_312), .ZN(n_1_1_845));
   NAND2_X1 i_1_1_1275 (.A1(n_1_1_848), .A2(n_1_1_847), .ZN(n_1_1_846));
   INV_X1 i_1_1_1276 (.A(n_1_1_546), .ZN(n_1_1_847));
   NAND3_X1 i_1_1_1277 (.A1(n_1_1_547), .A2(n_1_1_560), .A3(n_1_1_558), .ZN(
      n_1_1_546));
   INV_X1 i_1_1_1278 (.A(n_1_1_563), .ZN(n_1_1_848));
   NOR2_X1 i_1_1_1279 (.A1(n_1_1_850), .A2(n_1_1_849), .ZN(n_1_1_563));
   NOR2_X1 i_1_1_1280 (.A1(RAM_Data_RD_A[15]), .A2(n_1_1_625), .ZN(n_1_1_849));
   INV_X1 i_1_1_1281 (.A(Errortemp[15]), .ZN(n_1_1_625));
   AOI21_X1 i_1_1_1282 (.A(n_1_1_851), .B1(n_1_1_853), .B2(n_1_1_852), .ZN(
      n_1_1_850));
   OAI22_X1 i_1_1_1283 (.A1(n_1_1_641), .A2(Errortemp[15]), .B1(n_1_1_640), 
      .B2(Errortemp[14]), .ZN(n_1_1_851));
   INV_X1 i_1_1_1284 (.A(RAM_Data_RD_A[15]), .ZN(n_1_1_641));
   AOI22_X1 i_1_1_1285 (.A1(n_1_1_640), .A2(Errortemp[14]), .B1(n_1_1_639), 
      .B2(Errortemp[13]), .ZN(n_1_1_852));
   INV_X1 i_1_1_1286 (.A(RAM_Data_RD_A[14]), .ZN(n_1_1_640));
   OAI22_X1 i_1_1_1287 (.A1(n_1_1_855), .A2(n_1_1_854), .B1(n_1_1_639), .B2(
      Errortemp[13]), .ZN(n_1_1_853));
   NOR2_X1 i_1_1_1288 (.A1(RAM_Data_RD_A[12]), .A2(n_1_1_622), .ZN(n_1_1_854));
   INV_X1 i_1_1_1289 (.A(Errortemp[12]), .ZN(n_1_1_622));
   AOI21_X1 i_1_1_1290 (.A(n_1_1_856), .B1(n_1_1_858), .B2(n_1_1_857), .ZN(
      n_1_1_855));
   OAI22_X1 i_1_1_1291 (.A1(n_1_1_638), .A2(Errortemp[12]), .B1(n_1_1_637), 
      .B2(Errortemp[11]), .ZN(n_1_1_856));
   INV_X1 i_1_1_1292 (.A(RAM_Data_RD_A[12]), .ZN(n_1_1_638));
   AOI22_X1 i_1_1_1293 (.A1(n_1_1_637), .A2(Errortemp[11]), .B1(n_1_1_636), 
      .B2(Errortemp[10]), .ZN(n_1_1_857));
   INV_X1 i_1_1_1294 (.A(RAM_Data_RD_A[11]), .ZN(n_1_1_637));
   OAI221_X1 i_1_1_1295 (.A(n_1_1_859), .B1(n_1_1_636), .B2(Errortemp[10]), 
      .C1(n_1_1_861), .C2(n_1_1_860), .ZN(n_1_1_858));
   NAND2_X1 i_1_1_1296 (.A1(RAM_Data_RD_A[9]), .A2(n_1_1_619), .ZN(n_1_1_859));
   OAI22_X1 i_1_1_1297 (.A1(RAM_Data_RD_A[9]), .A2(n_1_1_619), .B1(
      RAM_Data_RD_A[8]), .B2(n_1_1_618), .ZN(n_1_1_860));
   INV_X1 i_1_1_1298 (.A(Errortemp[8]), .ZN(n_1_1_618));
   INV_X1 i_1_1_1299 (.A(Errortemp[9]), .ZN(n_1_1_619));
   AOI21_X1 i_1_1_1300 (.A(n_1_1_862), .B1(n_1_1_864), .B2(n_1_1_863), .ZN(
      n_1_1_861));
   OAI22_X1 i_1_1_1301 (.A1(n_1_1_634), .A2(Errortemp[8]), .B1(n_1_1_633), 
      .B2(Errortemp[7]), .ZN(n_1_1_862));
   INV_X1 i_1_1_1302 (.A(RAM_Data_RD_A[8]), .ZN(n_1_1_634));
   AOI22_X1 i_1_1_1303 (.A1(n_1_1_633), .A2(Errortemp[7]), .B1(n_1_1_632), 
      .B2(Errortemp[6]), .ZN(n_1_1_863));
   INV_X1 i_1_1_1304 (.A(RAM_Data_RD_A[7]), .ZN(n_1_1_633));
   OAI221_X1 i_1_1_1305 (.A(n_1_1_865), .B1(n_1_1_632), .B2(Errortemp[6]), 
      .C1(n_1_1_867), .C2(n_1_1_866), .ZN(n_1_1_864));
   NAND2_X1 i_1_1_1306 (.A1(RAM_Data_RD_A[5]), .A2(n_1_1_615), .ZN(n_1_1_865));
   OAI22_X1 i_1_1_1307 (.A1(RAM_Data_RD_A[5]), .A2(n_1_1_615), .B1(
      RAM_Data_RD_A[4]), .B2(n_1_1_614), .ZN(n_1_1_866));
   INV_X1 i_1_1_1308 (.A(Errortemp[4]), .ZN(n_1_1_614));
   INV_X1 i_1_1_1309 (.A(Errortemp[5]), .ZN(n_1_1_615));
   AOI21_X1 i_1_1_1310 (.A(n_1_1_868), .B1(n_1_1_870), .B2(n_1_1_869), .ZN(
      n_1_1_867));
   OAI22_X1 i_1_1_1311 (.A1(n_1_1_630), .A2(Errortemp[4]), .B1(n_1_1_629), 
      .B2(Errortemp[3]), .ZN(n_1_1_868));
   INV_X1 i_1_1_1312 (.A(RAM_Data_RD_A[4]), .ZN(n_1_1_630));
   AOI22_X1 i_1_1_1313 (.A1(n_1_1_629), .A2(Errortemp[3]), .B1(n_1_1_628), 
      .B2(Errortemp[2]), .ZN(n_1_1_869));
   INV_X1 i_1_1_1314 (.A(RAM_Data_RD_A[3]), .ZN(n_1_1_629));
   OR2_X1 i_1_1_1315 (.A1(n_1_1_871), .A2(n_1_1_872), .ZN(n_1_1_870));
   OAI22_X1 i_1_1_1316 (.A1(n_1_1_628), .A2(Errortemp[2]), .B1(n_1_1_627), 
      .B2(Errortemp[1]), .ZN(n_1_1_871));
   INV_X1 i_1_1_1317 (.A(RAM_Data_RD_A[2]), .ZN(n_1_1_628));
   AOI22_X1 i_1_1_1318 (.A1(n_1_1_627), .A2(Errortemp[1]), .B1(n_1_1_626), 
      .B2(Errortemp[0]), .ZN(n_1_1_872));
   INV_X1 i_1_1_1319 (.A(RAM_Data_RD_A[0]), .ZN(n_1_1_626));
   INV_X1 i_1_1_1320 (.A(RAM_Data_RD_A[1]), .ZN(n_1_1_627));
   INV_X1 i_1_1_1321 (.A(RAM_Data_RD_A[6]), .ZN(n_1_1_632));
   INV_X1 i_1_1_1322 (.A(RAM_Data_RD_A[10]), .ZN(n_1_1_636));
   INV_X1 i_1_1_1323 (.A(RAM_Data_RD_A[13]), .ZN(n_1_1_639));
   MUX2_X1 i_1_0_0 (.A(hstate[0]), .B(n_1_5), .S(n_1_7), .Z(n_1_81));
   MUX2_X1 i_1_0_1 (.A(hstate[1]), .B(n_1_6), .S(n_1_7), .Z(n_1_10));
   MUX2_X1 division_operation_reg_enable_mux_0 (.A(division_operation), .B(n_1_8), 
      .S(n_1_9), .Z(n_1_82));
   CLKGATETST_X1 clk_gate_htemp_reg (.CK(CLK), .E(n_235), .SE(1'b0), .GCK(n_2_0));
   DFF_X1 \htemp_reg[63]  (.D(n_132), .CK(n_2_0), .Q(htemp[63]), .QN());
   DFF_X1 \htemp_reg[62]  (.D(n_131), .CK(n_2_0), .Q(htemp[62]), .QN());
   DFF_X1 \htemp_reg[61]  (.D(n_130), .CK(n_2_0), .Q(htemp[61]), .QN());
   DFF_X1 \htemp_reg[60]  (.D(n_129), .CK(n_2_0), .Q(htemp[60]), .QN());
   DFF_X1 \htemp_reg[59]  (.D(n_128), .CK(n_2_0), .Q(htemp[59]), .QN());
   DFF_X1 \htemp_reg[58]  (.D(n_127), .CK(n_2_0), .Q(htemp[58]), .QN());
   DFF_X1 \htemp_reg[57]  (.D(n_126), .CK(n_2_0), .Q(htemp[57]), .QN());
   DFF_X1 \htemp_reg[56]  (.D(n_125), .CK(n_2_0), .Q(htemp[56]), .QN());
   DFF_X1 \htemp_reg[55]  (.D(n_124), .CK(n_2_0), .Q(htemp[55]), .QN());
   DFF_X1 \htemp_reg[54]  (.D(n_123), .CK(n_2_0), .Q(htemp[54]), .QN());
   DFF_X1 \htemp_reg[53]  (.D(n_122), .CK(n_2_0), .Q(htemp[53]), .QN());
   DFF_X1 \htemp_reg[52]  (.D(n_121), .CK(n_2_0), .Q(htemp[52]), .QN());
   DFF_X1 \htemp_reg[51]  (.D(n_120), .CK(n_2_0), .Q(htemp[51]), .QN());
   DFF_X1 \htemp_reg[50]  (.D(n_119), .CK(n_2_0), .Q(htemp[50]), .QN());
   DFF_X1 \htemp_reg[49]  (.D(n_118), .CK(n_2_0), .Q(htemp[49]), .QN());
   DFF_X1 \htemp_reg[48]  (.D(n_117), .CK(n_2_0), .Q(htemp[48]), .QN());
   DFF_X1 \htemp_reg[47]  (.D(n_116), .CK(n_2_0), .Q(htemp[47]), .QN());
   DFF_X1 \htemp_reg[46]  (.D(n_115), .CK(n_2_0), .Q(htemp[46]), .QN());
   DFF_X1 \htemp_reg[45]  (.D(n_114), .CK(n_2_0), .Q(htemp[45]), .QN());
   DFF_X1 \htemp_reg[44]  (.D(n_113), .CK(n_2_0), .Q(htemp[44]), .QN());
   DFF_X1 \htemp_reg[43]  (.D(n_112), .CK(n_2_0), .Q(htemp[43]), .QN());
   DFF_X1 \htemp_reg[42]  (.D(n_111), .CK(n_2_0), .Q(htemp[42]), .QN());
   DFF_X1 \htemp_reg[41]  (.D(n_110), .CK(n_2_0), .Q(htemp[41]), .QN());
   DFF_X1 \htemp_reg[40]  (.D(n_109), .CK(n_2_0), .Q(htemp[40]), .QN());
   DFF_X1 \htemp_reg[39]  (.D(n_108), .CK(n_2_0), .Q(htemp[39]), .QN());
   DFF_X1 \htemp_reg[38]  (.D(n_107), .CK(n_2_0), .Q(htemp[38]), .QN());
   DFF_X1 \htemp_reg[37]  (.D(n_106), .CK(n_2_0), .Q(htemp[37]), .QN());
   DFF_X1 \htemp_reg[36]  (.D(n_105), .CK(n_2_0), .Q(htemp[36]), .QN());
   DFF_X1 \htemp_reg[35]  (.D(n_104), .CK(n_2_0), .Q(htemp[35]), .QN());
   DFF_X1 \htemp_reg[34]  (.D(n_103), .CK(n_2_0), .Q(htemp[34]), .QN());
   DFF_X1 \htemp_reg[33]  (.D(n_102), .CK(n_2_0), .Q(htemp[33]), .QN());
   DFF_X1 \htemp_reg[32]  (.D(n_101), .CK(n_2_0), .Q(htemp[32]), .QN());
   DFF_X1 \htemp_reg[31]  (.D(n_100), .CK(n_2_0), .Q(htemp[31]), .QN());
   DFF_X1 \htemp_reg[30]  (.D(n_99), .CK(n_2_0), .Q(htemp[30]), .QN());
   DFF_X1 \htemp_reg[29]  (.D(n_98), .CK(n_2_0), .Q(htemp[29]), .QN());
   DFF_X1 \htemp_reg[28]  (.D(n_97), .CK(n_2_0), .Q(htemp[28]), .QN());
   DFF_X1 \htemp_reg[27]  (.D(n_96), .CK(n_2_0), .Q(htemp[27]), .QN());
   DFF_X1 \htemp_reg[26]  (.D(n_95), .CK(n_2_0), .Q(htemp[26]), .QN());
   DFF_X1 \htemp_reg[25]  (.D(n_94), .CK(n_2_0), .Q(htemp[25]), .QN());
   DFF_X1 \htemp_reg[24]  (.D(n_93), .CK(n_2_0), .Q(htemp[24]), .QN());
   DFF_X1 \htemp_reg[23]  (.D(n_92), .CK(n_2_0), .Q(htemp[23]), .QN());
   DFF_X1 \htemp_reg[22]  (.D(n_91), .CK(n_2_0), .Q(htemp[22]), .QN());
   DFF_X1 \htemp_reg[21]  (.D(n_90), .CK(n_2_0), .Q(htemp[21]), .QN());
   DFF_X1 \htemp_reg[20]  (.D(n_89), .CK(n_2_0), .Q(htemp[20]), .QN());
   DFF_X1 \htemp_reg[19]  (.D(n_88), .CK(n_2_0), .Q(htemp[19]), .QN());
   DFF_X1 \htemp_reg[18]  (.D(n_87), .CK(n_2_0), .Q(htemp[18]), .QN());
   DFF_X1 \htemp_reg[17]  (.D(n_86), .CK(n_2_0), .Q(htemp[17]), .QN());
   DFF_X1 \htemp_reg[16]  (.D(n_85), .CK(n_2_0), .Q(htemp[16]), .QN());
   CLKGATETST_X1 clk_gate_htemp_reg__47 (.CK(CLK), .E(n_234), .SE(1'b0), 
      .GCK(n_2_1));
   DFF_X1 \htemp_reg[15]  (.D(n_84), .CK(n_2_1), .Q(htemp[15]), .QN());
   DFF_X1 \htemp_reg[14]  (.D(n_83), .CK(n_2_1), .Q(htemp[14]), .QN());
   DFF_X1 \htemp_reg[13]  (.D(n_82), .CK(n_2_1), .Q(htemp[13]), .QN());
   DFF_X1 \htemp_reg[12]  (.D(n_81), .CK(n_2_1), .Q(htemp[12]), .QN());
   DFF_X1 \htemp_reg[11]  (.D(n_80), .CK(n_2_1), .Q(htemp[11]), .QN());
   DFF_X1 \htemp_reg[10]  (.D(n_79), .CK(n_2_1), .Q(htemp[10]), .QN());
   DFF_X1 \htemp_reg[9]  (.D(n_78), .CK(n_2_1), .Q(htemp[9]), .QN());
   DFF_X1 \htemp_reg[8]  (.D(n_77), .CK(n_2_1), .Q(htemp[8]), .QN());
   DFF_X1 \htemp_reg[7]  (.D(n_76), .CK(n_2_1), .Q(htemp[7]), .QN());
   DFF_X1 \htemp_reg[6]  (.D(n_75), .CK(n_2_1), .Q(htemp[6]), .QN());
   DFF_X1 \htemp_reg[5]  (.D(n_74), .CK(n_2_1), .Q(htemp[5]), .QN());
   DFF_X1 \htemp_reg[4]  (.D(n_73), .CK(n_2_1), .Q(htemp[4]), .QN());
   DFF_X1 \htemp_reg[3]  (.D(n_72), .CK(n_2_1), .Q(htemp[3]), .QN());
   DFF_X1 \htemp_reg[2]  (.D(n_71), .CK(n_2_1), .Q(htemp[2]), .QN());
   DFF_X1 \htemp_reg[1]  (.D(n_70), .CK(n_2_1), .Q(htemp[1]), .QN());
   DFF_X1 \htemp_reg[0]  (.D(n_69), .CK(n_2_1), .Q(htemp[0]), .QN());
   CLKGATETST_X1 clk_gate_Temp_reg__47 (.CK(CLK), .E(n_237), .SE(1'b0), .GCK(
      n_2_2));
   DFF_X1 \Temp_reg[15]  (.D(n_18), .CK(n_2_2), .Q(Temp[15]), .QN());
   DFF_X1 \Temp_reg[14]  (.D(n_17), .CK(n_2_2), .Q(Temp[14]), .QN());
   DFF_X1 \Temp_reg[13]  (.D(n_16), .CK(n_2_2), .Q(Temp[13]), .QN());
   DFF_X1 \Temp_reg[12]  (.D(n_15), .CK(n_2_2), .Q(Temp[12]), .QN());
   DFF_X1 \Temp_reg[11]  (.D(n_14), .CK(n_2_2), .Q(Temp[11]), .QN());
   DFF_X1 \Temp_reg[10]  (.D(n_13), .CK(n_2_2), .Q(Temp[10]), .QN());
   DFF_X1 \Temp_reg[9]  (.D(n_12), .CK(n_2_2), .Q(Temp[9]), .QN());
   DFF_X1 \Temp_reg[8]  (.D(n_11), .CK(n_2_2), .Q(Temp[8]), .QN());
   DFF_X1 \Temp_reg[7]  (.D(n_10), .CK(n_2_2), .Q(Temp[7]), .QN());
   DFF_X1 \Temp_reg[6]  (.D(n_9), .CK(n_2_2), .Q(Temp[6]), .QN());
   DFF_X1 \Temp_reg[5]  (.D(n_8), .CK(n_2_2), .Q(Temp[5]), .QN());
   DFF_X1 \Temp_reg[4]  (.D(n_7), .CK(n_2_2), .Q(Temp[4]), .QN());
   DFF_X1 \Temp_reg[3]  (.D(n_6), .CK(n_2_2), .Q(Temp[3]), .QN());
   DFF_X1 \Temp_reg[2]  (.D(n_5), .CK(n_2_2), .Q(Temp[2]), .QN());
   DFF_X1 \Temp_reg[1]  (.D(n_4), .CK(n_2_2), .Q(Temp[1]), .QN());
   DFF_X1 \Temp_reg[0]  (.D(n_3), .CK(n_2_2), .Q(Temp[0]), .QN());
   CLKGATETST_X1 clk_gate_RAM_Address_RD_A_reg (.CK(CLK), .E(n_198), .SE(1'b0), 
      .GCK(n_2_3));
   DFF_X1 \RAM_Address_RD_A_reg[12]  (.D(n_197), .CK(n_2_3), .Q(
      RAM_Address_RD_A[12]), .QN());
   DFF_X1 \RAM_Address_RD_A_reg[11]  (.D(n_196), .CK(n_2_3), .Q(
      RAM_Address_RD_A[11]), .QN());
   DFF_X1 \RAM_Address_RD_A_reg[10]  (.D(n_195), .CK(n_2_3), .Q(
      RAM_Address_RD_A[10]), .QN());
   DFF_X1 \RAM_Address_RD_A_reg[9]  (.D(n_194), .CK(n_2_3), .Q(
      RAM_Address_RD_A[9]), .QN());
   DFF_X1 \RAM_Address_RD_A_reg[8]  (.D(n_193), .CK(n_2_3), .Q(
      RAM_Address_RD_A[8]), .QN());
   DFF_X1 \RAM_Address_RD_A_reg[7]  (.D(n_192), .CK(n_2_3), .Q(
      RAM_Address_RD_A[7]), .QN());
   DFF_X1 \RAM_Address_RD_A_reg[6]  (.D(n_191), .CK(n_2_3), .Q(
      RAM_Address_RD_A[6]), .QN());
   DFF_X1 \RAM_Address_RD_A_reg[5]  (.D(n_190), .CK(n_2_3), .Q(
      RAM_Address_RD_A[5]), .QN());
   DFF_X1 \RAM_Address_RD_A_reg[4]  (.D(n_189), .CK(n_2_3), .Q(
      RAM_Address_RD_A[4]), .QN());
   DFF_X1 \RAM_Address_RD_A_reg[3]  (.D(n_188), .CK(n_2_3), .Q(
      RAM_Address_RD_A[3]), .QN());
   DFF_X1 \RAM_Address_RD_A_reg[2]  (.D(n_187), .CK(n_2_3), .Q(
      RAM_Address_RD_A[2]), .QN());
   DFF_X1 \RAM_Address_RD_A_reg[1]  (.D(n_186), .CK(n_2_3), .Q(
      RAM_Address_RD_A[1]), .QN());
   DFF_X1 \RAM_Address_RD_A_reg[0]  (.D(n_185), .CK(n_2_3), .Q(
      RAM_Address_RD_A[0]), .QN());
   DFF_X1 \in22_reg[15]  (.D(n_165), .CK(n_2_7), .Q(in22[15]), .QN());
   DFF_X1 \in22_reg[14]  (.D(n_164), .CK(n_2_7), .Q(in22[14]), .QN());
   DFF_X1 \in22_reg[13]  (.D(n_163), .CK(n_2_7), .Q(in22[13]), .QN());
   DFF_X1 \in22_reg[12]  (.D(n_162), .CK(n_2_7), .Q(in22[12]), .QN());
   DFF_X1 \in22_reg[11]  (.D(n_161), .CK(n_2_7), .Q(in22[11]), .QN());
   DFF_X1 \in22_reg[10]  (.D(n_160), .CK(n_2_7), .Q(in22[10]), .QN());
   DFF_X1 \in22_reg[9]  (.D(n_159), .CK(n_2_7), .Q(in22[9]), .QN());
   DFF_X1 \in22_reg[8]  (.D(n_158), .CK(n_2_7), .Q(in22[8]), .QN());
   DFF_X1 \in22_reg[7]  (.D(n_157), .CK(n_2_7), .Q(in22[7]), .QN());
   DFF_X1 \in22_reg[6]  (.D(n_156), .CK(n_2_7), .Q(in22[6]), .QN());
   DFF_X1 \in22_reg[5]  (.D(n_155), .CK(n_2_7), .Q(in22[5]), .QN());
   DFF_X1 \in22_reg[4]  (.D(n_154), .CK(n_2_7), .Q(in22[4]), .QN());
   DFF_X1 \in22_reg[3]  (.D(n_153), .CK(n_2_7), .Q(in22[3]), .QN());
   DFF_X1 \in22_reg[2]  (.D(n_152), .CK(n_2_7), .Q(in22[2]), .QN());
   DFF_X1 \in22_reg[1]  (.D(n_151), .CK(n_2_7), .Q(in22[1]), .QN());
   DFF_X1 \in22_reg[0]  (.D(n_150), .CK(n_2_7), .Q(in22[0]), .QN());
   DFF_X1 \in12_reg[15]  (.D(n_53), .CK(n_2_7), .Q(in12[15]), .QN());
   DFF_X1 \in12_reg[14]  (.D(n_52), .CK(n_2_7), .Q(in12[14]), .QN());
   DFF_X1 \in12_reg[13]  (.D(n_51), .CK(n_2_7), .Q(in12[13]), .QN());
   DFF_X1 \in12_reg[12]  (.D(n_50), .CK(n_2_7), .Q(in12[12]), .QN());
   DFF_X1 \in12_reg[11]  (.D(n_49), .CK(n_2_7), .Q(in12[11]), .QN());
   DFF_X1 \in12_reg[10]  (.D(n_48), .CK(n_2_7), .Q(in12[10]), .QN());
   DFF_X1 \in12_reg[9]  (.D(n_47), .CK(n_2_7), .Q(in12[9]), .QN());
   DFF_X1 \in12_reg[8]  (.D(n_46), .CK(n_2_7), .Q(in12[8]), .QN());
   DFF_X1 \in12_reg[7]  (.D(n_45), .CK(n_2_7), .Q(in12[7]), .QN());
   DFF_X1 \in12_reg[6]  (.D(n_44), .CK(n_2_7), .Q(in12[6]), .QN());
   DFF_X1 \in12_reg[5]  (.D(n_43), .CK(n_2_7), .Q(in12[5]), .QN());
   DFF_X1 \in12_reg[4]  (.D(n_42), .CK(n_2_7), .Q(in12[4]), .QN());
   DFF_X1 \in12_reg[3]  (.D(n_41), .CK(n_2_7), .Q(in12[3]), .QN());
   DFF_X1 \in12_reg[2]  (.D(n_40), .CK(n_2_7), .Q(in12[2]), .QN());
   DFF_X1 \in12_reg[1]  (.D(n_39), .CK(n_2_7), .Q(in12[1]), .QN());
   DFF_X1 \in12_reg[0]  (.D(n_38), .CK(n_2_7), .Q(in12[0]), .QN());
   CLKGATETST_X1 clk_gate_divisor_reg (.CK(CLK), .E(n_242), .SE(1'b0), .GCK(
      n_2_4));
   DFF_X1 \divisor_reg[15]  (.D(n_149), .CK(n_2_4), .Q(divisor[15]), .QN());
   DFF_X1 \divisor_reg[14]  (.D(n_148), .CK(n_2_4), .Q(divisor[14]), .QN());
   DFF_X1 \divisor_reg[13]  (.D(n_147), .CK(n_2_4), .Q(divisor[13]), .QN());
   DFF_X1 \divisor_reg[12]  (.D(n_146), .CK(n_2_4), .Q(divisor[12]), .QN());
   DFF_X1 \divisor_reg[11]  (.D(n_145), .CK(n_2_4), .Q(divisor[11]), .QN());
   DFF_X1 \divisor_reg[10]  (.D(n_144), .CK(n_2_4), .Q(divisor[10]), .QN());
   DFF_X1 \divisor_reg[9]  (.D(n_143), .CK(n_2_4), .Q(divisor[9]), .QN());
   DFF_X1 \divisor_reg[8]  (.D(n_142), .CK(n_2_4), .Q(divisor[8]), .QN());
   DFF_X1 \divisor_reg[7]  (.D(n_141), .CK(n_2_4), .Q(divisor[7]), .QN());
   DFF_X1 \divisor_reg[6]  (.D(n_140), .CK(n_2_4), .Q(divisor[6]), .QN());
   DFF_X1 \divisor_reg[5]  (.D(n_139), .CK(n_2_4), .Q(divisor[5]), .QN());
   DFF_X1 \divisor_reg[4]  (.D(n_138), .CK(n_2_4), .Q(divisor[4]), .QN());
   DFF_X1 \divisor_reg[3]  (.D(n_137), .CK(n_2_4), .Q(divisor[3]), .QN());
   DFF_X1 \divisor_reg[2]  (.D(n_136), .CK(n_2_4), .Q(divisor[2]), .QN());
   DFF_X1 \divisor_reg[1]  (.D(n_135), .CK(n_2_4), .Q(divisor[1]), .QN());
   DFF_X1 \divisor_reg[0]  (.D(n_134), .CK(n_2_4), .Q(divisor[0]), .QN());
   CLKGATETST_X1 clk_gate_RAM_Address_RD_B_reg (.CK(CLK), .E(n_212), .SE(1'b0), 
      .GCK(n_2_5));
   DFF_X1 \RAM_Address_RD_B_reg[12]  (.D(n_211), .CK(n_2_5), .Q(
      RAM_Address_RD_B[12]), .QN());
   DFF_X1 \RAM_Address_RD_B_reg[11]  (.D(n_210), .CK(n_2_5), .Q(
      RAM_Address_RD_B[11]), .QN());
   DFF_X1 \RAM_Address_RD_B_reg[10]  (.D(n_209), .CK(n_2_5), .Q(
      RAM_Address_RD_B[10]), .QN());
   DFF_X1 \RAM_Address_RD_B_reg[9]  (.D(n_208), .CK(n_2_5), .Q(
      RAM_Address_RD_B[9]), .QN());
   DFF_X1 \RAM_Address_RD_B_reg[8]  (.D(n_207), .CK(n_2_5), .Q(
      RAM_Address_RD_B[8]), .QN());
   DFF_X1 \RAM_Address_RD_B_reg[7]  (.D(n_206), .CK(n_2_5), .Q(
      RAM_Address_RD_B[7]), .QN());
   DFF_X1 \RAM_Address_RD_B_reg[6]  (.D(n_205), .CK(n_2_5), .Q(
      RAM_Address_RD_B[6]), .QN());
   DFF_X1 \RAM_Address_RD_B_reg[5]  (.D(n_204), .CK(n_2_5), .Q(
      RAM_Address_RD_B[5]), .QN());
   DFF_X1 \RAM_Address_RD_B_reg[4]  (.D(n_203), .CK(n_2_5), .Q(
      RAM_Address_RD_B[4]), .QN());
   DFF_X1 \RAM_Address_RD_B_reg[3]  (.D(n_202), .CK(n_2_5), .Q(
      RAM_Address_RD_B[3]), .QN());
   DFF_X1 \RAM_Address_RD_B_reg[2]  (.D(n_201), .CK(n_2_5), .Q(
      RAM_Address_RD_B[2]), .QN());
   DFF_X1 \RAM_Address_RD_B_reg[1]  (.D(n_200), .CK(n_2_5), .Q(
      RAM_Address_RD_B[1]), .QN());
   DFF_X1 \RAM_Address_RD_B_reg[0]  (.D(n_199), .CK(n_2_5), .Q(
      RAM_Address_RD_B[0]), .QN());
   CLKGATETST_X1 clk_gate_RAM_Address_WR_reg (.CK(CLK), .E(n_309), .SE(1'b0), 
      .GCK(n_2_6));
   DFF_X1 \RAM_Address_WR_reg[12]  (.D(n_227), .CK(n_2_6), .Q(RAM_Address_WR[12]), 
      .QN());
   DFF_X1 \RAM_Address_WR_reg[11]  (.D(n_226), .CK(n_2_6), .Q(RAM_Address_WR[11]), 
      .QN());
   DFF_X1 \RAM_Address_WR_reg[10]  (.D(n_225), .CK(n_2_6), .Q(RAM_Address_WR[10]), 
      .QN());
   DFF_X1 \RAM_Address_WR_reg[9]  (.D(n_224), .CK(n_2_6), .Q(RAM_Address_WR[9]), 
      .QN());
   DFF_X1 \RAM_Address_WR_reg[8]  (.D(n_223), .CK(n_2_6), .Q(RAM_Address_WR[8]), 
      .QN());
   DFF_X1 \RAM_Address_WR_reg[7]  (.D(n_222), .CK(n_2_6), .Q(RAM_Address_WR[7]), 
      .QN());
   DFF_X1 \RAM_Address_WR_reg[6]  (.D(n_221), .CK(n_2_6), .Q(RAM_Address_WR[6]), 
      .QN());
   DFF_X1 \RAM_Address_WR_reg[5]  (.D(n_220), .CK(n_2_6), .Q(RAM_Address_WR[5]), 
      .QN());
   DFF_X1 \RAM_Address_WR_reg[4]  (.D(n_219), .CK(n_2_6), .Q(RAM_Address_WR[4]), 
      .QN());
   DFF_X1 \RAM_Address_WR_reg[3]  (.D(n_218), .CK(n_2_6), .Q(RAM_Address_WR[3]), 
      .QN());
   DFF_X1 \RAM_Address_WR_reg[2]  (.D(n_217), .CK(n_2_6), .Q(RAM_Address_WR[2]), 
      .QN());
   DFF_X1 \RAM_Address_WR_reg[1]  (.D(n_216), .CK(n_2_6), .Q(RAM_Address_WR[1]), 
      .QN());
   DFF_X1 \RAM_Address_WR_reg[0]  (.D(n_215), .CK(n_2_6), .Q(RAM_Address_WR[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_in22_reg (.CK(CLK), .E(n_233), .SE(1'b0), .GCK(n_2_7));
   DFF_X1 mult_enable_reg (.D(n_3_5), .CK(CLK), .Q(mult_enable), .QN());
   DFF_X1 reset_reg (.D(n_3_7), .CK(CLK), .Q(reset), .QN());
   DFF_X1 sub2_reg (.D(n_3_8), .CK(CLK), .Q(sub2), .QN());
   CLKGATETST_X1 clk_gate_NextState_reg (.CK(CLK), .E(n_184), .SE(1'b0), 
      .GCK(n_3_0));
   DFF_X1 \NextState_reg[3]  (.D(n_2), .CK(n_3_0), .Q(NextState[3]), .QN());
   DFF_X1 \NextState_reg[2]  (.D(n_232), .CK(n_3_0), .Q(NextState[2]), .QN());
   DFF_X1 \NextState_reg[1]  (.D(n_238), .CK(n_3_0), .Q(NextState[1]), .QN());
   DFF_X1 \NextState_reg[0]  (.D(n_1), .CK(n_3_0), .Q(NextState[0]), .QN());
   DFF_X1 \flag_reg[0]  (.D(n_3_10), .CK(CLK), .Q(n_311), .QN());
   DFF_X1 \flag_reg[1]  (.D(n_3_9), .CK(CLK), .Q(n_312), .QN());
   DFF_X1 sub1_reg (.D(n_3_11), .CK(CLK), .Q(sub1), .QN());
   CLKGATETST_X1 clk_gate_in21_reg (.CK(CLK), .E(n_236), .SE(1'b0), .GCK(n_3_1));
   DFF_X1 \in21_reg[15]  (.D(n_182), .CK(n_3_1), .Q(in21[15]), .QN());
   DFF_X1 \in21_reg[14]  (.D(n_181), .CK(n_3_1), .Q(in21[14]), .QN());
   DFF_X1 \in21_reg[13]  (.D(n_180), .CK(n_3_1), .Q(in21[13]), .QN());
   DFF_X1 \in21_reg[12]  (.D(n_179), .CK(n_3_1), .Q(in21[12]), .QN());
   DFF_X1 \in21_reg[11]  (.D(n_178), .CK(n_3_1), .Q(in21[11]), .QN());
   DFF_X1 \in21_reg[10]  (.D(n_177), .CK(n_3_1), .Q(in21[10]), .QN());
   DFF_X1 \in21_reg[9]  (.D(n_176), .CK(n_3_1), .Q(in21[9]), .QN());
   DFF_X1 \in21_reg[8]  (.D(n_175), .CK(n_3_1), .Q(in21[8]), .QN());
   DFF_X1 \in21_reg[7]  (.D(n_174), .CK(n_3_1), .Q(in21[7]), .QN());
   DFF_X1 \in21_reg[6]  (.D(n_173), .CK(n_3_1), .Q(in21[6]), .QN());
   DFF_X1 \in21_reg[5]  (.D(n_172), .CK(n_3_1), .Q(in21[5]), .QN());
   DFF_X1 \in21_reg[4]  (.D(n_171), .CK(n_3_1), .Q(in21[4]), .QN());
   DFF_X1 \in21_reg[3]  (.D(n_170), .CK(n_3_1), .Q(in21[3]), .QN());
   DFF_X1 \in21_reg[2]  (.D(n_169), .CK(n_3_1), .Q(in21[2]), .QN());
   DFF_X1 \in21_reg[1]  (.D(n_168), .CK(n_3_1), .Q(in21[1]), .QN());
   DFF_X1 \in21_reg[0]  (.D(n_167), .CK(n_3_1), .Q(in21[0]), .QN());
   DFF_X1 Step_Memory_WR_Enable_reg (.D(n_3_12), .CK(CLK), .Q(
      Step_Memory_WR_Enable), .QN());
   CLKGATETST_X1 clk_gate_count_reg (.CK(CLK), .E(n_67), .SE(1'b0), .GCK(n_3_2));
   DFF_X1 \count_reg[12]  (.D(n_66), .CK(n_3_2), .Q(count[12]), .QN());
   DFF_X1 \count_reg[11]  (.D(n_65), .CK(n_3_2), .Q(count[11]), .QN());
   DFF_X1 \count_reg[10]  (.D(n_64), .CK(n_3_2), .Q(count[10]), .QN());
   DFF_X1 \count_reg[9]  (.D(n_63), .CK(n_3_2), .Q(count[9]), .QN());
   DFF_X1 \count_reg[8]  (.D(n_62), .CK(n_3_2), .Q(count[8]), .QN());
   DFF_X1 \count_reg[7]  (.D(n_61), .CK(n_3_2), .Q(count[7]), .QN());
   DFF_X1 \count_reg[6]  (.D(n_60), .CK(n_3_2), .Q(count[6]), .QN());
   DFF_X1 \count_reg[5]  (.D(n_59), .CK(n_3_2), .Q(count[5]), .QN());
   DFF_X1 \count_reg[4]  (.D(n_58), .CK(n_3_2), .Q(count[4]), .QN());
   DFF_X1 \count_reg[3]  (.D(n_57), .CK(n_3_2), .Q(count[3]), .QN());
   DFF_X1 \count_reg[2]  (.D(n_56), .CK(n_3_2), .Q(count[2]), .QN());
   DFF_X1 \count_reg[1]  (.D(n_55), .CK(n_3_2), .Q(count[1]), .QN());
   DFF_X1 \count_reg[0]  (.D(n_54), .CK(n_3_2), .Q(count[0]), .QN());
   CLKGATETST_X1 clk_gate_RAM_Data_WR_reg (.CK(CLK), .E(n_308), .SE(1'b0), 
      .GCK(n_3_6));
   DFF_X1 \RAM_Data_WR_reg[63]  (.D(n_307), .CK(n_3_6), .Q(RAM_Data_WR[63]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[62]  (.D(n_306), .CK(n_3_6), .Q(RAM_Data_WR[62]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[61]  (.D(n_305), .CK(n_3_6), .Q(RAM_Data_WR[61]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[60]  (.D(n_304), .CK(n_3_6), .Q(RAM_Data_WR[60]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[59]  (.D(n_303), .CK(n_3_6), .Q(RAM_Data_WR[59]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[58]  (.D(n_302), .CK(n_3_6), .Q(RAM_Data_WR[58]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[57]  (.D(n_301), .CK(n_3_6), .Q(RAM_Data_WR[57]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[56]  (.D(n_300), .CK(n_3_6), .Q(RAM_Data_WR[56]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[55]  (.D(n_299), .CK(n_3_6), .Q(RAM_Data_WR[55]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[54]  (.D(n_298), .CK(n_3_6), .Q(RAM_Data_WR[54]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[53]  (.D(n_297), .CK(n_3_6), .Q(RAM_Data_WR[53]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[52]  (.D(n_296), .CK(n_3_6), .Q(RAM_Data_WR[52]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[51]  (.D(n_295), .CK(n_3_6), .Q(RAM_Data_WR[51]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[50]  (.D(n_294), .CK(n_3_6), .Q(RAM_Data_WR[50]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[49]  (.D(n_293), .CK(n_3_6), .Q(RAM_Data_WR[49]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[48]  (.D(n_292), .CK(n_3_6), .Q(RAM_Data_WR[48]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[47]  (.D(n_291), .CK(n_3_6), .Q(RAM_Data_WR[47]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[46]  (.D(n_290), .CK(n_3_6), .Q(RAM_Data_WR[46]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[45]  (.D(n_289), .CK(n_3_6), .Q(RAM_Data_WR[45]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[44]  (.D(n_288), .CK(n_3_6), .Q(RAM_Data_WR[44]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[43]  (.D(n_287), .CK(n_3_6), .Q(RAM_Data_WR[43]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[42]  (.D(n_286), .CK(n_3_6), .Q(RAM_Data_WR[42]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[41]  (.D(n_285), .CK(n_3_6), .Q(RAM_Data_WR[41]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[40]  (.D(n_284), .CK(n_3_6), .Q(RAM_Data_WR[40]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[39]  (.D(n_283), .CK(n_3_6), .Q(RAM_Data_WR[39]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[38]  (.D(n_282), .CK(n_3_6), .Q(RAM_Data_WR[38]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[37]  (.D(n_281), .CK(n_3_6), .Q(RAM_Data_WR[37]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[36]  (.D(n_280), .CK(n_3_6), .Q(RAM_Data_WR[36]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[35]  (.D(n_279), .CK(n_3_6), .Q(RAM_Data_WR[35]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[34]  (.D(n_278), .CK(n_3_6), .Q(RAM_Data_WR[34]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[33]  (.D(n_277), .CK(n_3_6), .Q(RAM_Data_WR[33]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[32]  (.D(n_276), .CK(n_3_6), .Q(RAM_Data_WR[32]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[31]  (.D(n_275), .CK(n_3_6), .Q(RAM_Data_WR[31]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[30]  (.D(n_274), .CK(n_3_6), .Q(RAM_Data_WR[30]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[29]  (.D(n_273), .CK(n_3_6), .Q(RAM_Data_WR[29]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[28]  (.D(n_272), .CK(n_3_6), .Q(RAM_Data_WR[28]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[27]  (.D(n_271), .CK(n_3_6), .Q(RAM_Data_WR[27]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[26]  (.D(n_270), .CK(n_3_6), .Q(RAM_Data_WR[26]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[25]  (.D(n_269), .CK(n_3_6), .Q(RAM_Data_WR[25]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[24]  (.D(n_268), .CK(n_3_6), .Q(RAM_Data_WR[24]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[23]  (.D(n_267), .CK(n_3_6), .Q(RAM_Data_WR[23]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[22]  (.D(n_266), .CK(n_3_6), .Q(RAM_Data_WR[22]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[21]  (.D(n_265), .CK(n_3_6), .Q(RAM_Data_WR[21]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[20]  (.D(n_264), .CK(n_3_6), .Q(RAM_Data_WR[20]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[19]  (.D(n_263), .CK(n_3_6), .Q(RAM_Data_WR[19]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[18]  (.D(n_262), .CK(n_3_6), .Q(RAM_Data_WR[18]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[17]  (.D(n_261), .CK(n_3_6), .Q(RAM_Data_WR[17]), 
      .QN());
   CLKGATETST_X1 clk_gate_RAM_Data_WR_reg__46 (.CK(CLK), .E(n_310), .SE(1'b0), 
      .GCK(n_3_3));
   DFF_X1 \RAM_Data_WR_reg[16]  (.D(n_214), .CK(n_3_3), .Q(RAM_Data_WR[16]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[15]  (.D(n_213), .CK(n_3_3), .Q(RAM_Data_WR[15]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[14]  (.D(n_260), .CK(n_3_3), .Q(RAM_Data_WR[14]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[13]  (.D(n_259), .CK(n_3_3), .Q(RAM_Data_WR[13]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[12]  (.D(n_258), .CK(n_3_3), .Q(RAM_Data_WR[12]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[11]  (.D(n_257), .CK(n_3_3), .Q(RAM_Data_WR[11]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[10]  (.D(n_256), .CK(n_3_3), .Q(RAM_Data_WR[10]), 
      .QN());
   DFF_X1 \RAM_Data_WR_reg[9]  (.D(n_255), .CK(n_3_3), .Q(RAM_Data_WR[9]), .QN());
   DFF_X1 \RAM_Data_WR_reg[8]  (.D(n_254), .CK(n_3_3), .Q(RAM_Data_WR[8]), .QN());
   DFF_X1 \RAM_Data_WR_reg[7]  (.D(n_253), .CK(n_3_3), .Q(RAM_Data_WR[7]), .QN());
   DFF_X1 \RAM_Data_WR_reg[6]  (.D(n_252), .CK(n_3_3), .Q(RAM_Data_WR[6]), .QN());
   DFF_X1 \RAM_Data_WR_reg[5]  (.D(n_251), .CK(n_3_3), .Q(RAM_Data_WR[5]), .QN());
   DFF_X1 \RAM_Data_WR_reg[4]  (.D(n_250), .CK(n_3_3), .Q(RAM_Data_WR[4]), .QN());
   DFF_X1 \RAM_Data_WR_reg[3]  (.D(n_249), .CK(n_3_3), .Q(RAM_Data_WR[3]), .QN());
   DFF_X1 \RAM_Data_WR_reg[2]  (.D(n_248), .CK(n_3_3), .Q(RAM_Data_WR[2]), .QN());
   DFF_X1 \RAM_Data_WR_reg[1]  (.D(n_247), .CK(n_3_3), .Q(RAM_Data_WR[1]), .QN());
   DFF_X1 \RAM_Data_WR_reg[0]  (.D(n_246), .CK(n_3_3), .Q(RAM_Data_WR[0]), .QN());
   DFF_X1 Euler_Enable_reg (.D(n_3_13), .CK(CLK), .Q(Euler_Enable), .QN());
   CLKGATETST_X1 clk_gate_Errortemp_reg__47 (.CK(CLK), .E(n_166), .SE(1'b0), 
      .GCK(n_3_4));
   DFF_X1 \Errortemp_reg[15]  (.D(n_37), .CK(n_3_4), .Q(Errortemp[15]), .QN());
   DFF_X1 \Errortemp_reg[14]  (.D(n_36), .CK(n_3_4), .Q(Errortemp[14]), .QN());
   DFF_X1 \Errortemp_reg[13]  (.D(n_35), .CK(n_3_4), .Q(Errortemp[13]), .QN());
   DFF_X1 \Errortemp_reg[12]  (.D(n_34), .CK(n_3_4), .Q(Errortemp[12]), .QN());
   DFF_X1 \Errortemp_reg[11]  (.D(n_33), .CK(n_3_4), .Q(Errortemp[11]), .QN());
   DFF_X1 \Errortemp_reg[10]  (.D(n_32), .CK(n_3_4), .Q(Errortemp[10]), .QN());
   DFF_X1 \Errortemp_reg[9]  (.D(n_31), .CK(n_3_4), .Q(Errortemp[9]), .QN());
   DFF_X1 \Errortemp_reg[8]  (.D(n_30), .CK(n_3_4), .Q(Errortemp[8]), .QN());
   DFF_X1 \Errortemp_reg[7]  (.D(n_29), .CK(n_3_4), .Q(Errortemp[7]), .QN());
   DFF_X1 \Errortemp_reg[6]  (.D(n_28), .CK(n_3_4), .Q(Errortemp[6]), .QN());
   DFF_X1 \Errortemp_reg[5]  (.D(n_27), .CK(n_3_4), .Q(Errortemp[5]), .QN());
   DFF_X1 \Errortemp_reg[4]  (.D(n_26), .CK(n_3_4), .Q(Errortemp[4]), .QN());
   DFF_X1 \Errortemp_reg[3]  (.D(n_25), .CK(n_3_4), .Q(Errortemp[3]), .QN());
   DFF_X1 \Errortemp_reg[2]  (.D(n_24), .CK(n_3_4), .Q(Errortemp[2]), .QN());
   DFF_X1 \Errortemp_reg[1]  (.D(n_23), .CK(n_3_4), .Q(Errortemp[1]), .QN());
   DFF_X1 \Errortemp_reg[0]  (.D(n_22), .CK(n_3_4), .Q(Errortemp[0]), .QN());
   DFF_X1 Error_Flag_reg (.D(n_3_14), .CK(CLK), .Q(Error_Flag), .QN());
   MUX2_X1 mult_enable_reg_enable_mux_0 (.A(mult_enable), .B(n_133), .S(n_241), 
      .Z(n_3_5));
   NAND2_X1 reset_reg_enable_mux_0 (.A1(reset_reg_enable_mux_n_1), .A2(
      reset_reg_enable_mux_n_0), .ZN(n_3_7));
   NAND2_X1 reset_reg_enable_mux_1 (.A1(n_240), .A2(n_68), .ZN(
      reset_reg_enable_mux_n_0));
   NAND2_X1 reset_reg_enable_mux_2 (.A1(reset_reg_enable_mux_n_2), .A2(reset), 
      .ZN(reset_reg_enable_mux_n_1));
   INV_X1 reset_reg_enable_mux_3 (.A(n_240), .ZN(reset_reg_enable_mux_n_2));
   MUX2_X1 sub2_reg_enable_mux_0 (.A(sub2), .B(n_183), .S(n_239), .Z(n_3_8));
   MUX2_X1 i_3_0_0 (.A(n_311), .B(n_20), .S(n_243), .Z(n_3_10));
   MUX2_X1 i_3_0_1 (.A(n_312), .B(n_21), .S(n_243), .Z(n_3_9));
   MUX2_X1 sub1_reg_enable_mux_0 (.A(sub1), .B(n_19), .S(n_244), .Z(n_3_11));
   MUX2_X1 Step_Memory_WR_Enable_reg_enable_mux_0 (.A(Step_Memory_WR_Enable), 
      .B(n_0), .S(n_245), .Z(n_3_12));
   MUX2_X1 Euler_Enable_reg_enable_mux_0 (.A(Euler_Enable), .B(n_228), .S(n_229), 
      .Z(n_3_13));
   MUX2_X1 Error_Flag_reg_enable_mux_0 (.A(Error_Flag), .B(n_230), .S(n_231), 
      .Z(n_3_14));
   add_sub_cla__4_802 adder1 (.sub(sub1), .in1(in11), .in2(in21), .cin(), 
      .out(adder_out1), .cout(), .invalid(invalid1));
   add_sub_cla adder2 (.sub(sub2), .in1(in12), .in2(in22), .cin(), .out(
      adder_out2), .cout(), .invalid(invalid2));
   Division_CSA Division (.reset(reset), .clk(CLK), .dividend(dividend), 
      .divisor(divisor), .Q({uc_0, Q[14], uc_1, Q[12], Q[11], Q[10], Q[9], Q[8], 
      Q[7], Q[6], Q[5], Q[4], Q[3], Q[2], Q[1], Q[0]}), .ready(ready), .overFlow(
      div_overflow), .divideByZero(divideByZero));
   multiplier_16bit multiplier (.first_operand(first_operand), .second_operand(
      second_operand), .out(out), .enable(mult_enable), .overflow(mult_overflow));
   NOR2_X1 i_0_0_0 (.A1(n_311), .A2(n_312), .ZN(n_313));
   INV_X1 i_0_0_1 (.A(n_311), .ZN(n_0_0_0));
   AND2_X1 i_0_0_2 (.A1(n_0_0_0), .A2(n_312), .ZN(n_314));
   NOR2_X1 i_0_0_3 (.A1(n_0_0_0), .A2(n_312), .ZN(n_315));
endmodule
