/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 16:31:18 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3549782253 */

module datapath__0_28(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_0 (.A(B[0]), .B(p_0[0]), .CO(n_0), .S(p_1[0]));
   FA_X1 i_1 (.A(B[1]), .B(p_0[1]), .CI(n_0), .CO(n_1), .S(p_1[1]));
   FA_X1 i_2 (.A(B[2]), .B(p_0[2]), .CI(n_1), .CO(n_2), .S(p_1[2]));
   FA_X1 i_3 (.A(B[3]), .B(p_0[3]), .CI(n_2), .CO(n_3), .S(p_1[3]));
   FA_X1 i_4 (.A(B[4]), .B(p_0[4]), .CI(n_3), .CO(n_4), .S(p_1[4]));
   FA_X1 i_5 (.A(B[5]), .B(p_0[5]), .CI(n_4), .CO(n_5), .S(p_1[5]));
   FA_X1 i_6 (.A(B[6]), .B(p_0[6]), .CI(n_5), .CO(n_6), .S(p_1[6]));
   FA_X1 i_7 (.A(B[7]), .B(p_0[7]), .CI(n_6), .CO(n_7), .S(p_1[7]));
   FA_X1 i_8 (.A(B[8]), .B(p_0[8]), .CI(n_7), .CO(n_8), .S(p_1[8]));
   FA_X1 i_9 (.A(B[9]), .B(p_0[9]), .CI(n_8), .CO(n_9), .S(p_1[9]));
   FA_X1 i_10 (.A(B[10]), .B(p_0[10]), .CI(n_9), .CO(n_10), .S(p_1[10]));
   FA_X1 i_11 (.A(B[11]), .B(p_0[11]), .CI(n_10), .CO(n_11), .S(p_1[11]));
   FA_X1 i_12 (.A(B[15]), .B(p_0[14]), .CI(n_11), .CO(n_12), .S(p_1[12]));
   FA_X1 i_13 (.A(B[15]), .B(p_0[14]), .CI(n_12), .CO(n_13), .S(p_1[13]));
   FA_X1 i_14 (.A(B[15]), .B(p_0[14]), .CI(n_13), .CO(n_14), .S(p_1[14]));
   XNOR2_X1 i_15 (.A(B[15]), .B(p_0[15]), .ZN(n_15));
   XNOR2_X1 i_16 (.A(n_15), .B(n_14), .ZN(p_1[15]));
endmodule

module datapath__0_33(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[14]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[14]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[14]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[14]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_34(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(p_0[13]), .B2(n_15), .ZN(p_2[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_2[15]));
   NAND2_X1 i_16 (.A1(p_0[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_1[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_1[14]), .ZN(n_16));
endmodule

module datapath__0_39(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[13]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[13]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[13]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_40(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(p_0[13]), .B2(n_15), .ZN(p_2[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_2[15]));
   NAND2_X1 i_16 (.A1(p_0[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_1[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_1[14]), .ZN(n_16));
endmodule

module datapath__0_45(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[12]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[12]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[12]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[12]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_46(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(p_0[13]), .B2(n_15), .ZN(p_2[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_2[15]));
   NAND2_X1 i_16 (.A1(p_0[13]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_1[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_1[14]), .ZN(n_16));
endmodule

module booth_16bit_multiplier(A, B, product);
   input [15:0]A;
   input [15:0]B;
   output [31:0]product;

   wire n_0_174;
   wire n_0_2;
   wire n_0_175;
   wire n_0_3;
   wire n_0_176;
   wire n_0_4;
   wire n_0_177;
   wire n_0_5;
   wire n_0_178;
   wire n_0_6;
   wire n_0_179;
   wire n_0_7;
   wire n_0_180;
   wire n_0_8;
   wire n_0_181;
   wire n_0_9;
   wire n_0_182;
   wire n_0_10;
   wire n_0_183;
   wire n_0_11;
   wire n_0_184;
   wire n_0_12;
   wire n_0_185;
   wire n_0_13;
   wire n_0_186;
   wire n_0_14;
   wire n_0_187;
   wire n_0_0;
   wire n_0_188;
   wire n_0_1;
   wire n_0_189;
   wire n_0_15;
   wire n_0_190;
   wire n_0_16;
   wire n_0_191;
   wire n_0_17;
   wire n_0_192;
   wire n_0_18;
   wire n_0_193;
   wire n_0_19;
   wire n_0_194;
   wire n_0_20;
   wire n_0_195;
   wire n_0_21;
   wire n_0_196;
   wire n_0_22;
   wire n_0_197;
   wire n_0_23;
   wire n_0_198;
   wire n_0_24;
   wire n_0_199;
   wire n_0_25;
   wire n_0_200;
   wire n_0_26;
   wire n_0_201;
   wire n_0_27;
   wire n_0_202;
   wire n_0_28;
   wire n_0_203;
   wire n_0_29;
   wire n_0_204;
   wire n_0_30;
   wire n_0_205;
   wire n_0_31;
   wire n_0_206;
   wire n_0_32;
   wire n_0_207;
   wire n_0_33;
   wire n_0_208;
   wire n_0_34;
   wire n_0_209;
   wire n_0_35;
   wire n_0_210;
   wire n_0_36;
   wire n_0_211;
   wire n_0_37;
   wire n_0_212;
   wire n_0_38;
   wire n_0_213;
   wire n_0_39;
   wire n_0_214;
   wire n_0_40;
   wire n_0_215;
   wire n_0_41;
   wire n_0_216;
   wire n_0_42;
   wire n_0_217;
   wire n_0_43;
   wire n_0_218;
   wire n_0_44;
   wire n_0_219;
   wire n_0_45;
   wire n_0_220;
   wire n_0_46;
   wire n_0_221;
   wire n_0_47;
   wire n_0_222;
   wire n_0_48;
   wire n_0_223;
   wire n_0_49;
   wire n_0_224;
   wire n_0_50;
   wire n_0_225;
   wire n_0_51;
   wire n_0_226;
   wire n_0_52;
   wire n_0_227;
   wire n_0_53;
   wire n_0_228;
   wire n_0_54;
   wire n_0_229;
   wire n_0_55;
   wire n_0_230;
   wire n_0_56;
   wire n_0_231;
   wire n_0_57;
   wire n_0_232;
   wire n_0_58;
   wire n_0_233;
   wire n_0_59;
   wire n_0_234;
   wire n_0_60;
   wire n_0_235;
   wire n_0_61;
   wire n_0_236;
   wire n_0_62;
   wire n_0_237;
   wire n_0_63;
   wire n_0_238;
   wire n_0_64;
   wire n_0_239;
   wire n_0_65;
   wire n_0_240;
   wire n_0_66;
   wire n_0_241;
   wire n_0_67;
   wire n_0_242;
   wire n_0_68;
   wire n_0_243;
   wire n_0_69;
   wire n_0_244;
   wire n_0_70;
   wire n_0_245;
   wire n_0_71;
   wire n_0_246;
   wire n_0_72;
   wire n_0_247;
   wire n_0_73;
   wire n_0_248;
   wire n_0_74;
   wire n_0_249;
   wire n_0_75;
   wire n_0_250;
   wire n_0_76;
   wire n_0_251;
   wire n_0_77;
   wire n_0_252;
   wire n_0_78;
   wire n_0_253;
   wire n_0_79;
   wire n_0_254;
   wire n_0_80;
   wire n_0_255;
   wire n_0_81;
   wire n_0_256;
   wire n_0_82;
   wire n_0_257;
   wire n_0_83;
   wire n_0_258;
   wire n_0_84;
   wire n_0_259;
   wire n_0_85;
   wire n_0_260;
   wire n_0_86;
   wire n_0_261;
   wire n_0_87;
   wire n_0_262;
   wire n_0_88;
   wire n_0_263;
   wire n_0_89;
   wire n_0_264;
   wire n_0_90;
   wire n_0_265;
   wire n_0_91;
   wire n_0_266;
   wire n_0_92;
   wire n_0_267;
   wire n_0_93;
   wire n_0_268;
   wire n_0_94;
   wire n_0_269;
   wire n_0_95;
   wire n_0_270;
   wire n_0_96;
   wire n_0_271;
   wire n_0_97;
   wire n_0_272;
   wire n_0_98;
   wire n_0_273;
   wire n_0_99;
   wire n_0_274;
   wire n_0_100;
   wire n_0_275;
   wire n_0_101;
   wire n_0_276;
   wire n_0_102;
   wire n_0_277;
   wire n_0_103;
   wire n_0_278;
   wire n_0_104;
   wire n_0_279;
   wire n_0_105;
   wire n_0_280;
   wire n_0_106;
   wire n_0_281;
   wire n_0_107;
   wire n_0_282;
   wire n_0_108;
   wire n_0_283;
   wire n_0_109;
   wire n_0_284;
   wire n_0_110;
   wire n_0_285;
   wire n_0_111;
   wire n_0_286;
   wire n_0_112;
   wire n_0_287;
   wire n_0_113;
   wire n_0_288;
   wire n_0_114;
   wire n_0_289;
   wire n_0_115;
   wire n_0_290;
   wire n_0_116;
   wire n_0_291;
   wire n_0_117;
   wire n_0_292;
   wire n_0_118;
   wire n_0_293;
   wire n_0_119;
   wire n_0_294;
   wire n_0_120;
   wire n_0_295;
   wire n_0_121;
   wire n_0_296;
   wire n_0_122;
   wire n_0_297;
   wire n_0_123;
   wire n_0_298;
   wire n_0_124;
   wire n_0_299;
   wire n_0_125;
   wire n_0_300;
   wire n_0_126;
   wire n_0_301;
   wire n_0_127;
   wire n_0_302;
   wire n_0_128;
   wire n_0_303;
   wire n_0_129;
   wire n_0_304;
   wire n_0_130;
   wire n_0_305;
   wire n_0_131;
   wire n_0_306;
   wire n_0_132;
   wire n_0_307;
   wire n_0_133;
   wire n_0_308;
   wire n_0_134;
   wire n_0_309;
   wire n_0_135;
   wire n_0_310;
   wire n_0_136;
   wire n_0_311;
   wire n_0_137;
   wire n_0_312;
   wire n_0_138;
   wire n_0_313;
   wire n_0_139;
   wire n_0_314;
   wire n_0_140;
   wire n_0_315;
   wire n_0_141;
   wire n_0_316;
   wire n_0_142;
   wire n_0_317;
   wire n_0_143;
   wire n_0_318;
   wire n_0_144;
   wire n_0_319;
   wire n_0_145;
   wire n_0_320;
   wire n_0_146;
   wire n_0_321;
   wire n_0_147;
   wire n_0_322;
   wire n_0_148;
   wire n_0_323;
   wire n_0_149;
   wire n_0_324;
   wire n_0_150;
   wire n_0_325;
   wire n_0_151;
   wire n_0_326;
   wire n_0_152;
   wire n_0_327;
   wire n_0_153;
   wire n_0_328;
   wire n_0_154;
   wire n_0_329;
   wire n_0_155;
   wire n_0_330;
   wire n_0_156;
   wire n_0_331;
   wire n_0_157;
   wire n_0_332;
   wire n_0_158;
   wire n_0_333;
   wire n_0_159;
   wire n_0_334;
   wire n_0_160;
   wire n_0_335;
   wire n_0_161;
   wire n_0_336;
   wire n_0_162;
   wire n_0_337;
   wire n_0_163;
   wire n_0_338;
   wire n_0_164;
   wire n_0_339;
   wire n_0_165;
   wire n_0_340;
   wire n_0_166;
   wire n_0_341;
   wire n_0_167;
   wire n_0_342;
   wire n_0_168;
   wire n_0_343;
   wire n_0_169;
   wire n_0_344;
   wire n_0_170;
   wire n_0_345;
   wire n_0_171;
   wire n_0_346;
   wire n_0_172;
   wire n_0_347;
   wire n_0_173;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_0_419;
   wire n_0_420;
   wire n_0_421;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_425;
   wire n_0_426;
   wire n_0_427;
   wire n_0_428;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_436;
   wire n_0_437;
   wire n_0_438;
   wire n_0_439;
   wire n_0_440;
   wire n_0_441;
   wire n_0_442;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_458;
   wire n_0_459;
   wire n_0_460;
   wire n_0_461;
   wire n_0_462;
   wire n_0_463;
   wire n_0_464;
   wire n_0_465;
   wire n_0_466;
   wire n_0_467;
   wire n_0_468;
   wire n_0_469;
   wire n_0_470;
   wire n_0_471;
   wire n_0_472;
   wire n_0_473;
   wire n_0_474;
   wire n_0_475;
   wire n_0_476;
   wire n_0_477;
   wire n_0_478;
   wire n_0_479;
   wire n_0_480;
   wire n_0_481;
   wire n_0_482;
   wire n_0_483;
   wire n_0_484;
   wire n_0_485;
   wire n_0_486;
   wire n_0_487;
   wire n_0_488;
   wire n_0_489;
   wire n_0_490;
   wire n_0_491;
   wire n_0_492;
   wire n_0_493;
   wire n_0_494;
   wire n_0_495;
   wire n_0_496;
   wire n_0_497;
   wire n_0_498;
   wire n_0_499;
   wire n_0_500;
   wire n_0_501;
   wire n_0_502;
   wire n_0_503;
   wire n_0_504;
   wire n_0_505;
   wire n_0_506;
   wire n_0_507;
   wire n_0_508;
   wire n_0_509;
   wire n_0_510;
   wire n_0_511;
   wire n_0_512;
   wire n_0_513;
   wire n_0_514;
   wire n_0_515;
   wire n_0_516;
   wire n_0_517;
   wire n_0_518;
   wire n_0_519;
   wire n_0_520;
   wire n_0_521;
   wire n_0_522;
   wire n_0_523;
   wire n_0_524;
   wire n_0_525;
   wire n_0_526;
   wire n_0_527;
   wire n_0_528;
   wire n_0_529;
   wire n_0_530;
   wire n_0_531;
   wire n_0_532;
   wire n_0_533;
   wire n_0_534;
   wire n_0_535;
   wire n_0_536;
   wire n_0_537;
   wire n_0_538;
   wire n_0_539;
   wire n_0_540;
   wire n_0_541;
   wire n_0_542;
   wire n_0_543;
   wire n_0_544;
   wire n_0_545;
   wire n_0_546;
   wire n_0_547;
   wire n_0_548;
   wire n_0_549;
   wire n_0_550;
   wire n_0_551;
   wire n_0_552;
   wire n_0_553;
   wire n_0_554;
   wire n_0_555;
   wire n_0_556;
   wire n_0_557;
   wire n_0_558;
   wire n_0_559;
   wire n_0_560;
   wire n_0_561;
   wire n_0_562;
   wire n_0_563;
   wire n_0_564;
   wire n_0_565;
   wire n_0_566;
   wire n_0_567;
   wire n_0_568;
   wire n_0_569;
   wire n_0_570;
   wire n_0_571;
   wire n_0_572;
   wire n_0_573;
   wire n_0_574;
   wire n_0_575;
   wire n_0_576;
   wire n_0_577;
   wire n_0_578;
   wire n_0_579;
   wire n_0_580;
   wire n_0_581;
   wire n_0_582;
   wire n_0_583;
   wire n_0_584;
   wire n_0_585;
   wire n_0_586;
   wire n_0_587;
   wire n_0_588;
   wire n_0_589;
   wire n_0_590;
   wire n_0_591;
   wire n_0_592;
   wire n_0_593;
   wire n_0_594;
   wire n_0_595;
   wire n_0_596;
   wire n_0_597;
   wire n_0_598;
   wire n_0_599;
   wire n_0_600;
   wire n_0_601;
   wire n_0_602;
   wire n_0_603;
   wire n_0_604;
   wire n_0_605;
   wire n_0_606;
   wire n_0_607;
   wire n_0_608;
   wire n_0_609;
   wire n_0_610;
   wire n_0_611;
   wire n_0_612;
   wire n_0_613;
   wire n_0_614;
   wire n_0_615;
   wire n_0_616;
   wire n_0_617;
   wire n_0_618;
   wire n_0_619;
   wire n_0_620;
   wire n_0_621;
   wire n_0_622;
   wire n_0_623;
   wire n_0_624;
   wire n_0_625;
   wire n_0_626;
   wire n_0_627;
   wire n_0_628;
   wire n_0_629;
   wire n_0_630;
   wire n_0_631;
   wire n_0_632;
   wire n_0_633;
   wire n_0_634;
   wire n_0_635;
   wire n_0_636;
   wire n_0_637;
   wire n_0_638;
   wire n_0_639;
   wire n_0_640;
   wire n_0_641;
   wire n_0_642;
   wire n_0_643;
   wire n_0_644;
   wire n_0_645;
   wire n_0_646;
   wire n_0_647;
   wire n_0_648;
   wire n_0_649;
   wire n_0_650;
   wire n_0_651;
   wire n_0_652;
   wire n_0_653;
   wire n_0_654;
   wire n_0_655;
   wire n_0_656;
   wire n_0_657;
   wire n_0_658;
   wire n_0_659;
   wire n_0_660;
   wire n_0_661;
   wire n_0_662;
   wire n_0_663;
   wire n_0_664;
   wire n_0_665;
   wire n_0_666;
   wire n_0_667;
   wire n_0_668;
   wire n_0_669;
   wire n_0_670;
   wire n_0_671;
   wire n_0_672;
   wire n_0_673;
   wire n_0_674;
   wire n_0_675;
   wire n_0_676;
   wire n_0_677;
   wire n_0_678;
   wire n_0_679;
   wire n_0_680;
   wire n_0_681;
   wire n_0_682;
   wire n_0_683;
   wire n_0_684;
   wire n_0_685;
   wire n_0_686;
   wire n_0_687;
   wire n_0_688;
   wire n_0_689;

   datapath__0_28 i_2 (.B({B[12], uc_0, uc_1, uc_2, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({n_157, n_170, uc_3, 
      uc_4, n_169, n_168, n_167, n_166, n_165, n_164, n_163, n_162, n_161, n_160, 
      n_159, n_158}), .p_1({n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, 
      n_6, n_5, n_4, n_3, n_2, n_1, n_0}));
   datapath__0_33 i_5 (.B({uc_5, B[12], uc_6, uc_7, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_8, n_156, n_155, 
      n_154, n_153, n_152, n_151, n_150, n_149, n_148, n_147, n_146, n_145, 
      n_144, n_143, n_142}), .p_1({n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
      n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16}));
   datapath__0_34 i_6 (.p_0({uc_9, uc_10, n_170, n_169, n_168, n_167, n_166, 
      n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, B[0]}), .p_1({
      uc_11, n_156, n_155, n_154, n_153, n_152, n_151, n_150, n_149, n_148, 
      n_147, n_146, n_145, n_144, n_143, n_142}), .p_2({n_47, n_46, n_45, n_44, 
      n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32}));
   datapath__0_39 i_9 (.B({uc_12, uc_13, B[12], uc_14, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_15, n_141, 
      n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, n_132, n_131, 
      n_130, n_129, n_128, n_127}), .p_1({n_63, n_62, n_61, n_60, n_59, n_58, 
      n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48}));
   datapath__0_40 i_10 (.p_0({uc_16, uc_17, n_170, n_169, n_168, n_167, n_166, 
      n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, B[0]}), .p_1({
      uc_18, n_141, n_140, n_139, n_138, n_137, n_136, n_135, n_134, n_133, 
      n_132, n_131, n_130, n_129, n_128, n_127}), .p_2({n_79, n_78, n_77, n_76, 
      n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64}));
   datapath__0_45 i_13 (.B({uc_19, uc_20, uc_21, B[12], B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_22, n_126, 
      n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, n_117, n_116, 
      n_115, n_114, n_113, n_112}), .p_1({n_95, n_94, n_93, n_92, n_91, n_90, 
      n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80}));
   datapath__0_46 i_14 (.p_0({uc_23, uc_24, n_170, n_169, n_168, n_167, n_166, 
      n_165, n_164, n_163, n_162, n_161, n_160, n_159, n_158, B[0]}), .p_1({
      uc_25, n_126, n_125, n_124, n_123, n_122, n_121, n_120, n_119, n_118, 
      n_117, n_116, n_115, n_114, n_113, n_112}), .p_2({n_111, n_110, n_109, 
      n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
      n_97, n_96}));
   FA_X1 i_0_0 (.A(B[1]), .B(n_0_355), .CI(n_0_166), .CO(n_0_2), .S(n_0_174));
   FA_X1 i_0_1 (.A(B[2]), .B(n_0_362), .CI(n_0_2), .CO(n_0_3), .S(n_0_175));
   FA_X1 i_0_2 (.A(B[3]), .B(n_0_371), .CI(n_0_3), .CO(n_0_4), .S(n_0_176));
   FA_X1 i_0_3 (.A(B[4]), .B(n_0_382), .CI(n_0_4), .CO(n_0_5), .S(n_0_177));
   FA_X1 i_0_4 (.A(B[5]), .B(n_0_395), .CI(n_0_5), .CO(n_0_6), .S(n_0_178));
   FA_X1 i_0_5 (.A(B[6]), .B(n_0_410), .CI(n_0_6), .CO(n_0_7), .S(n_0_179));
   FA_X1 i_0_6 (.A(B[7]), .B(n_0_427), .CI(n_0_7), .CO(n_0_8), .S(n_0_180));
   FA_X1 i_0_7 (.A(B[8]), .B(n_0_444), .CI(n_0_8), .CO(n_0_9), .S(n_0_181));
   FA_X1 i_0_8 (.A(B[9]), .B(n_0_461), .CI(n_0_9), .CO(n_0_10), .S(n_0_182));
   FA_X1 i_0_9 (.A(B[10]), .B(n_0_478), .CI(n_0_10), .CO(n_0_11), .S(n_0_183));
   FA_X1 i_0_10 (.A(B[11]), .B(n_0_495), .CI(n_0_11), .CO(n_0_12), .S(n_0_184));
   FA_X1 i_0_11 (.A(B[12]), .B(n_0_512), .CI(n_0_12), .CO(n_0_13), .S(n_0_185));
   FA_X1 i_0_12 (.A(B[12]), .B(n_0_529), .CI(n_0_13), .CO(n_0_14), .S(n_0_186));
   FA_X1 i_0_13 (.A(n_158), .B(n_0_355), .CI(n_0_166), .CO(n_0_0), .S(n_0_187));
   FA_X1 i_0_14 (.A(n_159), .B(n_0_362), .CI(n_0_0), .CO(n_0_1), .S(n_0_188));
   FA_X1 i_0_15 (.A(n_160), .B(n_0_371), .CI(n_0_1), .CO(n_0_15), .S(n_0_189));
   FA_X1 i_0_16 (.A(n_161), .B(n_0_382), .CI(n_0_15), .CO(n_0_16), .S(n_0_190));
   FA_X1 i_0_17 (.A(n_162), .B(n_0_395), .CI(n_0_16), .CO(n_0_17), .S(n_0_191));
   FA_X1 i_0_18 (.A(n_163), .B(n_0_410), .CI(n_0_17), .CO(n_0_18), .S(n_0_192));
   FA_X1 i_0_19 (.A(n_164), .B(n_0_427), .CI(n_0_18), .CO(n_0_19), .S(n_0_193));
   FA_X1 i_0_20 (.A(n_165), .B(n_0_444), .CI(n_0_19), .CO(n_0_20), .S(n_0_194));
   FA_X1 i_0_21 (.A(n_166), .B(n_0_461), .CI(n_0_20), .CO(n_0_21), .S(n_0_195));
   FA_X1 i_0_22 (.A(n_167), .B(n_0_478), .CI(n_0_21), .CO(n_0_22), .S(n_0_196));
   FA_X1 i_0_23 (.A(n_168), .B(n_0_495), .CI(n_0_22), .CO(n_0_23), .S(n_0_197));
   FA_X1 i_0_24 (.A(n_169), .B(n_0_512), .CI(n_0_23), .CO(n_0_24), .S(n_0_198));
   FA_X1 i_0_25 (.A(n_170), .B(n_0_529), .CI(n_0_24), .CO(n_0_25), .S(n_0_199));
   FA_X1 i_0_26 (.A(B[1]), .B(n_0_360), .CI(n_0_167), .CO(n_0_26), .S(n_0_200));
   FA_X1 i_0_27 (.A(B[2]), .B(n_0_369), .CI(n_0_26), .CO(n_0_27), .S(n_0_201));
   FA_X1 i_0_28 (.A(B[3]), .B(n_0_380), .CI(n_0_27), .CO(n_0_28), .S(n_0_202));
   FA_X1 i_0_29 (.A(B[4]), .B(n_0_393), .CI(n_0_28), .CO(n_0_29), .S(n_0_203));
   FA_X1 i_0_30 (.A(B[5]), .B(n_0_408), .CI(n_0_29), .CO(n_0_30), .S(n_0_204));
   FA_X1 i_0_31 (.A(B[6]), .B(n_0_425), .CI(n_0_30), .CO(n_0_31), .S(n_0_205));
   FA_X1 i_0_32 (.A(B[7]), .B(n_0_442), .CI(n_0_31), .CO(n_0_32), .S(n_0_206));
   FA_X1 i_0_33 (.A(B[8]), .B(n_0_459), .CI(n_0_32), .CO(n_0_33), .S(n_0_207));
   FA_X1 i_0_34 (.A(B[9]), .B(n_0_476), .CI(n_0_33), .CO(n_0_34), .S(n_0_208));
   FA_X1 i_0_35 (.A(B[10]), .B(n_0_493), .CI(n_0_34), .CO(n_0_35), .S(n_0_209));
   FA_X1 i_0_36 (.A(B[11]), .B(n_0_510), .CI(n_0_35), .CO(n_0_36), .S(n_0_210));
   FA_X1 i_0_37 (.A(B[12]), .B(n_0_527), .CI(n_0_36), .CO(n_0_37), .S(n_0_211));
   FA_X1 i_0_38 (.A(B[12]), .B(n_0_544), .CI(n_0_37), .CO(n_0_38), .S(n_0_212));
   FA_X1 i_0_39 (.A(n_158), .B(n_0_360), .CI(n_0_167), .CO(n_0_39), .S(n_0_213));
   FA_X1 i_0_40 (.A(n_159), .B(n_0_369), .CI(n_0_39), .CO(n_0_40), .S(n_0_214));
   FA_X1 i_0_41 (.A(n_160), .B(n_0_380), .CI(n_0_40), .CO(n_0_41), .S(n_0_215));
   FA_X1 i_0_42 (.A(n_161), .B(n_0_393), .CI(n_0_41), .CO(n_0_42), .S(n_0_216));
   FA_X1 i_0_43 (.A(n_162), .B(n_0_408), .CI(n_0_42), .CO(n_0_43), .S(n_0_217));
   FA_X1 i_0_44 (.A(n_163), .B(n_0_425), .CI(n_0_43), .CO(n_0_44), .S(n_0_218));
   FA_X1 i_0_45 (.A(n_164), .B(n_0_442), .CI(n_0_44), .CO(n_0_45), .S(n_0_219));
   FA_X1 i_0_46 (.A(n_165), .B(n_0_459), .CI(n_0_45), .CO(n_0_46), .S(n_0_220));
   FA_X1 i_0_47 (.A(n_166), .B(n_0_476), .CI(n_0_46), .CO(n_0_47), .S(n_0_221));
   FA_X1 i_0_48 (.A(n_167), .B(n_0_493), .CI(n_0_47), .CO(n_0_48), .S(n_0_222));
   FA_X1 i_0_49 (.A(n_168), .B(n_0_510), .CI(n_0_48), .CO(n_0_49), .S(n_0_223));
   FA_X1 i_0_50 (.A(n_169), .B(n_0_527), .CI(n_0_49), .CO(n_0_50), .S(n_0_224));
   FA_X1 i_0_51 (.A(n_170), .B(n_0_544), .CI(n_0_50), .CO(n_0_51), .S(n_0_225));
   FA_X1 i_0_52 (.A(B[1]), .B(n_0_367), .CI(n_0_168), .CO(n_0_52), .S(n_0_226));
   FA_X1 i_0_53 (.A(B[2]), .B(n_0_378), .CI(n_0_52), .CO(n_0_53), .S(n_0_227));
   FA_X1 i_0_54 (.A(B[3]), .B(n_0_391), .CI(n_0_53), .CO(n_0_54), .S(n_0_228));
   FA_X1 i_0_55 (.A(B[4]), .B(n_0_406), .CI(n_0_54), .CO(n_0_55), .S(n_0_229));
   FA_X1 i_0_56 (.A(B[5]), .B(n_0_423), .CI(n_0_55), .CO(n_0_56), .S(n_0_230));
   FA_X1 i_0_57 (.A(B[6]), .B(n_0_440), .CI(n_0_56), .CO(n_0_57), .S(n_0_231));
   FA_X1 i_0_58 (.A(B[7]), .B(n_0_457), .CI(n_0_57), .CO(n_0_58), .S(n_0_232));
   FA_X1 i_0_59 (.A(B[8]), .B(n_0_474), .CI(n_0_58), .CO(n_0_59), .S(n_0_233));
   FA_X1 i_0_60 (.A(B[9]), .B(n_0_491), .CI(n_0_59), .CO(n_0_60), .S(n_0_234));
   FA_X1 i_0_61 (.A(B[10]), .B(n_0_508), .CI(n_0_60), .CO(n_0_61), .S(n_0_235));
   FA_X1 i_0_62 (.A(B[11]), .B(n_0_525), .CI(n_0_61), .CO(n_0_62), .S(n_0_236));
   FA_X1 i_0_63 (.A(B[12]), .B(n_0_542), .CI(n_0_62), .CO(n_0_63), .S(n_0_237));
   FA_X1 i_0_64 (.A(n_158), .B(n_0_367), .CI(n_0_168), .CO(n_0_64), .S(n_0_238));
   FA_X1 i_0_65 (.A(n_159), .B(n_0_378), .CI(n_0_64), .CO(n_0_65), .S(n_0_239));
   FA_X1 i_0_66 (.A(n_160), .B(n_0_391), .CI(n_0_65), .CO(n_0_66), .S(n_0_240));
   FA_X1 i_0_67 (.A(n_161), .B(n_0_406), .CI(n_0_66), .CO(n_0_67), .S(n_0_241));
   FA_X1 i_0_68 (.A(n_162), .B(n_0_423), .CI(n_0_67), .CO(n_0_68), .S(n_0_242));
   FA_X1 i_0_69 (.A(n_163), .B(n_0_440), .CI(n_0_68), .CO(n_0_69), .S(n_0_243));
   FA_X1 i_0_70 (.A(n_164), .B(n_0_457), .CI(n_0_69), .CO(n_0_70), .S(n_0_244));
   FA_X1 i_0_71 (.A(n_165), .B(n_0_474), .CI(n_0_70), .CO(n_0_71), .S(n_0_245));
   FA_X1 i_0_72 (.A(n_166), .B(n_0_491), .CI(n_0_71), .CO(n_0_72), .S(n_0_246));
   FA_X1 i_0_73 (.A(n_167), .B(n_0_508), .CI(n_0_72), .CO(n_0_73), .S(n_0_247));
   FA_X1 i_0_74 (.A(n_168), .B(n_0_525), .CI(n_0_73), .CO(n_0_74), .S(n_0_248));
   FA_X1 i_0_75 (.A(n_169), .B(n_0_542), .CI(n_0_74), .CO(n_0_75), .S(n_0_249));
   FA_X1 i_0_76 (.A(B[1]), .B(n_0_376), .CI(n_0_169), .CO(n_0_76), .S(n_0_250));
   FA_X1 i_0_77 (.A(B[2]), .B(n_0_389), .CI(n_0_76), .CO(n_0_77), .S(n_0_251));
   FA_X1 i_0_78 (.A(B[3]), .B(n_0_404), .CI(n_0_77), .CO(n_0_78), .S(n_0_252));
   FA_X1 i_0_79 (.A(B[4]), .B(n_0_421), .CI(n_0_78), .CO(n_0_79), .S(n_0_253));
   FA_X1 i_0_80 (.A(B[5]), .B(n_0_438), .CI(n_0_79), .CO(n_0_80), .S(n_0_254));
   FA_X1 i_0_81 (.A(B[6]), .B(n_0_455), .CI(n_0_80), .CO(n_0_81), .S(n_0_255));
   FA_X1 i_0_82 (.A(B[7]), .B(n_0_472), .CI(n_0_81), .CO(n_0_82), .S(n_0_256));
   FA_X1 i_0_83 (.A(B[8]), .B(n_0_489), .CI(n_0_82), .CO(n_0_83), .S(n_0_257));
   FA_X1 i_0_84 (.A(B[9]), .B(n_0_506), .CI(n_0_83), .CO(n_0_84), .S(n_0_258));
   FA_X1 i_0_85 (.A(B[10]), .B(n_0_523), .CI(n_0_84), .CO(n_0_85), .S(n_0_259));
   FA_X1 i_0_86 (.A(B[11]), .B(n_0_540), .CI(n_0_85), .CO(n_0_86), .S(n_0_260));
   FA_X1 i_0_87 (.A(n_158), .B(n_0_376), .CI(n_0_169), .CO(n_0_87), .S(n_0_261));
   FA_X1 i_0_88 (.A(n_159), .B(n_0_389), .CI(n_0_87), .CO(n_0_88), .S(n_0_262));
   FA_X1 i_0_89 (.A(n_160), .B(n_0_404), .CI(n_0_88), .CO(n_0_89), .S(n_0_263));
   FA_X1 i_0_90 (.A(n_161), .B(n_0_421), .CI(n_0_89), .CO(n_0_90), .S(n_0_264));
   FA_X1 i_0_91 (.A(n_162), .B(n_0_438), .CI(n_0_90), .CO(n_0_91), .S(n_0_265));
   FA_X1 i_0_92 (.A(n_163), .B(n_0_455), .CI(n_0_91), .CO(n_0_92), .S(n_0_266));
   FA_X1 i_0_93 (.A(n_164), .B(n_0_472), .CI(n_0_92), .CO(n_0_93), .S(n_0_267));
   FA_X1 i_0_94 (.A(n_165), .B(n_0_489), .CI(n_0_93), .CO(n_0_94), .S(n_0_268));
   FA_X1 i_0_95 (.A(n_166), .B(n_0_506), .CI(n_0_94), .CO(n_0_95), .S(n_0_269));
   FA_X1 i_0_96 (.A(n_167), .B(n_0_523), .CI(n_0_95), .CO(n_0_96), .S(n_0_270));
   FA_X1 i_0_97 (.A(n_168), .B(n_0_540), .CI(n_0_96), .CO(n_0_97), .S(n_0_271));
   FA_X1 i_0_98 (.A(B[1]), .B(n_0_387), .CI(n_0_170), .CO(n_0_98), .S(n_0_272));
   FA_X1 i_0_99 (.A(B[2]), .B(n_0_402), .CI(n_0_98), .CO(n_0_99), .S(n_0_273));
   FA_X1 i_0_100 (.A(B[3]), .B(n_0_419), .CI(n_0_99), .CO(n_0_100), .S(n_0_274));
   FA_X1 i_0_101 (.A(B[4]), .B(n_0_436), .CI(n_0_100), .CO(n_0_101), .S(n_0_275));
   FA_X1 i_0_102 (.A(B[5]), .B(n_0_453), .CI(n_0_101), .CO(n_0_102), .S(n_0_276));
   FA_X1 i_0_103 (.A(B[6]), .B(n_0_470), .CI(n_0_102), .CO(n_0_103), .S(n_0_277));
   FA_X1 i_0_104 (.A(B[7]), .B(n_0_487), .CI(n_0_103), .CO(n_0_104), .S(n_0_278));
   FA_X1 i_0_105 (.A(B[8]), .B(n_0_504), .CI(n_0_104), .CO(n_0_105), .S(n_0_279));
   FA_X1 i_0_106 (.A(B[9]), .B(n_0_521), .CI(n_0_105), .CO(n_0_106), .S(n_0_280));
   FA_X1 i_0_107 (.A(B[10]), .B(n_0_538), .CI(n_0_106), .CO(n_0_107), .S(n_0_281));
   FA_X1 i_0_108 (.A(n_158), .B(n_0_387), .CI(n_0_170), .CO(n_0_108), .S(n_0_282));
   FA_X1 i_0_109 (.A(n_159), .B(n_0_402), .CI(n_0_108), .CO(n_0_109), .S(n_0_283));
   FA_X1 i_0_110 (.A(n_160), .B(n_0_419), .CI(n_0_109), .CO(n_0_110), .S(n_0_284));
   FA_X1 i_0_111 (.A(n_161), .B(n_0_436), .CI(n_0_110), .CO(n_0_111), .S(n_0_285));
   FA_X1 i_0_112 (.A(n_162), .B(n_0_453), .CI(n_0_111), .CO(n_0_112), .S(n_0_286));
   FA_X1 i_0_113 (.A(n_163), .B(n_0_470), .CI(n_0_112), .CO(n_0_113), .S(n_0_287));
   FA_X1 i_0_114 (.A(n_164), .B(n_0_487), .CI(n_0_113), .CO(n_0_114), .S(n_0_288));
   FA_X1 i_0_115 (.A(n_165), .B(n_0_504), .CI(n_0_114), .CO(n_0_115), .S(n_0_289));
   FA_X1 i_0_116 (.A(n_166), .B(n_0_521), .CI(n_0_115), .CO(n_0_116), .S(n_0_290));
   FA_X1 i_0_117 (.A(n_167), .B(n_0_538), .CI(n_0_116), .CO(n_0_117), .S(n_0_291));
   FA_X1 i_0_118 (.A(B[1]), .B(n_0_400), .CI(n_0_171), .CO(n_0_118), .S(n_0_292));
   FA_X1 i_0_119 (.A(B[2]), .B(n_0_417), .CI(n_0_118), .CO(n_0_119), .S(n_0_293));
   FA_X1 i_0_120 (.A(B[3]), .B(n_0_434), .CI(n_0_119), .CO(n_0_120), .S(n_0_294));
   FA_X1 i_0_121 (.A(B[4]), .B(n_0_451), .CI(n_0_120), .CO(n_0_121), .S(n_0_295));
   FA_X1 i_0_122 (.A(B[5]), .B(n_0_468), .CI(n_0_121), .CO(n_0_122), .S(n_0_296));
   FA_X1 i_0_123 (.A(B[6]), .B(n_0_485), .CI(n_0_122), .CO(n_0_123), .S(n_0_297));
   FA_X1 i_0_124 (.A(B[7]), .B(n_0_502), .CI(n_0_123), .CO(n_0_124), .S(n_0_298));
   FA_X1 i_0_125 (.A(B[8]), .B(n_0_519), .CI(n_0_124), .CO(n_0_125), .S(n_0_299));
   FA_X1 i_0_126 (.A(B[9]), .B(n_0_536), .CI(n_0_125), .CO(n_0_126), .S(n_0_300));
   FA_X1 i_0_127 (.A(n_158), .B(n_0_400), .CI(n_0_171), .CO(n_0_127), .S(n_0_301));
   FA_X1 i_0_128 (.A(n_159), .B(n_0_417), .CI(n_0_127), .CO(n_0_128), .S(n_0_302));
   FA_X1 i_0_129 (.A(n_160), .B(n_0_434), .CI(n_0_128), .CO(n_0_129), .S(n_0_303));
   FA_X1 i_0_130 (.A(n_161), .B(n_0_451), .CI(n_0_129), .CO(n_0_130), .S(n_0_304));
   FA_X1 i_0_131 (.A(n_162), .B(n_0_468), .CI(n_0_130), .CO(n_0_131), .S(n_0_305));
   FA_X1 i_0_132 (.A(n_163), .B(n_0_485), .CI(n_0_131), .CO(n_0_132), .S(n_0_306));
   FA_X1 i_0_133 (.A(n_164), .B(n_0_502), .CI(n_0_132), .CO(n_0_133), .S(n_0_307));
   FA_X1 i_0_134 (.A(n_165), .B(n_0_519), .CI(n_0_133), .CO(n_0_134), .S(n_0_308));
   FA_X1 i_0_135 (.A(n_166), .B(n_0_536), .CI(n_0_134), .CO(n_0_135), .S(n_0_309));
   FA_X1 i_0_136 (.A(B[1]), .B(n_0_415), .CI(n_0_172), .CO(n_0_136), .S(n_0_310));
   FA_X1 i_0_137 (.A(B[2]), .B(n_0_432), .CI(n_0_136), .CO(n_0_137), .S(n_0_311));
   FA_X1 i_0_138 (.A(B[3]), .B(n_0_449), .CI(n_0_137), .CO(n_0_138), .S(n_0_312));
   FA_X1 i_0_139 (.A(B[4]), .B(n_0_466), .CI(n_0_138), .CO(n_0_139), .S(n_0_313));
   FA_X1 i_0_140 (.A(B[5]), .B(n_0_483), .CI(n_0_139), .CO(n_0_140), .S(n_0_314));
   FA_X1 i_0_141 (.A(B[6]), .B(n_0_500), .CI(n_0_140), .CO(n_0_141), .S(n_0_315));
   FA_X1 i_0_142 (.A(B[7]), .B(n_0_517), .CI(n_0_141), .CO(n_0_142), .S(n_0_316));
   FA_X1 i_0_143 (.A(B[8]), .B(n_0_534), .CI(n_0_142), .CO(n_0_143), .S(n_0_317));
   FA_X1 i_0_144 (.A(n_158), .B(n_0_415), .CI(n_0_172), .CO(n_0_144), .S(n_0_318));
   FA_X1 i_0_145 (.A(n_159), .B(n_0_432), .CI(n_0_144), .CO(n_0_145), .S(n_0_319));
   FA_X1 i_0_146 (.A(n_160), .B(n_0_449), .CI(n_0_145), .CO(n_0_146), .S(n_0_320));
   FA_X1 i_0_147 (.A(n_161), .B(n_0_466), .CI(n_0_146), .CO(n_0_147), .S(n_0_321));
   FA_X1 i_0_148 (.A(n_162), .B(n_0_483), .CI(n_0_147), .CO(n_0_148), .S(n_0_322));
   FA_X1 i_0_149 (.A(n_163), .B(n_0_500), .CI(n_0_148), .CO(n_0_149), .S(n_0_323));
   FA_X1 i_0_150 (.A(n_164), .B(n_0_517), .CI(n_0_149), .CO(n_0_150), .S(n_0_324));
   FA_X1 i_0_151 (.A(n_165), .B(n_0_534), .CI(n_0_150), .CO(n_0_151), .S(n_0_325));
   FA_X1 i_0_152 (.A(B[1]), .B(n_0_430), .CI(n_0_173), .CO(n_0_152), .S(n_0_326));
   FA_X1 i_0_153 (.A(B[2]), .B(n_0_447), .CI(n_0_152), .CO(n_0_153), .S(n_0_327));
   FA_X1 i_0_154 (.A(B[3]), .B(n_0_464), .CI(n_0_153), .CO(n_0_154), .S(n_0_328));
   FA_X1 i_0_155 (.A(B[4]), .B(n_0_481), .CI(n_0_154), .CO(n_0_155), .S(n_0_329));
   FA_X1 i_0_156 (.A(B[5]), .B(n_0_498), .CI(n_0_155), .CO(n_0_156), .S(n_0_330));
   FA_X1 i_0_157 (.A(B[6]), .B(n_0_515), .CI(n_0_156), .CO(n_0_157), .S(n_0_331));
   FA_X1 i_0_158 (.A(B[7]), .B(n_0_532), .CI(n_0_157), .CO(n_0_158), .S(n_0_332));
   FA_X1 i_0_159 (.A(n_158), .B(n_0_430), .CI(n_0_173), .CO(n_0_159), .S(n_0_333));
   FA_X1 i_0_160 (.A(n_159), .B(n_0_447), .CI(n_0_159), .CO(n_0_160), .S(n_0_334));
   FA_X1 i_0_161 (.A(n_160), .B(n_0_464), .CI(n_0_160), .CO(n_0_161), .S(n_0_335));
   FA_X1 i_0_162 (.A(n_161), .B(n_0_481), .CI(n_0_161), .CO(n_0_162), .S(n_0_336));
   FA_X1 i_0_163 (.A(n_162), .B(n_0_498), .CI(n_0_162), .CO(n_0_163), .S(n_0_337));
   FA_X1 i_0_164 (.A(n_163), .B(n_0_515), .CI(n_0_163), .CO(n_0_164), .S(n_0_338));
   FA_X1 i_0_165 (.A(n_164), .B(n_0_532), .CI(n_0_164), .CO(n_0_165), .S(n_0_339));
   HA_X1 i_0_166 (.A(B[0]), .B(n_0_350), .CO(n_0_166), .S(n_0_340));
   HA_X1 i_0_167 (.A(B[0]), .B(n_0_353), .CO(n_0_167), .S(n_0_341));
   HA_X1 i_0_168 (.A(B[0]), .B(n_0_358), .CO(n_0_168), .S(n_0_342));
   HA_X1 i_0_169 (.A(B[0]), .B(n_0_365), .CO(n_0_169), .S(n_0_343));
   HA_X1 i_0_170 (.A(B[0]), .B(n_0_374), .CO(n_0_170), .S(n_0_344));
   HA_X1 i_0_171 (.A(B[0]), .B(n_0_385), .CO(n_0_171), .S(n_0_345));
   HA_X1 i_0_172 (.A(B[0]), .B(n_0_398), .CO(n_0_172), .S(n_0_346));
   HA_X1 i_0_173 (.A(B[0]), .B(n_0_413), .CO(n_0_173), .S(n_0_347));
   INV_X1 i_0_174 (.A(n_0_348), .ZN(product[4]));
   AOI222_X1 i_0_175 (.A1(n_80), .A2(n_0_556), .B1(n_96), .B2(n_0_557), .C1(
      n_112), .C2(n_0_555), .ZN(n_0_348));
   OAI21_X1 i_0_176 (.A(n_0_349), .B1(n_0_545), .B2(n_0_351), .ZN(product[5]));
   NAND2_X1 i_0_177 (.A1(n_0_340), .A2(n_0_545), .ZN(n_0_349));
   INV_X1 i_0_178 (.A(n_0_351), .ZN(n_0_350));
   AOI222_X1 i_0_179 (.A1(n_81), .A2(n_0_556), .B1(n_97), .B2(n_0_557), .C1(
      n_113), .C2(n_0_555), .ZN(n_0_351));
   INV_X1 i_0_180 (.A(n_0_352), .ZN(product[6]));
   OAI22_X1 i_0_181 (.A1(n_0_559), .A2(n_0_353), .B1(n_0_341), .B2(n_0_558), 
      .ZN(n_0_352));
   OAI21_X1 i_0_182 (.A(n_0_354), .B1(n_0_545), .B2(n_0_356), .ZN(n_0_353));
   AOI22_X1 i_0_183 (.A1(n_0_187), .A2(n_0_551), .B1(n_0_174), .B2(n_0_548), 
      .ZN(n_0_354));
   INV_X1 i_0_184 (.A(n_0_356), .ZN(n_0_355));
   AOI222_X1 i_0_185 (.A1(n_82), .A2(n_0_556), .B1(n_98), .B2(n_0_557), .C1(
      n_114), .C2(n_0_555), .ZN(n_0_356));
   OAI21_X1 i_0_186 (.A(n_0_357), .B1(n_0_564), .B2(n_0_359), .ZN(product[7]));
   NAND2_X1 i_0_187 (.A1(n_0_342), .A2(n_0_564), .ZN(n_0_357));
   INV_X1 i_0_188 (.A(n_0_359), .ZN(n_0_358));
   AOI222_X1 i_0_189 (.A1(n_0_213), .A2(n_0_562), .B1(n_0_200), .B2(n_0_560), 
      .C1(n_0_558), .C2(n_0_360), .ZN(n_0_359));
   OAI21_X1 i_0_190 (.A(n_0_361), .B1(n_0_545), .B2(n_0_363), .ZN(n_0_360));
   AOI22_X1 i_0_191 (.A1(n_0_188), .A2(n_0_551), .B1(n_0_175), .B2(n_0_548), 
      .ZN(n_0_361));
   INV_X1 i_0_192 (.A(n_0_363), .ZN(n_0_362));
   AOI222_X1 i_0_193 (.A1(n_83), .A2(n_0_556), .B1(n_99), .B2(n_0_557), .C1(
      n_115), .C2(n_0_555), .ZN(n_0_363));
   INV_X1 i_0_194 (.A(n_0_364), .ZN(product[8]));
   OAI22_X1 i_0_195 (.A1(n_0_570), .A2(n_0_365), .B1(n_0_343), .B2(n_0_569), 
      .ZN(n_0_364));
   OAI21_X1 i_0_196 (.A(n_0_366), .B1(n_0_564), .B2(n_0_368), .ZN(n_0_365));
   AOI22_X1 i_0_197 (.A1(n_0_226), .A2(n_0_565), .B1(n_0_238), .B2(n_0_567), 
      .ZN(n_0_366));
   INV_X1 i_0_198 (.A(n_0_368), .ZN(n_0_367));
   AOI222_X1 i_0_199 (.A1(n_0_214), .A2(n_0_562), .B1(n_0_201), .B2(n_0_560), 
      .C1(n_0_558), .C2(n_0_369), .ZN(n_0_368));
   OAI21_X1 i_0_200 (.A(n_0_370), .B1(n_0_545), .B2(n_0_372), .ZN(n_0_369));
   AOI22_X1 i_0_201 (.A1(n_0_189), .A2(n_0_551), .B1(n_0_176), .B2(n_0_548), 
      .ZN(n_0_370));
   INV_X1 i_0_202 (.A(n_0_372), .ZN(n_0_371));
   AOI222_X1 i_0_203 (.A1(n_84), .A2(n_0_556), .B1(n_100), .B2(n_0_557), 
      .C1(n_116), .C2(n_0_555), .ZN(n_0_372));
   OAI21_X1 i_0_204 (.A(n_0_373), .B1(n_0_575), .B2(n_0_375), .ZN(product[9]));
   NAND2_X1 i_0_205 (.A1(n_0_344), .A2(n_0_575), .ZN(n_0_373));
   INV_X1 i_0_206 (.A(n_0_375), .ZN(n_0_374));
   AOI222_X1 i_0_207 (.A1(n_0_261), .A2(n_0_573), .B1(n_0_250), .B2(n_0_571), 
      .C1(n_0_569), .C2(n_0_376), .ZN(n_0_375));
   OAI21_X1 i_0_208 (.A(n_0_377), .B1(n_0_564), .B2(n_0_379), .ZN(n_0_376));
   AOI22_X1 i_0_209 (.A1(n_0_239), .A2(n_0_567), .B1(n_0_227), .B2(n_0_565), 
      .ZN(n_0_377));
   INV_X1 i_0_210 (.A(n_0_379), .ZN(n_0_378));
   AOI222_X1 i_0_211 (.A1(n_0_202), .A2(n_0_560), .B1(n_0_215), .B2(n_0_562), 
      .C1(n_0_558), .C2(n_0_380), .ZN(n_0_379));
   OAI21_X1 i_0_212 (.A(n_0_381), .B1(n_0_545), .B2(n_0_383), .ZN(n_0_380));
   AOI22_X1 i_0_213 (.A1(n_0_177), .A2(n_0_548), .B1(n_0_190), .B2(n_0_551), 
      .ZN(n_0_381));
   INV_X1 i_0_214 (.A(n_0_383), .ZN(n_0_382));
   AOI222_X1 i_0_215 (.A1(n_85), .A2(n_0_556), .B1(n_101), .B2(n_0_557), 
      .C1(n_117), .C2(n_0_555), .ZN(n_0_383));
   INV_X1 i_0_216 (.A(n_0_384), .ZN(product[10]));
   OAI22_X1 i_0_217 (.A1(n_0_581), .A2(n_0_385), .B1(n_0_345), .B2(n_0_580), 
      .ZN(n_0_384));
   OAI21_X1 i_0_218 (.A(n_0_386), .B1(n_0_575), .B2(n_0_388), .ZN(n_0_385));
   AOI22_X1 i_0_219 (.A1(n_0_272), .A2(n_0_578), .B1(n_0_282), .B2(n_0_576), 
      .ZN(n_0_386));
   INV_X1 i_0_220 (.A(n_0_388), .ZN(n_0_387));
   AOI222_X1 i_0_221 (.A1(n_0_251), .A2(n_0_571), .B1(n_0_262), .B2(n_0_573), 
      .C1(n_0_569), .C2(n_0_389), .ZN(n_0_388));
   OAI21_X1 i_0_222 (.A(n_0_390), .B1(n_0_564), .B2(n_0_392), .ZN(n_0_389));
   AOI22_X1 i_0_223 (.A1(n_0_240), .A2(n_0_567), .B1(n_0_228), .B2(n_0_565), 
      .ZN(n_0_390));
   INV_X1 i_0_224 (.A(n_0_392), .ZN(n_0_391));
   AOI222_X1 i_0_225 (.A1(n_0_203), .A2(n_0_560), .B1(n_0_216), .B2(n_0_562), 
      .C1(n_0_558), .C2(n_0_393), .ZN(n_0_392));
   OAI21_X1 i_0_226 (.A(n_0_394), .B1(n_0_545), .B2(n_0_396), .ZN(n_0_393));
   AOI22_X1 i_0_227 (.A1(n_0_178), .A2(n_0_548), .B1(n_0_191), .B2(n_0_551), 
      .ZN(n_0_394));
   INV_X1 i_0_228 (.A(n_0_396), .ZN(n_0_395));
   AOI222_X1 i_0_229 (.A1(n_86), .A2(n_0_556), .B1(n_102), .B2(n_0_557), 
      .C1(n_118), .C2(n_0_555), .ZN(n_0_396));
   OAI21_X1 i_0_230 (.A(n_0_397), .B1(n_0_586), .B2(n_0_399), .ZN(product[11]));
   NAND2_X1 i_0_231 (.A1(n_0_346), .A2(n_0_586), .ZN(n_0_397));
   INV_X1 i_0_232 (.A(n_0_399), .ZN(n_0_398));
   AOI222_X1 i_0_233 (.A1(n_0_301), .A2(n_0_584), .B1(n_0_292), .B2(n_0_582), 
      .C1(n_0_580), .C2(n_0_400), .ZN(n_0_399));
   OAI21_X1 i_0_234 (.A(n_0_401), .B1(n_0_575), .B2(n_0_403), .ZN(n_0_400));
   AOI22_X1 i_0_235 (.A1(n_0_283), .A2(n_0_576), .B1(n_0_273), .B2(n_0_578), 
      .ZN(n_0_401));
   INV_X1 i_0_236 (.A(n_0_403), .ZN(n_0_402));
   AOI222_X1 i_0_237 (.A1(n_0_263), .A2(n_0_573), .B1(n_0_252), .B2(n_0_571), 
      .C1(n_0_569), .C2(n_0_404), .ZN(n_0_403));
   OAI21_X1 i_0_238 (.A(n_0_405), .B1(n_0_564), .B2(n_0_407), .ZN(n_0_404));
   AOI22_X1 i_0_239 (.A1(n_0_241), .A2(n_0_567), .B1(n_0_229), .B2(n_0_565), 
      .ZN(n_0_405));
   INV_X1 i_0_240 (.A(n_0_407), .ZN(n_0_406));
   AOI222_X1 i_0_241 (.A1(n_0_204), .A2(n_0_560), .B1(n_0_217), .B2(n_0_562), 
      .C1(n_0_558), .C2(n_0_408), .ZN(n_0_407));
   OAI21_X1 i_0_242 (.A(n_0_409), .B1(n_0_545), .B2(n_0_411), .ZN(n_0_408));
   AOI22_X1 i_0_243 (.A1(n_0_192), .A2(n_0_551), .B1(n_0_179), .B2(n_0_548), 
      .ZN(n_0_409));
   INV_X1 i_0_244 (.A(n_0_411), .ZN(n_0_410));
   AOI222_X1 i_0_245 (.A1(n_87), .A2(n_0_556), .B1(n_103), .B2(n_0_557), 
      .C1(n_119), .C2(n_0_555), .ZN(n_0_411));
   OAI21_X1 i_0_246 (.A(n_0_412), .B1(n_0_677), .B2(n_0_591), .ZN(product[12]));
   NAND2_X1 i_0_247 (.A1(n_0_591), .A2(n_0_413), .ZN(n_0_412));
   OAI21_X1 i_0_248 (.A(n_0_414), .B1(n_0_586), .B2(n_0_416), .ZN(n_0_413));
   AOI22_X1 i_0_249 (.A1(n_0_318), .A2(n_0_589), .B1(n_0_310), .B2(n_0_587), 
      .ZN(n_0_414));
   INV_X1 i_0_250 (.A(n_0_416), .ZN(n_0_415));
   AOI222_X1 i_0_251 (.A1(n_0_302), .A2(n_0_584), .B1(n_0_293), .B2(n_0_582), 
      .C1(n_0_580), .C2(n_0_417), .ZN(n_0_416));
   OAI21_X1 i_0_252 (.A(n_0_418), .B1(n_0_575), .B2(n_0_420), .ZN(n_0_417));
   AOI22_X1 i_0_253 (.A1(n_0_284), .A2(n_0_576), .B1(n_0_274), .B2(n_0_578), 
      .ZN(n_0_418));
   INV_X1 i_0_254 (.A(n_0_420), .ZN(n_0_419));
   AOI222_X1 i_0_255 (.A1(n_0_264), .A2(n_0_573), .B1(n_0_253), .B2(n_0_571), 
      .C1(n_0_569), .C2(n_0_421), .ZN(n_0_420));
   OAI21_X1 i_0_256 (.A(n_0_422), .B1(n_0_564), .B2(n_0_424), .ZN(n_0_421));
   AOI22_X1 i_0_257 (.A1(n_0_242), .A2(n_0_567), .B1(n_0_230), .B2(n_0_565), 
      .ZN(n_0_422));
   INV_X1 i_0_258 (.A(n_0_424), .ZN(n_0_423));
   AOI222_X1 i_0_259 (.A1(n_0_218), .A2(n_0_562), .B1(n_0_205), .B2(n_0_560), 
      .C1(n_0_558), .C2(n_0_425), .ZN(n_0_424));
   OAI21_X1 i_0_260 (.A(n_0_426), .B1(n_0_545), .B2(n_0_428), .ZN(n_0_425));
   AOI22_X1 i_0_261 (.A1(n_0_180), .A2(n_0_548), .B1(n_0_193), .B2(n_0_551), 
      .ZN(n_0_426));
   INV_X1 i_0_262 (.A(n_0_428), .ZN(n_0_427));
   AOI222_X1 i_0_263 (.A1(n_88), .A2(n_0_556), .B1(n_104), .B2(n_0_557), 
      .C1(n_120), .C2(n_0_555), .ZN(n_0_428));
   INV_X1 i_0_264 (.A(n_0_429), .ZN(product[13]));
   AOI222_X1 i_0_265 (.A1(n_0_333), .A2(n_0_593), .B1(n_0_326), .B2(n_0_592), 
      .C1(n_0_591), .C2(n_0_430), .ZN(n_0_429));
   OAI21_X1 i_0_266 (.A(n_0_431), .B1(n_0_586), .B2(n_0_433), .ZN(n_0_430));
   AOI22_X1 i_0_267 (.A1(n_0_319), .A2(n_0_589), .B1(n_0_311), .B2(n_0_587), 
      .ZN(n_0_431));
   INV_X1 i_0_268 (.A(n_0_433), .ZN(n_0_432));
   AOI222_X1 i_0_269 (.A1(n_0_303), .A2(n_0_584), .B1(n_0_294), .B2(n_0_582), 
      .C1(n_0_580), .C2(n_0_434), .ZN(n_0_433));
   OAI21_X1 i_0_270 (.A(n_0_435), .B1(n_0_575), .B2(n_0_437), .ZN(n_0_434));
   AOI22_X1 i_0_271 (.A1(n_0_285), .A2(n_0_576), .B1(n_0_275), .B2(n_0_578), 
      .ZN(n_0_435));
   INV_X1 i_0_272 (.A(n_0_437), .ZN(n_0_436));
   AOI222_X1 i_0_273 (.A1(n_0_265), .A2(n_0_573), .B1(n_0_254), .B2(n_0_571), 
      .C1(n_0_569), .C2(n_0_438), .ZN(n_0_437));
   OAI21_X1 i_0_274 (.A(n_0_439), .B1(n_0_564), .B2(n_0_441), .ZN(n_0_438));
   AOI22_X1 i_0_275 (.A1(n_0_243), .A2(n_0_567), .B1(n_0_231), .B2(n_0_565), 
      .ZN(n_0_439));
   INV_X1 i_0_276 (.A(n_0_441), .ZN(n_0_440));
   AOI222_X1 i_0_277 (.A1(n_0_219), .A2(n_0_562), .B1(n_0_206), .B2(n_0_560), 
      .C1(n_0_558), .C2(n_0_442), .ZN(n_0_441));
   OAI21_X1 i_0_278 (.A(n_0_443), .B1(n_0_545), .B2(n_0_445), .ZN(n_0_442));
   AOI22_X1 i_0_279 (.A1(n_0_194), .A2(n_0_551), .B1(n_0_181), .B2(n_0_548), 
      .ZN(n_0_443));
   INV_X1 i_0_280 (.A(n_0_445), .ZN(n_0_444));
   AOI222_X1 i_0_281 (.A1(n_89), .A2(n_0_556), .B1(n_105), .B2(n_0_557), 
      .C1(n_121), .C2(n_0_555), .ZN(n_0_445));
   INV_X1 i_0_282 (.A(n_0_446), .ZN(product[14]));
   AOI222_X1 i_0_283 (.A1(n_0_334), .A2(n_0_593), .B1(n_0_327), .B2(n_0_592), 
      .C1(n_0_591), .C2(n_0_447), .ZN(n_0_446));
   OAI21_X1 i_0_284 (.A(n_0_448), .B1(n_0_586), .B2(n_0_450), .ZN(n_0_447));
   AOI22_X1 i_0_285 (.A1(n_0_320), .A2(n_0_589), .B1(n_0_312), .B2(n_0_587), 
      .ZN(n_0_448));
   INV_X1 i_0_286 (.A(n_0_450), .ZN(n_0_449));
   AOI222_X1 i_0_287 (.A1(n_0_304), .A2(n_0_584), .B1(n_0_295), .B2(n_0_582), 
      .C1(n_0_580), .C2(n_0_451), .ZN(n_0_450));
   OAI21_X1 i_0_288 (.A(n_0_452), .B1(n_0_575), .B2(n_0_454), .ZN(n_0_451));
   AOI22_X1 i_0_289 (.A1(n_0_286), .A2(n_0_576), .B1(n_0_276), .B2(n_0_578), 
      .ZN(n_0_452));
   INV_X1 i_0_290 (.A(n_0_454), .ZN(n_0_453));
   AOI222_X1 i_0_291 (.A1(n_0_266), .A2(n_0_573), .B1(n_0_255), .B2(n_0_571), 
      .C1(n_0_569), .C2(n_0_455), .ZN(n_0_454));
   OAI21_X1 i_0_292 (.A(n_0_456), .B1(n_0_564), .B2(n_0_458), .ZN(n_0_455));
   AOI22_X1 i_0_293 (.A1(n_0_244), .A2(n_0_567), .B1(n_0_232), .B2(n_0_565), 
      .ZN(n_0_456));
   INV_X1 i_0_294 (.A(n_0_458), .ZN(n_0_457));
   AOI222_X1 i_0_295 (.A1(n_0_220), .A2(n_0_562), .B1(n_0_207), .B2(n_0_560), 
      .C1(n_0_558), .C2(n_0_459), .ZN(n_0_458));
   OAI21_X1 i_0_296 (.A(n_0_460), .B1(n_0_545), .B2(n_0_462), .ZN(n_0_459));
   AOI22_X1 i_0_297 (.A1(n_0_182), .A2(n_0_548), .B1(n_0_195), .B2(n_0_551), 
      .ZN(n_0_460));
   INV_X1 i_0_298 (.A(n_0_462), .ZN(n_0_461));
   AOI222_X1 i_0_299 (.A1(n_90), .A2(n_0_556), .B1(n_106), .B2(n_0_557), 
      .C1(n_122), .C2(n_0_555), .ZN(n_0_462));
   INV_X1 i_0_300 (.A(n_0_463), .ZN(product[15]));
   AOI222_X1 i_0_301 (.A1(n_0_335), .A2(n_0_593), .B1(n_0_328), .B2(n_0_592), 
      .C1(n_0_591), .C2(n_0_464), .ZN(n_0_463));
   OAI21_X1 i_0_302 (.A(n_0_465), .B1(n_0_586), .B2(n_0_467), .ZN(n_0_464));
   AOI22_X1 i_0_303 (.A1(n_0_321), .A2(n_0_589), .B1(n_0_313), .B2(n_0_587), 
      .ZN(n_0_465));
   INV_X1 i_0_304 (.A(n_0_467), .ZN(n_0_466));
   AOI222_X1 i_0_305 (.A1(n_0_305), .A2(n_0_584), .B1(n_0_296), .B2(n_0_582), 
      .C1(n_0_580), .C2(n_0_468), .ZN(n_0_467));
   OAI21_X1 i_0_306 (.A(n_0_469), .B1(n_0_575), .B2(n_0_471), .ZN(n_0_468));
   AOI22_X1 i_0_307 (.A1(n_0_287), .A2(n_0_576), .B1(n_0_277), .B2(n_0_578), 
      .ZN(n_0_469));
   INV_X1 i_0_308 (.A(n_0_471), .ZN(n_0_470));
   AOI222_X1 i_0_309 (.A1(n_0_267), .A2(n_0_573), .B1(n_0_256), .B2(n_0_571), 
      .C1(n_0_569), .C2(n_0_472), .ZN(n_0_471));
   OAI21_X1 i_0_310 (.A(n_0_473), .B1(n_0_564), .B2(n_0_475), .ZN(n_0_472));
   AOI22_X1 i_0_311 (.A1(n_0_245), .A2(n_0_567), .B1(n_0_233), .B2(n_0_565), 
      .ZN(n_0_473));
   INV_X1 i_0_312 (.A(n_0_475), .ZN(n_0_474));
   AOI222_X1 i_0_313 (.A1(n_0_221), .A2(n_0_562), .B1(n_0_208), .B2(n_0_560), 
      .C1(n_0_558), .C2(n_0_476), .ZN(n_0_475));
   OAI21_X1 i_0_314 (.A(n_0_477), .B1(n_0_545), .B2(n_0_479), .ZN(n_0_476));
   AOI22_X1 i_0_315 (.A1(n_0_183), .A2(n_0_548), .B1(n_0_196), .B2(n_0_551), 
      .ZN(n_0_477));
   INV_X1 i_0_316 (.A(n_0_479), .ZN(n_0_478));
   AOI222_X1 i_0_317 (.A1(n_91), .A2(n_0_556), .B1(n_107), .B2(n_0_557), 
      .C1(n_123), .C2(n_0_555), .ZN(n_0_479));
   INV_X1 i_0_318 (.A(n_0_480), .ZN(product[16]));
   AOI222_X1 i_0_319 (.A1(n_0_336), .A2(n_0_593), .B1(n_0_329), .B2(n_0_592), 
      .C1(n_0_591), .C2(n_0_481), .ZN(n_0_480));
   OAI21_X1 i_0_320 (.A(n_0_482), .B1(n_0_586), .B2(n_0_484), .ZN(n_0_481));
   AOI22_X1 i_0_321 (.A1(n_0_322), .A2(n_0_589), .B1(n_0_314), .B2(n_0_587), 
      .ZN(n_0_482));
   INV_X1 i_0_322 (.A(n_0_484), .ZN(n_0_483));
   AOI222_X1 i_0_323 (.A1(n_0_306), .A2(n_0_584), .B1(n_0_297), .B2(n_0_582), 
      .C1(n_0_580), .C2(n_0_485), .ZN(n_0_484));
   OAI21_X1 i_0_324 (.A(n_0_486), .B1(n_0_575), .B2(n_0_488), .ZN(n_0_485));
   AOI22_X1 i_0_325 (.A1(n_0_288), .A2(n_0_576), .B1(n_0_278), .B2(n_0_578), 
      .ZN(n_0_486));
   INV_X1 i_0_326 (.A(n_0_488), .ZN(n_0_487));
   AOI222_X1 i_0_327 (.A1(n_0_268), .A2(n_0_573), .B1(n_0_257), .B2(n_0_571), 
      .C1(n_0_569), .C2(n_0_489), .ZN(n_0_488));
   OAI21_X1 i_0_328 (.A(n_0_490), .B1(n_0_564), .B2(n_0_492), .ZN(n_0_489));
   AOI22_X1 i_0_329 (.A1(n_0_246), .A2(n_0_567), .B1(n_0_234), .B2(n_0_565), 
      .ZN(n_0_490));
   INV_X1 i_0_330 (.A(n_0_492), .ZN(n_0_491));
   AOI222_X1 i_0_331 (.A1(n_0_222), .A2(n_0_562), .B1(n_0_209), .B2(n_0_560), 
      .C1(n_0_558), .C2(n_0_493), .ZN(n_0_492));
   OAI21_X1 i_0_332 (.A(n_0_494), .B1(n_0_545), .B2(n_0_496), .ZN(n_0_493));
   AOI22_X1 i_0_333 (.A1(n_0_197), .A2(n_0_551), .B1(n_0_184), .B2(n_0_548), 
      .ZN(n_0_494));
   INV_X1 i_0_334 (.A(n_0_496), .ZN(n_0_495));
   AOI222_X1 i_0_335 (.A1(n_92), .A2(n_0_556), .B1(n_108), .B2(n_0_557), 
      .C1(n_124), .C2(n_0_555), .ZN(n_0_496));
   INV_X1 i_0_336 (.A(n_0_497), .ZN(product[17]));
   AOI222_X1 i_0_337 (.A1(n_0_337), .A2(n_0_593), .B1(n_0_330), .B2(n_0_592), 
      .C1(n_0_591), .C2(n_0_498), .ZN(n_0_497));
   OAI21_X1 i_0_338 (.A(n_0_499), .B1(n_0_586), .B2(n_0_501), .ZN(n_0_498));
   AOI22_X1 i_0_339 (.A1(n_0_323), .A2(n_0_589), .B1(n_0_315), .B2(n_0_587), 
      .ZN(n_0_499));
   INV_X1 i_0_340 (.A(n_0_501), .ZN(n_0_500));
   AOI222_X1 i_0_341 (.A1(n_0_307), .A2(n_0_584), .B1(n_0_298), .B2(n_0_582), 
      .C1(n_0_580), .C2(n_0_502), .ZN(n_0_501));
   OAI21_X1 i_0_342 (.A(n_0_503), .B1(n_0_575), .B2(n_0_505), .ZN(n_0_502));
   AOI22_X1 i_0_343 (.A1(n_0_289), .A2(n_0_576), .B1(n_0_279), .B2(n_0_578), 
      .ZN(n_0_503));
   INV_X1 i_0_344 (.A(n_0_505), .ZN(n_0_504));
   AOI222_X1 i_0_345 (.A1(n_0_269), .A2(n_0_573), .B1(n_0_258), .B2(n_0_571), 
      .C1(n_0_569), .C2(n_0_506), .ZN(n_0_505));
   OAI21_X1 i_0_346 (.A(n_0_507), .B1(n_0_564), .B2(n_0_509), .ZN(n_0_506));
   AOI22_X1 i_0_347 (.A1(n_0_247), .A2(n_0_567), .B1(n_0_235), .B2(n_0_565), 
      .ZN(n_0_507));
   INV_X1 i_0_348 (.A(n_0_509), .ZN(n_0_508));
   AOI222_X1 i_0_349 (.A1(n_0_210), .A2(n_0_560), .B1(n_0_223), .B2(n_0_562), 
      .C1(n_0_558), .C2(n_0_510), .ZN(n_0_509));
   OAI21_X1 i_0_350 (.A(n_0_511), .B1(n_0_545), .B2(n_0_513), .ZN(n_0_510));
   AOI22_X1 i_0_351 (.A1(n_0_185), .A2(n_0_548), .B1(n_0_198), .B2(n_0_551), 
      .ZN(n_0_511));
   INV_X1 i_0_352 (.A(n_0_513), .ZN(n_0_512));
   AOI222_X1 i_0_353 (.A1(n_93), .A2(n_0_556), .B1(n_109), .B2(n_0_557), 
      .C1(n_125), .C2(n_0_555), .ZN(n_0_513));
   INV_X1 i_0_354 (.A(n_0_514), .ZN(product[18]));
   AOI222_X1 i_0_355 (.A1(n_0_338), .A2(n_0_593), .B1(n_0_331), .B2(n_0_592), 
      .C1(n_0_591), .C2(n_0_515), .ZN(n_0_514));
   OAI21_X1 i_0_356 (.A(n_0_516), .B1(n_0_586), .B2(n_0_518), .ZN(n_0_515));
   AOI22_X1 i_0_357 (.A1(n_0_324), .A2(n_0_589), .B1(n_0_316), .B2(n_0_587), 
      .ZN(n_0_516));
   INV_X1 i_0_358 (.A(n_0_518), .ZN(n_0_517));
   AOI222_X1 i_0_359 (.A1(n_0_308), .A2(n_0_584), .B1(n_0_299), .B2(n_0_582), 
      .C1(n_0_580), .C2(n_0_519), .ZN(n_0_518));
   OAI21_X1 i_0_360 (.A(n_0_520), .B1(n_0_575), .B2(n_0_522), .ZN(n_0_519));
   AOI22_X1 i_0_361 (.A1(n_0_290), .A2(n_0_576), .B1(n_0_280), .B2(n_0_578), 
      .ZN(n_0_520));
   INV_X1 i_0_362 (.A(n_0_522), .ZN(n_0_521));
   AOI222_X1 i_0_363 (.A1(n_0_270), .A2(n_0_573), .B1(n_0_259), .B2(n_0_571), 
      .C1(n_0_569), .C2(n_0_523), .ZN(n_0_522));
   OAI21_X1 i_0_364 (.A(n_0_524), .B1(n_0_564), .B2(n_0_526), .ZN(n_0_523));
   AOI22_X1 i_0_365 (.A1(n_0_248), .A2(n_0_567), .B1(n_0_236), .B2(n_0_565), 
      .ZN(n_0_524));
   INV_X1 i_0_366 (.A(n_0_526), .ZN(n_0_525));
   AOI222_X1 i_0_367 (.A1(n_0_224), .A2(n_0_562), .B1(n_0_211), .B2(n_0_560), 
      .C1(n_0_558), .C2(n_0_527), .ZN(n_0_526));
   OAI21_X1 i_0_368 (.A(n_0_528), .B1(n_0_545), .B2(n_0_530), .ZN(n_0_527));
   AOI22_X1 i_0_369 (.A1(n_0_199), .A2(n_0_551), .B1(n_0_186), .B2(n_0_548), 
      .ZN(n_0_528));
   INV_X1 i_0_370 (.A(n_0_530), .ZN(n_0_529));
   AOI221_X1 i_0_371 (.A(n_0_554), .B1(n_94), .B2(n_0_556), .C1(n_110), .C2(
      n_0_557), .ZN(n_0_530));
   INV_X1 i_0_372 (.A(n_0_531), .ZN(product[19]));
   AOI222_X1 i_0_373 (.A1(n_0_339), .A2(n_0_593), .B1(n_0_332), .B2(n_0_592), 
      .C1(n_0_591), .C2(n_0_532), .ZN(n_0_531));
   OAI21_X1 i_0_374 (.A(n_0_533), .B1(n_0_586), .B2(n_0_535), .ZN(n_0_532));
   AOI22_X1 i_0_375 (.A1(n_0_325), .A2(n_0_589), .B1(n_0_317), .B2(n_0_587), 
      .ZN(n_0_533));
   INV_X1 i_0_376 (.A(n_0_535), .ZN(n_0_534));
   AOI222_X1 i_0_377 (.A1(n_0_309), .A2(n_0_584), .B1(n_0_300), .B2(n_0_582), 
      .C1(n_0_580), .C2(n_0_536), .ZN(n_0_535));
   OAI21_X1 i_0_378 (.A(n_0_537), .B1(n_0_575), .B2(n_0_539), .ZN(n_0_536));
   AOI22_X1 i_0_379 (.A1(n_0_281), .A2(n_0_578), .B1(n_0_291), .B2(n_0_576), 
      .ZN(n_0_537));
   INV_X1 i_0_380 (.A(n_0_539), .ZN(n_0_538));
   AOI222_X1 i_0_381 (.A1(n_0_271), .A2(n_0_573), .B1(n_0_260), .B2(n_0_571), 
      .C1(n_0_569), .C2(n_0_540), .ZN(n_0_539));
   OAI21_X1 i_0_382 (.A(n_0_541), .B1(n_0_564), .B2(n_0_543), .ZN(n_0_540));
   AOI22_X1 i_0_383 (.A1(n_0_249), .A2(n_0_567), .B1(n_0_237), .B2(n_0_565), 
      .ZN(n_0_541));
   INV_X1 i_0_384 (.A(n_0_543), .ZN(n_0_542));
   AOI222_X1 i_0_385 (.A1(n_0_225), .A2(n_0_562), .B1(n_0_212), .B2(n_0_560), 
      .C1(n_0_558), .C2(n_0_544), .ZN(n_0_543));
   XOR2_X1 i_0_386 (.A(n_0_553), .B(n_0_546), .Z(n_0_544));
   NAND2_X1 i_0_387 (.A1(n_0_552), .A2(n_0_549), .ZN(n_0_545));
   AOI22_X1 i_0_388 (.A1(n_0_551), .A2(n_0_550), .B1(n_0_548), .B2(n_0_547), 
      .ZN(n_0_546));
   XOR2_X1 i_0_389 (.A(B[12]), .B(n_0_14), .Z(n_0_547));
   INV_X1 i_0_390 (.A(n_0_549), .ZN(n_0_548));
   NAND2_X1 i_0_391 (.A1(n_0_683), .A2(A[4]), .ZN(n_0_549));
   XOR2_X1 i_0_392 (.A(n_0_25), .B(n_170), .Z(n_0_550));
   INV_X1 i_0_393 (.A(n_0_552), .ZN(n_0_551));
   NAND2_X1 i_0_394 (.A1(A[5]), .A2(n_0_682), .ZN(n_0_552));
   AOI221_X1 i_0_395 (.A(n_0_554), .B1(n_95), .B2(n_0_556), .C1(n_111), .C2(
      n_0_557), .ZN(n_0_553));
   AND2_X1 i_0_396 (.A1(n_126), .A2(n_0_555), .ZN(n_0_554));
   NOR2_X1 i_0_397 (.A1(n_0_557), .A2(n_0_556), .ZN(n_0_555));
   NOR2_X1 i_0_398 (.A1(A[4]), .A2(n_0_681), .ZN(n_0_556));
   NOR2_X1 i_0_399 (.A1(n_0_682), .A2(A[3]), .ZN(n_0_557));
   INV_X1 i_0_400 (.A(n_0_559), .ZN(n_0_558));
   NAND2_X1 i_0_401 (.A1(n_0_563), .A2(n_0_561), .ZN(n_0_559));
   INV_X1 i_0_402 (.A(n_0_561), .ZN(n_0_560));
   NAND2_X1 i_0_403 (.A1(n_0_684), .A2(A[5]), .ZN(n_0_561));
   INV_X1 i_0_404 (.A(n_0_563), .ZN(n_0_562));
   NAND2_X1 i_0_405 (.A1(A[6]), .A2(n_0_683), .ZN(n_0_563));
   NAND2_X1 i_0_406 (.A1(n_0_568), .A2(n_0_566), .ZN(n_0_564));
   INV_X1 i_0_407 (.A(n_0_566), .ZN(n_0_565));
   NAND2_X1 i_0_408 (.A1(n_0_685), .A2(A[6]), .ZN(n_0_566));
   INV_X1 i_0_409 (.A(n_0_568), .ZN(n_0_567));
   NAND2_X1 i_0_410 (.A1(A[7]), .A2(n_0_684), .ZN(n_0_568));
   INV_X1 i_0_411 (.A(n_0_570), .ZN(n_0_569));
   NAND2_X1 i_0_412 (.A1(n_0_574), .A2(n_0_572), .ZN(n_0_570));
   INV_X1 i_0_413 (.A(n_0_572), .ZN(n_0_571));
   NAND2_X1 i_0_414 (.A1(n_0_686), .A2(A[7]), .ZN(n_0_572));
   INV_X1 i_0_415 (.A(n_0_574), .ZN(n_0_573));
   NAND2_X1 i_0_416 (.A1(A[8]), .A2(n_0_685), .ZN(n_0_574));
   NAND2_X1 i_0_417 (.A1(n_0_579), .A2(n_0_577), .ZN(n_0_575));
   INV_X1 i_0_418 (.A(n_0_577), .ZN(n_0_576));
   NAND2_X1 i_0_419 (.A1(A[9]), .A2(n_0_686), .ZN(n_0_577));
   INV_X1 i_0_420 (.A(n_0_579), .ZN(n_0_578));
   NAND2_X1 i_0_421 (.A1(n_0_687), .A2(A[8]), .ZN(n_0_579));
   INV_X1 i_0_422 (.A(n_0_581), .ZN(n_0_580));
   NAND2_X1 i_0_423 (.A1(n_0_585), .A2(n_0_583), .ZN(n_0_581));
   INV_X1 i_0_424 (.A(n_0_583), .ZN(n_0_582));
   NAND2_X1 i_0_425 (.A1(n_0_688), .A2(A[9]), .ZN(n_0_583));
   INV_X1 i_0_426 (.A(n_0_585), .ZN(n_0_584));
   NAND2_X1 i_0_427 (.A1(A[10]), .A2(n_0_687), .ZN(n_0_585));
   NAND2_X1 i_0_428 (.A1(n_0_590), .A2(n_0_588), .ZN(n_0_586));
   INV_X1 i_0_429 (.A(n_0_588), .ZN(n_0_587));
   NAND2_X1 i_0_430 (.A1(n_0_689), .A2(A[10]), .ZN(n_0_588));
   INV_X1 i_0_431 (.A(n_0_590), .ZN(n_0_589));
   NAND2_X1 i_0_432 (.A1(A[11]), .A2(n_0_688), .ZN(n_0_590));
   NOR2_X1 i_0_433 (.A1(n_0_593), .A2(n_0_592), .ZN(n_0_591));
   NOR2_X1 i_0_434 (.A1(A[12]), .A2(n_0_689), .ZN(n_0_592));
   AND2_X1 i_0_435 (.A1(A[12]), .A2(n_0_689), .ZN(n_0_593));
   INV_X1 i_0_436 (.A(n_0_594), .ZN(product[3]));
   AOI222_X1 i_0_437 (.A1(n_48), .A2(n_0_612), .B1(n_64), .B2(n_0_613), .C1(
      n_127), .C2(n_0_611), .ZN(n_0_594));
   INV_X1 i_0_438 (.A(n_0_595), .ZN(n_112));
   AOI222_X1 i_0_439 (.A1(n_49), .A2(n_0_612), .B1(n_65), .B2(n_0_613), .C1(
      n_128), .C2(n_0_611), .ZN(n_0_595));
   INV_X1 i_0_440 (.A(n_0_596), .ZN(n_113));
   AOI222_X1 i_0_441 (.A1(n_50), .A2(n_0_612), .B1(n_66), .B2(n_0_613), .C1(
      n_129), .C2(n_0_611), .ZN(n_0_596));
   INV_X1 i_0_442 (.A(n_0_597), .ZN(n_114));
   AOI222_X1 i_0_443 (.A1(n_51), .A2(n_0_612), .B1(n_67), .B2(n_0_613), .C1(
      n_130), .C2(n_0_611), .ZN(n_0_597));
   INV_X1 i_0_444 (.A(n_0_598), .ZN(n_115));
   AOI222_X1 i_0_445 (.A1(n_52), .A2(n_0_612), .B1(n_68), .B2(n_0_613), .C1(
      n_131), .C2(n_0_611), .ZN(n_0_598));
   INV_X1 i_0_446 (.A(n_0_599), .ZN(n_116));
   AOI222_X1 i_0_447 (.A1(n_53), .A2(n_0_612), .B1(n_69), .B2(n_0_613), .C1(
      n_132), .C2(n_0_611), .ZN(n_0_599));
   INV_X1 i_0_448 (.A(n_0_600), .ZN(n_117));
   AOI222_X1 i_0_449 (.A1(n_54), .A2(n_0_612), .B1(n_70), .B2(n_0_613), .C1(
      n_133), .C2(n_0_611), .ZN(n_0_600));
   INV_X1 i_0_450 (.A(n_0_601), .ZN(n_118));
   AOI222_X1 i_0_451 (.A1(n_55), .A2(n_0_612), .B1(n_71), .B2(n_0_613), .C1(
      n_134), .C2(n_0_611), .ZN(n_0_601));
   INV_X1 i_0_452 (.A(n_0_602), .ZN(n_119));
   AOI222_X1 i_0_453 (.A1(n_56), .A2(n_0_612), .B1(n_72), .B2(n_0_613), .C1(
      n_135), .C2(n_0_611), .ZN(n_0_602));
   INV_X1 i_0_454 (.A(n_0_603), .ZN(n_120));
   AOI222_X1 i_0_455 (.A1(n_57), .A2(n_0_612), .B1(n_73), .B2(n_0_613), .C1(
      n_136), .C2(n_0_611), .ZN(n_0_603));
   INV_X1 i_0_456 (.A(n_0_604), .ZN(n_121));
   AOI222_X1 i_0_457 (.A1(n_58), .A2(n_0_612), .B1(n_74), .B2(n_0_613), .C1(
      n_137), .C2(n_0_611), .ZN(n_0_604));
   INV_X1 i_0_458 (.A(n_0_605), .ZN(n_122));
   AOI222_X1 i_0_459 (.A1(n_59), .A2(n_0_612), .B1(n_75), .B2(n_0_613), .C1(
      n_138), .C2(n_0_611), .ZN(n_0_605));
   INV_X1 i_0_460 (.A(n_0_606), .ZN(n_123));
   AOI222_X1 i_0_461 (.A1(n_60), .A2(n_0_612), .B1(n_76), .B2(n_0_613), .C1(
      n_139), .C2(n_0_611), .ZN(n_0_606));
   INV_X1 i_0_462 (.A(n_0_607), .ZN(n_124));
   AOI222_X1 i_0_463 (.A1(n_61), .A2(n_0_612), .B1(n_77), .B2(n_0_613), .C1(
      n_140), .C2(n_0_611), .ZN(n_0_607));
   INV_X1 i_0_464 (.A(n_0_608), .ZN(n_125));
   AOI221_X1 i_0_465 (.A(n_0_610), .B1(n_62), .B2(n_0_612), .C1(n_78), .C2(
      n_0_613), .ZN(n_0_608));
   INV_X1 i_0_466 (.A(n_0_609), .ZN(n_126));
   AOI221_X1 i_0_467 (.A(n_0_610), .B1(n_63), .B2(n_0_612), .C1(n_79), .C2(
      n_0_613), .ZN(n_0_609));
   AND2_X1 i_0_468 (.A1(n_141), .A2(n_0_611), .ZN(n_0_610));
   NOR2_X1 i_0_469 (.A1(n_0_613), .A2(n_0_612), .ZN(n_0_611));
   NOR2_X1 i_0_470 (.A1(A[3]), .A2(n_0_680), .ZN(n_0_612));
   NOR2_X1 i_0_471 (.A1(n_0_681), .A2(A[2]), .ZN(n_0_613));
   INV_X1 i_0_472 (.A(n_0_614), .ZN(product[2]));
   AOI222_X1 i_0_473 (.A1(n_16), .A2(n_0_633), .B1(n_32), .B2(n_0_632), .C1(
      n_142), .C2(n_0_631), .ZN(n_0_614));
   INV_X1 i_0_474 (.A(n_0_615), .ZN(n_127));
   AOI222_X1 i_0_475 (.A1(n_17), .A2(n_0_633), .B1(n_33), .B2(n_0_632), .C1(
      n_143), .C2(n_0_631), .ZN(n_0_615));
   INV_X1 i_0_476 (.A(n_0_616), .ZN(n_128));
   AOI222_X1 i_0_477 (.A1(n_18), .A2(n_0_633), .B1(n_34), .B2(n_0_632), .C1(
      n_144), .C2(n_0_631), .ZN(n_0_616));
   INV_X1 i_0_478 (.A(n_0_617), .ZN(n_129));
   AOI222_X1 i_0_479 (.A1(n_19), .A2(n_0_633), .B1(n_35), .B2(n_0_632), .C1(
      n_145), .C2(n_0_631), .ZN(n_0_617));
   INV_X1 i_0_480 (.A(n_0_618), .ZN(n_130));
   AOI222_X1 i_0_481 (.A1(n_20), .A2(n_0_633), .B1(n_36), .B2(n_0_632), .C1(
      n_146), .C2(n_0_631), .ZN(n_0_618));
   INV_X1 i_0_482 (.A(n_0_619), .ZN(n_131));
   AOI222_X1 i_0_483 (.A1(n_21), .A2(n_0_633), .B1(n_37), .B2(n_0_632), .C1(
      n_147), .C2(n_0_631), .ZN(n_0_619));
   INV_X1 i_0_484 (.A(n_0_620), .ZN(n_132));
   AOI222_X1 i_0_485 (.A1(n_22), .A2(n_0_633), .B1(n_38), .B2(n_0_632), .C1(
      n_148), .C2(n_0_631), .ZN(n_0_620));
   INV_X1 i_0_486 (.A(n_0_621), .ZN(n_133));
   AOI222_X1 i_0_487 (.A1(n_23), .A2(n_0_633), .B1(n_39), .B2(n_0_632), .C1(
      n_149), .C2(n_0_631), .ZN(n_0_621));
   INV_X1 i_0_488 (.A(n_0_622), .ZN(n_134));
   AOI222_X1 i_0_489 (.A1(n_24), .A2(n_0_633), .B1(n_40), .B2(n_0_632), .C1(
      n_150), .C2(n_0_631), .ZN(n_0_622));
   INV_X1 i_0_490 (.A(n_0_623), .ZN(n_135));
   AOI222_X1 i_0_491 (.A1(n_25), .A2(n_0_633), .B1(n_41), .B2(n_0_632), .C1(
      n_151), .C2(n_0_631), .ZN(n_0_623));
   INV_X1 i_0_492 (.A(n_0_624), .ZN(n_136));
   AOI222_X1 i_0_493 (.A1(n_26), .A2(n_0_633), .B1(n_42), .B2(n_0_632), .C1(
      n_152), .C2(n_0_631), .ZN(n_0_624));
   INV_X1 i_0_494 (.A(n_0_625), .ZN(n_137));
   AOI222_X1 i_0_495 (.A1(n_27), .A2(n_0_633), .B1(n_43), .B2(n_0_632), .C1(
      n_153), .C2(n_0_631), .ZN(n_0_625));
   INV_X1 i_0_496 (.A(n_0_626), .ZN(n_138));
   AOI222_X1 i_0_497 (.A1(n_28), .A2(n_0_633), .B1(n_44), .B2(n_0_632), .C1(
      n_154), .C2(n_0_631), .ZN(n_0_626));
   INV_X1 i_0_498 (.A(n_0_627), .ZN(n_139));
   AOI222_X1 i_0_499 (.A1(n_29), .A2(n_0_633), .B1(n_45), .B2(n_0_632), .C1(
      n_155), .C2(n_0_631), .ZN(n_0_627));
   INV_X1 i_0_500 (.A(n_0_628), .ZN(n_140));
   AOI221_X1 i_0_501 (.A(n_0_630), .B1(n_30), .B2(n_0_633), .C1(n_46), .C2(
      n_0_632), .ZN(n_0_628));
   INV_X1 i_0_502 (.A(n_0_629), .ZN(n_141));
   AOI221_X1 i_0_503 (.A(n_0_630), .B1(n_31), .B2(n_0_633), .C1(n_47), .C2(
      n_0_632), .ZN(n_0_629));
   AND2_X1 i_0_504 (.A1(n_156), .A2(n_0_631), .ZN(n_0_630));
   NOR2_X1 i_0_505 (.A1(n_0_633), .A2(n_0_632), .ZN(n_0_631));
   NOR2_X1 i_0_506 (.A1(n_0_680), .A2(A[1]), .ZN(n_0_632));
   NOR2_X1 i_0_507 (.A1(A[2]), .A2(n_0_679), .ZN(n_0_633));
   INV_X1 i_0_508 (.A(n_0_634), .ZN(product[1]));
   AOI222_X1 i_0_509 (.A1(n_0), .A2(n_0_653), .B1(B[0]), .B2(n_0_651), .C1(n_158), 
      .C2(n_0_650), .ZN(n_0_634));
   INV_X1 i_0_510 (.A(n_0_635), .ZN(n_142));
   AOI222_X1 i_0_511 (.A1(n_1), .A2(n_0_653), .B1(n_158), .B2(n_0_651), .C1(
      n_159), .C2(n_0_650), .ZN(n_0_635));
   INV_X1 i_0_512 (.A(n_0_636), .ZN(n_143));
   AOI222_X1 i_0_513 (.A1(n_2), .A2(n_0_653), .B1(n_159), .B2(n_0_651), .C1(
      n_160), .C2(n_0_650), .ZN(n_0_636));
   INV_X1 i_0_514 (.A(n_0_637), .ZN(n_144));
   AOI222_X1 i_0_515 (.A1(n_3), .A2(n_0_653), .B1(n_160), .B2(n_0_651), .C1(
      n_161), .C2(n_0_650), .ZN(n_0_637));
   INV_X1 i_0_516 (.A(n_0_638), .ZN(n_145));
   AOI222_X1 i_0_517 (.A1(n_4), .A2(n_0_653), .B1(n_161), .B2(n_0_651), .C1(
      n_162), .C2(n_0_650), .ZN(n_0_638));
   INV_X1 i_0_518 (.A(n_0_639), .ZN(n_146));
   AOI222_X1 i_0_519 (.A1(n_162), .A2(n_0_651), .B1(n_5), .B2(n_0_653), .C1(
      n_163), .C2(n_0_650), .ZN(n_0_639));
   INV_X1 i_0_520 (.A(n_0_640), .ZN(n_147));
   AOI222_X1 i_0_521 (.A1(n_6), .A2(n_0_653), .B1(n_163), .B2(n_0_651), .C1(
      n_164), .C2(n_0_650), .ZN(n_0_640));
   INV_X1 i_0_522 (.A(n_0_641), .ZN(n_148));
   AOI222_X1 i_0_523 (.A1(n_164), .A2(n_0_651), .B1(n_7), .B2(n_0_653), .C1(
      n_165), .C2(n_0_650), .ZN(n_0_641));
   INV_X1 i_0_524 (.A(n_0_642), .ZN(n_149));
   AOI222_X1 i_0_525 (.A1(n_8), .A2(n_0_653), .B1(n_165), .B2(n_0_651), .C1(
      n_166), .C2(n_0_650), .ZN(n_0_642));
   INV_X1 i_0_526 (.A(n_0_643), .ZN(n_150));
   AOI222_X1 i_0_527 (.A1(n_9), .A2(n_0_653), .B1(n_166), .B2(n_0_651), .C1(
      n_167), .C2(n_0_650), .ZN(n_0_643));
   INV_X1 i_0_528 (.A(n_0_644), .ZN(n_151));
   AOI222_X1 i_0_529 (.A1(n_10), .A2(n_0_653), .B1(n_167), .B2(n_0_651), 
      .C1(n_168), .C2(n_0_650), .ZN(n_0_644));
   INV_X1 i_0_530 (.A(n_0_645), .ZN(n_152));
   AOI222_X1 i_0_531 (.A1(n_11), .A2(n_0_653), .B1(n_168), .B2(n_0_651), 
      .C1(n_169), .C2(n_0_650), .ZN(n_0_645));
   INV_X1 i_0_532 (.A(n_0_646), .ZN(n_153));
   AOI222_X1 i_0_533 (.A1(A[1]), .A2(n_157), .B1(n_12), .B2(n_0_653), .C1(n_169), 
      .C2(n_0_651), .ZN(n_0_646));
   INV_X1 i_0_534 (.A(n_0_647), .ZN(n_154));
   AOI21_X1 i_0_535 (.A(n_0_652), .B1(n_13), .B2(n_0_653), .ZN(n_0_647));
   INV_X1 i_0_536 (.A(n_0_648), .ZN(n_155));
   AOI21_X1 i_0_537 (.A(n_0_652), .B1(n_14), .B2(n_0_653), .ZN(n_0_648));
   INV_X1 i_0_538 (.A(n_0_649), .ZN(n_156));
   AOI21_X1 i_0_539 (.A(n_0_652), .B1(n_15), .B2(n_0_653), .ZN(n_0_649));
   NOR2_X1 i_0_540 (.A1(n_0_678), .A2(n_0_653), .ZN(n_0_650));
   NOR2_X1 i_0_541 (.A1(n_0_679), .A2(A[0]), .ZN(n_0_651));
   NOR2_X1 i_0_542 (.A1(n_0_679), .A2(n_0_655), .ZN(n_0_652));
   NOR2_X1 i_0_543 (.A1(A[1]), .A2(n_0_678), .ZN(n_0_653));
   AND2_X1 i_0_544 (.A1(B[0]), .A2(A[0]), .ZN(product[0]));
   NOR2_X1 i_0_545 (.A1(n_0_678), .A2(n_0_655), .ZN(n_157));
   AOI21_X1 i_0_546 (.A(n_0_676), .B1(B[1]), .B2(B[0]), .ZN(n_158));
   AOI21_X1 i_0_547 (.A(n_0_674), .B1(B[2]), .B2(n_0_675), .ZN(n_159));
   AOI21_X1 i_0_548 (.A(n_0_672), .B1(B[3]), .B2(n_0_673), .ZN(n_160));
   AOI21_X1 i_0_549 (.A(n_0_670), .B1(B[4]), .B2(n_0_671), .ZN(n_161));
   AOI21_X1 i_0_550 (.A(n_0_668), .B1(B[5]), .B2(n_0_669), .ZN(n_162));
   AOI21_X1 i_0_551 (.A(n_0_666), .B1(B[6]), .B2(n_0_667), .ZN(n_163));
   AOI21_X1 i_0_552 (.A(n_0_664), .B1(B[7]), .B2(n_0_665), .ZN(n_164));
   AOI21_X1 i_0_553 (.A(n_0_662), .B1(B[8]), .B2(n_0_663), .ZN(n_165));
   AOI21_X1 i_0_554 (.A(n_0_660), .B1(B[9]), .B2(n_0_661), .ZN(n_166));
   AOI21_X1 i_0_555 (.A(n_0_658), .B1(B[10]), .B2(n_0_659), .ZN(n_167));
   AOI21_X1 i_0_556 (.A(n_0_656), .B1(B[11]), .B2(n_0_657), .ZN(n_168));
   INV_X1 i_0_557 (.A(n_0_654), .ZN(n_169));
   AOI21_X1 i_0_558 (.A(n_170), .B1(B[12]), .B2(n_0_656), .ZN(n_0_654));
   INV_X1 i_0_559 (.A(n_170), .ZN(n_0_655));
   NOR2_X1 i_0_560 (.A1(B[12]), .A2(n_0_656), .ZN(n_170));
   NOR2_X1 i_0_561 (.A1(B[11]), .A2(n_0_657), .ZN(n_0_656));
   INV_X1 i_0_562 (.A(n_0_658), .ZN(n_0_657));
   NOR2_X1 i_0_563 (.A1(B[10]), .A2(n_0_659), .ZN(n_0_658));
   INV_X1 i_0_564 (.A(n_0_660), .ZN(n_0_659));
   NOR2_X1 i_0_565 (.A1(B[9]), .A2(n_0_661), .ZN(n_0_660));
   INV_X1 i_0_566 (.A(n_0_662), .ZN(n_0_661));
   NOR2_X1 i_0_567 (.A1(B[8]), .A2(n_0_663), .ZN(n_0_662));
   INV_X1 i_0_568 (.A(n_0_664), .ZN(n_0_663));
   NOR2_X1 i_0_569 (.A1(B[7]), .A2(n_0_665), .ZN(n_0_664));
   INV_X1 i_0_570 (.A(n_0_666), .ZN(n_0_665));
   NOR2_X1 i_0_571 (.A1(B[6]), .A2(n_0_667), .ZN(n_0_666));
   INV_X1 i_0_572 (.A(n_0_668), .ZN(n_0_667));
   NOR2_X1 i_0_573 (.A1(B[5]), .A2(n_0_669), .ZN(n_0_668));
   INV_X1 i_0_574 (.A(n_0_670), .ZN(n_0_669));
   NOR2_X1 i_0_575 (.A1(B[4]), .A2(n_0_671), .ZN(n_0_670));
   INV_X1 i_0_576 (.A(n_0_672), .ZN(n_0_671));
   NOR2_X1 i_0_577 (.A1(B[3]), .A2(n_0_673), .ZN(n_0_672));
   INV_X1 i_0_578 (.A(n_0_674), .ZN(n_0_673));
   NOR2_X1 i_0_579 (.A1(B[2]), .A2(n_0_675), .ZN(n_0_674));
   INV_X1 i_0_580 (.A(n_0_676), .ZN(n_0_675));
   NOR2_X1 i_0_581 (.A1(B[1]), .A2(B[0]), .ZN(n_0_676));
   INV_X1 i_0_582 (.A(n_0_347), .ZN(n_0_677));
   INV_X1 i_0_583 (.A(A[0]), .ZN(n_0_678));
   INV_X1 i_0_584 (.A(A[1]), .ZN(n_0_679));
   INV_X1 i_0_585 (.A(A[2]), .ZN(n_0_680));
   INV_X1 i_0_586 (.A(A[3]), .ZN(n_0_681));
   INV_X1 i_0_587 (.A(A[4]), .ZN(n_0_682));
   INV_X1 i_0_588 (.A(A[5]), .ZN(n_0_683));
   INV_X1 i_0_589 (.A(A[6]), .ZN(n_0_684));
   INV_X1 i_0_590 (.A(A[7]), .ZN(n_0_685));
   INV_X1 i_0_591 (.A(A[8]), .ZN(n_0_686));
   INV_X1 i_0_592 (.A(A[9]), .ZN(n_0_687));
   INV_X1 i_0_593 (.A(A[10]), .ZN(n_0_688));
   INV_X1 i_0_594 (.A(A[11]), .ZN(n_0_689));
endmodule

module multiplier_16bit(first_operand, second_operand, out, enable, overflow);
   input [15:0]first_operand;
   input [15:0]second_operand;
   output [15:0]out;
   input enable;
   output overflow;

   wire [31:0]temp_result_wire;
   wire [15:0]second_operand_number;
   wire [15:0]first_operand_number;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;

   booth_16bit_multiplier mult (.A({uc_0, uc_1, uc_2, first_operand_number[12], 
      first_operand_number[11], first_operand_number[10], 
      first_operand_number[9], first_operand_number[8], first_operand_number[7], 
      first_operand_number[6], first_operand_number[5], first_operand_number[4], 
      first_operand_number[3], first_operand_number[2], first_operand_number[1], 
      first_operand_number[0]}), .B({uc_3, uc_4, uc_5, second_operand_number[12], 
      second_operand_number[11], second_operand_number[10], 
      second_operand_number[9], second_operand_number[8], 
      second_operand_number[7], second_operand_number[6], 
      second_operand_number[5], second_operand_number[4], 
      second_operand_number[3], second_operand_number[2], 
      second_operand_number[1], second_operand_number[0]}), .product({uc_6, uc_7, 
      uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, 
      temp_result_wire[19], temp_result_wire[18], temp_result_wire[17], 
      temp_result_wire[16], temp_result_wire[15], temp_result_wire[14], 
      temp_result_wire[13], temp_result_wire[12], temp_result_wire[11], 
      temp_result_wire[10], temp_result_wire[9], temp_result_wire[8], 
      temp_result_wire[7], temp_result_wire[6], temp_result_wire[5], 
      temp_result_wire[4], temp_result_wire[3], temp_result_wire[2], 
      temp_result_wire[1], temp_result_wire[0]}));
   DLH_X1 \out_reg[15]  (.D(n_15), .G(enable), .Q(out[15]));
   DLH_X1 \out_reg[14]  (.D(n_14), .G(enable), .Q(out[14]));
   DLH_X1 \out_reg[13]  (.D(n_13), .G(enable), .Q(out[13]));
   DLH_X1 \out_reg[12]  (.D(n_12), .G(enable), .Q(out[12]));
   DLH_X1 \out_reg[11]  (.D(n_11), .G(enable), .Q(out[11]));
   DLH_X1 \out_reg[10]  (.D(n_10), .G(enable), .Q(out[10]));
   DLH_X1 \out_reg[9]  (.D(n_9), .G(enable), .Q(out[9]));
   DLH_X1 \out_reg[8]  (.D(n_8), .G(enable), .Q(out[8]));
   DLH_X1 \out_reg[7]  (.D(n_7), .G(enable), .Q(out[7]));
   DLH_X1 \out_reg[6]  (.D(n_6), .G(enable), .Q(out[6]));
   DLH_X1 \out_reg[5]  (.D(n_5), .G(enable), .Q(out[5]));
   DLH_X1 \out_reg[4]  (.D(n_4), .G(enable), .Q(out[4]));
   DLH_X1 \out_reg[3]  (.D(n_3), .G(enable), .Q(out[3]));
   DLH_X1 \out_reg[2]  (.D(n_2), .G(enable), .Q(out[2]));
   DLH_X1 \out_reg[1]  (.D(n_1), .G(enable), .Q(out[1]));
   DLH_X1 \out_reg[0]  (.D(n_0), .G(enable), .Q(out[0]));
   DLH_X1 \second_operand_number_reg[12]  (.D(second_operand[12]), .G(enable), 
      .Q(second_operand_number[12]));
   DLH_X1 \second_operand_number_reg[11]  (.D(second_operand[11]), .G(enable), 
      .Q(second_operand_number[11]));
   DLH_X1 \second_operand_number_reg[10]  (.D(second_operand[10]), .G(enable), 
      .Q(second_operand_number[10]));
   DLH_X1 \second_operand_number_reg[9]  (.D(second_operand[9]), .G(enable), 
      .Q(second_operand_number[9]));
   DLH_X1 \second_operand_number_reg[8]  (.D(second_operand[8]), .G(enable), 
      .Q(second_operand_number[8]));
   DLH_X1 \second_operand_number_reg[7]  (.D(second_operand[7]), .G(enable), 
      .Q(second_operand_number[7]));
   DLH_X1 \second_operand_number_reg[6]  (.D(second_operand[6]), .G(enable), 
      .Q(second_operand_number[6]));
   DLH_X1 \second_operand_number_reg[5]  (.D(second_operand[5]), .G(enable), 
      .Q(second_operand_number[5]));
   DLH_X1 \second_operand_number_reg[4]  (.D(second_operand[4]), .G(enable), 
      .Q(second_operand_number[4]));
   DLH_X1 \second_operand_number_reg[3]  (.D(second_operand[3]), .G(enable), 
      .Q(second_operand_number[3]));
   DLH_X1 \second_operand_number_reg[2]  (.D(second_operand[2]), .G(enable), 
      .Q(second_operand_number[2]));
   DLH_X1 \second_operand_number_reg[1]  (.D(second_operand[1]), .G(enable), 
      .Q(second_operand_number[1]));
   DLH_X1 \second_operand_number_reg[0]  (.D(second_operand[0]), .G(enable), 
      .Q(second_operand_number[0]));
   DLH_X1 \first_operand_number_reg[12]  (.D(first_operand[12]), .G(enable), 
      .Q(first_operand_number[12]));
   DLH_X1 \first_operand_number_reg[11]  (.D(first_operand[11]), .G(enable), 
      .Q(first_operand_number[11]));
   DLH_X1 \first_operand_number_reg[10]  (.D(first_operand[10]), .G(enable), 
      .Q(first_operand_number[10]));
   DLH_X1 \first_operand_number_reg[9]  (.D(first_operand[9]), .G(enable), 
      .Q(first_operand_number[9]));
   DLH_X1 \first_operand_number_reg[8]  (.D(first_operand[8]), .G(enable), 
      .Q(first_operand_number[8]));
   DLH_X1 \first_operand_number_reg[7]  (.D(first_operand[7]), .G(enable), 
      .Q(first_operand_number[7]));
   DLH_X1 \first_operand_number_reg[6]  (.D(first_operand[6]), .G(enable), 
      .Q(first_operand_number[6]));
   DLH_X1 \first_operand_number_reg[5]  (.D(first_operand[5]), .G(enable), 
      .Q(first_operand_number[5]));
   DLH_X1 \first_operand_number_reg[4]  (.D(first_operand[4]), .G(enable), 
      .Q(first_operand_number[4]));
   DLH_X1 \first_operand_number_reg[3]  (.D(first_operand[3]), .G(enable), 
      .Q(first_operand_number[3]));
   DLH_X1 \first_operand_number_reg[2]  (.D(first_operand[2]), .G(enable), 
      .Q(first_operand_number[2]));
   DLH_X1 \first_operand_number_reg[1]  (.D(first_operand[1]), .G(enable), 
      .Q(first_operand_number[1]));
   DLH_X1 \first_operand_number_reg[0]  (.D(first_operand[0]), .G(enable), 
      .Q(first_operand_number[0]));
   MUX2_X1 i_0_0 (.A(temp_result_wire[0]), .B(temp_result_wire[4]), .S(n_0_41), 
      .Z(n_0_0));
   MUX2_X1 i_0_1 (.A(temp_result_wire[1]), .B(temp_result_wire[5]), .S(n_0_41), 
      .Z(n_0_1));
   MUX2_X1 i_0_2 (.A(temp_result_wire[2]), .B(temp_result_wire[6]), .S(n_0_41), 
      .Z(n_0_2));
   MUX2_X1 i_0_3 (.A(temp_result_wire[3]), .B(temp_result_wire[7]), .S(n_0_41), 
      .Z(n_0_3));
   MUX2_X1 i_0_4 (.A(temp_result_wire[4]), .B(temp_result_wire[8]), .S(n_0_41), 
      .Z(n_0_4));
   MUX2_X1 i_0_5 (.A(temp_result_wire[5]), .B(temp_result_wire[9]), .S(n_0_41), 
      .Z(n_0_5));
   MUX2_X1 i_0_6 (.A(temp_result_wire[6]), .B(temp_result_wire[10]), .S(n_0_41), 
      .Z(n_0_6));
   MUX2_X1 i_0_7 (.A(temp_result_wire[7]), .B(temp_result_wire[11]), .S(n_0_41), 
      .Z(n_0_7));
   MUX2_X1 i_0_8 (.A(temp_result_wire[8]), .B(temp_result_wire[12]), .S(n_0_41), 
      .Z(n_0_8));
   MUX2_X1 i_0_9 (.A(temp_result_wire[9]), .B(temp_result_wire[13]), .S(n_0_41), 
      .Z(n_0_9));
   MUX2_X1 i_0_10 (.A(temp_result_wire[10]), .B(temp_result_wire[14]), .S(n_0_41), 
      .Z(n_0_10));
   MUX2_X1 i_0_11 (.A(temp_result_wire[11]), .B(temp_result_wire[15]), .S(n_0_41), 
      .Z(n_0_11));
   MUX2_X1 i_0_12 (.A(temp_result_wire[12]), .B(temp_result_wire[16]), .S(n_0_41), 
      .Z(n_0_12));
   MUX2_X1 i_0_13 (.A(temp_result_wire[13]), .B(temp_result_wire[17]), .S(n_0_41), 
      .Z(n_0_13));
   MUX2_X1 i_0_14 (.A(temp_result_wire[14]), .B(temp_result_wire[18]), .S(n_0_41), 
      .Z(n_0_14));
   MUX2_X1 i_0_15 (.A(temp_result_wire[15]), .B(temp_result_wire[19]), .S(n_0_41), 
      .Z(n_0_15));
   MUX2_X1 i_0_16 (.A(n_0_0), .B(n_0_2), .S(n_0_40), .Z(n_0_16));
   MUX2_X1 i_0_17 (.A(n_0_1), .B(n_0_3), .S(n_0_40), .Z(n_0_17));
   MUX2_X1 i_0_18 (.A(n_0_2), .B(n_0_4), .S(n_0_40), .Z(n_0_18));
   MUX2_X1 i_0_19 (.A(n_0_3), .B(n_0_5), .S(n_0_40), .Z(n_0_19));
   MUX2_X1 i_0_20 (.A(n_0_4), .B(n_0_6), .S(n_0_40), .Z(n_0_20));
   MUX2_X1 i_0_21 (.A(n_0_5), .B(n_0_7), .S(n_0_40), .Z(n_0_21));
   MUX2_X1 i_0_22 (.A(n_0_6), .B(n_0_8), .S(n_0_40), .Z(n_0_22));
   MUX2_X1 i_0_23 (.A(n_0_7), .B(n_0_9), .S(n_0_40), .Z(n_0_23));
   MUX2_X1 i_0_24 (.A(n_0_8), .B(n_0_10), .S(n_0_40), .Z(n_0_24));
   MUX2_X1 i_0_25 (.A(n_0_9), .B(n_0_11), .S(n_0_40), .Z(n_0_25));
   MUX2_X1 i_0_26 (.A(n_0_10), .B(n_0_12), .S(n_0_40), .Z(n_0_26));
   MUX2_X1 i_0_27 (.A(n_0_11), .B(n_0_13), .S(n_0_40), .Z(n_0_27));
   MUX2_X1 i_0_28 (.A(n_0_12), .B(n_0_14), .S(n_0_40), .Z(n_0_28));
   MUX2_X1 i_0_29 (.A(n_0_13), .B(n_0_15), .S(n_0_40), .Z(n_0_29));
   MUX2_X1 i_0_30 (.A(n_0_16), .B(n_0_17), .S(n_0_39), .Z(n_0));
   MUX2_X1 i_0_31 (.A(n_0_17), .B(n_0_18), .S(n_0_39), .Z(n_1));
   MUX2_X1 i_0_32 (.A(n_0_18), .B(n_0_19), .S(n_0_39), .Z(n_2));
   MUX2_X1 i_0_33 (.A(n_0_19), .B(n_0_20), .S(n_0_39), .Z(n_3));
   MUX2_X1 i_0_34 (.A(n_0_20), .B(n_0_21), .S(n_0_39), .Z(n_4));
   MUX2_X1 i_0_35 (.A(n_0_21), .B(n_0_22), .S(n_0_39), .Z(n_5));
   MUX2_X1 i_0_36 (.A(n_0_22), .B(n_0_23), .S(n_0_39), .Z(n_6));
   MUX2_X1 i_0_37 (.A(n_0_23), .B(n_0_24), .S(n_0_39), .Z(n_7));
   MUX2_X1 i_0_38 (.A(n_0_24), .B(n_0_25), .S(n_0_39), .Z(n_8));
   MUX2_X1 i_0_39 (.A(n_0_25), .B(n_0_26), .S(n_0_39), .Z(n_9));
   MUX2_X1 i_0_40 (.A(n_0_26), .B(n_0_27), .S(n_0_39), .Z(n_10));
   MUX2_X1 i_0_41 (.A(n_0_27), .B(n_0_28), .S(n_0_39), .Z(n_11));
   MUX2_X1 i_0_42 (.A(n_0_28), .B(n_0_29), .S(n_0_39), .Z(n_12));
   INV_X1 i_0_43 (.A(second_operand[13]), .ZN(n_0_30));
   INV_X1 i_0_44 (.A(second_operand[14]), .ZN(n_0_31));
   OAI211_X1 i_0_45 (.A(n_0_30), .B(first_operand[13]), .C1(n_0_31), .C2(
      first_operand[14]), .ZN(n_0_32));
   INV_X1 i_0_46 (.A(first_operand[14]), .ZN(n_0_33));
   OAI21_X1 i_0_47 (.A(n_0_32), .B1(second_operand[14]), .B2(n_0_33), .ZN(n_0_34));
   INV_X1 i_0_48 (.A(second_operand[15]), .ZN(n_0_35));
   OAI21_X1 i_0_49 (.A(n_0_34), .B1(first_operand[15]), .B2(n_0_35), .ZN(n_0_36));
   INV_X1 i_0_50 (.A(first_operand[15]), .ZN(n_0_37));
   OAI21_X1 i_0_51 (.A(n_0_36), .B1(second_operand[15]), .B2(n_0_37), .ZN(n_0_38));
   MUX2_X1 i_0_52 (.A(first_operand[13]), .B(second_operand[13]), .S(n_0_38), 
      .Z(n_0_39));
   MUX2_X1 i_0_53 (.A(first_operand[14]), .B(second_operand[14]), .S(n_0_38), 
      .Z(n_0_40));
   MUX2_X1 i_0_54 (.A(first_operand[15]), .B(second_operand[15]), .S(n_0_38), 
      .Z(n_0_41));
   MUX2_X1 i_0_55 (.A(second_operand[13]), .B(first_operand[13]), .S(n_0_38), 
      .Z(n_13));
   MUX2_X1 i_0_56 (.A(second_operand[14]), .B(first_operand[14]), .S(n_0_38), 
      .Z(n_14));
   MUX2_X1 i_0_57 (.A(second_operand[15]), .B(first_operand[15]), .S(n_0_38), 
      .Z(n_15));
endmodule

module Division_CLHA(reset, clk, dividend, divisor, Q, ready, overFlow, 
      divideByZero);
   input reset;
   input clk;
   input [15:0]dividend;
   input [15:0]divisor;
   output [15:0]Q;
   output ready;
   output overFlow;
   output divideByZero;

   wire cla0_n_0;
   wire cla0_n_1;
   wire cla0_n_2;
   wire cla1_n_0;
   wire [15:0]negated_second_operand_number;
   wire [15:0]second_operand_number;
   wire [4:0]number_of_bits_in_dividend;
   wire sign;
   wire n_0_1;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_40;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_97;
   wire n_0_98;
   wire n_0_108;
   wire n_0_109;
   wire n_0_112;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_124;
   wire n_0_125;
   wire n_0_133;
   wire n_0_149;
   wire n_0_150;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_174;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_317;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_337;
   wire n_0_0;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_2;
   wire n_0_366;
   wire n_0_3;
   wire n_0_369;
   wire n_0_370;
   wire n_0_4;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_5;
   wire n_0_379;
   wire n_0_380;
   wire n_0_24;
   wire n_0_385;
   wire n_0_396;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_419;
   wire n_0_420;
   wire n_0_421;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_41;
   wire n_0_428;
   wire n_0_56;
   wire n_0_68;
   wire n_0_69;
   wire n_0_76;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_451;
   wire n_0_453;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_84;
   wire n_0_85;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_110;
   wire n_0_111;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_122;
   wire n_0_123;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_173;
   wire n_0_175;
   wire n_0_226;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_360;
   wire n_0_364;
   wire n_0_365;
   wire n_0_367;
   wire n_0_368;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_377;
   wire n_0_378;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_0_425;
   wire n_0_426;
   wire n_0_427;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_436;
   wire n_0_437;
   wire n_0_438;
   wire n_0_439;
   wire n_0_440;
   wire n_0_441;
   wire n_0_442;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_449;
   wire n_0_450;
   wire n_0_452;
   wire n_0_454;
   wire n_0_455;

   INV_X1 cla0_i_5 (.A(divisor[13]), .ZN(cla0_n_0));
   INV_X1 cla0_i_6 (.A(divisor[14]), .ZN(cla0_n_1));
   INV_X1 cla0_i_7 (.A(divisor[15]), .ZN(cla0_n_2));
   INV_X1 cla1_i_5 (.A(dividend[13]), .ZN(cla1_n_0));
   DFF_X1 divideByZero_reg (.D(n_116), .CK(n_6), .Q(divideByZero), .QN());
   DFF_X1 overFlow_reg (.D(n_128), .CK(clk), .Q(overFlow), .QN());
   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_85), .SE(1'b0), .GCK(n_0));
   DFF_X1 \Q_reg[14]  (.D(n_113), .CK(n_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_49), .CK(n_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_48), .CK(n_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_47), .CK(n_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_46), .CK(n_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_45), .CK(n_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_44), .CK(n_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_43), .CK(n_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_42), .CK(n_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_41), .CK(n_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_40), .CK(n_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_39), .CK(n_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_38), .CK(n_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_37), .CK(n_0), .Q(Q[0]), .QN());
   CLKGATETST_X1 clk_gate_A_reg (.CK(clk), .E(n_84), .SE(1'b0), .GCK(n_1));
   DFF_X1 \A_reg[31]  (.D(n_82), .CK(n_1), .Q(n_4), .QN());
   DFF_X1 \A_reg[30]  (.D(n_81), .CK(n_1), .Q(n_5), .QN());
   DFF_X1 \A_reg[29]  (.D(n_80), .CK(n_1), .Q(n_7), .QN());
   DFF_X1 \A_reg[28]  (.D(n_79), .CK(n_1), .Q(n_8), .QN());
   DFF_X1 \A_reg[27]  (.D(n_78), .CK(n_1), .Q(n_9), .QN());
   DFF_X1 \A_reg[26]  (.D(n_77), .CK(n_1), .Q(n_10), .QN());
   DFF_X1 \A_reg[25]  (.D(n_76), .CK(n_1), .Q(n_11), .QN());
   DFF_X1 \A_reg[24]  (.D(n_75), .CK(n_1), .Q(n_12), .QN());
   DFF_X1 \A_reg[23]  (.D(n_74), .CK(n_1), .Q(n_13), .QN());
   DFF_X1 \A_reg[22]  (.D(n_73), .CK(n_1), .Q(n_14), .QN());
   DFF_X1 \A_reg[21]  (.D(n_72), .CK(n_1), .Q(n_15), .QN());
   DFF_X1 \A_reg[20]  (.D(n_71), .CK(n_1), .Q(n_16), .QN());
   DFF_X1 \A_reg[19]  (.D(n_70), .CK(n_1), .Q(n_17), .QN());
   DFF_X1 \A_reg[18]  (.D(n_69), .CK(n_1), .Q(n_18), .QN());
   DFF_X1 \A_reg[17]  (.D(n_68), .CK(n_1), .Q(n_19), .QN());
   DFF_X1 \A_reg[16]  (.D(n_67), .CK(n_1), .Q(n_20), .QN());
   CLKGATETST_X1 clk_gate_A_reg__15 (.CK(clk), .E(n_83), .SE(1'b0), .GCK(n_2));
   DFF_X1 \A_reg[15]  (.D(n_66), .CK(n_2), .Q(n_21), .QN());
   DFF_X1 \A_reg[14]  (.D(n_127), .CK(n_2), .Q(n_22), .QN());
   DFF_X1 \A_reg[13]  (.D(n_65), .CK(n_2), .Q(n_23), .QN());
   DFF_X1 \A_reg[12]  (.D(n_64), .CK(n_2), .Q(n_24), .QN());
   DFF_X1 \A_reg[11]  (.D(n_63), .CK(n_2), .Q(n_25), .QN());
   DFF_X1 \A_reg[10]  (.D(n_62), .CK(n_2), .Q(n_26), .QN());
   DFF_X1 \A_reg[9]  (.D(n_61), .CK(n_2), .Q(n_27), .QN());
   DFF_X1 \A_reg[8]  (.D(n_60), .CK(n_2), .Q(n_28), .QN());
   DFF_X1 \A_reg[7]  (.D(n_126), .CK(n_2), .Q(n_29), .QN());
   DFF_X1 \A_reg[6]  (.D(n_59), .CK(n_2), .Q(n_30), .QN());
   DFF_X1 \A_reg[5]  (.D(n_58), .CK(n_2), .Q(n_31), .QN());
   DFF_X1 \A_reg[4]  (.D(n_124), .CK(n_2), .Q(n_32), .QN());
   DFF_X1 \A_reg[3]  (.D(n_57), .CK(n_2), .Q(n_33), .QN());
   DFF_X1 \A_reg[2]  (.D(n_56), .CK(n_2), .Q(n_34), .QN());
   DFF_X1 \A_reg[1]  (.D(n_55), .CK(n_2), .Q(n_35), .QN());
   DFF_X1 \A_reg[0]  (.D(n_54), .CK(n_2), .Q(n_36), .QN());
   DFF_X1 \negated_second_operand_number_reg[15]  (.D(n_104), .CK(n_6), .Q(
      negated_second_operand_number[15]), .QN());
   DFF_X1 \negated_second_operand_number_reg[14]  (.D(n_103), .CK(n_6), .Q(
      negated_second_operand_number[14]), .QN());
   DFF_X1 \negated_second_operand_number_reg[13]  (.D(n_102), .CK(n_6), .Q(
      negated_second_operand_number[13]), .QN());
   DFF_X1 \negated_second_operand_number_reg[12]  (.D(n_101), .CK(n_6), .Q(
      negated_second_operand_number[12]), .QN());
   DFF_X1 \negated_second_operand_number_reg[11]  (.D(n_100), .CK(n_6), .Q(
      negated_second_operand_number[11]), .QN());
   DFF_X1 \negated_second_operand_number_reg[10]  (.D(n_99), .CK(n_6), .Q(
      negated_second_operand_number[10]), .QN());
   DFF_X1 \negated_second_operand_number_reg[9]  (.D(n_98), .CK(n_6), .Q(
      negated_second_operand_number[9]), .QN());
   DFF_X1 \negated_second_operand_number_reg[8]  (.D(n_97), .CK(n_6), .Q(
      negated_second_operand_number[8]), .QN());
   DFF_X1 \negated_second_operand_number_reg[7]  (.D(n_96), .CK(n_6), .Q(
      negated_second_operand_number[7]), .QN());
   DFF_X1 \negated_second_operand_number_reg[6]  (.D(n_95), .CK(n_6), .Q(
      negated_second_operand_number[6]), .QN());
   DFF_X1 \negated_second_operand_number_reg[5]  (.D(n_94), .CK(n_6), .Q(
      negated_second_operand_number[5]), .QN());
   DFF_X1 \negated_second_operand_number_reg[4]  (.D(n_93), .CK(n_6), .Q(
      negated_second_operand_number[4]), .QN());
   DFF_X1 \negated_second_operand_number_reg[3]  (.D(n_92), .CK(n_6), .Q(
      negated_second_operand_number[3]), .QN());
   DFF_X1 \negated_second_operand_number_reg[2]  (.D(n_91), .CK(n_6), .Q(
      negated_second_operand_number[2]), .QN());
   DFF_X1 \negated_second_operand_number_reg[1]  (.D(n_90), .CK(n_6), .Q(
      negated_second_operand_number[1]), .QN());
   DFF_X1 \second_operand_number_reg[15]  (.D(n_123), .CK(n_6), .Q(
      second_operand_number[15]), .QN());
   DFF_X1 \second_operand_number_reg[14]  (.D(n_111), .CK(n_6), .Q(
      second_operand_number[14]), .QN());
   DFF_X1 \second_operand_number_reg[13]  (.D(n_122), .CK(n_6), .Q(
      second_operand_number[13]), .QN());
   DFF_X1 \second_operand_number_reg[12]  (.D(n_121), .CK(n_6), .Q(
      second_operand_number[12]), .QN());
   DFF_X1 \second_operand_number_reg[11]  (.D(n_120), .CK(n_6), .Q(
      second_operand_number[11]), .QN());
   DFF_X1 \second_operand_number_reg[10]  (.D(n_119), .CK(n_6), .Q(
      second_operand_number[10]), .QN());
   DFF_X1 \second_operand_number_reg[9]  (.D(n_118), .CK(n_6), .Q(
      second_operand_number[9]), .QN());
   DFF_X1 \second_operand_number_reg[8]  (.D(n_117), .CK(n_6), .Q(
      second_operand_number[8]), .QN());
   DFF_X1 \second_operand_number_reg[7]  (.D(n_110), .CK(n_6), .Q(
      second_operand_number[7]), .QN());
   DFF_X1 \second_operand_number_reg[6]  (.D(n_109), .CK(n_6), .Q(
      second_operand_number[6]), .QN());
   DFF_X1 \second_operand_number_reg[5]  (.D(n_108), .CK(n_6), .Q(
      second_operand_number[5]), .QN());
   DFF_X1 \second_operand_number_reg[4]  (.D(n_107), .CK(n_6), .Q(
      second_operand_number[4]), .QN());
   DFF_X1 \second_operand_number_reg[3]  (.D(n_106), .CK(n_6), .Q(
      second_operand_number[3]), .QN());
   DFF_X1 \second_operand_number_reg[2]  (.D(n_105), .CK(n_6), .Q(
      second_operand_number[2]), .QN());
   DFF_X1 \second_operand_number_reg[1]  (.D(n_89), .CK(n_6), .Q(
      second_operand_number[1]), .QN());
   DFF_X1 ready_reg (.D(n_129), .CK(clk), .Q(ready), .QN());
   CLKGATETST_X1 clk_gate_number_of_bits_in_dividend_reg (.CK(clk), .E(n_125), 
      .SE(1'b0), .GCK(n_3));
   DFF_X1 \number_of_bits_in_dividend_reg[4]  (.D(n_115), .CK(n_3), .Q(
      number_of_bits_in_dividend[4]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[3]  (.D(n_114), .CK(n_3), .Q(
      number_of_bits_in_dividend[3]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[2]  (.D(n_52), .CK(n_3), .Q(
      number_of_bits_in_dividend[2]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[1]  (.D(n_112), .CK(n_3), .Q(
      number_of_bits_in_dividend[1]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[0]  (.D(n_51), .CK(n_3), .Q(
      number_of_bits_in_dividend[0]), .QN());
   DFF_X1 sign_reg (.D(n_50), .CK(n_6), .Q(sign), .QN());
   CLKGATETST_X1 clk_gate_divideByZero_reg (.CK(clk), .E(reset), .SE(1'b0), 
      .GCK(n_6));
   DFF_X1 \negated_second_operand_number_reg[0]  (.D(n_88), .CK(n_6), .Q(
      negated_second_operand_number[0]), .QN());
   AND2_X1 i_0_0 (.A1(n_113), .A2(n_36), .ZN(n_37));
   NOR2_X1 i_0_1 (.A1(reset), .A2(n_0_16), .ZN(n_38));
   NOR2_X1 i_0_2 (.A1(reset), .A2(n_0_18), .ZN(n_39));
   NOR2_X1 i_0_3 (.A1(reset), .A2(n_0_22), .ZN(n_40));
   NOR2_X1 i_0_4 (.A1(reset), .A2(n_0_333), .ZN(n_41));
   NOR2_X1 i_0_5 (.A1(reset), .A2(n_0_28), .ZN(n_42));
   AND2_X1 i_0_6 (.A1(n_113), .A2(n_0_35), .ZN(n_43));
   NOR2_X1 i_0_7 (.A1(reset), .A2(n_0_393), .ZN(n_44));
   NOR2_X1 i_0_8 (.A1(reset), .A2(n_0_42), .ZN(n_45));
   NOR2_X1 i_0_9 (.A1(reset), .A2(n_0_49), .ZN(n_46));
   NOR2_X1 i_0_10 (.A1(reset), .A2(n_0_52), .ZN(n_47));
   NOR2_X1 i_0_11 (.A1(reset), .A2(n_0_62), .ZN(n_48));
   NOR2_X1 i_0_12 (.A1(reset), .A2(n_0_71), .ZN(n_49));
   XNOR2_X1 i_0_13 (.A(n_0_451), .B(dividend[12]), .ZN(n_50));
   NAND2_X1 i_0_14 (.A1(n_113), .A2(number_of_bits_in_dividend[0]), .ZN(n_51));
   NAND3_X1 i_0_15 (.A1(n_113), .A2(n_0_80), .A3(n_0_1), .ZN(n_52));
   OAI21_X1 i_0_16 (.A(number_of_bits_in_dividend[2]), .B1(
      number_of_bits_in_dividend[1]), .B2(number_of_bits_in_dividend[0]), 
      .ZN(n_0_1));
   NAND2_X1 i_0_17 (.A1(n_113), .A2(n_0_317), .ZN(n_53));
   OAI221_X1 i_0_18 (.A(n_0_14), .B1(n_0_10), .B2(n_0_229), .C1(n_0_6), .C2(
      n_0_230), .ZN(n_54));
   XNOR2_X1 i_0_19 (.A(negated_second_operand_number[15]), .B(n_0_7), .ZN(n_0_6));
   OAI21_X1 i_0_20 (.A(n_0_8), .B1(negated_second_operand_number[14]), .B2(n_5), 
      .ZN(n_0_7));
   NAND2_X1 i_0_21 (.A1(n_0_234), .A2(n_0_9), .ZN(n_0_8));
   NAND2_X1 i_0_22 (.A1(n_5), .A2(negated_second_operand_number[14]), .ZN(n_0_9));
   XNOR2_X1 i_0_23 (.A(second_operand_number[15]), .B(n_0_11), .ZN(n_0_10));
   OAI21_X1 i_0_24 (.A(n_0_12), .B1(n_0_274), .B2(n_0_13), .ZN(n_0_11));
   NAND2_X1 i_0_25 (.A1(n_5), .A2(second_operand_number[14]), .ZN(n_0_12));
   NOR2_X1 i_0_26 (.A1(n_5), .A2(second_operand_number[14]), .ZN(n_0_13));
   NAND2_X1 i_0_27 (.A1(n_36), .A2(n_0_434), .ZN(n_0_14));
   OAI21_X1 i_0_28 (.A(n_0_15), .B1(n_0_319), .B2(n_0_16), .ZN(n_55));
   NAND2_X1 i_0_29 (.A1(n_36), .A2(n_0_173), .ZN(n_0_15));
   XOR2_X1 i_0_30 (.A(n_35), .B(n_0_20), .Z(n_0_16));
   OAI21_X1 i_0_31 (.A(n_0_17), .B1(n_0_319), .B2(n_0_18), .ZN(n_56));
   NAND2_X1 i_0_32 (.A1(n_35), .A2(n_0_173), .ZN(n_0_17));
   XOR2_X1 i_0_33 (.A(n_34), .B(n_0_19), .Z(n_0_18));
   NAND2_X1 i_0_34 (.A1(n_0_336), .A2(sign), .ZN(n_0_19));
   NAND2_X1 i_0_35 (.A1(n_36), .A2(sign), .ZN(n_0_20));
   OAI21_X1 i_0_36 (.A(n_0_21), .B1(n_0_22), .B2(n_0_319), .ZN(n_57));
   NAND2_X1 i_0_37 (.A1(n_34), .A2(n_0_173), .ZN(n_0_21));
   XOR2_X1 i_0_38 (.A(n_33), .B(n_0_23), .Z(n_0_22));
   OAI21_X1 i_0_39 (.A(sign), .B1(n_0_336), .B2(n_34), .ZN(n_0_23));
   OAI221_X1 i_0_40 (.A(n_0_30), .B1(n_0_394), .B2(n_0_373), .C1(n_0_28), 
      .C2(n_0_319), .ZN(n_58));
   XOR2_X1 i_0_41 (.A(n_31), .B(n_0_29), .Z(n_0_28));
   NAND2_X1 i_0_42 (.A1(n_0_388), .A2(sign), .ZN(n_0_29));
   AOI21_X1 i_0_43 (.A(n_0_31), .B1(n_0_173), .B2(n_32), .ZN(n_0_30));
   NOR3_X1 i_0_44 (.A1(n_0_365), .A2(n_0_270), .A3(n_0_412), .ZN(n_0_31));
   OAI221_X1 i_0_45 (.A(n_0_34), .B1(n_0_32), .B2(n_0_360), .C1(n_0_383), 
      .C2(n_0_394), .ZN(n_59));
   AOI21_X1 i_0_46 (.A(n_0_33), .B1(n_0_384), .B2(n_0_386), .ZN(n_0_32));
   NOR3_X1 i_0_47 (.A1(n_0_270), .A2(n_0_386), .A3(n_0_373), .ZN(n_0_33));
   AOI22_X1 i_0_48 (.A1(n_0_35), .A2(n_0_434), .B1(n_0_173), .B2(n_31), .ZN(
      n_0_34));
   XNOR2_X1 i_0_49 (.A(n_30), .B(n_0_389), .ZN(n_0_35));
   OAI221_X1 i_0_50 (.A(n_0_40), .B1(n_0_398), .B2(n_0_47), .C1(n_0_42), 
      .C2(n_0_319), .ZN(n_60));
   AOI222_X1 i_0_51 (.A1(n_0_175), .A2(n_0_405), .B1(n_0_381), .B2(n_0_387), 
      .C1(n_29), .C2(n_0_173), .ZN(n_0_40));
   XOR2_X1 i_0_52 (.A(n_28), .B(n_0_43), .Z(n_0_42));
   NAND2_X1 i_0_53 (.A1(n_0_75), .A2(sign), .ZN(n_0_43));
   OAI21_X1 i_0_54 (.A(n_0_44), .B1(n_0_49), .B2(n_0_319), .ZN(n_61));
   AOI21_X1 i_0_55 (.A(n_0_45), .B1(n_0_55), .B2(n_0_364), .ZN(n_0_44));
   OAI221_X1 i_0_56 (.A(n_0_46), .B1(n_0_394), .B2(n_0_417), .C1(n_0_47), 
      .C2(n_0_412), .ZN(n_0_45));
   NAND2_X1 i_0_57 (.A1(n_28), .A2(n_0_173), .ZN(n_0_46));
   AOI21_X1 i_0_58 (.A(n_0_48), .B1(n_0_60), .B2(n_0_271), .ZN(n_0_47));
   NOR2_X1 i_0_59 (.A1(n_0_378), .A2(n_0_383), .ZN(n_0_48));
   XOR2_X1 i_0_60 (.A(n_27), .B(n_0_50), .Z(n_0_49));
   NAND2_X1 i_0_61 (.A1(n_0_74), .A2(sign), .ZN(n_0_50));
   OAI211_X1 i_0_62 (.A(n_0_51), .B(n_0_54), .C1(n_0_319), .C2(n_0_52), .ZN(n_62));
   AOI222_X1 i_0_63 (.A1(n_0_55), .A2(n_0_387), .B1(n_0_410), .B2(n_0_175), 
      .C1(n_27), .C2(n_0_173), .ZN(n_0_51));
   XOR2_X1 i_0_64 (.A(n_26), .B(n_0_53), .Z(n_0_52));
   OAI21_X1 i_0_65 (.A(sign), .B1(n_0_74), .B2(n_27), .ZN(n_0_53));
   NAND2_X1 i_0_66 (.A1(n_0_59), .A2(n_0_364), .ZN(n_0_54));
   OAI22_X1 i_0_67 (.A1(n_0_377), .A2(n_0_67), .B1(n_0_378), .B2(n_0_371), 
      .ZN(n_0_55));
   OAI221_X1 i_0_68 (.A(n_0_57), .B1(n_0_62), .B2(n_0_319), .C1(n_0_398), 
      .C2(n_0_66), .ZN(n_63));
   AOI221_X1 i_0_69 (.A(n_0_58), .B1(n_0_173), .B2(n_26), .C1(n_0_59), .C2(
      n_0_387), .ZN(n_0_57));
   NOR2_X1 i_0_70 (.A1(n_0_427), .A2(n_0_394), .ZN(n_0_58));
   MUX2_X1 i_0_71 (.A(n_0_60), .B(n_0_83), .S(n_0_271), .Z(n_0_59));
   OAI21_X1 i_0_72 (.A(n_0_61), .B1(n_0_308), .B2(n_0_365), .ZN(n_0_60));
   NAND2_X1 i_0_73 (.A1(n_0_308), .A2(n_0_405), .ZN(n_0_61));
   XOR2_X1 i_0_74 (.A(n_25), .B(n_0_63), .Z(n_0_62));
   NAND2_X1 i_0_75 (.A1(n_0_73), .A2(sign), .ZN(n_0_63));
   OAI211_X1 i_0_76 (.A(n_0_64), .B(n_0_70), .C1(n_0_71), .C2(n_0_319), .ZN(n_64));
   AOI221_X1 i_0_77 (.A(n_0_65), .B1(n_0_403), .B2(n_0_175), .C1(n_25), .C2(
      n_0_173), .ZN(n_0_64));
   NOR2_X1 i_0_78 (.A1(n_0_66), .A2(n_0_412), .ZN(n_0_65));
   MUX2_X1 i_0_79 (.A(n_0_67), .B(n_0_425), .S(n_0_271), .Z(n_0_66));
   MUX2_X1 i_0_80 (.A(n_0_373), .B(n_0_417), .S(n_0_308), .Z(n_0_67));
   NAND2_X1 i_0_81 (.A1(n_0_82), .A2(n_0_364), .ZN(n_0_70));
   XOR2_X1 i_0_82 (.A(n_24), .B(n_0_72), .Z(n_0_71));
   OAI21_X1 i_0_83 (.A(sign), .B1(n_0_73), .B2(n_25), .ZN(n_0_72));
   OR3_X1 i_0_84 (.A1(n_0_74), .A2(n_27), .A3(n_26), .ZN(n_0_73));
   OR2_X1 i_0_85 (.A1(n_0_75), .A2(n_28), .ZN(n_0_74));
   OR2_X1 i_0_86 (.A1(n_0_391), .A2(n_29), .ZN(n_0_75));
   OAI21_X1 i_0_87 (.A(n_0_81), .B1(n_0_413), .B2(n_0_398), .ZN(n_65));
   AOI21_X1 i_0_88 (.A(n_0_87), .B1(n_0_82), .B2(n_0_387), .ZN(n_0_81));
   MUX2_X1 i_0_89 (.A(n_0_83), .B(n_0_401), .S(n_0_271), .Z(n_0_82));
   AOI21_X1 i_0_90 (.A(n_0_86), .B1(n_0_383), .B2(n_0_309), .ZN(n_0_83));
   NOR2_X1 i_0_91 (.A1(n_0_410), .A2(n_0_309), .ZN(n_0_86));
   OAI21_X1 i_0_92 (.A(n_0_88), .B1(n_0_415), .B2(n_0_394), .ZN(n_0_87));
   AOI21_X1 i_0_93 (.A(n_0_434), .B1(n_0_173), .B2(n_24), .ZN(n_0_88));
   OAI221_X1 i_0_94 (.A(n_0_97), .B1(n_0_399), .B2(n_0_412), .C1(n_0_119), 
      .C2(n_0_398), .ZN(n_66));
   AOI21_X1 i_0_95 (.A(n_0_98), .B1(n_0_173), .B2(n_22), .ZN(n_0_97));
   NOR2_X1 i_0_96 (.A1(n_0_124), .A2(n_0_394), .ZN(n_0_98));
   OAI221_X1 i_0_97 (.A(n_0_133), .B1(n_0_108), .B2(n_0_398), .C1(n_0_412), 
      .C2(n_0_119), .ZN(n_67));
   OAI21_X1 i_0_98 (.A(n_0_112), .B1(n_0_109), .B2(n_0_377), .ZN(n_0_108));
   MUX2_X1 i_0_99 (.A(n_0_403), .B(n_0_149), .S(n_0_308), .Z(n_0_109));
   NAND2_X1 i_0_100 (.A1(n_0_377), .A2(n_0_407), .ZN(n_0_112));
   AOI21_X1 i_0_101 (.A(n_0_120), .B1(n_0_414), .B2(n_0_377), .ZN(n_0_119));
   OAI22_X1 i_0_102 (.A1(n_0_270), .A2(n_0_124), .B1(n_0_427), .B2(n_0_121), 
      .ZN(n_0_120));
   NAND2_X1 i_0_103 (.A1(n_0_271), .A2(n_0_309), .ZN(n_0_121));
   XOR2_X1 i_0_104 (.A(dividend[11]), .B(n_0_125), .Z(n_0_124));
   NAND2_X1 i_0_105 (.A1(n_0_150), .A2(dividend[12]), .ZN(n_0_125));
   AOI222_X1 i_0_106 (.A1(n_21), .A2(n_0_173), .B1(n_0_149), .B2(n_0_175), 
      .C1(n_0_320), .C2(n_19), .ZN(n_0_133));
   NOR3_X1 i_0_107 (.A1(n_0_438), .A2(n_0_150), .A3(dividend[11]), .ZN(n_0_149));
   OR2_X1 i_0_108 (.A1(n_0_430), .A2(dividend[10]), .ZN(n_0_150));
   INV_X1 i_0_109 (.A(n_0_158), .ZN(n_68));
   AOI22_X1 i_0_110 (.A1(n_18), .A2(n_0_320), .B1(n_0_159), .B2(n_0_173), 
      .ZN(n_0_158));
   XOR2_X1 i_0_111 (.A(n_20), .B(negated_second_operand_number[0]), .Z(n_0_159));
   INV_X1 i_0_112 (.A(n_0_160), .ZN(n_69));
   AOI22_X1 i_0_113 (.A1(n_0_161), .A2(n_0_173), .B1(n_17), .B2(n_0_320), 
      .ZN(n_0_160));
   XNOR2_X1 i_0_114 (.A(n_0_163), .B(n_0_162), .ZN(n_0_161));
   XNOR2_X1 i_0_115 (.A(n_19), .B(n_0_445), .ZN(n_0_162));
   MUX2_X1 i_0_116 (.A(negated_second_operand_number[1]), .B(
      second_operand_number[1]), .S(n_4), .Z(n_0_163));
   INV_X1 i_0_117 (.A(n_0_164), .ZN(n_70));
   AOI22_X1 i_0_118 (.A1(n_0_165), .A2(n_0_173), .B1(n_16), .B2(n_0_320), 
      .ZN(n_0_164));
   XNOR2_X1 i_0_119 (.A(n_18), .B(n_0_166), .ZN(n_0_165));
   OAI21_X1 i_0_120 (.A(n_0_167), .B1(n_0_168), .B2(n_4), .ZN(n_0_166));
   NAND2_X1 i_0_121 (.A1(n_4), .A2(n_0_169), .ZN(n_0_167));
   XOR2_X1 i_0_122 (.A(negated_second_operand_number[2]), .B(n_0_442), .Z(
      n_0_168));
   XNOR2_X1 i_0_123 (.A(second_operand_number[2]), .B(n_0_454), .ZN(n_0_169));
   INV_X1 i_0_124 (.A(n_0_170), .ZN(n_71));
   AOI22_X1 i_0_125 (.A1(n_0_171), .A2(n_0_173), .B1(n_15), .B2(n_0_320), 
      .ZN(n_0_170));
   XOR2_X1 i_0_126 (.A(n_17), .B(n_0_172), .Z(n_0_171));
   OAI21_X1 i_0_127 (.A(n_0_174), .B1(n_0_439), .B2(n_4), .ZN(n_0_172));
   NAND2_X1 i_0_128 (.A1(n_0_449), .A2(n_4), .ZN(n_0_174));
   OAI221_X1 i_0_129 (.A(n_0_180), .B1(n_0_178), .B2(n_0_229), .C1(n_0_176), 
      .C2(n_0_230), .ZN(n_72));
   XNOR2_X1 i_0_130 (.A(n_0_264), .B(n_0_177), .ZN(n_0_176));
   XNOR2_X1 i_0_131 (.A(n_16), .B(negated_second_operand_number[4]), .ZN(n_0_177));
   XNOR2_X1 i_0_132 (.A(n_0_304), .B(n_0_179), .ZN(n_0_178));
   XNOR2_X1 i_0_133 (.A(n_16), .B(second_operand_number[4]), .ZN(n_0_179));
   NAND2_X1 i_0_134 (.A1(n_14), .A2(n_0_320), .ZN(n_0_180));
   OAI221_X1 i_0_135 (.A(n_0_185), .B1(n_0_183), .B2(n_0_230), .C1(n_0_181), 
      .C2(n_0_229), .ZN(n_73));
   XNOR2_X1 i_0_136 (.A(n_0_301), .B(n_0_182), .ZN(n_0_181));
   XNOR2_X1 i_0_137 (.A(n_15), .B(second_operand_number[5]), .ZN(n_0_182));
   XNOR2_X1 i_0_138 (.A(n_0_261), .B(n_0_184), .ZN(n_0_183));
   XOR2_X1 i_0_139 (.A(n_15), .B(negated_second_operand_number[5]), .Z(n_0_184));
   NAND2_X1 i_0_140 (.A1(n_13), .A2(n_0_320), .ZN(n_0_185));
   OAI221_X1 i_0_141 (.A(n_0_190), .B1(n_0_188), .B2(n_0_229), .C1(n_0_186), 
      .C2(n_0_230), .ZN(n_74));
   XNOR2_X1 i_0_142 (.A(n_0_257), .B(n_0_187), .ZN(n_0_186));
   XNOR2_X1 i_0_143 (.A(n_14), .B(negated_second_operand_number[6]), .ZN(n_0_187));
   XNOR2_X1 i_0_144 (.A(n_0_298), .B(n_0_189), .ZN(n_0_188));
   XOR2_X1 i_0_145 (.A(n_14), .B(second_operand_number[6]), .Z(n_0_189));
   NAND2_X1 i_0_146 (.A1(n_12), .A2(n_0_320), .ZN(n_0_190));
   OAI221_X1 i_0_147 (.A(n_0_191), .B1(n_0_230), .B2(n_0_194), .C1(n_0_192), 
      .C2(n_0_229), .ZN(n_75));
   NAND2_X1 i_0_148 (.A1(n_11), .A2(n_0_320), .ZN(n_0_191));
   XNOR2_X1 i_0_149 (.A(n_0_295), .B(n_0_193), .ZN(n_0_192));
   XOR2_X1 i_0_150 (.A(n_13), .B(second_operand_number[7]), .Z(n_0_193));
   XNOR2_X1 i_0_151 (.A(n_0_255), .B(n_0_195), .ZN(n_0_194));
   XOR2_X1 i_0_152 (.A(n_13), .B(negated_second_operand_number[7]), .Z(n_0_195));
   INV_X1 i_0_153 (.A(n_0_196), .ZN(n_76));
   AOI22_X1 i_0_154 (.A1(n_0_197), .A2(n_0_173), .B1(n_10), .B2(n_0_320), 
      .ZN(n_0_196));
   XNOR2_X1 i_0_155 (.A(n_12), .B(n_0_198), .ZN(n_0_197));
   AOI21_X1 i_0_156 (.A(n_0_199), .B1(n_0_201), .B2(n_4), .ZN(n_0_198));
   NOR2_X1 i_0_157 (.A1(n_4), .A2(n_0_200), .ZN(n_0_199));
   XNOR2_X1 i_0_158 (.A(negated_second_operand_number[8]), .B(n_0_252), .ZN(
      n_0_200));
   XNOR2_X1 i_0_159 (.A(second_operand_number[8]), .B(n_0_291), .ZN(n_0_201));
   OAI221_X1 i_0_160 (.A(n_0_206), .B1(n_0_229), .B2(n_0_202), .C1(n_0_230), 
      .C2(n_0_204), .ZN(n_77));
   XNOR2_X1 i_0_161 (.A(n_0_289), .B(n_0_203), .ZN(n_0_202));
   XOR2_X1 i_0_162 (.A(n_11), .B(second_operand_number[9]), .Z(n_0_203));
   XNOR2_X1 i_0_163 (.A(n_0_249), .B(n_0_205), .ZN(n_0_204));
   XNOR2_X1 i_0_164 (.A(n_11), .B(negated_second_operand_number[9]), .ZN(n_0_205));
   NAND2_X1 i_0_165 (.A1(n_9), .A2(n_0_320), .ZN(n_0_206));
   OAI221_X1 i_0_166 (.A(n_0_211), .B1(n_0_207), .B2(n_0_230), .C1(n_0_229), 
      .C2(n_0_209), .ZN(n_78));
   XNOR2_X1 i_0_167 (.A(n_0_245), .B(n_0_208), .ZN(n_0_207));
   XNOR2_X1 i_0_168 (.A(n_10), .B(negated_second_operand_number[10]), .ZN(
      n_0_208));
   XNOR2_X1 i_0_169 (.A(n_0_285), .B(n_0_210), .ZN(n_0_209));
   XNOR2_X1 i_0_170 (.A(n_10), .B(second_operand_number[10]), .ZN(n_0_210));
   NAND2_X1 i_0_171 (.A1(n_8), .A2(n_0_320), .ZN(n_0_211));
   INV_X1 i_0_172 (.A(n_0_212), .ZN(n_79));
   AOI22_X1 i_0_173 (.A1(n_0_213), .A2(n_0_173), .B1(n_7), .B2(n_0_320), 
      .ZN(n_0_212));
   XNOR2_X1 i_0_174 (.A(n_9), .B(n_0_214), .ZN(n_0_213));
   AOI21_X1 i_0_175 (.A(n_0_215), .B1(n_0_217), .B2(n_4), .ZN(n_0_214));
   NOR2_X1 i_0_176 (.A1(n_4), .A2(n_0_216), .ZN(n_0_215));
   XNOR2_X1 i_0_177 (.A(negated_second_operand_number[11]), .B(n_0_243), 
      .ZN(n_0_216));
   XOR2_X1 i_0_178 (.A(second_operand_number[11]), .B(n_0_283), .Z(n_0_217));
   OAI221_X1 i_0_179 (.A(n_0_218), .B1(n_0_219), .B2(n_0_230), .C1(n_0_221), 
      .C2(n_0_229), .ZN(n_80));
   NAND2_X1 i_0_180 (.A1(n_5), .A2(n_0_320), .ZN(n_0_218));
   XNOR2_X1 i_0_181 (.A(n_0_240), .B(n_0_220), .ZN(n_0_219));
   XNOR2_X1 i_0_182 (.A(n_8), .B(negated_second_operand_number[12]), .ZN(n_0_220));
   XNOR2_X1 i_0_183 (.A(n_0_279), .B(n_0_222), .ZN(n_0_221));
   XNOR2_X1 i_0_184 (.A(n_8), .B(second_operand_number[12]), .ZN(n_0_222));
   OAI22_X1 i_0_185 (.A1(n_0_223), .A2(n_0_446), .B1(n_0_227), .B2(n_0_230), 
      .ZN(n_81));
   AOI21_X1 i_0_186 (.A(n_0_320), .B1(n_0_224), .B2(n_0_173), .ZN(n_0_223));
   XNOR2_X1 i_0_187 (.A(n_0_277), .B(n_0_225), .ZN(n_0_224));
   XNOR2_X1 i_0_188 (.A(n_7), .B(second_operand_number[13]), .ZN(n_0_225));
   XNOR2_X1 i_0_189 (.A(n_0_237), .B(n_0_228), .ZN(n_0_227));
   XOR2_X1 i_0_190 (.A(n_7), .B(negated_second_operand_number[13]), .Z(n_0_228));
   NOR3_X1 i_0_191 (.A1(reset), .A2(n_0_328), .A3(n_0_231), .ZN(n_82));
   NAND2_X1 i_0_192 (.A1(n_4), .A2(n_0_173), .ZN(n_0_229));
   NAND2_X1 i_0_193 (.A1(n_0_173), .A2(n_0_446), .ZN(n_0_230));
   XNOR2_X1 i_0_194 (.A(n_5), .B(n_0_232), .ZN(n_0_231));
   OAI21_X1 i_0_195 (.A(n_0_272), .B1(n_0_233), .B2(n_4), .ZN(n_0_232));
   XOR2_X1 i_0_196 (.A(negated_second_operand_number[14]), .B(n_0_234), .Z(
      n_0_233));
   OAI21_X1 i_0_197 (.A(n_0_235), .B1(negated_second_operand_number[13]), 
      .B2(n_7), .ZN(n_0_234));
   INV_X1 i_0_198 (.A(n_0_236), .ZN(n_0_235));
   AOI21_X1 i_0_199 (.A(n_0_237), .B1(negated_second_operand_number[13]), 
      .B2(n_7), .ZN(n_0_236));
   OAI21_X1 i_0_200 (.A(n_0_239), .B1(n_0_240), .B2(n_0_238), .ZN(n_0_237));
   NOR2_X1 i_0_201 (.A1(n_8), .A2(negated_second_operand_number[12]), .ZN(
      n_0_238));
   NAND2_X1 i_0_202 (.A1(n_8), .A2(negated_second_operand_number[12]), .ZN(
      n_0_239));
   OAI21_X1 i_0_203 (.A(n_0_241), .B1(negated_second_operand_number[11]), 
      .B2(n_9), .ZN(n_0_240));
   INV_X1 i_0_204 (.A(n_0_242), .ZN(n_0_241));
   AOI21_X1 i_0_205 (.A(n_0_243), .B1(negated_second_operand_number[11]), 
      .B2(n_9), .ZN(n_0_242));
   AOI21_X1 i_0_206 (.A(n_0_244), .B1(n_0_245), .B2(n_0_248), .ZN(n_0_243));
   NOR2_X1 i_0_207 (.A1(n_10), .A2(negated_second_operand_number[10]), .ZN(
      n_0_244));
   OAI21_X1 i_0_208 (.A(n_0_246), .B1(negated_second_operand_number[9]), 
      .B2(n_11), .ZN(n_0_245));
   NAND2_X1 i_0_209 (.A1(n_0_249), .A2(n_0_247), .ZN(n_0_246));
   NAND2_X1 i_0_210 (.A1(n_11), .A2(negated_second_operand_number[9]), .ZN(
      n_0_247));
   NAND2_X1 i_0_211 (.A1(n_10), .A2(negated_second_operand_number[10]), .ZN(
      n_0_248));
   AOI21_X1 i_0_212 (.A(n_0_250), .B1(negated_second_operand_number[8]), 
      .B2(n_12), .ZN(n_0_249));
   INV_X1 i_0_213 (.A(n_0_251), .ZN(n_0_250));
   OAI21_X1 i_0_214 (.A(n_0_252), .B1(negated_second_operand_number[8]), 
      .B2(n_12), .ZN(n_0_251));
   NOR2_X1 i_0_215 (.A1(n_0_254), .A2(n_0_253), .ZN(n_0_252));
   NOR2_X1 i_0_216 (.A1(n_13), .A2(negated_second_operand_number[7]), .ZN(
      n_0_253));
   AOI21_X1 i_0_217 (.A(n_0_255), .B1(negated_second_operand_number[7]), 
      .B2(n_13), .ZN(n_0_254));
   AOI21_X1 i_0_218 (.A(n_0_256), .B1(n_0_257), .B2(n_0_260), .ZN(n_0_255));
   NOR2_X1 i_0_219 (.A1(n_14), .A2(negated_second_operand_number[6]), .ZN(
      n_0_256));
   OAI21_X1 i_0_220 (.A(n_0_258), .B1(n_0_261), .B2(
      negated_second_operand_number[5]), .ZN(n_0_257));
   INV_X1 i_0_221 (.A(n_0_259), .ZN(n_0_258));
   AOI21_X1 i_0_222 (.A(n_15), .B1(negated_second_operand_number[5]), .B2(
      n_0_261), .ZN(n_0_259));
   NAND2_X1 i_0_223 (.A1(n_14), .A2(negated_second_operand_number[6]), .ZN(
      n_0_260));
   OAI21_X1 i_0_224 (.A(n_0_263), .B1(n_0_264), .B2(n_0_262), .ZN(n_0_261));
   NOR2_X1 i_0_225 (.A1(n_16), .A2(negated_second_operand_number[4]), .ZN(
      n_0_262));
   NAND2_X1 i_0_226 (.A1(n_16), .A2(negated_second_operand_number[4]), .ZN(
      n_0_263));
   OAI21_X1 i_0_227 (.A(n_0_265), .B1(negated_second_operand_number[3]), 
      .B2(n_17), .ZN(n_0_264));
   NAND2_X1 i_0_228 (.A1(n_0_440), .A2(n_0_266), .ZN(n_0_265));
   NAND2_X1 i_0_229 (.A1(n_17), .A2(negated_second_operand_number[3]), .ZN(
      n_0_266));
   NAND2_X1 i_0_230 (.A1(n_0_273), .A2(n_4), .ZN(n_0_272));
   XNOR2_X1 i_0_231 (.A(second_operand_number[14]), .B(n_0_274), .ZN(n_0_273));
   OAI21_X1 i_0_232 (.A(n_0_275), .B1(second_operand_number[13]), .B2(n_7), 
      .ZN(n_0_274));
   INV_X1 i_0_233 (.A(n_0_276), .ZN(n_0_275));
   AOI21_X1 i_0_234 (.A(n_0_277), .B1(second_operand_number[13]), .B2(n_7), 
      .ZN(n_0_276));
   AOI21_X1 i_0_235 (.A(n_0_278), .B1(n_0_279), .B2(n_0_282), .ZN(n_0_277));
   NOR2_X1 i_0_236 (.A1(n_8), .A2(second_operand_number[12]), .ZN(n_0_278));
   OAI21_X1 i_0_237 (.A(n_0_280), .B1(n_0_283), .B2(second_operand_number[11]), 
      .ZN(n_0_279));
   INV_X1 i_0_238 (.A(n_0_281), .ZN(n_0_280));
   AOI21_X1 i_0_239 (.A(n_9), .B1(n_0_283), .B2(second_operand_number[11]), 
      .ZN(n_0_281));
   NAND2_X1 i_0_240 (.A1(n_8), .A2(second_operand_number[12]), .ZN(n_0_282));
   AOI21_X1 i_0_241 (.A(n_0_284), .B1(n_0_285), .B2(n_0_288), .ZN(n_0_283));
   NOR2_X1 i_0_242 (.A1(n_10), .A2(second_operand_number[10]), .ZN(n_0_284));
   OAI21_X1 i_0_243 (.A(n_0_286), .B1(n_0_289), .B2(second_operand_number[9]), 
      .ZN(n_0_285));
   INV_X1 i_0_244 (.A(n_0_287), .ZN(n_0_286));
   AOI21_X1 i_0_245 (.A(n_11), .B1(n_0_289), .B2(second_operand_number[9]), 
      .ZN(n_0_287));
   NAND2_X1 i_0_246 (.A1(n_10), .A2(second_operand_number[10]), .ZN(n_0_288));
   AOI21_X1 i_0_247 (.A(n_0_290), .B1(n_0_291), .B2(n_0_294), .ZN(n_0_289));
   NOR2_X1 i_0_248 (.A1(n_12), .A2(second_operand_number[8]), .ZN(n_0_290));
   OAI21_X1 i_0_249 (.A(n_0_292), .B1(n_0_295), .B2(second_operand_number[7]), 
      .ZN(n_0_291));
   INV_X1 i_0_250 (.A(n_0_293), .ZN(n_0_292));
   AOI21_X1 i_0_251 (.A(n_13), .B1(n_0_295), .B2(second_operand_number[7]), 
      .ZN(n_0_293));
   NAND2_X1 i_0_252 (.A1(n_12), .A2(second_operand_number[8]), .ZN(n_0_294));
   NOR2_X1 i_0_253 (.A1(n_0_297), .A2(n_0_296), .ZN(n_0_295));
   NOR2_X1 i_0_254 (.A1(n_14), .A2(second_operand_number[6]), .ZN(n_0_296));
   AOI21_X1 i_0_255 (.A(n_0_298), .B1(second_operand_number[6]), .B2(n_14), 
      .ZN(n_0_297));
   AOI21_X1 i_0_256 (.A(n_0_299), .B1(n_0_300), .B2(n_0_301), .ZN(n_0_298));
   NOR2_X1 i_0_257 (.A1(n_15), .A2(second_operand_number[5]), .ZN(n_0_299));
   NAND2_X1 i_0_258 (.A1(n_15), .A2(second_operand_number[5]), .ZN(n_0_300));
   AOI21_X1 i_0_259 (.A(n_0_302), .B1(second_operand_number[4]), .B2(n_16), 
      .ZN(n_0_301));
   NOR2_X1 i_0_260 (.A1(n_0_304), .A2(n_0_303), .ZN(n_0_302));
   NOR2_X1 i_0_261 (.A1(n_16), .A2(second_operand_number[4]), .ZN(n_0_303));
   OAI21_X1 i_0_262 (.A(n_0_305), .B1(second_operand_number[3]), .B2(n_17), 
      .ZN(n_0_304));
   NAND2_X1 i_0_263 (.A1(n_0_450), .A2(n_0_306), .ZN(n_0_305));
   NAND2_X1 i_0_264 (.A1(n_17), .A2(second_operand_number[3]), .ZN(n_0_306));
   OAI21_X1 i_0_367 (.A(n_0_321), .B1(n_0_331), .B2(ready), .ZN(n_83));
   NAND2_X1 i_0_368 (.A1(ready), .A2(n_0_321), .ZN(n_84));
   OAI21_X1 i_0_371 (.A(n_113), .B1(n_0_317), .B2(n_0_331), .ZN(n_85));
   NOR2_X1 i_0_372 (.A1(reset), .A2(n_0_332), .ZN(n_86));
   OAI21_X1 i_0_373 (.A(n_113), .B1(n_0_317), .B2(n_0_332), .ZN(n_87));
   OR2_X1 i_0_265 (.A1(n_0_329), .A2(ready), .ZN(n_0_317));
   NOR2_X1 i_0_381 (.A1(n_0_145), .A2(n_0_447), .ZN(n_88));
   OAI21_X1 i_0_382 (.A(n_0_324), .B1(n_0_145), .B2(n_0_423), .ZN(n_89));
   OAI21_X1 i_0_383 (.A(n_0_324), .B1(n_0_322), .B2(n_0_145), .ZN(n_90));
   XNOR2_X1 i_0_384 (.A(n_0_448), .B(n_0_323), .ZN(n_0_322));
   NAND2_X1 i_0_385 (.A1(n_0_451), .A2(divisor[0]), .ZN(n_0_323));
   NAND3_X1 i_0_386 (.A1(divisor[0]), .A2(n_0_25), .A3(n_0_145), .ZN(n_0_324));
   NOR2_X1 i_0_387 (.A1(n_0_342), .A2(n_0_325), .ZN(n_91));
   NOR3_X1 i_0_388 (.A1(n_0_385), .A2(n_0_346), .A3(n_0_344), .ZN(n_0_325));
   XNOR2_X1 i_0_389 (.A(n_106), .B(n_0_342), .ZN(n_92));
   XOR2_X1 i_0_390 (.A(n_107), .B(n_0_341), .Z(n_93));
   XOR2_X1 i_0_391 (.A(n_108), .B(n_0_0), .Z(n_94));
   NOR2_X1 i_0_392 (.A1(n_0_100), .A2(n_0_326), .ZN(n_95));
   INV_X1 i_0_266 (.A(n_0_327), .ZN(n_0_326));
   OAI21_X1 i_0_267 (.A(n_109), .B1(n_108), .B2(n_0_0), .ZN(n_0_327));
   XNOR2_X1 i_0_268 (.A(n_110), .B(n_0_100), .ZN(n_96));
   XOR2_X1 i_0_396 (.A(n_117), .B(n_0_99), .Z(n_97));
   XNOR2_X1 i_0_269 (.A(n_118), .B(n_0_337), .ZN(n_98));
   XNOR2_X1 i_0_398 (.A(n_119), .B(n_0_96), .ZN(n_99));
   XOR2_X1 i_0_399 (.A(n_120), .B(n_0_95), .Z(n_100));
   XOR2_X1 i_0_400 (.A(n_121), .B(n_0_94), .Z(n_101));
   XOR2_X1 i_0_401 (.A(n_122), .B(n_0_93), .Z(n_102));
   XNOR2_X1 i_0_402 (.A(n_111), .B(n_0_92), .ZN(n_103));
   XOR2_X1 i_0_403 (.A(n_0_89), .B(n_123), .Z(n_104));
   NOR2_X1 i_0_270 (.A1(n_0_99), .A2(n_117), .ZN(n_0_337));
   OR2_X1 i_0_271 (.A1(n_107), .A2(n_0_341), .ZN(n_0_0));
   OR2_X1 i_0_272 (.A1(n_0_343), .A2(n_106), .ZN(n_0_341));
   INV_X1 i_0_419 (.A(n_0_343), .ZN(n_0_342));
   OAI21_X1 i_0_273 (.A(n_0_346), .B1(n_0_344), .B2(n_0_385), .ZN(n_0_343));
   NOR2_X1 i_0_274 (.A1(divisor[0]), .A2(n_0_345), .ZN(n_0_344));
   NOR2_X1 i_0_275 (.A1(n_0_145), .A2(n_0_448), .ZN(n_0_345));
   INV_X1 i_0_276 (.A(n_105), .ZN(n_0_346));
   OAI221_X1 i_0_277 (.A(n_0_347), .B1(n_0_369), .B2(n_0_145), .C1(n_0_144), 
      .C2(n_0_351), .ZN(n_105));
   NAND3_X1 i_0_278 (.A1(n_0_145), .A2(n_0_422), .A3(n_0_25), .ZN(n_0_347));
   OAI21_X1 i_0_279 (.A(n_0_348), .B1(n_0_453), .B2(n_0_145), .ZN(n_106));
   OAI211_X1 i_0_280 (.A(n_0_349), .B(n_0_145), .C1(n_0_76), .C2(n_0_350), 
      .ZN(n_0_348));
   NAND2_X1 i_0_281 (.A1(n_0_76), .A2(n_0_352), .ZN(n_0_349));
   OAI21_X1 i_0_282 (.A(n_0_351), .B1(n_0_369), .B2(n_0_396), .ZN(n_0_350));
   NAND2_X1 i_0_283 (.A1(divisor[0]), .A2(n_0_358), .ZN(n_0_351));
   OAI222_X1 i_0_284 (.A1(n_0_144), .A2(n_0_354), .B1(n_0_352), .B2(n_0_146), 
      .C1(n_0_379), .C2(n_0_145), .ZN(n_107));
   AOI22_X1 i_0_285 (.A1(n_0_422), .A2(n_0_358), .B1(n_0_25), .B2(n_0_375), 
      .ZN(n_0_352));
   OAI221_X1 i_0_286 (.A(n_0_353), .B1(n_0_113), .B2(n_0_145), .C1(n_0_144), 
      .C2(n_0_357), .ZN(n_108));
   OAI21_X1 i_0_287 (.A(n_0_147), .B1(n_0_356), .B2(n_0_355), .ZN(n_0_353));
   NOR2_X1 i_0_288 (.A1(n_0_356), .A2(n_0_355), .ZN(n_0_354));
   NOR3_X1 i_0_289 (.A1(n_0_151), .A2(n_0_143), .A3(n_0_369), .ZN(n_0_355));
   NOR2_X1 i_0_290 (.A1(n_0_362), .A2(n_0_148), .ZN(n_0_356));
   OAI222_X1 i_0_291 (.A1(n_0_361), .A2(n_0_144), .B1(n_0_145), .B2(n_0_123), 
      .C1(n_0_357), .C2(n_0_146), .ZN(n_109));
   AOI21_X1 i_0_292 (.A(n_0_359), .B1(n_0_358), .B2(n_0_375), .ZN(n_0_357));
   NOR2_X1 i_0_293 (.A1(n_0_151), .A2(n_0_143), .ZN(n_0_358));
   NOR2_X1 i_0_294 (.A1(n_0_2), .A2(n_0_148), .ZN(n_0_359));
   OAI222_X1 i_0_295 (.A1(n_0_361), .A2(n_0_146), .B1(n_0_101), .B2(n_0_144), 
      .C1(n_0_145), .C2(n_0_117), .ZN(n_110));
   MUX2_X1 i_0_296 (.A(n_0_362), .B(n_0_3), .S(n_0_151), .Z(n_0_361));
   OAI21_X1 i_0_297 (.A(n_0_363), .B1(n_0_142), .B2(divisor[0]), .ZN(n_0_362));
   NAND2_X1 i_0_298 (.A1(n_0_142), .A2(n_0_379), .ZN(n_0_363));
   OAI21_X1 i_0_299 (.A(n_0_366), .B1(n_0_422), .B2(n_0_142), .ZN(n_0_2));
   NAND2_X1 i_0_300 (.A1(n_0_142), .A2(n_0_113), .ZN(n_0_366));
   MUX2_X1 i_0_301 (.A(n_0_369), .B(n_0_123), .S(n_0_142), .Z(n_0_3));
   XOR2_X1 i_0_302 (.A(divisor[2]), .B(n_0_370), .Z(n_0_369));
   NAND2_X1 i_0_303 (.A1(n_0_421), .A2(divisor[12]), .ZN(n_0_370));
   OAI21_X1 i_0_304 (.A(n_0_374), .B1(n_0_375), .B2(n_0_142), .ZN(n_0_4));
   NAND2_X1 i_0_305 (.A1(n_0_142), .A2(n_0_117), .ZN(n_0_374));
   XNOR2_X1 i_0_306 (.A(divisor[3]), .B(n_0_376), .ZN(n_0_375));
   NAND2_X1 i_0_307 (.A1(n_0_420), .A2(divisor[12]), .ZN(n_0_376));
   MUX2_X1 i_0_465 (.A(n_0_379), .B(n_0_141), .S(n_0_142), .Z(n_0_5));
   XOR2_X1 i_0_308 (.A(divisor[4]), .B(n_0_380), .Z(n_0_379));
   OAI21_X1 i_0_309 (.A(divisor[12]), .B1(n_0_420), .B2(divisor[3]), .ZN(n_0_380));
   NAND2_X1 i_0_310 (.A1(n_0_419), .A2(divisor[12]), .ZN(n_0_24));
   NOR2_X1 i_0_311 (.A1(n_0_25), .A2(n_0_313), .ZN(n_0_385));
   INV_X1 i_0_479 (.A(n_0_90), .ZN(n_111));
   NAND2_X1 i_0_312 (.A1(n_0_151), .A2(n_0_142), .ZN(n_0_396));
   NOR2_X1 i_0_313 (.A1(n_0_143), .A2(n_0_148), .ZN(n_0_25));
   OAI21_X1 i_0_490 (.A(divisor[12]), .B1(n_0_139), .B2(divisor[9]), .ZN(n_0_26));
   NOR2_X1 i_0_494 (.A1(n_0_140), .A2(n_0_451), .ZN(n_0_27));
   NAND2_X1 i_0_499 (.A1(n_0_139), .A2(divisor[12]), .ZN(n_0_36));
   NOR2_X1 i_0_314 (.A1(n_0_138), .A2(n_0_451), .ZN(n_0_37));
   OAI21_X1 i_0_315 (.A(divisor[12]), .B1(n_0_39), .B2(divisor[6]), .ZN(n_0_38));
   OR2_X1 i_0_316 (.A1(n_0_419), .A2(divisor[5]), .ZN(n_0_39));
   OR3_X1 i_0_317 (.A1(n_0_420), .A2(divisor[3]), .A3(divisor[4]), .ZN(n_0_419));
   OR2_X1 i_0_318 (.A1(n_0_421), .A2(divisor[2]), .ZN(n_0_420));
   NAND2_X1 i_0_319 (.A1(n_0_448), .A2(n_0_447), .ZN(n_0_421));
   INV_X1 i_0_320 (.A(n_0_423), .ZN(n_0_422));
   XNOR2_X1 i_0_321 (.A(n_0_448), .B(n_0_424), .ZN(n_0_423));
   NAND2_X1 i_0_322 (.A1(divisor[12]), .A2(divisor[0]), .ZN(n_0_424));
   OAI21_X1 i_0_517 (.A(n_0_428), .B1(n_0_69), .B2(n_0_318), .ZN(n_0_41));
   NAND2_X1 i_0_518 (.A1(dividend[14]), .A2(cla0_n_1), .ZN(n_0_428));
   XNOR2_X1 i_0_519 (.A(n_0_340), .B(cla0_n_2), .ZN(n_0_56));
   XNOR2_X1 i_0_522 (.A(n_0_339), .B(cla0_n_1), .ZN(n_0_68));
   NOR2_X1 i_0_523 (.A1(dividend[13]), .A2(cla0_n_0), .ZN(n_0_69));
   XOR2_X1 i_0_323 (.A(dividend[13]), .B(cla0_n_0), .Z(n_0_76));
   INV_X1 i_0_324 (.A(n_4), .ZN(n_0_446));
   INV_X1 i_0_325 (.A(divisor[0]), .ZN(n_0_447));
   INV_X1 i_0_326 (.A(divisor[1]), .ZN(n_0_448));
   INV_X1 i_0_327 (.A(divisor[12]), .ZN(n_0_451));
   INV_X1 i_0_328 (.A(n_0_375), .ZN(n_0_453));
   OAI211_X1 i_0_329 (.A(n_0_77), .B(n_113), .C1(number_of_bits_in_dividend[1]), 
      .C2(number_of_bits_in_dividend[0]), .ZN(n_112));
   NAND2_X1 i_0_330 (.A1(number_of_bits_in_dividend[1]), .A2(
      number_of_bits_in_dividend[0]), .ZN(n_0_77));
   INV_X1 i_0_331 (.A(reset), .ZN(n_113));
   INV_X1 i_0_332 (.A(n_0_78), .ZN(n_114));
   AOI211_X1 i_0_333 (.A(reset), .B(n_0_79), .C1(number_of_bits_in_dividend[3]), 
      .C2(n_0_80), .ZN(n_0_78));
   NOR2_X1 i_0_334 (.A1(number_of_bits_in_dividend[3]), .A2(n_0_80), .ZN(n_0_79));
   OR3_X1 i_0_335 (.A1(number_of_bits_in_dividend[2]), .A2(
      number_of_bits_in_dividend[0]), .A3(number_of_bits_in_dividend[1]), 
      .ZN(n_0_80));
   OR2_X1 i_0_336 (.A1(n_116), .A2(n_0_84), .ZN(n_115));
   AOI211_X1 i_0_337 (.A(n_0_85), .B(reset), .C1(number_of_bits_in_dividend[4]), 
      .C2(n_0_79), .ZN(n_0_84));
   NOR2_X1 i_0_338 (.A1(number_of_bits_in_dividend[4]), .A2(n_0_79), .ZN(n_0_85));
   NOR3_X1 i_0_339 (.A1(n_113), .A2(n_123), .A3(n_0_89), .ZN(n_116));
   NAND2_X1 i_0_340 (.A1(n_0_92), .A2(n_0_90), .ZN(n_0_89));
   INV_X1 i_0_341 (.A(n_0_91), .ZN(n_0_90));
   OAI22_X1 i_0_342 (.A1(n_0_146), .A2(n_0_114), .B1(n_0_144), .B2(n_0_131), 
      .ZN(n_0_91));
   NOR2_X1 i_0_343 (.A1(n_122), .A2(n_0_93), .ZN(n_0_92));
   OR2_X1 i_0_344 (.A1(n_121), .A2(n_0_94), .ZN(n_0_93));
   OR2_X1 i_0_345 (.A1(n_120), .A2(n_0_95), .ZN(n_0_94));
   NAND2_X1 i_0_346 (.A1(n_0_105), .A2(n_0_96), .ZN(n_0_95));
   NOR3_X1 i_0_347 (.A1(n_117), .A2(n_0_99), .A3(n_118), .ZN(n_0_96));
   NAND2_X1 i_0_348 (.A1(n_0_152), .A2(n_0_100), .ZN(n_0_99));
   NOR3_X1 i_0_349 (.A1(n_109), .A2(n_0_0), .A3(n_108), .ZN(n_0_100));
   OAI222_X1 i_0_350 (.A1(n_0_146), .A2(n_0_101), .B1(n_0_144), .B2(n_0_103), 
      .C1(n_0_145), .C2(n_0_141), .ZN(n_117));
   INV_X1 i_0_351 (.A(n_0_102), .ZN(n_0_101));
   OAI22_X1 i_0_352 (.A1(n_0_2), .A2(n_0_151), .B1(n_0_4), .B2(n_0_148), 
      .ZN(n_0_102));
   OAI222_X1 i_0_353 (.A1(n_0_144), .A2(n_0_106), .B1(n_0_145), .B2(n_0_129), 
      .C1(n_0_146), .C2(n_0_103), .ZN(n_118));
   INV_X1 i_0_354 (.A(n_0_104), .ZN(n_0_103));
   OAI22_X1 i_0_355 (.A1(n_0_3), .A2(n_0_151), .B1(n_0_5), .B2(n_0_148), 
      .ZN(n_0_104));
   INV_X1 i_0_356 (.A(n_119), .ZN(n_0_105));
   OAI222_X1 i_0_357 (.A1(n_0_144), .A2(n_0_107), .B1(n_0_145), .B2(n_0_134), 
      .C1(n_0_146), .C2(n_0_106), .ZN(n_119));
   AOI22_X1 i_0_358 (.A1(n_0_156), .A2(n_0_148), .B1(n_0_151), .B2(n_0_111), 
      .ZN(n_0_106));
   OAI222_X1 i_0_359 (.A1(n_0_146), .A2(n_0_107), .B1(n_0_144), .B2(n_0_110), 
      .C1(n_0_145), .C2(n_0_130), .ZN(n_120));
   AOI22_X1 i_0_360 (.A1(n_0_153), .A2(n_0_148), .B1(n_0_151), .B2(n_0_122), 
      .ZN(n_0_107));
   OAI222_X1 i_0_361 (.A1(n_0_146), .A2(n_0_110), .B1(n_0_145), .B2(n_0_137), 
      .C1(n_0_144), .C2(n_0_118), .ZN(n_121));
   AOI22_X1 i_0_362 (.A1(n_0_148), .A2(n_0_111), .B1(n_0_151), .B2(n_0_116), 
      .ZN(n_0_110));
   OAI22_X1 i_0_363 (.A1(n_0_142), .A2(n_0_113), .B1(n_0_143), .B2(n_0_129), 
      .ZN(n_0_111));
   XOR2_X1 i_0_364 (.A(divisor[5]), .B(n_0_24), .Z(n_0_113));
   OAI22_X1 i_0_365 (.A1(n_0_146), .A2(n_0_118), .B1(n_0_144), .B2(n_0_114), 
      .ZN(n_122));
   AOI21_X1 i_0_366 (.A(n_0_115), .B1(n_0_148), .B2(n_0_116), .ZN(n_0_114));
   NOR2_X1 i_0_369 (.A1(n_0_135), .A2(n_0_129), .ZN(n_0_115));
   OAI22_X1 i_0_370 (.A1(n_0_142), .A2(n_0_117), .B1(n_0_143), .B2(n_0_130), 
      .ZN(n_0_116));
   XOR2_X1 i_0_374 (.A(divisor[7]), .B(n_0_38), .Z(n_0_117));
   AOI22_X1 i_0_375 (.A1(n_0_151), .A2(n_0_136), .B1(n_0_148), .B2(n_0_122), 
      .ZN(n_0_118));
   OAI22_X1 i_0_376 (.A1(n_0_142), .A2(n_0_123), .B1(n_0_143), .B2(n_0_134), 
      .ZN(n_0_122));
   XOR2_X1 i_0_377 (.A(divisor[6]), .B(n_0_126), .Z(n_0_123));
   NAND2_X1 i_0_378 (.A1(divisor[12]), .A2(n_0_39), .ZN(n_0_126));
   OAI33_X1 i_0_379 (.A1(n_0_76), .A2(n_0_313), .A3(n_0_131), .B1(n_0_144), 
      .B2(n_0_142), .B3(n_0_127), .ZN(n_123));
   INV_X1 i_0_380 (.A(n_0_128), .ZN(n_0_127));
   OAI22_X1 i_0_393 (.A1(n_0_148), .A2(n_0_130), .B1(n_0_151), .B2(n_0_129), 
      .ZN(n_0_128));
   XOR2_X1 i_0_394 (.A(divisor[9]), .B(n_0_36), .Z(n_0_129));
   XOR2_X1 i_0_395 (.A(n_0_155), .B(n_0_37), .Z(n_0_130));
   AOI21_X1 i_0_397 (.A(n_0_132), .B1(n_0_148), .B2(n_0_136), .ZN(n_0_131));
   NOR2_X1 i_0_404 (.A1(n_0_135), .A2(n_0_134), .ZN(n_0_132));
   XOR2_X1 i_0_405 (.A(divisor[10]), .B(n_0_26), .Z(n_0_134));
   NAND2_X1 i_0_406 (.A1(n_0_151), .A2(n_0_143), .ZN(n_0_135));
   OAI22_X1 i_0_407 (.A1(n_0_142), .A2(n_0_141), .B1(n_0_143), .B2(n_0_137), 
      .ZN(n_0_136));
   NAND3_X1 i_0_408 (.A1(divisor[12]), .A2(n_0_155), .A3(n_0_138), .ZN(n_0_137));
   NOR3_X1 i_0_409 (.A1(divisor[9]), .A2(n_0_139), .A3(divisor[10]), .ZN(n_0_138));
   NAND2_X1 i_0_410 (.A1(n_0_154), .A2(n_0_140), .ZN(n_0_139));
   NOR3_X1 i_0_411 (.A1(divisor[6]), .A2(n_0_39), .A3(divisor[7]), .ZN(n_0_140));
   XOR2_X1 i_0_412 (.A(n_0_154), .B(n_0_27), .Z(n_0_141));
   INV_X1 i_0_413 (.A(n_0_143), .ZN(n_0_142));
   XOR2_X1 i_0_414 (.A(n_0_56), .B(n_0_41), .Z(n_0_143));
   NAND2_X1 i_0_415 (.A1(n_0_76), .A2(n_0_145), .ZN(n_0_144));
   OAI21_X1 i_0_416 (.A(n_0_146), .B1(n_0_313), .B2(n_0_25), .ZN(n_0_145));
   INV_X1 i_0_417 (.A(n_0_147), .ZN(n_0_146));
   NOR2_X1 i_0_418 (.A1(n_0_76), .A2(n_0_313), .ZN(n_0_147));
   INV_X1 i_0_420 (.A(n_0_151), .ZN(n_0_148));
   XOR2_X1 i_0_421 (.A(n_0_69), .B(n_0_68), .Z(n_0_151));
   INV_X1 i_0_422 (.A(n_110), .ZN(n_0_152));
   INV_X1 i_0_423 (.A(n_0_5), .ZN(n_0_153));
   INV_X1 i_0_424 (.A(divisor[8]), .ZN(n_0_154));
   INV_X1 i_0_425 (.A(divisor[11]), .ZN(n_0_155));
   INV_X1 i_0_426 (.A(n_0_4), .ZN(n_0_156));
   OAI21_X1 i_0_427 (.A(n_0_157), .B1(n_0_333), .B2(n_0_319), .ZN(n_124));
   AOI22_X1 i_0_428 (.A1(dividend[0]), .A2(n_0_175), .B1(n_33), .B2(n_0_173), 
      .ZN(n_0_157));
   NOR2_X1 i_0_429 (.A1(reset), .A2(n_0_328), .ZN(n_0_173));
   NOR2_X1 i_0_430 (.A1(n_113), .A2(n_0_226), .ZN(n_0_175));
   INV_X1 i_0_431 (.A(n_0_267), .ZN(n_0_226));
   OAI21_X1 i_0_432 (.A(n_0_313), .B1(n_0_270), .B2(n_0_268), .ZN(n_0_267));
   INV_X1 i_0_433 (.A(n_0_269), .ZN(n_0_268));
   AOI21_X1 i_0_434 (.A(n_0_311), .B1(divisor[13]), .B2(cla1_n_0), .ZN(n_0_269));
   NAND2_X1 i_0_435 (.A1(n_0_308), .A2(n_0_271), .ZN(n_0_270));
   XNOR2_X1 i_0_436 (.A(n_0_311), .B(n_0_307), .ZN(n_0_271));
   OAI22_X1 i_0_437 (.A1(n_0_339), .A2(divisor[14]), .B1(dividend[14]), .B2(
      n_0_338), .ZN(n_0_307));
   INV_X1 i_0_438 (.A(n_0_309), .ZN(n_0_308));
   XOR2_X1 i_0_439 (.A(n_0_312), .B(n_0_310), .Z(n_0_309));
   OAI22_X1 i_0_440 (.A1(dividend[14]), .A2(n_0_338), .B1(n_0_315), .B2(n_0_311), 
      .ZN(n_0_310));
   NOR2_X1 i_0_441 (.A1(divisor[13]), .A2(cla1_n_0), .ZN(n_0_311));
   XOR2_X1 i_0_442 (.A(n_0_340), .B(divisor[15]), .Z(n_0_312));
   OAI22_X1 i_0_443 (.A1(dividend[15]), .A2(cla0_n_2), .B1(n_0_315), .B2(n_0_314), 
      .ZN(n_0_313));
   OAI22_X1 i_0_444 (.A1(n_0_318), .A2(n_0_316), .B1(n_0_340), .B2(divisor[15]), 
      .ZN(n_0_314));
   NOR2_X1 i_0_445 (.A1(n_0_339), .A2(divisor[14]), .ZN(n_0_315));
   NAND2_X1 i_0_446 (.A1(dividend[13]), .A2(cla0_n_0), .ZN(n_0_316));
   NOR2_X1 i_0_447 (.A1(dividend[14]), .A2(cla0_n_1), .ZN(n_0_318));
   NAND2_X1 i_0_448 (.A1(n_0_332), .A2(n_0_320), .ZN(n_0_319));
   NOR2_X1 i_0_449 (.A1(ready), .A2(n_125), .ZN(n_0_320));
   INV_X1 i_0_450 (.A(n_0_321), .ZN(n_125));
   NOR2_X1 i_0_451 (.A1(reset), .A2(n_0_329), .ZN(n_0_321));
   INV_X1 i_0_452 (.A(n_0_329), .ZN(n_0_328));
   NAND4_X1 i_0_453 (.A1(number_of_bits_in_dividend[2]), .A2(
      number_of_bits_in_dividend[1]), .A3(number_of_bits_in_dividend[0]), 
      .A4(n_0_330), .ZN(n_0_329));
   AND2_X1 i_0_454 (.A1(number_of_bits_in_dividend[4]), .A2(
      number_of_bits_in_dividend[3]), .ZN(n_0_330));
   INV_X1 i_0_455 (.A(n_0_332), .ZN(n_0_331));
   NOR4_X1 i_0_456 (.A1(n_21), .A2(n_22), .A3(n_23), .A4(n_24), .ZN(n_0_332));
   XOR2_X1 i_0_457 (.A(n_32), .B(n_0_334), .Z(n_0_333));
   NAND2_X1 i_0_458 (.A1(sign), .A2(n_0_335), .ZN(n_0_334));
   OR3_X1 i_0_459 (.A1(n_34), .A2(n_0_336), .A3(n_33), .ZN(n_0_335));
   OR2_X1 i_0_460 (.A1(n_35), .A2(n_36), .ZN(n_0_336));
   INV_X1 i_0_461 (.A(divisor[14]), .ZN(n_0_338));
   INV_X1 i_0_462 (.A(dividend[14]), .ZN(n_0_339));
   INV_X1 i_0_463 (.A(dividend[15]), .ZN(n_0_340));
   NAND2_X1 i_0_464 (.A1(n_0_226), .A2(reset), .ZN(n_0_360));
   NOR2_X1 i_0_466 (.A1(n_0_360), .A2(n_0_268), .ZN(n_0_364));
   INV_X1 i_0_467 (.A(dividend[0]), .ZN(n_0_365));
   OR3_X1 i_0_468 (.A1(dividend[2]), .A2(dividend[1]), .A3(dividend[0]), 
      .ZN(n_0_367));
   NAND2_X1 i_0_469 (.A1(n_0_367), .A2(dividend[12]), .ZN(n_0_368));
   XOR2_X1 i_0_470 (.A(n_0_368), .B(dividend[3]), .Z(n_0_371));
   NAND2_X1 i_0_471 (.A1(dividend[12]), .A2(dividend[0]), .ZN(n_0_372));
   XOR2_X1 i_0_472 (.A(n_0_372), .B(dividend[1]), .Z(n_0_373));
   INV_X1 i_0_473 (.A(n_0_271), .ZN(n_0_377));
   NAND2_X1 i_0_474 (.A1(n_0_377), .A2(n_0_308), .ZN(n_0_378));
   OAI22_X1 i_0_475 (.A1(n_0_371), .A2(n_0_270), .B1(n_0_378), .B2(n_0_373), 
      .ZN(n_0_381));
   OAI21_X1 i_0_476 (.A(dividend[12]), .B1(dividend[1]), .B2(dividend[0]), 
      .ZN(n_0_382));
   XOR2_X1 i_0_477 (.A(n_0_382), .B(dividend[2]), .Z(n_0_383));
   OAI22_X1 i_0_478 (.A1(n_0_383), .A2(n_0_270), .B1(n_0_378), .B2(n_0_365), 
      .ZN(n_0_384));
   INV_X1 i_0_480 (.A(n_0_268), .ZN(n_0_386));
   NOR2_X1 i_0_481 (.A1(n_0_360), .A2(n_0_386), .ZN(n_0_387));
   OR2_X1 i_0_482 (.A1(n_32), .A2(n_0_335), .ZN(n_0_388));
   OAI21_X1 i_0_483 (.A(sign), .B1(n_0_388), .B2(n_31), .ZN(n_0_389));
   INV_X1 i_0_484 (.A(n_30), .ZN(n_0_390));
   NAND2_X1 i_0_485 (.A1(n_0_389), .A2(n_0_390), .ZN(n_0_391));
   NAND2_X1 i_0_486 (.A1(n_0_391), .A2(sign), .ZN(n_0_392));
   XOR2_X1 i_0_487 (.A(n_29), .B(n_0_392), .Z(n_0_393));
   NAND2_X1 i_0_488 (.A1(reset), .A2(n_0_267), .ZN(n_0_394));
   AOI222_X1 i_0_489 (.A1(n_0_381), .A2(n_0_364), .B1(n_0_384), .B2(n_0_387), 
      .C1(n_0_173), .C2(n_30), .ZN(n_0_395));
   OAI221_X1 i_0_491 (.A(n_0_395), .B1(n_0_319), .B2(n_0_393), .C1(n_0_394), 
      .C2(n_0_371), .ZN(n_126));
   OAI221_X1 i_0_492 (.A(n_0_397), .B1(n_0_399), .B2(n_0_398), .C1(n_0_413), 
      .C2(n_0_412), .ZN(n_127));
   AOI221_X1 i_0_493 (.A(n_0_434), .B1(n_0_175), .B2(n_0_408), .C1(n_0_173), 
      .C2(n_23), .ZN(n_0_397));
   NAND3_X1 i_0_495 (.A1(reset), .A2(n_0_386), .A3(n_0_226), .ZN(n_0_398));
   AOI21_X1 i_0_496 (.A(n_0_400), .B1(n_0_377), .B2(n_0_401), .ZN(n_0_399));
   NOR2_X1 i_0_497 (.A1(n_0_377), .A2(n_0_407), .ZN(n_0_400));
   INV_X1 i_0_498 (.A(n_0_402), .ZN(n_0_401));
   OAI22_X1 i_0_500 (.A1(n_0_436), .A2(n_0_403), .B1(n_0_308), .B2(n_0_405), 
      .ZN(n_0_402));
   XNOR2_X1 i_0_501 (.A(dividend[8]), .B(n_0_404), .ZN(n_0_403));
   NAND2_X1 i_0_502 (.A1(dividend[12]), .A2(n_0_431), .ZN(n_0_404));
   XNOR2_X1 i_0_503 (.A(dividend[4]), .B(n_0_406), .ZN(n_0_405));
   OAI21_X1 i_0_504 (.A(dividend[12]), .B1(n_0_367), .B2(dividend[3]), .ZN(
      n_0_406));
   OAI22_X1 i_0_505 (.A1(n_0_309), .A2(n_0_408), .B1(n_0_308), .B2(n_0_410), 
      .ZN(n_0_407));
   XNOR2_X1 i_0_506 (.A(dividend[10]), .B(n_0_409), .ZN(n_0_408));
   NAND2_X1 i_0_507 (.A1(dividend[12]), .A2(n_0_430), .ZN(n_0_409));
   XNOR2_X1 i_0_508 (.A(dividend[6]), .B(n_0_411), .ZN(n_0_410));
   NAND2_X1 i_0_509 (.A1(dividend[12]), .A2(n_0_432), .ZN(n_0_411));
   NAND3_X1 i_0_510 (.A1(n_0_313), .A2(n_0_268), .A3(reset), .ZN(n_0_412));
   OAI22_X1 i_0_511 (.A1(n_0_435), .A2(n_0_414), .B1(n_0_271), .B2(n_0_426), 
      .ZN(n_0_413));
   OAI22_X1 i_0_512 (.A1(n_0_436), .A2(n_0_415), .B1(n_0_308), .B2(n_0_417), 
      .ZN(n_0_414));
   XOR2_X1 i_0_513 (.A(dividend[9]), .B(n_0_416), .Z(n_0_415));
   OAI21_X1 i_0_514 (.A(dividend[12]), .B1(dividend[8]), .B2(n_0_431), .ZN(
      n_0_416));
   XNOR2_X1 i_0_515 (.A(dividend[5]), .B(n_0_418), .ZN(n_0_417));
   NOR2_X1 i_0_516 (.A1(n_0_438), .A2(n_0_433), .ZN(n_0_418));
   INV_X1 i_0_520 (.A(n_0_426), .ZN(n_0_425));
   OAI22_X1 i_0_521 (.A1(n_0_436), .A2(n_0_427), .B1(n_0_308), .B2(n_0_371), 
      .ZN(n_0_426));
   XOR2_X1 i_0_524 (.A(dividend[7]), .B(n_0_429), .Z(n_0_427));
   OAI21_X1 i_0_525 (.A(dividend[12]), .B1(dividend[6]), .B2(n_0_432), .ZN(
      n_0_429));
   OR3_X1 i_0_526 (.A1(dividend[8]), .A2(n_0_431), .A3(dividend[9]), .ZN(n_0_430));
   OR3_X1 i_0_527 (.A1(dividend[6]), .A2(n_0_432), .A3(dividend[7]), .ZN(n_0_431));
   NAND2_X1 i_0_528 (.A1(n_0_437), .A2(n_0_433), .ZN(n_0_432));
   NOR3_X1 i_0_529 (.A1(n_0_367), .A2(dividend[3]), .A3(dividend[4]), .ZN(
      n_0_433));
   NOR3_X1 i_0_530 (.A1(n_125), .A2(n_0_331), .A3(ready), .ZN(n_0_434));
   INV_X1 i_0_531 (.A(n_0_271), .ZN(n_0_435));
   INV_X1 i_0_532 (.A(n_0_308), .ZN(n_0_436));
   INV_X1 i_0_533 (.A(dividend[5]), .ZN(n_0_437));
   INV_X1 i_0_534 (.A(dividend[12]), .ZN(n_0_438));
   XOR2_X1 i_0_535 (.A(negated_second_operand_number[3]), .B(n_0_440), .Z(
      n_0_439));
   OAI22_X1 i_0_536 (.A1(n_18), .A2(negated_second_operand_number[2]), .B1(
      n_0_442), .B2(n_0_441), .ZN(n_0_440));
   AND2_X1 i_0_537 (.A1(n_18), .A2(negated_second_operand_number[2]), .ZN(
      n_0_441));
   NOR2_X1 i_0_538 (.A1(n_0_444), .A2(n_0_443), .ZN(n_0_442));
   AOI21_X1 i_0_539 (.A(negated_second_operand_number[1]), .B1(n_19), .B2(
      n_0_445), .ZN(n_0_443));
   NOR2_X1 i_0_540 (.A1(n_19), .A2(n_0_445), .ZN(n_0_444));
   AND2_X1 i_0_541 (.A1(n_20), .A2(negated_second_operand_number[0]), .ZN(
      n_0_445));
   XNOR2_X1 i_0_542 (.A(second_operand_number[3]), .B(n_0_450), .ZN(n_0_449));
   AOI22_X1 i_0_543 (.A1(second_operand_number[2]), .A2(n_18), .B1(n_0_454), 
      .B2(n_0_452), .ZN(n_0_450));
   OR2_X1 i_0_544 (.A1(second_operand_number[2]), .A2(n_18), .ZN(n_0_452));
   NOR2_X1 i_0_545 (.A1(n_0_444), .A2(n_0_455), .ZN(n_0_454));
   AOI21_X1 i_0_546 (.A(second_operand_number[1]), .B1(n_0_445), .B2(n_19), 
      .ZN(n_0_455));
   MUX2_X1 overFlow_reg_enable_mux_0 (.A(overFlow), .B(n_86), .S(n_87), .Z(n_128));
   MUX2_X1 ready_reg_enable_mux_0 (.A(ready), .B(n_113), .S(n_53), .Z(n_129));
endmodule

module Interpolation(RST, CLK, Interpolation_Enable, Interpolation_Intialize, 
      Interpolation_Memory_WR_Enable, Interpolation_RAM_RD1_Data, 
      Interpolation_RAM_RD2_Data, Interpolation_RAM_WR_Data, 
      Interpolation_RAM_RD1_Address, Interpolation_RAM_RD2_Address, 
      Interpolation_RAM_WR_Address, Interpolation_Done, Intialization_Done, 
      Error, intialization_state, interpolation_state);
   input RST;
   input CLK;
   input Interpolation_Enable;
   input Interpolation_Intialize;
   output Interpolation_Memory_WR_Enable;
   input [63:0]Interpolation_RAM_RD1_Data;
   input [63:0]Interpolation_RAM_RD2_Data;
   output [63:0]Interpolation_RAM_WR_Data;
   output [12:0]Interpolation_RAM_RD1_Address;
   output [12:0]Interpolation_RAM_RD2_Address;
   output [12:0]Interpolation_RAM_WR_Address;
   output Interpolation_Done;
   output Intialization_Done;
   output Error;
   output [3:0]intialization_state;
   output [3:0]interpolation_state;

   wire [63:0]UN;
   wire [63:0]Temp;
   wire [12:0]UZ_ADD;
   wire [12:0]TZ_ADD;
   wire n_0_0;
   wire [3:0]current_intialization_state;
   wire n_0_1;
   wire [3:0]current_interpolation_state;
   wire [15:0]adder_sub1_In1;
   wire [15:0]adder_sub1_In2;
   wire n_0_2;
   wire n_0_3;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_10;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_11;
   wire n_0_0_7;
   wire n_0_12;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_13;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_14;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_15;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_16;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_17;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_18;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_19;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_20;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_21;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_22;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_23;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_24;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_25;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_26;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_27;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_28;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_29;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_30;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_36;
   wire n_0_0_166;
   wire n_0_37;
   wire n_0_0_167;
   wire n_0_38;
   wire n_0_0_168;
   wire n_0_39;
   wire n_0_0_169;
   wire n_0_40;
   wire n_0_0_170;
   wire n_0_41;
   wire n_0_0_171;
   wire n_0_42;
   wire n_0_0_172;
   wire n_0_43;
   wire n_0_0_173;
   wire n_0_44;
   wire n_0_0_174;
   wire n_0_45;
   wire n_0_0_175;
   wire n_0_46;
   wire n_0_0_176;
   wire n_0_47;
   wire n_0_0_177;
   wire n_0_48;
   wire n_0_0_178;
   wire n_0_49;
   wire n_0_0_179;
   wire n_0_50;
   wire n_0_0_180;
   wire n_0_51;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_52;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_53;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_54;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_55;
   wire n_0_0_204;
   wire n_0_56;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_57;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_58;
   wire n_0_0_209;
   wire n_0_59;
   wire n_0_0_210;
   wire n_0_60;
   wire n_0_0_211;
   wire n_0_61;
   wire n_0_0_212;
   wire n_0_62;
   wire n_0_0_213;
   wire n_0_63;
   wire n_0_0_214;
   wire n_0_64;
   wire n_0_0_215;
   wire n_0_65;
   wire n_0_0_216;
   wire n_0_66;
   wire n_0_0_217;
   wire n_0_67;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_68;
   wire n_0_0_244;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_84;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_85;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_87;
   wire n_0_89;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_88;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_90;
   wire n_0_91;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_92;
   wire n_0_93;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_0_366;
   wire n_0_0_367;
   wire n_0_0_368;
   wire n_0_0_369;
   wire n_0_0_370;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_86;
   wire n_0_0_371;
   wire n_0_0_372;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_377;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_0_383;
   wire n_0_0_384;
   wire n_0_0_385;
   wire n_0_0_386;
   wire n_0_0_387;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_0_391;
   wire n_0_0_392;
   wire n_0_0_393;
   wire n_0_0_394;
   wire n_0_0_395;
   wire n_0_0_396;
   wire n_0_0_397;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_0_402;
   wire n_0_0_403;
   wire n_0_0_404;
   wire n_0_0_405;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_0_408;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire [15:0]adder_sub3_In2;
   wire [15:0]adder_sub3_In1;
   wire [15:0]div1_divisor;
   wire [15:0]div1_dividend;
   wire n_1_0;
   wire mult1_enable;
   wire [15:0]mult1_second_operand;
   wire [15:0]mult1_first_operand;
   wire div1_reset;
   wire [15:0]adder_sub2_In1;
   wire [15:0]adder_sub2_In2;
   wire Start_Intialization;
   wire Start_Interpolation;
   wire n_1_1;
   wire [2:0]Count2;
   wire n_1_2;
   wire n_1_3;
   wire Div_Count;
   wire n_1_14;
   wire [4:0]USIZE;
   wire [7:0]U_CURRENT_SIZE;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire adder_sub1_Sub;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_15;
   wire n_1_13;
   wire n_1_12;
   wire n_1_16;
   wire [15:0]mult1_out;
   wire div1_divideByZero;
   wire div1_overFlow;
   wire div1_ready;
   wire [15:0]div1_Q;
   wire [15:0]adder_sub1_Out;
   wire adder_sub1_i_0_n_0;
   wire adder_sub1_i_0_n_1;
   wire adder_sub1_i_0_n_2;
   wire adder_sub1_i_0_n_3;
   wire adder_sub1_i_0_n_4;
   wire adder_sub1_i_0_n_5;
   wire adder_sub1_i_0_n_6;
   wire adder_sub1_i_0_n_7;
   wire adder_sub1_i_0_n_8;
   wire adder_sub1_i_0_n_9;
   wire adder_sub1_i_0_n_10;
   wire adder_sub1_i_0_n_11;
   wire adder_sub1_i_0_n_12;
   wire adder_sub1_i_0_n_13;
   wire adder_sub1_i_0_n_14;
   wire adder_sub1_i_0_n_67;
   wire adder_sub1_i_0_n_68;
   wire adder_sub1_i_0_n_69;
   wire adder_sub1_i_0_n_70;
   wire adder_sub1_i_0_n_74;
   wire adder_sub1_i_0_n_75;
   wire adder_sub1_i_0_n_76;
   wire adder_sub1_i_0_n_80;
   wire adder_sub1_i_0_n_81;
   wire adder_sub1_i_0_n_82;
   wire adder_sub1_i_0_n_83;
   wire adder_sub1_i_0_n_86;
   wire adder_sub1_i_0_n_87;
   wire adder_sub1_i_0_n_88;
   wire adder_sub1_i_0_n_89;
   wire adder_sub1_i_0_n_90;
   wire adder_sub1_i_0_n_92;
   wire adder_sub1_i_0_n_93;
   wire adder_sub1_i_0_n_94;
   wire adder_sub1_i_0_n_95;
   wire adder_sub1_i_0_n_96;
   wire adder_sub1_i_0_n_97;
   wire adder_sub1_i_0_n_98;
   wire adder_sub1_i_0_n_100;
   wire adder_sub1_i_0_n_101;
   wire adder_sub1_i_0_n_102;
   wire adder_sub1_i_0_n_103;
   wire adder_sub1_i_0_n_105;
   wire adder_sub1_i_0_n_106;
   wire adder_sub1_i_0_n_107;
   wire adder_sub1_i_0_n_108;
   wire adder_sub1_i_0_n_109;
   wire adder_sub1_i_0_n_110;
   wire adder_sub1_i_0_n_111;
   wire adder_sub1_i_0_n_114;
   wire adder_sub1_i_0_n_115;
   wire adder_sub1_i_0_n_116;
   wire adder_sub1_i_0_n_117;
   wire adder_sub1_i_0_n_119;
   wire adder_sub1_i_0_n_120;
   wire adder_sub1_i_0_n_121;
   wire adder_sub1_i_0_n_124;
   wire adder_sub1_i_0_n_125;
   wire adder_sub1_i_0_n_126;
   wire adder_sub1_i_0_n_127;
   wire adder_sub1_i_0_n_128;
   wire adder_sub1_i_0_n_130;
   wire adder_sub1_i_0_n_131;
   wire adder_sub1_i_0_n_132;
   wire adder_sub1_i_0_n_133;
   wire adder_sub1_i_0_n_134;
   wire adder_sub1_i_0_n_135;
   wire adder_sub1_i_0_n_136;
   wire adder_sub1_i_0_n_137;
   wire adder_sub1_i_0_n_138;
   wire adder_sub1_i_0_n_139;
   wire adder_sub1_i_0_n_140;
   wire adder_sub1_i_0_n_141;
   wire adder_sub1_i_0_n_142;
   wire adder_sub1_i_0_n_143;
   wire adder_sub1_i_0_n_144;
   wire adder_sub1_i_0_n_145;
   wire adder_sub1_i_0_n_146;
   wire adder_sub1_i_0_n_147;
   wire adder_sub1_i_0_n_148;
   wire adder_sub1_i_0_n_149;
   wire adder_sub1_i_0_n_150;
   wire adder_sub1_i_0_n_151;
   wire adder_sub1_i_0_n_152;
   wire adder_sub1_i_0_n_153;
   wire adder_sub1_i_0_n_161;
   wire adder_sub1_i_0_n_162;
   wire adder_sub1_i_0_n_163;
   wire adder_sub1_i_0_n_164;
   wire adder_sub1_i_0_n_166;
   wire adder_sub1_i_0_n_167;
   wire adder_sub1_i_0_n_168;
   wire adder_sub1_i_0_n_169;
   wire adder_sub1_i_0_n_170;
   wire adder_sub1_i_0_n_171;
   wire adder_sub1_i_0_n_190;
   wire adder_sub1_i_0_n_198;
   wire adder_sub1_i_0_n_15;
   wire adder_sub1_i_0_n_16;
   wire adder_sub1_i_0_n_17;
   wire adder_sub1_i_0_n_18;
   wire adder_sub1_i_0_n_19;
   wire adder_sub1_i_0_n_20;
   wire adder_sub1_i_0_n_21;
   wire adder_sub1_i_0_n_22;
   wire adder_sub1_i_0_n_23;
   wire adder_sub1_i_0_n_24;
   wire adder_sub1_i_0_n_25;
   wire adder_sub1_i_0_n_26;
   wire adder_sub1_i_0_n_27;
   wire adder_sub1_i_0_n_28;
   wire adder_sub1_i_0_n_29;
   wire adder_sub1_i_0_n_30;
   wire adder_sub1_i_0_n_31;
   wire adder_sub1_i_0_n_32;
   wire adder_sub1_i_0_n_33;
   wire adder_sub1_i_0_n_34;
   wire adder_sub1_i_0_n_35;
   wire adder_sub1_i_0_n_36;
   wire adder_sub1_i_0_n_37;
   wire adder_sub1_i_0_n_38;
   wire adder_sub1_i_0_n_39;
   wire adder_sub1_i_0_n_40;
   wire adder_sub1_i_0_n_41;
   wire adder_sub1_i_0_n_42;
   wire adder_sub1_i_0_n_43;
   wire adder_sub1_i_0_n_44;
   wire adder_sub1_i_0_n_45;
   wire adder_sub1_i_0_n_46;
   wire adder_sub1_i_0_n_47;
   wire adder_sub1_i_0_n_48;
   wire adder_sub1_i_0_n_49;
   wire adder_sub1_i_0_n_50;
   wire adder_sub1_i_0_n_51;
   wire adder_sub1_i_0_n_52;
   wire adder_sub1_i_0_n_53;
   wire adder_sub1_i_0_n_54;
   wire adder_sub1_i_0_n_55;
   wire adder_sub1_i_0_n_56;
   wire adder_sub1_i_0_n_57;
   wire adder_sub1_i_0_n_58;
   wire adder_sub1_i_0_n_59;
   wire adder_sub1_i_0_n_60;
   wire adder_sub1_i_0_n_61;
   wire adder_sub1_i_0_n_62;
   wire adder_sub1_i_0_n_63;
   wire adder_sub1_i_0_n_64;
   wire adder_sub1_i_0_n_65;
   wire adder_sub1_i_0_n_66;
   wire adder_sub1_i_0_n_71;
   wire adder_sub1_i_0_n_72;
   wire adder_sub1_i_0_n_73;
   wire adder_sub1_i_0_n_77;
   wire adder_sub1_i_0_n_78;
   wire adder_sub1_i_0_n_79;
   wire adder_sub1_i_0_n_84;
   wire adder_sub1_i_0_n_85;
   wire adder_sub1_i_0_n_91;
   wire adder_sub1_i_0_n_99;
   wire adder_sub1_i_0_n_104;
   wire adder_sub1_i_0_n_112;
   wire adder_sub1_i_0_n_113;
   wire adder_sub1_i_0_n_118;
   wire adder_sub1_i_0_n_122;
   wire adder_sub1_i_0_n_123;
   wire adder_sub1_i_0_n_129;
   wire adder_sub1_i_0_n_154;
   wire adder_sub1_i_0_n_155;
   wire adder_sub1_i_0_n_156;
   wire adder_sub1_i_0_n_157;
   wire adder_sub1_i_0_n_158;
   wire adder_sub1_i_0_n_159;
   wire adder_sub1_i_0_n_160;
   wire adder_sub1_i_0_n_165;
   wire adder_sub1_i_0_n_172;
   wire adder_sub1_i_0_n_173;
   wire adder_sub1_i_0_n_174;
   wire adder_sub1_i_0_n_175;
   wire adder_sub1_i_0_n_176;
   wire adder_sub1_i_0_n_177;
   wire adder_sub1_i_0_n_178;
   wire adder_sub1_i_0_n_179;
   wire adder_sub1_i_0_n_180;
   wire adder_sub1_i_0_n_181;
   wire adder_sub1_i_0_n_182;
   wire adder_sub1_i_0_n_183;
   wire adder_sub1_i_0_n_184;
   wire adder_sub1_i_0_n_185;
   wire adder_sub1_i_0_n_186;
   wire adder_sub1_i_0_n_187;
   wire adder_sub1_i_0_n_188;
   wire adder_sub1_i_0_n_189;
   wire adder_sub1_i_0_n_191;
   wire adder_sub1_i_0_n_192;
   wire adder_sub1_i_0_n_193;
   wire adder_sub1_i_0_n_194;
   wire adder_sub1_i_0_n_195;
   wire adder_sub1_i_0_n_196;
   wire adder_sub1_i_0_n_197;
   wire adder_sub1_i_0_n_199;
   wire adder_sub1_i_0_n_200;
   wire adder_sub2_i_0_n_2;
   wire adder_sub2_i_0_n_4;
   wire adder_sub2_i_0_n_5;
   wire adder_sub2_i_0_n_6;
   wire adder_sub2_i_0_n_7;
   wire adder_sub2_i_0_n_8;
   wire adder_sub2_i_0_n_9;
   wire adder_sub2_i_0_n_10;
   wire adder_sub2_i_0_n_11;
   wire adder_sub2_i_0_n_12;
   wire adder_sub2_i_0_n_13;
   wire adder_sub2_i_0_n_14;
   wire adder_sub2_i_0_n_26;
   wire adder_sub2_i_0_n_0;
   wire adder_sub2_i_0_n_1;
   wire adder_sub2_i_0_n_3;
   wire adder_sub2_i_0_n_15;
   wire adder_sub2_i_0_n_16;
   wire adder_sub2_i_0_n_17;
   wire adder_sub2_i_0_n_18;
   wire adder_sub2_i_0_n_19;
   wire adder_sub2_i_0_n_20;
   wire adder_sub2_i_0_n_21;
   wire adder_sub2_i_0_n_22;
   wire adder_sub2_i_0_n_23;
   wire adder_sub2_i_0_n_24;
   wire adder_sub2_i_0_n_25;
   wire adder_sub2_i_0_n_27;
   wire adder_sub2_i_0_n_28;
   wire n_2_0_0;
   wire n_2_0_1;

   assign Interpolation_RAM_WR_Data[63] = 1'b0;
   assign Interpolation_RAM_WR_Data[62] = 1'b0;
   assign Interpolation_RAM_WR_Data[61] = 1'b0;
   assign Interpolation_RAM_WR_Data[60] = 1'b0;
   assign Interpolation_RAM_WR_Data[59] = 1'b0;
   assign Interpolation_RAM_WR_Data[58] = 1'b0;
   assign Interpolation_RAM_WR_Data[57] = 1'b0;
   assign Interpolation_RAM_WR_Data[56] = 1'b0;
   assign Interpolation_RAM_WR_Data[55] = 1'b0;
   assign Interpolation_RAM_WR_Data[54] = 1'b0;
   assign Interpolation_RAM_WR_Data[53] = 1'b0;
   assign Interpolation_RAM_WR_Data[52] = 1'b0;
   assign Interpolation_RAM_WR_Data[51] = 1'b0;
   assign Interpolation_RAM_WR_Data[50] = 1'b0;
   assign Interpolation_RAM_WR_Data[49] = 1'b0;
   assign Interpolation_RAM_WR_Data[48] = 1'b0;
   assign Interpolation_RAM_WR_Data[47] = 1'b0;
   assign Interpolation_RAM_WR_Data[46] = 1'b0;
   assign Interpolation_RAM_WR_Data[45] = 1'b0;
   assign Interpolation_RAM_WR_Data[44] = 1'b0;
   assign Interpolation_RAM_WR_Data[43] = 1'b0;
   assign Interpolation_RAM_WR_Data[42] = 1'b0;
   assign Interpolation_RAM_WR_Data[41] = 1'b0;
   assign Interpolation_RAM_WR_Data[40] = 1'b0;
   assign Interpolation_RAM_WR_Data[39] = 1'b0;
   assign Interpolation_RAM_WR_Data[38] = 1'b0;
   assign Interpolation_RAM_WR_Data[37] = 1'b0;
   assign Interpolation_RAM_WR_Data[36] = 1'b0;
   assign Interpolation_RAM_WR_Data[35] = 1'b0;
   assign Interpolation_RAM_WR_Data[34] = 1'b0;
   assign Interpolation_RAM_WR_Data[33] = 1'b0;
   assign Interpolation_RAM_WR_Data[32] = 1'b0;
   assign Interpolation_RAM_WR_Data[31] = 1'b0;
   assign Interpolation_RAM_WR_Data[30] = 1'b0;
   assign Interpolation_RAM_WR_Data[29] = 1'b0;
   assign Interpolation_RAM_WR_Data[28] = 1'b0;
   assign Interpolation_RAM_WR_Data[27] = 1'b0;
   assign Interpolation_RAM_WR_Data[26] = 1'b0;
   assign Interpolation_RAM_WR_Data[25] = 1'b0;
   assign Interpolation_RAM_WR_Data[24] = 1'b0;
   assign Interpolation_RAM_WR_Data[23] = 1'b0;
   assign Interpolation_RAM_WR_Data[22] = 1'b0;
   assign Interpolation_RAM_WR_Data[21] = 1'b0;
   assign Interpolation_RAM_WR_Data[20] = 1'b0;
   assign Interpolation_RAM_WR_Data[19] = 1'b0;
   assign Interpolation_RAM_WR_Data[18] = 1'b0;
   assign Interpolation_RAM_WR_Data[17] = 1'b0;
   assign Interpolation_RAM_WR_Data[16] = 1'b0;

   DFF_X1 \UN_reg[15]  (.D(n_0_51), .CK(CLK), .Q(UN[15]), .QN());
   DFF_X1 \UN_reg[14]  (.D(n_0_50), .CK(CLK), .Q(UN[14]), .QN());
   DFF_X1 \UN_reg[13]  (.D(n_0_49), .CK(CLK), .Q(UN[13]), .QN());
   DFF_X1 \UN_reg[12]  (.D(n_0_48), .CK(CLK), .Q(UN[12]), .QN());
   DFF_X1 \UN_reg[11]  (.D(n_0_47), .CK(CLK), .Q(UN[11]), .QN());
   DFF_X1 \UN_reg[10]  (.D(n_0_46), .CK(CLK), .Q(UN[10]), .QN());
   DFF_X1 \UN_reg[9]  (.D(n_0_45), .CK(CLK), .Q(UN[9]), .QN());
   DFF_X1 \UN_reg[8]  (.D(n_0_44), .CK(CLK), .Q(UN[8]), .QN());
   DFF_X1 \UN_reg[7]  (.D(n_0_43), .CK(CLK), .Q(UN[7]), .QN());
   DFF_X1 \UN_reg[6]  (.D(n_0_42), .CK(CLK), .Q(UN[6]), .QN());
   DFF_X1 \UN_reg[5]  (.D(n_0_41), .CK(CLK), .Q(UN[5]), .QN());
   DFF_X1 \UN_reg[4]  (.D(n_0_40), .CK(CLK), .Q(UN[4]), .QN());
   DFF_X1 \UN_reg[3]  (.D(n_0_39), .CK(CLK), .Q(UN[3]), .QN());
   DFF_X1 \UN_reg[2]  (.D(n_0_38), .CK(CLK), .Q(UN[2]), .QN());
   DFF_X1 \UN_reg[1]  (.D(n_0_37), .CK(CLK), .Q(UN[1]), .QN());
   DFF_X1 \UN_reg[0]  (.D(n_0_36), .CK(CLK), .Q(UN[0]), .QN());
   DFF_X1 \intialization_state_reg[3]  (.D(n_0_86), .CK(CLK), .Q(
      intialization_state[3]), .QN());
   DFF_X1 \intialization_state_reg[2]  (.D(n_0_6), .CK(CLK), .Q(
      intialization_state[2]), .QN());
   DFF_X1 \intialization_state_reg[1]  (.D(n_0_5), .CK(CLK), .Q(
      intialization_state[1]), .QN());
   DFF_X1 \intialization_state_reg[0]  (.D(n_0_4), .CK(CLK), .Q(
      intialization_state[0]), .QN());
   DFF_X1 \Temp_reg[15]  (.D(n_0_83), .CK(CLK), .Q(Temp[15]), .QN());
   DFF_X1 \Temp_reg[14]  (.D(n_0_82), .CK(CLK), .Q(Temp[14]), .QN());
   DFF_X1 \Temp_reg[13]  (.D(n_0_81), .CK(CLK), .Q(Temp[13]), .QN());
   DFF_X1 \Temp_reg[12]  (.D(n_0_80), .CK(CLK), .Q(Temp[12]), .QN());
   DFF_X1 \Temp_reg[11]  (.D(n_0_79), .CK(CLK), .Q(Temp[11]), .QN());
   DFF_X1 \Temp_reg[10]  (.D(n_0_78), .CK(CLK), .Q(Temp[10]), .QN());
   DFF_X1 \Temp_reg[9]  (.D(n_0_77), .CK(CLK), .Q(Temp[9]), .QN());
   DFF_X1 \Temp_reg[8]  (.D(n_0_76), .CK(CLK), .Q(Temp[8]), .QN());
   DFF_X1 \Temp_reg[7]  (.D(n_0_75), .CK(CLK), .Q(Temp[7]), .QN());
   DFF_X1 \Temp_reg[6]  (.D(n_0_74), .CK(CLK), .Q(Temp[6]), .QN());
   DFF_X1 \Temp_reg[5]  (.D(n_0_73), .CK(CLK), .Q(Temp[5]), .QN());
   DFF_X1 \Temp_reg[4]  (.D(n_0_72), .CK(CLK), .Q(Temp[4]), .QN());
   DFF_X1 \Temp_reg[3]  (.D(n_0_71), .CK(CLK), .Q(Temp[3]), .QN());
   DFF_X1 \Temp_reg[2]  (.D(n_0_70), .CK(CLK), .Q(Temp[2]), .QN());
   DFF_X1 \Temp_reg[1]  (.D(n_0_69), .CK(CLK), .Q(Temp[1]), .QN());
   DFF_X1 \Temp_reg[0]  (.D(n_0_68), .CK(CLK), .Q(Temp[0]), .QN());
   DFF_X1 Intialization_Done_reg (.D(n_0_94), .CK(CLK), .Q(Intialization_Done), 
      .QN());
   DFF_X1 Interpolation_Done_reg (.D(n_0_95), .CK(CLK), .Q(Interpolation_Done), 
      .QN());
   DFF_X1 \UZ_ADD_reg[12]  (.D(n_93), .CK(n_0_2), .Q(UZ_ADD[12]), .QN());
   DFF_X1 \UZ_ADD_reg[11]  (.D(n_91), .CK(n_0_2), .Q(UZ_ADD[11]), .QN());
   DFF_X1 \UZ_ADD_reg[10]  (.D(n_89), .CK(n_0_2), .Q(UZ_ADD[10]), .QN());
   DFF_X1 \UZ_ADD_reg[9]  (.D(n_87), .CK(n_0_2), .Q(UZ_ADD[9]), .QN());
   DFF_X1 \UZ_ADD_reg[8]  (.D(n_85), .CK(n_0_2), .Q(UZ_ADD[8]), .QN());
   DFF_X1 \UZ_ADD_reg[7]  (.D(n_83), .CK(n_0_2), .Q(UZ_ADD[7]), .QN());
   DFF_X1 \UZ_ADD_reg[6]  (.D(n_0_34), .CK(n_0_2), .Q(UZ_ADD[6]), .QN());
   DFF_X1 \UZ_ADD_reg[5]  (.D(n_0_33), .CK(n_0_2), .Q(UZ_ADD[5]), .QN());
   DFF_X1 \UZ_ADD_reg[4]  (.D(n_77), .CK(n_0_2), .Q(UZ_ADD[4]), .QN());
   DFF_X1 \UZ_ADD_reg[3]  (.D(n_75), .CK(n_0_2), .Q(UZ_ADD[3]), .QN());
   DFF_X1 \UZ_ADD_reg[2]  (.D(n_0_32), .CK(n_0_2), .Q(UZ_ADD[2]), .QN());
   DFF_X1 \UZ_ADD_reg[1]  (.D(n_0_31), .CK(n_0_2), .Q(UZ_ADD[1]), .QN());
   DFF_X1 \UZ_ADD_reg[0]  (.D(n_5), .CK(n_0_2), .Q(UZ_ADD[0]), .QN());
   DFF_X1 \TZ_ADD_reg[12]  (.D(n_162), .CK(n_0_2), .Q(TZ_ADD[12]), .QN());
   DFF_X1 \TZ_ADD_reg[11]  (.D(n_161), .CK(n_0_2), .Q(TZ_ADD[11]), .QN());
   DFF_X1 \TZ_ADD_reg[10]  (.D(n_160), .CK(n_0_2), .Q(TZ_ADD[10]), .QN());
   DFF_X1 \TZ_ADD_reg[9]  (.D(n_159), .CK(n_0_2), .Q(TZ_ADD[9]), .QN());
   DFF_X1 \TZ_ADD_reg[8]  (.D(n_158), .CK(n_0_2), .Q(TZ_ADD[8]), .QN());
   DFF_X1 \TZ_ADD_reg[7]  (.D(n_157), .CK(n_0_2), .Q(TZ_ADD[7]), .QN());
   DFF_X1 \TZ_ADD_reg[6]  (.D(n_156), .CK(n_0_2), .Q(TZ_ADD[6]), .QN());
   DFF_X1 \TZ_ADD_reg[5]  (.D(n_155), .CK(n_0_2), .Q(TZ_ADD[5]), .QN());
   DFF_X1 \TZ_ADD_reg[4]  (.D(n_154), .CK(n_0_2), .Q(TZ_ADD[4]), .QN());
   DFF_X1 \TZ_ADD_reg[3]  (.D(n_153), .CK(n_0_2), .Q(TZ_ADD[3]), .QN());
   DFF_X1 \TZ_ADD_reg[2]  (.D(n_0_88), .CK(n_0_2), .Q(TZ_ADD[2]), .QN());
   DFF_X1 \TZ_ADD_reg[1]  (.D(n_151), .CK(n_0_2), .Q(TZ_ADD[1]), .QN());
   DFF_X1 \TZ_ADD_reg[0]  (.D(n_150), .CK(n_0_2), .Q(TZ_ADD[0]), .QN());
   CLKGATETST_X1 clk_gate_current_intialization_state_reg (.CK(CLK), .E(n_0_84), 
      .SE(1'b0), .GCK(n_0_0));
   DFF_X1 \current_intialization_state_reg[3]  (.D(n_0_14), .CK(n_0_0), .Q(
      current_intialization_state[3]), .QN());
   DFF_X1 \current_intialization_state_reg[2]  (.D(n_0_13), .CK(n_0_0), .Q(
      current_intialization_state[2]), .QN());
   DFF_X1 \current_intialization_state_reg[1]  (.D(n_0_12), .CK(n_0_0), .Q(
      current_intialization_state[1]), .QN());
   DFF_X1 \current_intialization_state_reg[0]  (.D(n_0_11), .CK(n_0_0), .Q(
      current_intialization_state[0]), .QN());
   CLKGATETST_X1 clk_gate_current_interpolation_state_reg (.CK(CLK), .E(n_0_85), 
      .SE(1'b0), .GCK(n_0_1));
   DFF_X1 \current_interpolation_state_reg[3]  (.D(n_0_10), .CK(n_0_1), .Q(
      current_interpolation_state[3]), .QN());
   DFF_X1 \current_interpolation_state_reg[2]  (.D(n_0_9), .CK(n_0_1), .Q(
      current_interpolation_state[2]), .QN());
   DFF_X1 \current_interpolation_state_reg[1]  (.D(n_0_8), .CK(n_0_1), .Q(
      current_interpolation_state[1]), .QN());
   DFF_X1 \current_interpolation_state_reg[0]  (.D(n_0_7), .CK(n_0_1), .Q(
      current_interpolation_state[0]), .QN());
   DFF_X1 \adder_sub1_In1_reg[15]  (.D(n_0_30), .CK(n_0_3), .Q(
      adder_sub1_In1[15]), .QN());
   DFF_X1 \adder_sub1_In1_reg[14]  (.D(n_0_29), .CK(n_0_3), .Q(
      adder_sub1_In1[14]), .QN());
   DFF_X1 \adder_sub1_In1_reg[13]  (.D(n_0_28), .CK(n_0_3), .Q(
      adder_sub1_In1[13]), .QN());
   DFF_X1 \adder_sub1_In1_reg[12]  (.D(n_0_27), .CK(n_0_3), .Q(
      adder_sub1_In1[12]), .QN());
   DFF_X1 \adder_sub1_In1_reg[11]  (.D(n_0_26), .CK(n_0_3), .Q(
      adder_sub1_In1[11]), .QN());
   DFF_X1 \adder_sub1_In1_reg[10]  (.D(n_0_25), .CK(n_0_3), .Q(
      adder_sub1_In1[10]), .QN());
   DFF_X1 \adder_sub1_In1_reg[9]  (.D(n_0_24), .CK(n_0_3), .Q(adder_sub1_In1[9]), 
      .QN());
   DFF_X1 \adder_sub1_In1_reg[8]  (.D(n_0_23), .CK(n_0_3), .Q(adder_sub1_In1[8]), 
      .QN());
   DFF_X1 \adder_sub1_In1_reg[7]  (.D(n_0_22), .CK(n_0_3), .Q(adder_sub1_In1[7]), 
      .QN());
   DFF_X1 \adder_sub1_In1_reg[6]  (.D(n_0_21), .CK(n_0_3), .Q(adder_sub1_In1[6]), 
      .QN());
   DFF_X1 \adder_sub1_In1_reg[5]  (.D(n_0_20), .CK(n_0_3), .Q(adder_sub1_In1[5]), 
      .QN());
   DFF_X1 \adder_sub1_In1_reg[4]  (.D(n_0_19), .CK(n_0_3), .Q(adder_sub1_In1[4]), 
      .QN());
   DFF_X1 \adder_sub1_In1_reg[3]  (.D(n_0_18), .CK(n_0_3), .Q(adder_sub1_In1[3]), 
      .QN());
   DFF_X1 \adder_sub1_In1_reg[2]  (.D(n_0_17), .CK(n_0_3), .Q(adder_sub1_In1[2]), 
      .QN());
   DFF_X1 \adder_sub1_In1_reg[1]  (.D(n_0_16), .CK(n_0_3), .Q(adder_sub1_In1[1]), 
      .QN());
   DFF_X1 \adder_sub1_In1_reg[0]  (.D(n_0_15), .CK(n_0_3), .Q(adder_sub1_In1[0]), 
      .QN());
   DFF_X1 \adder_sub1_In2_reg[15]  (.D(n_0_67), .CK(n_0_3), .Q(
      adder_sub1_In2[15]), .QN());
   DFF_X1 \adder_sub1_In2_reg[14]  (.D(n_0_66), .CK(n_0_3), .Q(
      adder_sub1_In2[14]), .QN());
   DFF_X1 \adder_sub1_In2_reg[13]  (.D(n_0_65), .CK(n_0_3), .Q(
      adder_sub1_In2[13]), .QN());
   DFF_X1 \adder_sub1_In2_reg[12]  (.D(n_0_64), .CK(n_0_3), .Q(
      adder_sub1_In2[12]), .QN());
   DFF_X1 \adder_sub1_In2_reg[11]  (.D(n_0_63), .CK(n_0_3), .Q(
      adder_sub1_In2[11]), .QN());
   DFF_X1 \adder_sub1_In2_reg[10]  (.D(n_0_62), .CK(n_0_3), .Q(
      adder_sub1_In2[10]), .QN());
   DFF_X1 \adder_sub1_In2_reg[9]  (.D(n_0_61), .CK(n_0_3), .Q(adder_sub1_In2[9]), 
      .QN());
   DFF_X1 \adder_sub1_In2_reg[8]  (.D(n_0_60), .CK(n_0_3), .Q(adder_sub1_In2[8]), 
      .QN());
   DFF_X1 \adder_sub1_In2_reg[7]  (.D(n_0_59), .CK(n_0_3), .Q(adder_sub1_In2[7]), 
      .QN());
   DFF_X1 \adder_sub1_In2_reg[6]  (.D(n_0_58), .CK(n_0_3), .Q(adder_sub1_In2[6]), 
      .QN());
   DFF_X1 \adder_sub1_In2_reg[5]  (.D(n_0_57), .CK(n_0_3), .Q(adder_sub1_In2[5]), 
      .QN());
   DFF_X1 \adder_sub1_In2_reg[4]  (.D(n_0_56), .CK(n_0_3), .Q(adder_sub1_In2[4]), 
      .QN());
   DFF_X1 \adder_sub1_In2_reg[3]  (.D(n_0_55), .CK(n_0_3), .Q(adder_sub1_In2[3]), 
      .QN());
   DFF_X1 \adder_sub1_In2_reg[2]  (.D(n_0_54), .CK(n_0_3), .Q(adder_sub1_In2[2]), 
      .QN());
   DFF_X1 \adder_sub1_In2_reg[1]  (.D(n_0_53), .CK(n_0_3), .Q(adder_sub1_In2[1]), 
      .QN());
   DFF_X1 \adder_sub1_In2_reg[0]  (.D(n_0_52), .CK(n_0_3), .Q(adder_sub1_In2[0]), 
      .QN());
   DFF_X1 Interpolation_Memory_WR_Enable_reg (.D(n_0_96), .CK(CLK), .Q(
      Interpolation_Memory_WR_Enable), .QN());
   CLKGATETST_X1 clk_gate_UZ_ADD_reg (.CK(CLK), .E(n_0_35), .SE(1'b0), .GCK(
      n_0_2));
   CLKGATETST_X1 clk_gate_adder_sub1_In1_reg (.CK(CLK), .E(n_4), .SE(1'b0), 
      .GCK(n_0_3));
   AND3_X1 i_0_0_0 (.A1(n_177), .A2(n_0_0_360), .A3(n_0_0_356), .ZN(n_0));
   AND3_X1 i_0_0_1 (.A1(n_0_0_394), .A2(n_177), .A3(n_0_0_255), .ZN(n_0_7));
   OAI33_X1 i_0_0_2 (.A1(n_0_0_260), .A2(n_0_0_3), .A3(RST), .B1(n_0_0_1), 
      .B2(n_0_0_349), .B3(n_0_0_359), .ZN(n_0_8));
   NOR2_X1 i_0_0_3 (.A1(n_0_0_1), .A2(n_0_0_0), .ZN(n_0_9));
   XNOR2_X1 i_0_0_4 (.A(n_0_0_396), .B(n_0_0_358), .ZN(n_0_0_0));
   NAND2_X1 i_0_0_5 (.A1(n_0_0_397), .A2(n_177), .ZN(n_0_0_1));
   AOI21_X1 i_0_0_6 (.A(RST), .B1(n_0_0_354), .B2(n_0_0_2), .ZN(n_0_10));
   NAND2_X1 i_0_0_7 (.A1(n_0_0_259), .A2(n_0_0_3), .ZN(n_0_0_2));
   AOI211_X1 i_0_0_8 (.A(n_176), .B(n_175), .C1(n_0_0_6), .C2(n_0_0_4), .ZN(
      n_0_0_3));
   OAI222_X1 i_0_0_9 (.A1(n_0_0_5), .A2(n_191), .B1(n_0_0_372), .B2(n_192), 
      .C1(n_193), .C2(n_0_0_373), .ZN(n_0_0_4));
   OAI21_X1 i_0_0_10 (.A(n_172), .B1(n_173), .B2(n_0_0_399), .ZN(n_0_0_5));
   NAND2_X1 i_0_0_11 (.A1(n_0_0_373), .A2(n_193), .ZN(n_0_0_6));
   NOR3_X1 i_0_0_12 (.A1(RST), .A2(n_0_0_407), .A3(n_0_0_363), .ZN(n_1));
   NOR4_X1 i_0_0_13 (.A1(RST), .A2(current_intialization_state[0]), .A3(n_0_0_8), 
      .A4(n_0_0_7), .ZN(n_0_11));
   AOI211_X1 i_0_0_14 (.A(current_intialization_state[1]), .B(n_0_0_393), 
      .C1(div1_ready), .C2(Div_Count), .ZN(n_0_0_7));
   AOI211_X1 i_0_0_15 (.A(RST), .B(n_0_0_8), .C1(n_0_0_314), .C2(n_0_0_378), 
      .ZN(n_0_12));
   NOR2_X1 i_0_0_16 (.A1(n_0_0_9), .A2(n_0_0_393), .ZN(n_0_0_8));
   NOR2_X1 i_0_0_17 (.A1(current_intialization_state[2]), .A2(n_0_0_14), 
      .ZN(n_0_0_9));
   NOR2_X1 i_0_0_18 (.A1(RST), .A2(n_0_0_10), .ZN(n_0_13));
   AOI22_X1 i_0_0_19 (.A1(n_0_0_301), .A2(n_0_0_14), .B1(n_0_0_11), .B2(
      n_0_0_393), .ZN(n_0_0_10));
   XNOR2_X1 i_0_0_20 (.A(current_intialization_state[2]), .B(n_0_0_364), 
      .ZN(n_0_0_11));
   NOR2_X1 i_0_0_21 (.A1(RST), .A2(n_0_0_12), .ZN(n_0_14));
   AOI21_X1 i_0_0_22 (.A(n_0_0_351), .B1(n_0_0_13), .B2(n_0_0_364), .ZN(n_0_0_12));
   NOR3_X1 i_0_0_23 (.A1(n_0_0_14), .A2(n_0_0_368), .A3(n_0_0_253), .ZN(n_0_0_13));
   AOI21_X1 i_0_0_24 (.A(n_0_0_391), .B1(n_0_0_16), .B2(n_0_0_15), .ZN(n_0_0_14));
   AOI211_X1 i_0_0_25 (.A(USIZE[4]), .B(USIZE[3]), .C1(USIZE[2]), .C2(n_0_0_403), 
      .ZN(n_0_0_15));
   OAI21_X1 i_0_0_26 (.A(n_0_0_17), .B1(n_0_0_403), .B2(USIZE[2]), .ZN(n_0_0_16));
   OAI21_X1 i_0_0_27 (.A(n_0_0_18), .B1(adder_sub1_Out[1]), .B2(n_0_0_406), 
      .ZN(n_0_0_17));
   OAI211_X1 i_0_0_28 (.A(USIZE[0]), .B(n_0_0_401), .C1(n_0_0_402), .C2(USIZE[1]), 
      .ZN(n_0_0_18));
   NAND2_X1 i_0_0_29 (.A1(n_0_0_367), .A2(n_0_0_350), .ZN(n_2));
   OAI21_X1 i_0_0_30 (.A(n_0_0_19), .B1(n_0_0_224), .B2(RST), .ZN(n_3));
   NAND3_X1 i_0_0_31 (.A1(current_intialization_state[1]), .A2(n_0_0_340), 
      .A3(n_0_0_326), .ZN(n_0_0_19));
   NAND3_X1 i_0_0_32 (.A1(n_0_0_326), .A2(n_0_0_224), .A3(n_0_0_20), .ZN(n_4));
   OAI21_X1 i_0_0_33 (.A(n_0_0_377), .B1(n_0_0_340), .B2(n_0_0_278), .ZN(
      n_0_0_20));
   AOI21_X1 i_0_0_34 (.A(n_0_0_27), .B1(n_0_0_21), .B2(n_0_0_90), .ZN(n_0_15));
   AOI221_X1 i_0_0_35 (.A(n_0_0_22), .B1(n_0_0_158), .B2(UN[0]), .C1(UZ_ADD[0]), 
      .C2(n_0_0_133), .ZN(n_0_0_21));
   AOI21_X1 i_0_0_36 (.A(n_0_0_58), .B1(n_0_0_24), .B2(n_0_0_23), .ZN(n_0_0_22));
   AOI22_X1 i_0_0_37 (.A1(UZ_ADD[0]), .A2(n_0_0_136), .B1(n_0_0_57), .B2(
      Interpolation_RAM_RD2_Data[0]), .ZN(n_0_0_23));
   OAI21_X1 i_0_0_38 (.A(n_0_0_25), .B1(n_0_0_333), .B2(
      Interpolation_RAM_RD2_Data[0]), .ZN(n_0_0_24));
   INV_X1 i_0_0_39 (.A(n_0_0_26), .ZN(n_0_0_25));
   AOI22_X1 i_0_0_40 (.A1(Interpolation_RAM_RD1_Data[0]), .A2(n_0_0_313), 
      .B1(n_0_0_278), .B2(Count2[0]), .ZN(n_0_0_26));
   AOI21_X1 i_0_0_41 (.A(n_0_0_28), .B1(n_0_0_152), .B2(
      Interpolation_RAM_RD2_Data[0]), .ZN(n_0_0_27));
   AOI211_X1 i_0_0_42 (.A(n_0_0_47), .B(n_0_0_29), .C1(n_0_0_33), .C2(n_0_0_409), 
      .ZN(n_0_0_28));
   AOI221_X1 i_0_0_43 (.A(n_0_0_30), .B1(n_0_0_313), .B2(
      Interpolation_RAM_RD1_Data[0]), .C1(UZ_ADD[0]), .C2(n_0_0_317), .ZN(
      n_0_0_29));
   AOI22_X1 i_0_0_44 (.A1(n_0_0_337), .A2(n_0_0_31), .B1(n_0_0_194), .B2(
      Interpolation_Intialize), .ZN(n_0_0_30));
   AOI22_X1 i_0_0_45 (.A1(n_0_0_32), .A2(n_0_0_34), .B1(n_0_0_278), .B2(
      Count2[0]), .ZN(n_0_0_31));
   NOR2_X1 i_0_0_46 (.A1(n_0_0_194), .A2(n_0_0_33), .ZN(n_0_0_32));
   NAND2_X1 i_0_0_47 (.A1(n_0_0_339), .A2(Interpolation_RAM_RD2_Data[0]), 
      .ZN(n_0_0_33));
   OAI21_X1 i_0_0_48 (.A(n_0_0_225), .B1(n_0_0_376), .B2(
      current_intialization_state[0]), .ZN(n_0_0_34));
   AOI21_X1 i_0_0_49 (.A(n_0_0_39), .B1(n_0_0_35), .B2(n_0_0_338), .ZN(n_0_16));
   AOI221_X1 i_0_0_50 (.A(n_0_0_36), .B1(n_0_0_158), .B2(UN[1]), .C1(UZ_ADD[1]), 
      .C2(n_0_0_133), .ZN(n_0_0_35));
   NOR2_X1 i_0_0_51 (.A1(n_0_0_58), .A2(n_0_0_37), .ZN(n_0_0_36));
   AOI221_X1 i_0_0_52 (.A(n_0_0_38), .B1(n_0_0_57), .B2(
      Interpolation_RAM_RD2_Data[1]), .C1(UZ_ADD[1]), .C2(n_0_0_136), .ZN(
      n_0_0_37));
   AOI22_X1 i_0_0_53 (.A1(n_0_0_379), .A2(n_0_0_141), .B1(n_0_0_43), .B2(
      n_0_0_42), .ZN(n_0_0_38));
   AOI22_X1 i_0_0_54 (.A1(n_0_0_223), .A2(n_0_0_40), .B1(n_0_0_152), .B2(
      Interpolation_RAM_RD2_Data[1]), .ZN(n_0_0_39));
   AOI21_X1 i_0_0_55 (.A(n_0_0_48), .B1(n_0_0_41), .B2(n_0_0_42), .ZN(n_0_0_40));
   AOI221_X1 i_0_0_56 (.A(n_0_0_154), .B1(n_0_0_50), .B2(Count2[1]), .C1(
      n_0_0_317), .C2(UZ_ADD[1]), .ZN(n_0_0_41));
   NAND2_X1 i_0_0_57 (.A1(Interpolation_RAM_RD1_Data[1]), .A2(n_0_0_313), 
      .ZN(n_0_0_42));
   NAND2_X1 i_0_0_58 (.A1(Count2[1]), .A2(n_0_0_278), .ZN(n_0_0_43));
   AOI22_X1 i_0_0_59 (.A1(n_0_0_44), .A2(n_0_0_45), .B1(n_0_0_51), .B2(n_0_0_338), 
      .ZN(n_0_17));
   AOI21_X1 i_0_0_60 (.A(n_0_0_46), .B1(n_0_0_152), .B2(
      Interpolation_RAM_RD2_Data[2]), .ZN(n_0_0_44));
   NAND3_X1 i_0_0_61 (.A1(UZ_ADD[2]), .A2(n_0_0_317), .A3(n_0_0_223), .ZN(
      n_0_0_45));
   AOI211_X1 i_0_0_62 (.A(n_0_0_409), .B(n_0_0_47), .C1(n_0_0_49), .C2(n_0_0_337), 
      .ZN(n_0_0_46));
   OR2_X1 i_0_0_63 (.A1(RST), .A2(n_0_0_48), .ZN(n_0_0_47));
   NOR3_X1 i_0_0_64 (.A1(n_0_0_389), .A2(n_0_0_246), .A3(n_0_0_340), .ZN(
      n_0_0_48));
   AOI22_X1 i_0_0_65 (.A1(Interpolation_RAM_RD1_Data[2]), .A2(n_0_0_313), 
      .B1(n_0_0_50), .B2(Count2[2]), .ZN(n_0_0_49));
   AOI21_X1 i_0_0_66 (.A(n_0_0_277), .B1(n_0_0_194), .B2(Interpolation_Intialize), 
      .ZN(n_0_0_50));
   AOI221_X1 i_0_0_67 (.A(n_0_0_52), .B1(n_0_0_158), .B2(UN[2]), .C1(UZ_ADD[2]), 
      .C2(n_0_0_133), .ZN(n_0_0_51));
   AOI21_X1 i_0_0_68 (.A(n_0_0_58), .B1(n_0_0_54), .B2(n_0_0_53), .ZN(n_0_0_52));
   AOI22_X1 i_0_0_69 (.A1(UZ_ADD[2]), .A2(n_0_0_136), .B1(n_0_0_57), .B2(
      Interpolation_RAM_RD2_Data[2]), .ZN(n_0_0_53));
   OAI21_X1 i_0_0_70 (.A(n_0_0_55), .B1(n_0_0_333), .B2(
      Interpolation_RAM_RD2_Data[2]), .ZN(n_0_0_54));
   INV_X1 i_0_0_71 (.A(n_0_0_56), .ZN(n_0_0_55));
   AOI22_X1 i_0_0_72 (.A1(Interpolation_RAM_RD1_Data[2]), .A2(n_0_0_313), 
      .B1(n_0_0_278), .B2(Count2[2]), .ZN(n_0_0_56));
   OAI21_X1 i_0_0_73 (.A(n_0_0_220), .B1(n_0_0_308), .B2(n_0_0_333), .ZN(
      n_0_0_57));
   AOI21_X1 i_0_0_74 (.A(n_0_0_61), .B1(n_0_0_60), .B2(n_0_0_59), .ZN(n_0_0_58));
   AOI21_X1 i_0_0_75 (.A(n_0_0_332), .B1(n_0_0_334), .B2(n_0_0_407), .ZN(
      n_0_0_59));
   OAI21_X1 i_0_0_76 (.A(n_0_0_312), .B1(n_0_0_141), .B2(Interpolation_Intialize), 
      .ZN(n_0_0_60));
   AOI21_X1 i_0_0_77 (.A(n_0_0_329), .B1(n_0_0_307), .B2(n_0_0_220), .ZN(
      n_0_0_61));
   AOI21_X1 i_0_0_78 (.A(n_0_0_67), .B1(n_0_0_63), .B2(n_0_0_62), .ZN(n_0_18));
   AOI21_X1 i_0_0_79 (.A(n_0_0_64), .B1(n_0_0_91), .B2(
      Interpolation_RAM_RD2_Data[3]), .ZN(n_0_0_62));
   AOI221_X1 i_0_0_80 (.A(n_0_0_337), .B1(n_0_0_158), .B2(UN[3]), .C1(n_0_0_133), 
      .C2(UZ_ADD[3]), .ZN(n_0_0_63));
   AOI21_X1 i_0_0_81 (.A(n_0_0_65), .B1(n_0_0_66), .B2(n_0_0_162), .ZN(n_0_0_64));
   OAI21_X1 i_0_0_82 (.A(n_0_0_139), .B1(n_0_0_333), .B2(
      Interpolation_RAM_RD2_Data[3]), .ZN(n_0_0_65));
   AOI22_X1 i_0_0_83 (.A1(Interpolation_RAM_RD1_Data[3]), .A2(n_0_0_313), 
      .B1(n_0_0_136), .B2(UZ_ADD[3]), .ZN(n_0_0_66));
   AOI22_X1 i_0_0_84 (.A1(Interpolation_RAM_RD2_Data[3]), .A2(n_0_0_152), 
      .B1(n_0_0_68), .B2(n_0_0_223), .ZN(n_0_0_67));
   NAND2_X1 i_0_0_85 (.A1(n_0_0_69), .A2(n_0_0_337), .ZN(n_0_0_68));
   AOI22_X1 i_0_0_86 (.A1(UZ_ADD[3]), .A2(n_0_0_317), .B1(n_0_0_313), .B2(
      Interpolation_RAM_RD1_Data[3]), .ZN(n_0_0_69));
   OAI211_X1 i_0_0_87 (.A(n_0_0_73), .B(n_0_0_70), .C1(n_0_0_71), .C2(n_0_0_335), 
      .ZN(n_0_19));
   AOI222_X1 i_0_0_88 (.A1(UZ_ADD[4]), .A2(n_0_0_129), .B1(n_0_0_126), .B2(
      Interpolation_RAM_RD1_Data[4]), .C1(n_0_0_119), .C2(UN[4]), .ZN(n_0_0_70));
   AOI21_X1 i_0_0_89 (.A(n_0_0_72), .B1(n_0_0_133), .B2(UZ_ADD[4]), .ZN(n_0_0_71));
   NOR3_X1 i_0_0_90 (.A1(n_0_0_332), .A2(n_0_0_75), .A3(n_0_0_141), .ZN(n_0_0_72));
   OAI21_X1 i_0_0_91 (.A(Interpolation_RAM_RD2_Data[4]), .B1(n_0_0_150), 
      .B2(n_0_0_74), .ZN(n_0_0_73));
   AOI21_X1 i_0_0_92 (.A(n_0_0_410), .B1(n_0_0_75), .B2(n_0_0_220), .ZN(n_0_0_74));
   AOI221_X1 i_0_0_93 (.A(n_0_0_163), .B1(n_0_0_136), .B2(UZ_ADD[4]), .C1(
      Interpolation_RAM_RD1_Data[4]), .C2(n_0_0_313), .ZN(n_0_0_75));
   NAND2_X1 i_0_0_94 (.A1(n_0_0_81), .A2(n_0_0_76), .ZN(n_0_20));
   AOI221_X1 i_0_0_95 (.A(n_0_0_77), .B1(n_0_0_150), .B2(
      Interpolation_RAM_RD2_Data[5]), .C1(UZ_ADD[5]), .C2(n_0_0_129), .ZN(
      n_0_0_76));
   AOI21_X1 i_0_0_96 (.A(n_0_0_335), .B1(n_0_0_79), .B2(n_0_0_78), .ZN(n_0_0_77));
   OAI211_X1 i_0_0_97 (.A(Interpolation_RAM_RD2_Data[5]), .B(n_0_0_139), 
      .C1(n_0_0_137), .C2(n_0_0_82), .ZN(n_0_0_78));
   AOI211_X1 i_0_0_98 (.A(n_0_0_332), .B(n_0_0_80), .C1(n_0_0_133), .C2(
      UZ_ADD[5]), .ZN(n_0_0_79));
   NOR2_X1 i_0_0_99 (.A1(n_0_0_83), .A2(n_0_0_141), .ZN(n_0_0_80));
   AOI22_X1 i_0_0_100 (.A1(Interpolation_RAM_RD1_Data[5]), .A2(n_0_0_126), 
      .B1(n_0_0_119), .B2(UN[5]), .ZN(n_0_0_81));
   INV_X1 i_0_0_101 (.A(n_0_0_83), .ZN(n_0_0_82));
   AOI22_X1 i_0_0_102 (.A1(Interpolation_RAM_RD1_Data[5]), .A2(n_0_0_313), 
      .B1(n_0_0_136), .B2(UZ_ADD[5]), .ZN(n_0_0_83));
   AOI21_X1 i_0_0_103 (.A(n_0_0_87), .B1(n_0_0_84), .B2(n_0_0_335), .ZN(n_0_21));
   AOI22_X1 i_0_0_104 (.A1(Interpolation_RAM_RD2_Data[6]), .A2(n_0_0_152), 
      .B1(n_0_0_85), .B2(n_0_0_223), .ZN(n_0_0_84));
   INV_X1 i_0_0_105 (.A(n_0_0_86), .ZN(n_0_0_85));
   AOI22_X1 i_0_0_106 (.A1(UZ_ADD[6]), .A2(n_0_0_317), .B1(n_0_0_313), .B2(
      Interpolation_RAM_RD1_Data[6]), .ZN(n_0_0_86));
   AOI21_X1 i_0_0_107 (.A(n_0_0_88), .B1(n_0_0_91), .B2(
      Interpolation_RAM_RD2_Data[6]), .ZN(n_0_0_87));
   OAI211_X1 i_0_0_108 (.A(n_0_0_90), .B(n_0_0_89), .C1(n_0_0_93), .C2(n_0_0_92), 
      .ZN(n_0_0_88));
   AOI22_X1 i_0_0_109 (.A1(UN[6]), .A2(n_0_0_158), .B1(n_0_0_133), .B2(UZ_ADD[6]), 
      .ZN(n_0_0_89));
   NOR2_X1 i_0_0_110 (.A1(n_0_0_357), .A2(n_0_0_344), .ZN(n_0_0_90));
   NOR3_X1 i_0_0_111 (.A1(n_0_0_332), .A2(n_0_0_158), .A3(n_0_0_220), .ZN(
      n_0_0_91));
   OAI21_X1 i_0_0_112 (.A(n_0_0_139), .B1(n_0_0_333), .B2(
      Interpolation_RAM_RD2_Data[6]), .ZN(n_0_0_92));
   AOI221_X1 i_0_0_113 (.A(n_0_0_163), .B1(n_0_0_136), .B2(UZ_ADD[6]), .C1(
      Interpolation_RAM_RD1_Data[6]), .C2(n_0_0_313), .ZN(n_0_0_93));
   NAND2_X1 i_0_0_114 (.A1(n_0_0_95), .A2(n_0_0_94), .ZN(n_0_22));
   AOI222_X1 i_0_0_115 (.A1(UZ_ADD[7]), .A2(n_0_0_124), .B1(n_0_0_123), .B2(
      n_0_0_96), .C1(Interpolation_RAM_RD2_Data[7]), .C2(n_0_0_219), .ZN(
      n_0_0_94));
   AOI22_X1 i_0_0_116 (.A1(Interpolation_RAM_RD1_Data[7]), .A2(n_0_0_126), 
      .B1(n_0_0_119), .B2(UN[7]), .ZN(n_0_0_95));
   AOI21_X1 i_0_0_117 (.A(n_0_0_97), .B1(n_0_0_98), .B2(n_0_0_162), .ZN(n_0_0_96));
   NOR2_X1 i_0_0_118 (.A1(n_0_0_333), .A2(Interpolation_RAM_RD2_Data[7]), 
      .ZN(n_0_0_97));
   AOI22_X1 i_0_0_119 (.A1(Interpolation_RAM_RD1_Data[7]), .A2(n_0_0_313), 
      .B1(n_0_0_136), .B2(UZ_ADD[7]), .ZN(n_0_0_98));
   NAND2_X1 i_0_0_120 (.A1(n_0_0_100), .A2(n_0_0_99), .ZN(n_0_23));
   AOI222_X1 i_0_0_121 (.A1(n_0_0_101), .A2(n_0_0_336), .B1(
      Interpolation_RAM_RD2_Data[8]), .B2(n_0_0_150), .C1(n_0_0_129), .C2(
      UZ_ADD[8]), .ZN(n_0_0_99));
   AOI22_X1 i_0_0_122 (.A1(Interpolation_RAM_RD1_Data[8]), .A2(n_0_0_126), 
      .B1(n_0_0_119), .B2(UN[8]), .ZN(n_0_0_100));
   OAI21_X1 i_0_0_123 (.A(n_0_0_102), .B1(n_0_0_103), .B2(n_0_0_104), .ZN(
      n_0_0_101));
   AOI21_X1 i_0_0_124 (.A(n_0_0_332), .B1(n_0_0_133), .B2(UZ_ADD[8]), .ZN(
      n_0_0_102));
   AOI221_X1 i_0_0_125 (.A(n_0_0_137), .B1(n_0_0_136), .B2(UZ_ADD[8]), .C1(
      Interpolation_RAM_RD1_Data[8]), .C2(n_0_0_313), .ZN(n_0_0_103));
   AOI21_X1 i_0_0_126 (.A(n_0_0_140), .B1(n_0_0_139), .B2(
      Interpolation_RAM_RD2_Data[8]), .ZN(n_0_0_104));
   OAI211_X1 i_0_0_127 (.A(n_0_0_106), .B(n_0_0_105), .C1(n_0_0_107), .C2(
      n_0_0_335), .ZN(n_0_24));
   AOI22_X1 i_0_0_128 (.A1(Interpolation_RAM_RD2_Data[9]), .A2(n_0_0_150), 
      .B1(n_0_0_126), .B2(Interpolation_RAM_RD1_Data[9]), .ZN(n_0_0_105));
   NAND2_X1 i_0_0_129 (.A1(UZ_ADD[9]), .A2(n_0_0_129), .ZN(n_0_0_106));
   AOI221_X1 i_0_0_130 (.A(n_0_0_108), .B1(n_0_0_158), .B2(UN[9]), .C1(UZ_ADD[9]), 
      .C2(n_0_0_133), .ZN(n_0_0_107));
   NOR2_X1 i_0_0_131 (.A1(n_0_0_110), .A2(n_0_0_109), .ZN(n_0_0_108));
   AOI221_X1 i_0_0_132 (.A(n_0_0_137), .B1(n_0_0_136), .B2(UZ_ADD[9]), .C1(
      Interpolation_RAM_RD1_Data[9]), .C2(n_0_0_313), .ZN(n_0_0_109));
   AOI21_X1 i_0_0_133 (.A(n_0_0_140), .B1(n_0_0_139), .B2(
      Interpolation_RAM_RD2_Data[9]), .ZN(n_0_0_110));
   NAND4_X1 i_0_0_134 (.A1(n_0_0_113), .A2(n_0_0_111), .A3(n_0_0_112), .A4(
      n_0_0_116), .ZN(n_0_25));
   AOI22_X1 i_0_0_135 (.A1(n_0_0_219), .A2(Interpolation_RAM_RD2_Data[10]), 
      .B1(UN[10]), .B2(n_0_0_119), .ZN(n_0_0_111));
   NAND3_X1 i_0_0_136 (.A1(Interpolation_RAM_RD1_Data[10]), .A2(n_0_0_313), 
      .A3(n_0_0_130), .ZN(n_0_0_112));
   OAI211_X1 i_0_0_137 (.A(n_0_0_123), .B(n_0_0_114), .C1(
      Interpolation_RAM_RD2_Data[10]), .C2(n_0_0_333), .ZN(n_0_0_113));
   NAND2_X1 i_0_0_138 (.A1(n_0_0_115), .A2(n_0_0_162), .ZN(n_0_0_114));
   AOI22_X1 i_0_0_139 (.A1(Interpolation_RAM_RD1_Data[10]), .A2(n_0_0_313), 
      .B1(n_0_0_136), .B2(UZ_ADD[10]), .ZN(n_0_0_115));
   NAND2_X1 i_0_0_140 (.A1(n_0_0_124), .A2(UZ_ADD[10]), .ZN(n_0_0_116));
   NAND2_X1 i_0_0_141 (.A1(n_0_0_118), .A2(n_0_0_117), .ZN(n_0_26));
   AOI222_X1 i_0_0_142 (.A1(UZ_ADD[11]), .A2(n_0_0_124), .B1(n_0_0_123), 
      .B2(n_0_0_120), .C1(Interpolation_RAM_RD2_Data[11]), .C2(n_0_0_219), 
      .ZN(n_0_0_117));
   AOI22_X1 i_0_0_143 (.A1(Interpolation_RAM_RD1_Data[11]), .A2(n_0_0_126), 
      .B1(n_0_0_119), .B2(UN[11]), .ZN(n_0_0_118));
   NOR2_X1 i_0_0_144 (.A1(n_0_0_335), .A2(n_0_0_157), .ZN(n_0_0_119));
   AOI21_X1 i_0_0_145 (.A(n_0_0_121), .B1(n_0_0_122), .B2(n_0_0_162), .ZN(
      n_0_0_120));
   NOR2_X1 i_0_0_146 (.A1(n_0_0_333), .A2(Interpolation_RAM_RD2_Data[11]), 
      .ZN(n_0_0_121));
   AOI22_X1 i_0_0_147 (.A1(Interpolation_RAM_RD1_Data[11]), .A2(n_0_0_313), 
      .B1(n_0_0_136), .B2(UZ_ADD[11]), .ZN(n_0_0_122));
   AND2_X1 i_0_0_148 (.A1(n_0_0_336), .A2(n_0_0_139), .ZN(n_0_0_123));
   OAI21_X1 i_0_0_149 (.A(n_0_0_128), .B1(n_0_0_132), .B2(n_0_0_335), .ZN(
      n_0_0_124));
   OAI211_X1 i_0_0_150 (.A(n_0_0_127), .B(n_0_0_125), .C1(n_0_0_131), .C2(
      n_0_0_335), .ZN(n_0_27));
   AOI22_X1 i_0_0_151 (.A1(Interpolation_RAM_RD2_Data[12]), .A2(n_0_0_150), 
      .B1(n_0_0_126), .B2(Interpolation_RAM_RD1_Data[12]), .ZN(n_0_0_125));
   NOR3_X1 i_0_0_152 (.A1(n_0_0_154), .A2(RST), .A3(n_0_0_312), .ZN(n_0_0_126));
   NAND2_X1 i_0_0_153 (.A1(UZ_ADD[12]), .A2(n_0_0_129), .ZN(n_0_0_127));
   INV_X1 i_0_0_154 (.A(n_0_0_129), .ZN(n_0_0_128));
   AND2_X1 i_0_0_155 (.A1(n_0_0_317), .A2(n_0_0_130), .ZN(n_0_0_129));
   NOR2_X1 i_0_0_156 (.A1(n_0_0_154), .A2(RST), .ZN(n_0_0_130));
   AOI221_X1 i_0_0_157 (.A(n_0_0_134), .B1(n_0_0_133), .B2(UZ_ADD[12]), .C1(
      UN[12]), .C2(n_0_0_158), .ZN(n_0_0_131));
   INV_X1 i_0_0_158 (.A(n_0_0_133), .ZN(n_0_0_132));
   NOR2_X1 i_0_0_159 (.A1(n_0_0_329), .A2(n_0_0_339), .ZN(n_0_0_133));
   NOR2_X1 i_0_0_160 (.A1(n_0_0_138), .A2(n_0_0_135), .ZN(n_0_0_134));
   AOI221_X1 i_0_0_161 (.A(n_0_0_137), .B1(n_0_0_136), .B2(UZ_ADD[12]), .C1(
      Interpolation_RAM_RD1_Data[12]), .C2(n_0_0_313), .ZN(n_0_0_135));
   NOR2_X1 i_0_0_162 (.A1(n_0_0_334), .A2(n_0_0_307), .ZN(n_0_0_136));
   NAND2_X1 i_0_0_163 (.A1(n_0_0_220), .A2(n_0_0_162), .ZN(n_0_0_137));
   AOI21_X1 i_0_0_164 (.A(n_0_0_140), .B1(n_0_0_139), .B2(
      Interpolation_RAM_RD2_Data[12]), .ZN(n_0_0_138));
   NOR3_X1 i_0_0_165 (.A1(n_0_0_332), .A2(n_0_0_283), .A3(n_0_0_158), .ZN(
      n_0_0_139));
   NOR3_X1 i_0_0_166 (.A1(n_0_0_141), .A2(n_0_0_221), .A3(n_0_0_332), .ZN(
      n_0_0_140));
   OAI21_X1 i_0_0_167 (.A(n_0_0_333), .B1(n_0_0_376), .B2(
      current_intialization_state[1]), .ZN(n_0_0_141));
   OAI21_X1 i_0_0_168 (.A(n_0_0_142), .B1(n_0_0_144), .B2(n_0_0_143), .ZN(n_0_28));
   AOI22_X1 i_0_0_169 (.A1(Interpolation_RAM_RD1_Data[13]), .A2(n_0_0_153), 
      .B1(n_0_0_149), .B2(Interpolation_RAM_RD2_Data[13]), .ZN(n_0_0_142));
   OAI221_X1 i_0_0_170 (.A(n_0_0_159), .B1(n_0_0_157), .B2(UN[13]), .C1(
      n_0_0_161), .C2(Interpolation_RAM_RD2_Data[13]), .ZN(n_0_0_143));
   AOI221_X1 i_0_0_171 (.A(n_0_0_334), .B1(n_0_0_221), .B2(
      Interpolation_RAM_RD2_Data[13]), .C1(n_0_0_160), .C2(
      Interpolation_RAM_RD1_Data[13]), .ZN(n_0_0_144));
   OAI21_X1 i_0_0_172 (.A(n_0_0_145), .B1(n_0_0_147), .B2(n_0_0_146), .ZN(n_0_29));
   AOI22_X1 i_0_0_173 (.A1(Interpolation_RAM_RD1_Data[14]), .A2(n_0_0_153), 
      .B1(n_0_0_149), .B2(Interpolation_RAM_RD2_Data[14]), .ZN(n_0_0_145));
   OAI221_X1 i_0_0_174 (.A(n_0_0_159), .B1(n_0_0_157), .B2(UN[14]), .C1(
      n_0_0_161), .C2(Interpolation_RAM_RD2_Data[14]), .ZN(n_0_0_146));
   AOI221_X1 i_0_0_175 (.A(n_0_0_334), .B1(n_0_0_221), .B2(
      Interpolation_RAM_RD2_Data[14]), .C1(n_0_0_160), .C2(
      Interpolation_RAM_RD1_Data[14]), .ZN(n_0_0_147));
   OAI21_X1 i_0_0_176 (.A(n_0_0_148), .B1(n_0_0_156), .B2(n_0_0_155), .ZN(n_0_30));
   AOI22_X1 i_0_0_177 (.A1(Interpolation_RAM_RD1_Data[15]), .A2(n_0_0_153), 
      .B1(n_0_0_149), .B2(Interpolation_RAM_RD2_Data[15]), .ZN(n_0_0_148));
   AOI21_X1 i_0_0_178 (.A(n_0_0_151), .B1(n_0_0_249), .B2(n_0_0_338), .ZN(
      n_0_0_149));
   NOR2_X1 i_0_0_179 (.A1(n_0_0_338), .A2(n_0_0_151), .ZN(n_0_0_150));
   INV_X1 i_0_0_180 (.A(n_0_0_152), .ZN(n_0_0_151));
   AOI21_X1 i_0_0_181 (.A(RST), .B1(n_0_0_224), .B2(n_0_0_220), .ZN(n_0_0_152));
   AOI211_X1 i_0_0_182 (.A(n_0_0_312), .B(RST), .C1(n_0_0_154), .C2(n_0_0_249), 
      .ZN(n_0_0_153));
   NAND2_X1 i_0_0_183 (.A1(n_0_0_337), .A2(n_0_0_224), .ZN(n_0_0_154));
   OAI221_X1 i_0_0_184 (.A(n_0_0_159), .B1(n_0_0_157), .B2(UN[15]), .C1(
      n_0_0_161), .C2(Interpolation_RAM_RD2_Data[15]), .ZN(n_0_0_155));
   AOI221_X1 i_0_0_185 (.A(n_0_0_334), .B1(n_0_0_221), .B2(
      Interpolation_RAM_RD2_Data[15]), .C1(n_0_0_160), .C2(
      Interpolation_RAM_RD1_Data[15]), .ZN(n_0_0_156));
   OAI21_X1 i_0_0_186 (.A(n_0_0_334), .B1(n_0_0_312), .B2(n_0_0_407), .ZN(
      n_0_0_157));
   NOR2_X1 i_0_0_187 (.A1(n_0_0_185), .A2(n_0_0_333), .ZN(n_0_0_158));
   NOR3_X1 i_0_0_188 (.A1(n_0_0_194), .A2(n_0_0_332), .A3(RST), .ZN(n_0_0_159));
   AOI211_X1 i_0_0_189 (.A(n_0_0_298), .B(n_0_0_312), .C1(n_0_0_345), .C2(
      n_0_0_346), .ZN(n_0_0_160));
   NAND2_X1 i_0_0_190 (.A1(n_0_0_334), .A2(n_0_0_185), .ZN(n_0_0_161));
   NAND2_X1 i_0_0_191 (.A1(n_0_0_334), .A2(n_0_0_313), .ZN(n_0_0_162));
   NOR2_X1 i_0_0_192 (.A1(n_0_0_333), .A2(n_0_0_312), .ZN(n_0_0_163));
   NAND2_X1 i_0_0_193 (.A1(n_0_0_401), .A2(n_177), .ZN(n_5));
   NAND2_X1 i_0_0_194 (.A1(n_0_0_402), .A2(n_177), .ZN(n_0_31));
   NAND2_X1 i_0_0_195 (.A1(n_0_0_403), .A2(n_177), .ZN(n_0_32));
   NAND2_X1 i_0_0_196 (.A1(n_0_0_404), .A2(n_177), .ZN(n_0_33));
   NAND2_X1 i_0_0_197 (.A1(n_0_0_405), .A2(n_177), .ZN(n_0_34));
   NAND2_X1 i_0_0_198 (.A1(n_177), .A2(n_0_0_374), .ZN(n_0_35));
   OAI22_X1 i_0_0_199 (.A1(n_0_0_287), .A2(n_0_0_165), .B1(n_0_0_164), .B2(
      n_0_0_398), .ZN(n_6));
   NOR3_X1 i_0_0_200 (.A1(RST), .A2(Interpolation_Enable), .A3(n_0_0_287), 
      .ZN(n_7));
   OAI22_X1 i_0_0_201 (.A1(n_0_0_290), .A2(n_0_0_165), .B1(n_0_0_164), .B2(
      n_0_0_399), .ZN(n_8));
   NOR3_X1 i_0_0_202 (.A1(RST), .A2(Interpolation_Enable), .A3(n_0_0_290), 
      .ZN(n_9));
   OAI22_X1 i_0_0_203 (.A1(n_0_0_296), .A2(n_0_0_165), .B1(n_0_0_164), .B2(
      n_0_0_400), .ZN(n_10));
   NAND3_X1 i_0_0_204 (.A1(n_0_0_259), .A2(n_0_0_356), .A3(n_177), .ZN(n_0_0_164));
   NAND2_X1 i_0_0_205 (.A1(n_0_0_258), .A2(n_0_0_361), .ZN(n_0_0_165));
   NOR3_X1 i_0_0_206 (.A1(RST), .A2(Interpolation_Enable), .A3(n_0_0_296), 
      .ZN(n_11));
   INV_X1 i_0_0_207 (.A(n_0_0_166), .ZN(n_0_36));
   AOI22_X1 i_0_0_208 (.A1(UN[0]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[0]), .ZN(n_0_0_166));
   INV_X1 i_0_0_209 (.A(n_0_0_167), .ZN(n_0_37));
   AOI22_X1 i_0_0_210 (.A1(UN[1]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[1]), .ZN(n_0_0_167));
   INV_X1 i_0_0_211 (.A(n_0_0_168), .ZN(n_0_38));
   AOI22_X1 i_0_0_212 (.A1(UN[2]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[2]), .ZN(n_0_0_168));
   INV_X1 i_0_0_213 (.A(n_0_0_169), .ZN(n_0_39));
   AOI22_X1 i_0_0_214 (.A1(UN[3]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[3]), .ZN(n_0_0_169));
   INV_X1 i_0_0_215 (.A(n_0_0_170), .ZN(n_0_40));
   AOI22_X1 i_0_0_216 (.A1(UN[4]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[4]), .ZN(n_0_0_170));
   INV_X1 i_0_0_217 (.A(n_0_0_171), .ZN(n_0_41));
   AOI22_X1 i_0_0_218 (.A1(UN[5]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[5]), .ZN(n_0_0_171));
   INV_X1 i_0_0_219 (.A(n_0_0_172), .ZN(n_0_42));
   AOI22_X1 i_0_0_220 (.A1(UN[6]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[6]), .ZN(n_0_0_172));
   INV_X1 i_0_0_221 (.A(n_0_0_173), .ZN(n_0_43));
   AOI22_X1 i_0_0_222 (.A1(UN[7]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[7]), .ZN(n_0_0_173));
   INV_X1 i_0_0_223 (.A(n_0_0_174), .ZN(n_0_44));
   AOI22_X1 i_0_0_224 (.A1(UN[8]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[8]), .ZN(n_0_0_174));
   INV_X1 i_0_0_225 (.A(n_0_0_175), .ZN(n_0_45));
   AOI22_X1 i_0_0_226 (.A1(UN[9]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[9]), .ZN(n_0_0_175));
   INV_X1 i_0_0_227 (.A(n_0_0_176), .ZN(n_0_46));
   AOI22_X1 i_0_0_228 (.A1(UN[10]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[10]), .ZN(n_0_0_176));
   INV_X1 i_0_0_229 (.A(n_0_0_177), .ZN(n_0_47));
   AOI22_X1 i_0_0_230 (.A1(UN[11]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[11]), .ZN(n_0_0_177));
   INV_X1 i_0_0_231 (.A(n_0_0_178), .ZN(n_0_48));
   AOI22_X1 i_0_0_232 (.A1(UN[12]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[12]), .ZN(n_0_0_178));
   INV_X1 i_0_0_233 (.A(n_0_0_179), .ZN(n_0_49));
   AOI22_X1 i_0_0_234 (.A1(UN[13]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[13]), .ZN(n_0_0_179));
   INV_X1 i_0_0_235 (.A(n_0_0_180), .ZN(n_0_50));
   AOI22_X1 i_0_0_236 (.A1(UN[14]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[14]), .ZN(n_0_0_180));
   INV_X1 i_0_0_237 (.A(n_0_0_181), .ZN(n_0_51));
   AOI22_X1 i_0_0_238 (.A1(UN[15]), .A2(n_0_0_183), .B1(n_0_0_182), .B2(
      Interpolation_RAM_RD2_Data[15]), .ZN(n_0_0_181));
   NOR2_X1 i_0_0_239 (.A1(RST), .A2(n_0_0_184), .ZN(n_0_0_182));
   NOR2_X1 i_0_0_240 (.A1(n_50), .A2(n_0_0_185), .ZN(n_0_0_183));
   NOR2_X1 i_0_0_241 (.A1(n_0_0_248), .A2(n_0_0_185), .ZN(n_0_0_184));
   NOR2_X1 i_0_0_242 (.A1(n_0_0_312), .A2(n_0_0_407), .ZN(n_0_0_185));
   OAI21_X1 i_0_0_243 (.A(n_0_0_195), .B1(n_0_0_186), .B2(RST), .ZN(n_0_52));
   AOI22_X1 i_0_0_244 (.A1(n_0_0_194), .A2(n_0_0_192), .B1(n_0_0_188), .B2(
      n_0_0_187), .ZN(n_0_0_186));
   OAI211_X1 i_0_0_245 (.A(n_0_0_395), .B(n_0_0_344), .C1(n_0_0_194), .C2(
      n_0_0_381), .ZN(n_0_0_187));
   NAND2_X1 i_0_0_246 (.A1(n_0_0_189), .A2(n_0_0_225), .ZN(n_0_0_188));
   AOI221_X1 i_0_0_247 (.A(n_0_0_191), .B1(n_0_0_190), .B2(n_0_0_192), .C1(
      n_0_0_250), .C2(mult1_out[0]), .ZN(n_0_0_189));
   OAI21_X1 i_0_0_248 (.A(n_0_0_297), .B1(n_0_0_330), .B2(n_0_0_357), .ZN(
      n_0_0_190));
   NOR3_X1 i_0_0_249 (.A1(n_0_0_287), .A2(n_0_0_305), .A3(n_0_0_331), .ZN(
      n_0_0_191));
   NAND2_X1 i_0_0_250 (.A1(n_0_0_193), .A2(n_0_0_277), .ZN(n_0_0_192));
   AOI22_X1 i_0_0_251 (.A1(Interpolation_RAM_RD2_Data[0]), .A2(n_0_0_313), 
      .B1(n_0_0_308), .B2(n_0_0_319), .ZN(n_0_0_193));
   NAND2_X1 i_0_0_252 (.A1(n_0_0_356), .A2(n_0_0_342), .ZN(n_0_0_194));
   NAND3_X1 i_0_0_253 (.A1(Interpolation_RAM_RD1_Data[0]), .A2(n_0_0_326), 
      .A3(n_0_0_221), .ZN(n_0_0_195));
   OAI211_X1 i_0_0_254 (.A(n_0_0_198), .B(n_0_0_196), .C1(n_0_0_289), .C2(
      n_0_0_199), .ZN(n_0_53));
   OAI211_X1 i_0_0_255 (.A(n_0_0_197), .B(n_0_0_326), .C1(n_0_0_224), .C2(
      n_0_0_221), .ZN(n_0_0_196));
   OAI222_X1 i_0_0_256 (.A1(n_0_0_380), .A2(n_0_0_339), .B1(n_0_0_321), .B2(
      n_0_0_307), .C1(n_0_0_312), .C2(n_0_0_379), .ZN(n_0_0_197));
   AOI22_X1 i_0_0_257 (.A1(n_0_0_219), .A2(Interpolation_RAM_RD1_Data[1]), 
      .B1(mult1_out[1]), .B2(n_134), .ZN(n_0_0_198));
   OAI211_X1 i_0_0_258 (.A(n_0_0_200), .B(n_0_0_201), .C1(n_0_0_294), .C2(
      n_0_0_199), .ZN(n_0_54));
   NAND4_X1 i_0_0_259 (.A1(n_0_0_332), .A2(n_0_0_388), .A3(n_177), .A4(
      Start_Interpolation), .ZN(n_0_0_199));
   AOI21_X1 i_0_0_260 (.A(n_0_0_202), .B1(n_134), .B2(mult1_out[2]), .ZN(
      n_0_0_200));
   NAND2_X1 i_0_0_261 (.A1(n_0_0_219), .A2(Interpolation_RAM_RD1_Data[2]), 
      .ZN(n_0_0_201));
   AOI211_X1 i_0_0_262 (.A(n_0_0_203), .B(n_0_0_325), .C1(n_0_0_409), .C2(
      n_0_0_220), .ZN(n_0_0_202));
   AOI22_X1 i_0_0_263 (.A1(Interpolation_RAM_RD2_Data[2]), .A2(n_0_0_313), 
      .B1(n_0_0_308), .B2(n_0_0_322), .ZN(n_0_0_203));
   INV_X1 i_0_0_264 (.A(n_0_0_204), .ZN(n_0_55));
   AOI222_X1 i_0_0_265 (.A1(Interpolation_RAM_RD1_Data[3]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[3]), .C1(mult1_out[3]), 
      .C2(n_134), .ZN(n_0_0_204));
   NAND2_X1 i_0_0_266 (.A1(n_0_0_205), .A2(n_0_0_206), .ZN(n_0_56));
   AOI222_X1 i_0_0_267 (.A1(Interpolation_RAM_RD1_Data[4]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[4]), .C1(mult1_out[4]), 
      .C2(n_134), .ZN(n_0_0_205));
   NAND3_X1 i_0_0_268 (.A1(U_CURRENT_SIZE[4]), .A2(n_0_0_315), .A3(n_0_0_224), 
      .ZN(n_0_0_206));
   NAND2_X1 i_0_0_269 (.A1(n_0_0_207), .A2(n_0_0_208), .ZN(n_0_57));
   AOI222_X1 i_0_0_270 (.A1(Interpolation_RAM_RD1_Data[5]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[5]), .C1(mult1_out[5]), 
      .C2(n_134), .ZN(n_0_0_207));
   NAND3_X1 i_0_0_271 (.A1(U_CURRENT_SIZE[5]), .A2(n_0_0_315), .A3(n_0_0_224), 
      .ZN(n_0_0_208));
   INV_X1 i_0_0_272 (.A(n_0_0_209), .ZN(n_0_58));
   AOI222_X1 i_0_0_273 (.A1(Interpolation_RAM_RD1_Data[6]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[6]), .C1(mult1_out[6]), 
      .C2(n_134), .ZN(n_0_0_209));
   INV_X1 i_0_0_274 (.A(n_0_0_210), .ZN(n_0_59));
   AOI222_X1 i_0_0_275 (.A1(Interpolation_RAM_RD1_Data[7]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[7]), .C1(mult1_out[7]), 
      .C2(n_134), .ZN(n_0_0_210));
   INV_X1 i_0_0_276 (.A(n_0_0_211), .ZN(n_0_60));
   AOI222_X1 i_0_0_277 (.A1(Interpolation_RAM_RD1_Data[8]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[8]), .C1(mult1_out[8]), 
      .C2(n_134), .ZN(n_0_0_211));
   INV_X1 i_0_0_278 (.A(n_0_0_212), .ZN(n_0_61));
   AOI222_X1 i_0_0_279 (.A1(Interpolation_RAM_RD1_Data[9]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[9]), .C1(mult1_out[9]), 
      .C2(n_134), .ZN(n_0_0_212));
   INV_X1 i_0_0_280 (.A(n_0_0_213), .ZN(n_0_62));
   AOI222_X1 i_0_0_281 (.A1(Interpolation_RAM_RD1_Data[10]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[10]), .C1(mult1_out[10]), 
      .C2(n_134), .ZN(n_0_0_213));
   INV_X1 i_0_0_282 (.A(n_0_0_214), .ZN(n_0_63));
   AOI222_X1 i_0_0_283 (.A1(Interpolation_RAM_RD1_Data[11]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[11]), .C1(mult1_out[11]), 
      .C2(n_134), .ZN(n_0_0_214));
   INV_X1 i_0_0_284 (.A(n_0_0_215), .ZN(n_0_64));
   AOI222_X1 i_0_0_285 (.A1(Interpolation_RAM_RD1_Data[12]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[12]), .C1(mult1_out[12]), 
      .C2(n_134), .ZN(n_0_0_215));
   INV_X1 i_0_0_286 (.A(n_0_0_216), .ZN(n_0_65));
   AOI222_X1 i_0_0_287 (.A1(Interpolation_RAM_RD1_Data[13]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[13]), .C1(mult1_out[13]), 
      .C2(n_134), .ZN(n_0_0_216));
   INV_X1 i_0_0_288 (.A(n_0_0_217), .ZN(n_0_66));
   AOI222_X1 i_0_0_289 (.A1(Interpolation_RAM_RD1_Data[14]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[14]), .C1(mult1_out[14]), 
      .C2(n_134), .ZN(n_0_0_217));
   INV_X1 i_0_0_290 (.A(n_0_0_218), .ZN(n_0_67));
   AOI222_X1 i_0_0_291 (.A1(Interpolation_RAM_RD1_Data[15]), .A2(n_0_0_219), 
      .B1(n_0_0_222), .B2(Interpolation_RAM_RD2_Data[15]), .C1(mult1_out[15]), 
      .C2(n_134), .ZN(n_0_0_218));
   OAI22_X1 i_0_0_292 (.A1(n_0_0_325), .A2(n_0_0_220), .B1(n_0_0_224), .B2(RST), 
      .ZN(n_0_0_219));
   NAND3_X1 i_0_0_293 (.A1(n_0_0_340), .A2(n_0_0_392), .A3(
      current_intialization_state[1]), .ZN(n_0_0_220));
   NOR2_X1 i_0_0_294 (.A1(n_0_0_376), .A2(n_0_0_314), .ZN(n_0_0_221));
   NOR3_X1 i_0_0_295 (.A1(n_0_0_325), .A2(n_0_0_312), .A3(n_0_0_409), .ZN(
      n_0_0_222));
   NOR2_X1 i_0_0_296 (.A1(RST), .A2(n_0_0_409), .ZN(n_0_0_223));
   OR2_X1 i_0_0_297 (.A1(n_0_0_225), .A2(n_0_0_357), .ZN(n_0_0_224));
   NAND3_X1 i_0_0_298 (.A1(n_0_0_344), .A2(n_0_0_395), .A3(
      current_interpolation_state[0]), .ZN(n_0_0_225));
   NOR2_X1 i_0_0_299 (.A1(n_0_0_380), .A2(RST), .ZN(n_12));
   AND2_X1 i_0_0_300 (.A1(n_177), .A2(U_CURRENT_SIZE[4]), .ZN(n_13));
   AND2_X1 i_0_0_301 (.A1(n_177), .A2(U_CURRENT_SIZE[5]), .ZN(n_14));
   OAI21_X1 i_0_0_302 (.A(n_177), .B1(n_0_0_339), .B2(n_0_0_407), .ZN(n_15));
   NOR2_X1 i_0_0_303 (.A1(n_0_0_381), .A2(RST), .ZN(n_16));
   NOR2_X1 i_0_0_304 (.A1(n_0_0_382), .A2(RST), .ZN(n_17));
   AND2_X1 i_0_0_305 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[2]), .ZN(n_18));
   AND2_X1 i_0_0_306 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[3]), .ZN(n_19));
   AND2_X1 i_0_0_307 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[4]), .ZN(n_20));
   AND2_X1 i_0_0_308 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[5]), .ZN(n_21));
   AND2_X1 i_0_0_309 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[6]), .ZN(n_22));
   AND2_X1 i_0_0_310 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[7]), .ZN(n_23));
   AND2_X1 i_0_0_311 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[8]), .ZN(n_24));
   AND2_X1 i_0_0_312 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[9]), .ZN(n_25));
   AND2_X1 i_0_0_313 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[10]), .ZN(n_26));
   AND2_X1 i_0_0_314 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[11]), .ZN(n_27));
   AND2_X1 i_0_0_315 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[12]), .ZN(n_28));
   AND2_X1 i_0_0_316 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[13]), .ZN(n_29));
   AND2_X1 i_0_0_317 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[14]), .ZN(n_30));
   AND2_X1 i_0_0_318 (.A1(n_177), .A2(Interpolation_RAM_RD1_Data[15]), .ZN(n_31));
   NAND2_X1 i_0_0_319 (.A1(n_0_0_227), .A2(n_0_0_226), .ZN(n_32));
   NAND2_X1 i_0_0_320 (.A1(adder_sub1_Out[0]), .A2(n_0_0_243), .ZN(n_0_0_226));
   NAND3_X1 i_0_0_321 (.A1(n_177), .A2(n_0_0_247), .A3(Temp[0]), .ZN(n_0_0_227));
   INV_X1 i_0_0_322 (.A(n_0_0_228), .ZN(n_33));
   AOI22_X1 i_0_0_323 (.A1(adder_sub1_Out[1]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_52), .ZN(n_0_0_228));
   INV_X1 i_0_0_324 (.A(n_0_0_229), .ZN(n_34));
   AOI22_X1 i_0_0_325 (.A1(adder_sub1_Out[2]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_53), .ZN(n_0_0_229));
   INV_X1 i_0_0_326 (.A(n_0_0_230), .ZN(n_35));
   AOI22_X1 i_0_0_327 (.A1(adder_sub1_Out[3]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_54), .ZN(n_0_0_230));
   INV_X1 i_0_0_328 (.A(n_0_0_231), .ZN(n_36));
   AOI22_X1 i_0_0_329 (.A1(adder_sub1_Out[4]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_55), .ZN(n_0_0_231));
   INV_X1 i_0_0_330 (.A(n_0_0_232), .ZN(n_37));
   AOI22_X1 i_0_0_331 (.A1(adder_sub1_Out[5]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_56), .ZN(n_0_0_232));
   INV_X1 i_0_0_332 (.A(n_0_0_233), .ZN(n_38));
   AOI22_X1 i_0_0_333 (.A1(adder_sub1_Out[6]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_57), .ZN(n_0_0_233));
   INV_X1 i_0_0_334 (.A(n_0_0_234), .ZN(n_39));
   AOI22_X1 i_0_0_335 (.A1(adder_sub1_Out[7]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_58), .ZN(n_0_0_234));
   INV_X1 i_0_0_336 (.A(n_0_0_235), .ZN(n_40));
   AOI22_X1 i_0_0_337 (.A1(adder_sub1_Out[8]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_59), .ZN(n_0_0_235));
   INV_X1 i_0_0_338 (.A(n_0_0_236), .ZN(n_41));
   AOI22_X1 i_0_0_339 (.A1(adder_sub1_Out[9]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_60), .ZN(n_0_0_236));
   INV_X1 i_0_0_340 (.A(n_0_0_237), .ZN(n_42));
   AOI22_X1 i_0_0_341 (.A1(adder_sub1_Out[10]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_61), .ZN(n_0_0_237));
   INV_X1 i_0_0_342 (.A(n_0_0_238), .ZN(n_43));
   AOI22_X1 i_0_0_343 (.A1(adder_sub1_Out[11]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_62), .ZN(n_0_0_238));
   INV_X1 i_0_0_344 (.A(n_0_0_239), .ZN(n_44));
   AOI22_X1 i_0_0_345 (.A1(adder_sub1_Out[12]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_63), .ZN(n_0_0_239));
   INV_X1 i_0_0_346 (.A(n_0_0_240), .ZN(n_45));
   AOI22_X1 i_0_0_347 (.A1(adder_sub1_Out[13]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_64), .ZN(n_0_0_240));
   INV_X1 i_0_0_348 (.A(n_0_0_241), .ZN(n_46));
   AOI22_X1 i_0_0_349 (.A1(adder_sub1_Out[14]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_65), .ZN(n_0_0_241));
   INV_X1 i_0_0_350 (.A(n_0_0_242), .ZN(n_47));
   AOI22_X1 i_0_0_351 (.A1(adder_sub1_Out[15]), .A2(n_0_0_243), .B1(n_0_0_247), 
      .B2(n_66), .ZN(n_0_0_242));
   NOR2_X1 i_0_0_352 (.A1(n_0_0_247), .A2(RST), .ZN(n_0_0_243));
   AOI21_X1 i_0_0_353 (.A(n_0_0_244), .B1(n_0_0_245), .B2(n_0_0_401), .ZN(n_0_68));
   OAI21_X1 i_0_0_354 (.A(n_177), .B1(n_0_0_245), .B2(Temp[0]), .ZN(n_0_0_244));
   MUX2_X1 i_0_0_355 (.A(n_52), .B(n_71), .S(n_0_0_245), .Z(n_0_69));
   MUX2_X1 i_0_0_356 (.A(n_53), .B(n_73), .S(n_0_0_245), .Z(n_0_70));
   MUX2_X1 i_0_0_357 (.A(n_54), .B(n_75), .S(n_0_0_245), .Z(n_0_71));
   MUX2_X1 i_0_0_358 (.A(n_55), .B(n_77), .S(n_0_0_245), .Z(n_0_72));
   MUX2_X1 i_0_0_359 (.A(n_56), .B(n_79), .S(n_0_0_245), .Z(n_0_73));
   MUX2_X1 i_0_0_360 (.A(n_57), .B(n_81), .S(n_0_0_245), .Z(n_0_74));
   MUX2_X1 i_0_0_361 (.A(n_58), .B(n_83), .S(n_0_0_245), .Z(n_0_75));
   MUX2_X1 i_0_0_362 (.A(n_59), .B(n_85), .S(n_0_0_245), .Z(n_0_76));
   MUX2_X1 i_0_0_363 (.A(n_60), .B(n_87), .S(n_0_0_245), .Z(n_0_77));
   MUX2_X1 i_0_0_364 (.A(n_61), .B(n_89), .S(n_0_0_245), .Z(n_0_78));
   MUX2_X1 i_0_0_365 (.A(n_62), .B(n_91), .S(n_0_0_245), .Z(n_0_79));
   MUX2_X1 i_0_0_366 (.A(n_63), .B(n_93), .S(n_0_0_245), .Z(n_0_80));
   MUX2_X1 i_0_0_367 (.A(n_64), .B(n_95), .S(n_0_0_245), .Z(n_0_81));
   MUX2_X1 i_0_0_368 (.A(n_65), .B(n_97), .S(n_0_0_245), .Z(n_0_82));
   MUX2_X1 i_0_0_369 (.A(n_66), .B(n_99), .S(n_0_0_245), .Z(n_0_83));
   NAND2_X1 i_0_0_370 (.A1(n_0_0_247), .A2(n_0_0_246), .ZN(n_0_0_245));
   NAND2_X1 i_0_0_371 (.A1(n_0_0_298), .A2(n_0_0_356), .ZN(n_0_0_246));
   OR3_X1 i_0_0_372 (.A1(n_0_0_407), .A2(n_0_0_376), .A3(n_0_0_364), .ZN(
      n_0_0_247));
   NOR3_X1 i_0_0_373 (.A1(n_0_0_394), .A2(n_0_0_249), .A3(RST), .ZN(n_48));
   OR2_X1 i_0_0_374 (.A1(n_50), .A2(n_0_0_250), .ZN(n_49));
   OR2_X1 i_0_0_375 (.A1(RST), .A2(n_0_0_248), .ZN(n_50));
   NOR3_X1 i_0_0_376 (.A1(n_0_0_394), .A2(n_0_0_249), .A3(n_0_0_357), .ZN(
      n_0_0_248));
   NAND2_X1 i_0_0_377 (.A1(current_interpolation_state[2]), .A2(n_0_0_345), 
      .ZN(n_0_0_249));
   NOR2_X1 i_0_0_378 (.A1(n_0_0_333), .A2(n_0_0_357), .ZN(n_0_0_250));
   OR2_X1 i_0_0_379 (.A1(RST), .A2(Temp[0]), .ZN(n_51));
   AND2_X1 i_0_0_380 (.A1(n_177), .A2(Temp[1]), .ZN(n_52));
   AND2_X1 i_0_0_381 (.A1(n_177), .A2(Temp[2]), .ZN(n_53));
   AND2_X1 i_0_0_382 (.A1(n_177), .A2(Temp[3]), .ZN(n_54));
   AND2_X1 i_0_0_383 (.A1(n_177), .A2(Temp[4]), .ZN(n_55));
   AND2_X1 i_0_0_384 (.A1(n_177), .A2(Temp[5]), .ZN(n_56));
   AND2_X1 i_0_0_385 (.A1(n_177), .A2(Temp[6]), .ZN(n_57));
   AND2_X1 i_0_0_386 (.A1(n_177), .A2(Temp[7]), .ZN(n_58));
   AND2_X1 i_0_0_387 (.A1(n_177), .A2(Temp[8]), .ZN(n_59));
   AND2_X1 i_0_0_388 (.A1(n_177), .A2(Temp[9]), .ZN(n_60));
   AND2_X1 i_0_0_389 (.A1(n_177), .A2(Temp[10]), .ZN(n_61));
   AND2_X1 i_0_0_390 (.A1(n_177), .A2(Temp[11]), .ZN(n_62));
   AND2_X1 i_0_0_391 (.A1(n_177), .A2(Temp[12]), .ZN(n_63));
   AND2_X1 i_0_0_392 (.A1(n_177), .A2(Temp[13]), .ZN(n_64));
   AND2_X1 i_0_0_393 (.A1(n_177), .A2(Temp[14]), .ZN(n_65));
   AND2_X1 i_0_0_394 (.A1(n_177), .A2(Temp[15]), .ZN(n_66));
   NOR2_X1 i_0_0_395 (.A1(RST), .A2(Div_Count), .ZN(n_67));
   OAI21_X1 i_0_0_396 (.A(n_177), .B1(n_0_0_383), .B2(n_0_0_367), .ZN(n_68));
   AOI22_X1 i_0_0_397 (.A1(n_0_86), .A2(n_0_0_251), .B1(n_177), .B2(n_0_0_407), 
      .ZN(n_0_84));
   INV_X1 i_0_0_398 (.A(n_0_0_252), .ZN(n_0_0_251));
   AOI21_X1 i_0_0_399 (.A(current_intialization_state[2]), .B1(n_0_0_366), 
      .B2(n_0_0_253), .ZN(n_0_0_252));
   AOI211_X1 i_0_0_400 (.A(current_intialization_state[1]), .B(
      current_intialization_state[0]), .C1(Div_Count), .C2(div1_ready), .ZN(
      n_0_0_253));
   INV_X1 i_0_0_401 (.A(n_0_0_254), .ZN(n_0_85));
   AOI21_X1 i_0_0_402 (.A(RST), .B1(n_0_0_356), .B2(n_0_0_255), .ZN(n_0_0_254));
   OAI21_X1 i_0_0_403 (.A(current_interpolation_state[3]), .B1(
      current_interpolation_state[2]), .B2(current_interpolation_state[1]), 
      .ZN(n_0_0_255));
   AOI221_X1 i_0_0_404 (.A(RST), .B1(n_0_0_259), .B2(n_0_0_356), .C1(n_0_0_353), 
      .C2(n_0_0_277), .ZN(n_0_87));
   NAND3_X1 i_0_0_405 (.A1(n_0_0_279), .A2(n_0_0_258), .A3(n_0_0_256), .ZN(
      n_0_89));
   NAND3_X1 i_0_0_406 (.A1(n_0_0_377), .A2(n_0_0_257), .A3(n_0_0_369), .ZN(
      n_0_0_256));
   NAND2_X1 i_0_0_407 (.A1(n_0_0_378), .A2(n_0_0_314), .ZN(n_0_0_257));
   NAND2_X1 i_0_0_408 (.A1(n_0_0_259), .A2(n_0_0_356), .ZN(n_0_0_258));
   INV_X1 i_0_0_409 (.A(n_0_0_260), .ZN(n_0_0_259));
   NAND3_X1 i_0_0_410 (.A1(current_interpolation_state[3]), .A2(n_0_0_349), 
      .A3(n_0_0_396), .ZN(n_0_0_260));
   INV_X1 i_0_0_411 (.A(n_0_0_261), .ZN(n_69));
   AOI22_X1 i_0_0_412 (.A1(div1_Q[0]), .A2(n_0_0_279), .B1(n_0_0_262), .B2(
      adder_sub1_Out[0]), .ZN(n_0_0_261));
   NOR2_X1 i_0_0_413 (.A1(n_0_0_353), .A2(RST), .ZN(n_0_0_262));
   INV_X1 i_0_0_414 (.A(n_0_0_263), .ZN(n_70));
   AOI22_X1 i_0_0_415 (.A1(div1_Q[1]), .A2(n_0_0_279), .B1(n_71), .B2(n_0_0_408), 
      .ZN(n_0_0_263));
   NOR2_X1 i_0_0_416 (.A1(n_0_0_402), .A2(RST), .ZN(n_71));
   INV_X1 i_0_0_417 (.A(n_0_0_264), .ZN(n_72));
   AOI22_X1 i_0_0_418 (.A1(div1_Q[2]), .A2(n_0_0_279), .B1(n_73), .B2(n_0_0_408), 
      .ZN(n_0_0_264));
   NOR2_X1 i_0_0_419 (.A1(n_0_0_403), .A2(RST), .ZN(n_73));
   INV_X1 i_0_0_420 (.A(n_0_0_265), .ZN(n_74));
   AOI22_X1 i_0_0_421 (.A1(div1_Q[3]), .A2(n_0_0_279), .B1(n_75), .B2(n_0_0_408), 
      .ZN(n_0_0_265));
   AND2_X1 i_0_0_422 (.A1(n_177), .A2(adder_sub1_Out[3]), .ZN(n_75));
   INV_X1 i_0_0_423 (.A(n_0_0_266), .ZN(n_76));
   AOI22_X1 i_0_0_424 (.A1(div1_Q[4]), .A2(n_0_0_279), .B1(n_77), .B2(n_0_0_408), 
      .ZN(n_0_0_266));
   AND2_X1 i_0_0_425 (.A1(n_177), .A2(adder_sub1_Out[4]), .ZN(n_77));
   INV_X1 i_0_0_426 (.A(n_0_0_267), .ZN(n_78));
   AOI22_X1 i_0_0_427 (.A1(div1_Q[5]), .A2(n_0_0_279), .B1(n_79), .B2(n_0_0_408), 
      .ZN(n_0_0_267));
   NOR2_X1 i_0_0_428 (.A1(n_0_0_404), .A2(RST), .ZN(n_79));
   INV_X1 i_0_0_429 (.A(n_0_0_268), .ZN(n_80));
   AOI22_X1 i_0_0_430 (.A1(div1_Q[6]), .A2(n_0_0_279), .B1(n_81), .B2(n_0_0_408), 
      .ZN(n_0_0_268));
   NOR2_X1 i_0_0_431 (.A1(n_0_0_405), .A2(RST), .ZN(n_81));
   INV_X1 i_0_0_432 (.A(n_0_0_269), .ZN(n_82));
   AOI22_X1 i_0_0_433 (.A1(div1_Q[7]), .A2(n_0_0_279), .B1(n_83), .B2(n_0_0_408), 
      .ZN(n_0_0_269));
   AND2_X1 i_0_0_434 (.A1(n_177), .A2(adder_sub1_Out[7]), .ZN(n_83));
   INV_X1 i_0_0_435 (.A(n_0_0_270), .ZN(n_84));
   AOI22_X1 i_0_0_436 (.A1(div1_Q[8]), .A2(n_0_0_279), .B1(n_85), .B2(n_0_0_408), 
      .ZN(n_0_0_270));
   AND2_X1 i_0_0_437 (.A1(n_177), .A2(adder_sub1_Out[8]), .ZN(n_85));
   INV_X1 i_0_0_438 (.A(n_0_0_271), .ZN(n_86));
   AOI22_X1 i_0_0_439 (.A1(div1_Q[9]), .A2(n_0_0_279), .B1(n_87), .B2(n_0_0_408), 
      .ZN(n_0_0_271));
   AND2_X1 i_0_0_440 (.A1(n_177), .A2(adder_sub1_Out[9]), .ZN(n_87));
   INV_X1 i_0_0_441 (.A(n_0_0_272), .ZN(n_88));
   AOI22_X1 i_0_0_442 (.A1(div1_Q[10]), .A2(n_0_0_279), .B1(n_89), .B2(n_0_0_408), 
      .ZN(n_0_0_272));
   AND2_X1 i_0_0_443 (.A1(n_177), .A2(adder_sub1_Out[10]), .ZN(n_89));
   INV_X1 i_0_0_444 (.A(n_0_0_273), .ZN(n_90));
   AOI22_X1 i_0_0_445 (.A1(div1_Q[11]), .A2(n_0_0_279), .B1(n_91), .B2(n_0_0_408), 
      .ZN(n_0_0_273));
   AND2_X1 i_0_0_446 (.A1(n_177), .A2(adder_sub1_Out[11]), .ZN(n_91));
   INV_X1 i_0_0_447 (.A(n_0_0_274), .ZN(n_92));
   AOI22_X1 i_0_0_448 (.A1(div1_Q[12]), .A2(n_0_0_279), .B1(n_93), .B2(n_0_0_408), 
      .ZN(n_0_0_274));
   AND2_X1 i_0_0_449 (.A1(n_177), .A2(adder_sub1_Out[12]), .ZN(n_93));
   INV_X1 i_0_0_450 (.A(n_0_0_275), .ZN(n_94));
   AOI22_X1 i_0_0_451 (.A1(div1_Q[14]), .A2(n_0_0_279), .B1(n_95), .B2(n_0_0_408), 
      .ZN(n_0_0_275));
   AND2_X1 i_0_0_452 (.A1(n_177), .A2(adder_sub1_Out[13]), .ZN(n_95));
   INV_X1 i_0_0_453 (.A(n_0_0_276), .ZN(n_96));
   AOI22_X1 i_0_0_454 (.A1(div1_Q[14]), .A2(n_0_0_279), .B1(n_97), .B2(n_0_0_408), 
      .ZN(n_0_0_276));
   AND2_X1 i_0_0_455 (.A1(n_177), .A2(adder_sub1_Out[14]), .ZN(n_97));
   AND2_X1 i_0_0_456 (.A1(n_0_0_408), .A2(n_99), .ZN(n_98));
   AND2_X1 i_0_0_457 (.A1(n_177), .A2(adder_sub1_Out[15]), .ZN(n_99));
   OAI21_X1 i_0_0_458 (.A(n_0_0_279), .B1(n_0_0_277), .B2(n_0_0_407), .ZN(n_100));
   NAND3_X1 i_0_0_459 (.A1(n_0_0_369), .A2(n_0_0_391), .A3(
      current_intialization_state[0]), .ZN(n_0_0_277));
   NOR2_X1 i_0_0_460 (.A1(n_0_0_378), .A2(n_0_0_368), .ZN(n_0_0_278));
   INV_X1 i_0_0_461 (.A(n_0_0_279), .ZN(n_101));
   NOR2_X1 i_0_0_462 (.A1(RST), .A2(n_0_0_408), .ZN(n_0_0_279));
   OAI211_X1 i_0_0_463 (.A(n_0_0_281), .B(n_0_0_280), .C1(RST), .C2(n_0_0_341), 
      .ZN(n_102));
   NAND3_X1 i_0_0_464 (.A1(n_0_0_348), .A2(n_0_0_283), .A3(n_0_4), .ZN(n_0_0_280));
   NAND2_X1 i_0_0_465 (.A1(adder_sub1_Out[0]), .A2(n_0_0_284), .ZN(n_0_0_281));
   AOI21_X1 i_0_0_466 (.A(RST), .B1(n_0_0_282), .B2(n_0_0_341), .ZN(n_103));
   AOI22_X1 i_0_0_467 (.A1(adder_sub1_Out[1]), .A2(n_0_0_285), .B1(n_0_0_283), 
      .B2(n_0_0_348), .ZN(n_0_0_282));
   NOR2_X1 i_0_0_468 (.A1(n_0_0_376), .A2(current_intialization_state[1]), 
      .ZN(n_0_0_283));
   AND2_X1 i_0_0_469 (.A1(adder_sub1_Out[2]), .A2(n_0_0_284), .ZN(n_104));
   AND2_X1 i_0_0_470 (.A1(adder_sub1_Out[3]), .A2(n_0_0_284), .ZN(n_105));
   AND2_X1 i_0_0_471 (.A1(adder_sub1_Out[4]), .A2(n_0_0_284), .ZN(n_106));
   AND2_X1 i_0_0_472 (.A1(adder_sub1_Out[5]), .A2(n_0_0_284), .ZN(n_107));
   AND2_X1 i_0_0_473 (.A1(adder_sub1_Out[6]), .A2(n_0_0_284), .ZN(n_108));
   AND2_X1 i_0_0_474 (.A1(adder_sub1_Out[7]), .A2(n_0_0_284), .ZN(n_109));
   AND2_X1 i_0_0_475 (.A1(adder_sub1_Out[8]), .A2(n_0_0_284), .ZN(n_110));
   AND2_X1 i_0_0_476 (.A1(adder_sub1_Out[9]), .A2(n_0_0_284), .ZN(n_111));
   AND2_X1 i_0_0_477 (.A1(adder_sub1_Out[10]), .A2(n_0_0_284), .ZN(n_112));
   AND2_X1 i_0_0_478 (.A1(adder_sub1_Out[11]), .A2(n_0_0_284), .ZN(n_113));
   AND2_X1 i_0_0_479 (.A1(adder_sub1_Out[12]), .A2(n_0_0_284), .ZN(n_114));
   AND3_X1 i_0_0_480 (.A1(n_177), .A2(n_0_0_341), .A3(n_0_0_285), .ZN(n_0_0_284));
   OAI21_X1 i_0_0_481 (.A(n_0_0_348), .B1(n_0_0_352), .B2(n_0_0_378), .ZN(
      n_0_0_285));
   NAND2_X1 i_0_0_482 (.A1(n_177), .A2(n_0_0_386), .ZN(n_0_88));
   OAI211_X1 i_0_0_483 (.A(n_0_0_323), .B(n_0_0_286), .C1(n_0_0_287), .C2(
      n_0_0_304), .ZN(n_115));
   NAND2_X1 i_0_0_484 (.A1(TZ_ADD[0]), .A2(n_0_0_315), .ZN(n_0_0_286));
   AOI22_X1 i_0_0_485 (.A1(n_0_0_300), .A2(n_0_0_319), .B1(adder_sub1_Out[0]), 
      .B2(n_0_0_303), .ZN(n_0_0_287));
   OAI21_X1 i_0_0_486 (.A(n_0_0_288), .B1(n_0_0_289), .B2(n_0_0_304), .ZN(n_116));
   NAND2_X1 i_0_0_487 (.A1(TZ_ADD[1]), .A2(n_0_0_315), .ZN(n_0_0_288));
   AOI22_X1 i_0_0_488 (.A1(n_0_0_291), .A2(n_0_0_297), .B1(n_0_0_303), .B2(
      adder_sub1_Out[1]), .ZN(n_0_0_289));
   AOI21_X1 i_0_0_489 (.A(n_0_0_291), .B1(n_0_0_303), .B2(adder_sub1_Out[1]), 
      .ZN(n_0_0_290));
   INV_X1 i_0_0_490 (.A(n_0_0_292), .ZN(n_0_0_291));
   NAND3_X1 i_0_0_491 (.A1(n_0_0_389), .A2(n_0_0_300), .A3(Count2[1]), .ZN(
      n_0_0_292));
   OAI221_X1 i_0_0_492 (.A(n_0_0_293), .B1(n_0_0_294), .B2(n_0_0_304), .C1(
      current_intialization_state[1]), .C2(n_0_0_323), .ZN(n_117));
   NAND2_X1 i_0_0_493 (.A1(TZ_ADD[2]), .A2(n_0_0_315), .ZN(n_0_0_293));
   INV_X1 i_0_0_494 (.A(n_0_0_295), .ZN(n_0_0_294));
   OAI21_X1 i_0_0_495 (.A(n_0_0_302), .B1(n_0_0_299), .B2(n_0_0_298), .ZN(
      n_0_0_295));
   AND2_X1 i_0_0_496 (.A1(n_0_0_302), .A2(n_0_0_299), .ZN(n_0_0_296));
   INV_X1 i_0_0_497 (.A(n_0_0_298), .ZN(n_0_0_297));
   NOR2_X1 i_0_0_498 (.A1(n_0_0_355), .A2(n_0_0_346), .ZN(n_0_0_298));
   NAND2_X1 i_0_0_499 (.A1(n_0_0_300), .A2(n_0_0_322), .ZN(n_0_0_299));
   OAI211_X1 i_0_0_500 (.A(Start_Intialization), .B(n_0_0_301), .C1(n_0_0_365), 
      .C2(current_intialization_state[1]), .ZN(n_0_0_300));
   NOR2_X1 i_0_0_501 (.A1(n_0_0_368), .A2(current_intialization_state[0]), 
      .ZN(n_0_0_301));
   NAND2_X1 i_0_0_502 (.A1(adder_sub1_Out[2]), .A2(n_0_0_303), .ZN(n_0_0_302));
   NOR3_X1 i_0_0_503 (.A1(n_0_0_407), .A2(n_0_0_368), .A3(n_0_0_314), .ZN(
      n_0_0_303));
   NAND3_X1 i_0_0_504 (.A1(Start_Interpolation), .A2(n_0_0_361), .A3(n_0_0_329), 
      .ZN(n_0_0_304));
   NAND2_X1 i_0_0_505 (.A1(n_0_0_388), .A2(Start_Interpolation), .ZN(n_0_0_305));
   AND2_X1 i_0_0_506 (.A1(TZ_ADD[3]), .A2(n_0_0_315), .ZN(n_118));
   OAI21_X1 i_0_0_507 (.A(n_0_0_306), .B1(n_0_0_323), .B2(
      current_intialization_state[1]), .ZN(n_119));
   NAND2_X1 i_0_0_508 (.A1(TZ_ADD[4]), .A2(n_0_0_315), .ZN(n_0_0_306));
   NAND2_X1 i_0_0_509 (.A1(n_0_0_324), .A2(n_0_0_391), .ZN(n_0_0_307));
   NOR3_X1 i_0_0_510 (.A1(n_0_0_352), .A2(current_intialization_state[0]), 
      .A3(current_intialization_state[1]), .ZN(n_0_0_308));
   NAND2_X1 i_0_0_511 (.A1(n_0_0_323), .A2(n_0_0_309), .ZN(n_120));
   NAND2_X1 i_0_0_512 (.A1(TZ_ADD[5]), .A2(n_0_0_315), .ZN(n_0_0_309));
   INV_X1 i_0_0_513 (.A(n_0_0_310), .ZN(n_121));
   AOI22_X1 i_0_0_514 (.A1(TZ_ADD[6]), .A2(n_0_0_315), .B1(n_0_0_313), .B2(
      n_0_0_326), .ZN(n_0_0_310));
   AND2_X1 i_0_0_515 (.A1(TZ_ADD[7]), .A2(n_0_0_315), .ZN(n_122));
   INV_X1 i_0_0_516 (.A(n_0_0_311), .ZN(n_123));
   AOI22_X1 i_0_0_517 (.A1(TZ_ADD[8]), .A2(n_0_0_315), .B1(n_0_0_313), .B2(
      n_0_0_326), .ZN(n_0_0_311));
   NAND2_X1 i_0_0_518 (.A1(current_intialization_state[1]), .A2(n_0_0_324), 
      .ZN(n_0_0_312));
   NOR2_X1 i_0_0_519 (.A1(n_0_0_352), .A2(n_0_0_314), .ZN(n_0_0_313));
   NAND2_X1 i_0_0_520 (.A1(n_0_0_390), .A2(current_intialization_state[1]), 
      .ZN(n_0_0_314));
   AND2_X1 i_0_0_521 (.A1(TZ_ADD[9]), .A2(n_0_0_315), .ZN(n_124));
   AND2_X1 i_0_0_522 (.A1(TZ_ADD[10]), .A2(n_0_0_315), .ZN(n_125));
   AND2_X1 i_0_0_523 (.A1(TZ_ADD[11]), .A2(n_0_0_315), .ZN(n_126));
   AND2_X1 i_0_0_524 (.A1(TZ_ADD[12]), .A2(n_0_0_315), .ZN(n_127));
   NOR2_X1 i_0_0_525 (.A1(n_0_0_339), .A2(n_0_0_325), .ZN(n_0_0_315));
   OAI21_X1 i_0_0_526 (.A(n_0_0_326), .B1(n_0_0_316), .B2(n_0_0_407), .ZN(n_128));
   NOR2_X1 i_0_0_527 (.A1(n_0_0_324), .A2(n_0_0_317), .ZN(n_0_0_316));
   NOR3_X1 i_0_0_528 (.A1(current_intialization_state[3]), .A2(
      current_intialization_state[1]), .A3(current_intialization_state[0]), 
      .ZN(n_0_0_317));
   NOR2_X1 i_0_0_529 (.A1(RST), .A2(n_0_0_318), .ZN(n_129));
   AOI221_X1 i_0_0_530 (.A(n_0_0_327), .B1(n_0_0_324), .B2(n_0_0_319), .C1(
      n_0_0_320), .C2(n_0_0_389), .ZN(n_0_0_318));
   AND2_X1 i_0_0_531 (.A1(n_0_0_389), .A2(Count2[0]), .ZN(n_0_0_319));
   NOR3_X1 i_0_0_532 (.A1(n_0_0_376), .A2(n_0_0_337), .A3(n_0_0_370), .ZN(
      n_0_0_320));
   OAI22_X1 i_0_0_533 (.A1(n_0_0_335), .A2(n_0_0_333), .B1(n_0_0_323), .B2(
      n_0_0_321), .ZN(n_130));
   NAND2_X1 i_0_0_534 (.A1(n_0_0_389), .A2(Count2[1]), .ZN(n_0_0_321));
   OAI33_X1 i_0_0_535 (.A1(n_0_0_323), .A2(Interpolation_Intialize), .A3(
      n_0_0_384), .B1(n_0_0_331), .B2(RST), .B3(n_0_0_357), .ZN(n_131));
   NOR2_X1 i_0_0_536 (.A1(n_0_0_384), .A2(Interpolation_Intialize), .ZN(
      n_0_0_322));
   NAND2_X1 i_0_0_537 (.A1(n_0_0_326), .A2(n_0_0_324), .ZN(n_0_0_323));
   NOR2_X1 i_0_0_538 (.A1(n_0_0_352), .A2(current_intialization_state[0]), 
      .ZN(n_0_0_324));
   OAI21_X1 i_0_0_539 (.A(n_177), .B1(n_0_0_337), .B2(n_0_0_328), .ZN(n_0_0_325));
   NOR2_X1 i_0_0_540 (.A1(RST), .A2(n_0_0_327), .ZN(n_0_0_326));
   NOR2_X1 i_0_0_541 (.A1(n_0_0_335), .A2(n_0_0_328), .ZN(n_132));
   NOR2_X1 i_0_0_542 (.A1(n_0_0_337), .A2(n_0_0_328), .ZN(n_0_0_327));
   NAND2_X1 i_0_0_543 (.A1(n_0_0_330), .A2(n_0_0_346), .ZN(n_0_0_328));
   NAND2_X1 i_0_0_544 (.A1(n_0_0_333), .A2(n_0_0_331), .ZN(n_0_0_329));
   AOI21_X1 i_0_0_545 (.A(n_0_0_355), .B1(current_interpolation_state[0]), 
      .B2(current_interpolation_state[2]), .ZN(n_0_0_330));
   NOR2_X1 i_0_0_546 (.A1(n_0_0_335), .A2(n_0_0_331), .ZN(n_133));
   NAND2_X1 i_0_0_547 (.A1(n_0_0_359), .A2(n_0_0_344), .ZN(n_0_0_331));
   NOR2_X1 i_0_0_548 (.A1(n_0_0_358), .A2(n_0_0_343), .ZN(n_0_0_332));
   NOR2_X1 i_0_0_549 (.A1(n_0_0_335), .A2(n_0_0_333), .ZN(n_134));
   NAND4_X1 i_0_0_550 (.A1(n_0_0_397), .A2(n_0_0_394), .A3(
      current_interpolation_state[1]), .A4(current_interpolation_state[2]), 
      .ZN(n_0_0_333));
   NOR3_X1 i_0_0_551 (.A1(n_0_0_396), .A2(n_0_0_355), .A3(
      current_interpolation_state[0]), .ZN(n_0_0_334));
   NAND2_X1 i_0_0_552 (.A1(n_0_0_338), .A2(n_177), .ZN(n_0_0_335));
   NOR2_X1 i_0_0_553 (.A1(n_0_0_337), .A2(RST), .ZN(n_0_0_336));
   OAI21_X1 i_0_0_554 (.A(n_0_0_356), .B1(n_0_0_359), .B2(n_0_0_343), .ZN(
      n_0_0_337));
   AOI21_X1 i_0_0_555 (.A(n_0_0_357), .B1(n_0_0_344), .B2(n_0_0_358), .ZN(
      n_0_0_338));
   OAI211_X1 i_0_0_556 (.A(n_0_0_347), .B(n_0_0_348), .C1(n_0_0_407), .C2(
      n_0_0_339), .ZN(n_135));
   NAND3_X1 i_0_0_557 (.A1(n_0_0_370), .A2(n_0_0_392), .A3(n_0_0_393), .ZN(
      n_0_0_339));
   NOR2_X1 i_0_0_558 (.A1(current_intialization_state[3]), .A2(
      current_intialization_state[0]), .ZN(n_0_0_340));
   AOI21_X1 i_0_0_559 (.A(RST), .B1(n_0_0_385), .B2(n_0_0_341), .ZN(n_136));
   AND2_X1 i_0_0_560 (.A1(n_0_0_341), .A2(n_151), .ZN(n_137));
   AND2_X1 i_0_0_561 (.A1(n_0_0_341), .A2(n_152), .ZN(n_138));
   AND2_X1 i_0_0_562 (.A1(n_0_0_341), .A2(n_153), .ZN(n_139));
   AND2_X1 i_0_0_563 (.A1(n_0_0_341), .A2(n_154), .ZN(n_140));
   AND2_X1 i_0_0_564 (.A1(n_0_0_341), .A2(n_155), .ZN(n_141));
   AND2_X1 i_0_0_565 (.A1(n_0_0_341), .A2(n_156), .ZN(n_142));
   AND2_X1 i_0_0_566 (.A1(n_0_0_341), .A2(n_157), .ZN(n_143));
   AND2_X1 i_0_0_567 (.A1(n_0_0_341), .A2(n_158), .ZN(n_144));
   AND2_X1 i_0_0_568 (.A1(n_0_0_341), .A2(n_159), .ZN(n_145));
   AND2_X1 i_0_0_569 (.A1(n_0_0_341), .A2(n_160), .ZN(n_146));
   AND2_X1 i_0_0_570 (.A1(n_0_0_341), .A2(n_161), .ZN(n_147));
   AND2_X1 i_0_0_571 (.A1(n_0_0_341), .A2(n_162), .ZN(n_148));
   NAND3_X1 i_0_0_572 (.A1(n_0_0_356), .A2(n_0_0_349), .A3(n_0_0_344), .ZN(
      n_0_0_341));
   NAND2_X1 i_0_0_573 (.A1(n_0_0_349), .A2(n_0_0_344), .ZN(n_0_0_342));
   NAND2_X1 i_0_0_574 (.A1(n_0_0_397), .A2(n_0_0_396), .ZN(n_0_0_343));
   NOR2_X1 i_0_0_575 (.A1(current_interpolation_state[3]), .A2(
      current_interpolation_state[2]), .ZN(n_0_0_344));
   NOR2_X1 i_0_0_576 (.A1(current_interpolation_state[3]), .A2(
      current_interpolation_state[1]), .ZN(n_0_0_345));
   NAND2_X1 i_0_0_577 (.A1(n_0_0_396), .A2(n_0_0_394), .ZN(n_0_0_346));
   NAND2_X1 i_0_0_578 (.A1(n_0_0_347), .A2(n_0_0_348), .ZN(n_149));
   NOR2_X1 i_0_0_579 (.A1(RST), .A2(n_0_0_375), .ZN(n_0_0_347));
   NAND3_X1 i_0_0_580 (.A1(n_0_0_349), .A2(n_0_0_356), .A3(n_0_0_397), .ZN(
      n_0_0_348));
   NOR2_X1 i_0_0_581 (.A1(current_interpolation_state[1]), .A2(
      current_interpolation_state[0]), .ZN(n_0_0_349));
   NOR2_X1 i_0_0_582 (.A1(n_0_0_385), .A2(RST), .ZN(n_150));
   AND2_X1 i_0_0_583 (.A1(n_177), .A2(n_179), .ZN(n_151));
   NOR2_X1 i_0_0_584 (.A1(n_0_0_386), .A2(RST), .ZN(n_152));
   AND2_X1 i_0_0_585 (.A1(n_177), .A2(n_189), .ZN(n_153));
   AND2_X1 i_0_0_586 (.A1(n_177), .A2(n_180), .ZN(n_154));
   AND2_X1 i_0_0_587 (.A1(n_177), .A2(n_190), .ZN(n_155));
   AND2_X1 i_0_0_588 (.A1(n_177), .A2(n_181), .ZN(n_156));
   AND2_X1 i_0_0_589 (.A1(n_177), .A2(n_182), .ZN(n_157));
   AND2_X1 i_0_0_590 (.A1(n_177), .A2(n_183), .ZN(n_158));
   AND2_X1 i_0_0_591 (.A1(n_177), .A2(n_184), .ZN(n_159));
   AND2_X1 i_0_0_592 (.A1(n_177), .A2(n_185), .ZN(n_160));
   AND2_X1 i_0_0_593 (.A1(n_177), .A2(n_186), .ZN(n_161));
   AND2_X1 i_0_0_594 (.A1(n_177), .A2(n_187), .ZN(n_162));
   NAND2_X1 i_0_0_595 (.A1(n_0_0_353), .A2(n_0_0_350), .ZN(n_163));
   INV_X1 i_0_0_596 (.A(n_0_0_350), .ZN(n_164));
   AOI21_X1 i_0_0_597 (.A(RST), .B1(n_0_0_351), .B2(n_0_0_377), .ZN(n_0_0_350));
   OAI21_X1 i_0_0_598 (.A(n_177), .B1(n_0_0_364), .B2(n_0_0_352), .ZN(n_165));
   NOR2_X1 i_0_0_599 (.A1(n_0_0_364), .A2(n_0_0_352), .ZN(n_0_0_351));
   NAND2_X1 i_0_0_600 (.A1(n_0_0_393), .A2(current_intialization_state[2]), 
      .ZN(n_0_0_352));
   OR2_X1 i_0_0_601 (.A1(n_0_0_354), .A2(n_0_0_357), .ZN(n_0_0_353));
   NAND3_X1 i_0_0_602 (.A1(n_0_0_359), .A2(n_0_0_397), .A3(
      current_interpolation_state[2]), .ZN(n_0_0_354));
   NAND2_X1 i_0_0_603 (.A1(n_0_0_397), .A2(current_interpolation_state[1]), 
      .ZN(n_0_0_355));
   NAND2_X1 i_0_0_604 (.A1(n_0_0_388), .A2(n_0_0_387), .ZN(n_0_0_356));
   NOR2_X1 i_0_0_605 (.A1(Interpolation_Enable), .A2(Start_Interpolation), 
      .ZN(n_0_0_357));
   NAND2_X1 i_0_0_606 (.A1(current_interpolation_state[1]), .A2(
      current_interpolation_state[0]), .ZN(n_0_0_358));
   NOR2_X1 i_0_0_607 (.A1(n_0_0_395), .A2(n_0_0_394), .ZN(n_0_0_359));
   NOR2_X1 i_0_0_608 (.A1(n_0_0_360), .A2(RST), .ZN(n_0_90));
   OAI21_X1 i_0_0_609 (.A(n_0_0_361), .B1(n_0_0_360), .B2(n_0_0_387), .ZN(n_0_91));
   NAND4_X1 i_0_0_610 (.A1(n_0_0_396), .A2(n_0_0_395), .A3(
      current_interpolation_state[0]), .A4(current_interpolation_state[3]), 
      .ZN(n_0_0_360));
   NOR2_X1 i_0_0_611 (.A1(RST), .A2(Interpolation_Enable), .ZN(n_0_0_361));
   NOR3_X1 i_0_0_612 (.A1(n_0_0_368), .A2(n_0_0_364), .A3(RST), .ZN(n_0_92));
   INV_X1 i_0_0_613 (.A(n_0_0_362), .ZN(n_0_93));
   AOI211_X1 i_0_0_614 (.A(RST), .B(Interpolation_Intialize), .C1(n_0_0_363), 
      .C2(Start_Intialization), .ZN(n_0_0_362));
   NOR2_X1 i_0_0_615 (.A1(n_0_0_368), .A2(n_0_0_364), .ZN(n_0_0_363));
   NAND2_X1 i_0_0_616 (.A1(current_intialization_state[1]), .A2(
      current_intialization_state[0]), .ZN(n_0_0_364));
   NOR2_X1 i_0_0_617 (.A1(RST), .A2(n_0_0_366), .ZN(n_166));
   OAI21_X1 i_0_0_618 (.A(n_177), .B1(n_0_0_367), .B2(n_0_0_366), .ZN(n_167));
   INV_X1 i_0_0_619 (.A(n_0_0_366), .ZN(n_0_0_365));
   NOR2_X1 i_0_0_620 (.A1(div1_divideByZero), .A2(div1_overFlow), .ZN(n_0_0_366));
   NAND3_X1 i_0_0_621 (.A1(n_0_0_377), .A2(n_0_0_370), .A3(n_0_0_369), .ZN(
      n_0_0_367));
   NAND2_X1 i_0_0_622 (.A1(n_0_0_392), .A2(current_intialization_state[3]), 
      .ZN(n_0_0_368));
   NOR2_X1 i_0_0_623 (.A1(n_0_0_393), .A2(current_intialization_state[2]), 
      .ZN(n_0_0_369));
   NOR2_X1 i_0_0_624 (.A1(current_intialization_state[1]), .A2(
      current_intialization_state[0]), .ZN(n_0_0_370));
   NOR2_X1 i_0_0_625 (.A1(n_0_0_390), .A2(RST), .ZN(n_0_4));
   NOR2_X1 i_0_0_626 (.A1(n_0_0_391), .A2(RST), .ZN(n_0_5));
   NOR2_X1 i_0_0_627 (.A1(n_0_0_392), .A2(RST), .ZN(n_0_6));
   NOR2_X1 i_0_0_628 (.A1(n_0_0_393), .A2(RST), .ZN(n_0_86));
   NOR2_X1 i_0_0_629 (.A1(n_0_0_394), .A2(RST), .ZN(n_168));
   NOR2_X1 i_0_0_630 (.A1(n_0_0_395), .A2(RST), .ZN(n_169));
   NOR2_X1 i_0_0_631 (.A1(n_0_0_396), .A2(RST), .ZN(n_170));
   NOR2_X1 i_0_0_632 (.A1(n_0_0_397), .A2(RST), .ZN(n_171));
   OAI21_X1 i_0_0_633 (.A(n_0_0_371), .B1(n_0_0_374), .B2(n_0_0_381), .ZN(n_172));
   NAND2_X1 i_0_0_634 (.A1(n_0_0_374), .A2(USIZE[0]), .ZN(n_0_0_371));
   INV_X1 i_0_0_635 (.A(n_0_0_372), .ZN(n_173));
   MUX2_X1 i_0_0_636 (.A(n_0_0_382), .B(n_0_0_406), .S(n_0_0_374), .Z(n_0_0_372));
   INV_X1 i_0_0_637 (.A(n_174), .ZN(n_0_0_373));
   MUX2_X1 i_0_0_638 (.A(Interpolation_RAM_RD1_Data[2]), .B(USIZE[2]), .S(
      n_0_0_374), .Z(n_174));
   MUX2_X1 i_0_0_639 (.A(Interpolation_RAM_RD1_Data[3]), .B(USIZE[3]), .S(
      n_0_0_374), .Z(n_175));
   MUX2_X1 i_0_0_640 (.A(Interpolation_RAM_RD1_Data[4]), .B(USIZE[4]), .S(
      n_0_0_374), .Z(n_176));
   NAND2_X1 i_0_0_641 (.A1(n_0_0_375), .A2(n_0_0_392), .ZN(n_0_0_374));
   NOR3_X1 i_0_0_642 (.A1(n_0_0_378), .A2(n_0_0_407), .A3(
      current_intialization_state[3]), .ZN(n_0_0_375));
   NAND2_X1 i_0_0_643 (.A1(n_0_0_393), .A2(n_0_0_392), .ZN(n_0_0_376));
   OR2_X1 i_0_0_644 (.A1(Start_Intialization), .A2(Interpolation_Intialize), 
      .ZN(n_0_0_377));
   NAND2_X1 i_0_0_645 (.A1(n_0_0_391), .A2(current_intialization_state[0]), 
      .ZN(n_0_0_378));
   INV_X1 i_0_0_646 (.A(Interpolation_RAM_RD2_Data[1]), .ZN(n_0_0_379));
   INV_X1 i_0_0_647 (.A(U_CURRENT_SIZE[1]), .ZN(n_0_0_380));
   INV_X1 i_0_0_648 (.A(Interpolation_RAM_RD1_Data[0]), .ZN(n_0_0_381));
   INV_X1 i_0_0_649 (.A(Interpolation_RAM_RD1_Data[1]), .ZN(n_0_0_382));
   INV_X1 i_0_0_650 (.A(div1_ready), .ZN(n_0_0_383));
   INV_X1 i_0_0_651 (.A(Count2[2]), .ZN(n_0_0_384));
   INV_X1 i_0_0_652 (.A(n_178), .ZN(n_0_0_385));
   INV_X1 i_0_0_653 (.A(n_188), .ZN(n_0_0_386));
   INV_X1 i_0_0_654 (.A(Start_Interpolation), .ZN(n_0_0_387));
   INV_X1 i_0_0_655 (.A(Interpolation_Enable), .ZN(n_0_0_388));
   INV_X1 i_0_0_656 (.A(Interpolation_Intialize), .ZN(n_0_0_389));
   INV_X1 i_0_0_657 (.A(current_intialization_state[0]), .ZN(n_0_0_390));
   INV_X1 i_0_0_658 (.A(current_intialization_state[1]), .ZN(n_0_0_391));
   INV_X1 i_0_0_659 (.A(current_intialization_state[2]), .ZN(n_0_0_392));
   INV_X1 i_0_0_660 (.A(current_intialization_state[3]), .ZN(n_0_0_393));
   INV_X1 i_0_0_661 (.A(RST), .ZN(n_177));
   INV_X1 i_0_0_662 (.A(current_interpolation_state[0]), .ZN(n_0_0_394));
   INV_X1 i_0_0_663 (.A(current_interpolation_state[1]), .ZN(n_0_0_395));
   INV_X1 i_0_0_664 (.A(current_interpolation_state[2]), .ZN(n_0_0_396));
   INV_X1 i_0_0_665 (.A(current_interpolation_state[3]), .ZN(n_0_0_397));
   INV_X1 i_0_0_666 (.A(n_191), .ZN(n_0_0_398));
   INV_X1 i_0_0_667 (.A(n_192), .ZN(n_0_0_399));
   INV_X1 i_0_0_668 (.A(n_193), .ZN(n_0_0_400));
   INV_X1 i_0_0_669 (.A(adder_sub1_Out[0]), .ZN(n_0_0_401));
   INV_X1 i_0_0_670 (.A(adder_sub1_Out[1]), .ZN(n_0_0_402));
   INV_X1 i_0_0_671 (.A(adder_sub1_Out[2]), .ZN(n_0_0_403));
   INV_X1 i_0_0_672 (.A(adder_sub1_Out[5]), .ZN(n_0_0_404));
   INV_X1 i_0_0_673 (.A(adder_sub1_Out[6]), .ZN(n_0_0_405));
   INV_X1 i_0_0_674 (.A(USIZE[1]), .ZN(n_0_0_406));
   INV_X1 i_0_0_675 (.A(n_0_0_377), .ZN(n_0_0_407));
   INV_X1 i_0_0_676 (.A(n_0_0_353), .ZN(n_0_0_408));
   INV_X1 i_0_0_677 (.A(n_0_0_224), .ZN(n_0_0_409));
   INV_X1 i_0_0_678 (.A(n_0_0_123), .ZN(n_0_0_410));
   MUX2_X1 Intialization_Done_reg_enable_mux_0 (.A(Intialization_Done), .B(
      n_0_92), .S(n_0_93), .Z(n_0_94));
   MUX2_X1 Interpolation_Done_reg_enable_mux_0 (.A(Interpolation_Done), .B(
      n_0_90), .S(n_0_91), .Z(n_0_95));
   MUX2_X1 Interpolation_Memory_WR_Enable_reg_enable_mux_0 (.A(
      Interpolation_Memory_WR_Enable), .B(n_0_87), .S(n_0_89), .Z(n_0_96));
   DFF_X1 \adder_sub3_In2_reg[0]  (.D(n_177), .CK(n_1_4), .Q(adder_sub3_In2[0]), 
      .QN());
   DFF_X1 \adder_sub3_In1_reg[2]  (.D(n_11), .CK(n_1_4), .Q(adder_sub3_In1[2]), 
      .QN());
   DFF_X1 \adder_sub3_In1_reg[1]  (.D(n_9), .CK(n_1_4), .Q(adder_sub3_In1[1]), 
      .QN());
   DFF_X1 \adder_sub3_In1_reg[0]  (.D(n_7), .CK(n_1_4), .Q(adder_sub3_In1[0]), 
      .QN());
   DFF_X1 \div1_divisor_reg[15]  (.D(n_66), .CK(n_1_5), .Q(div1_divisor[15]), 
      .QN());
   DFF_X1 \div1_divisor_reg[14]  (.D(n_65), .CK(n_1_5), .Q(div1_divisor[14]), 
      .QN());
   DFF_X1 \div1_divisor_reg[13]  (.D(n_64), .CK(n_1_5), .Q(div1_divisor[13]), 
      .QN());
   DFF_X1 \div1_divisor_reg[12]  (.D(n_63), .CK(n_1_5), .Q(div1_divisor[12]), 
      .QN());
   DFF_X1 \div1_divisor_reg[11]  (.D(n_62), .CK(n_1_5), .Q(div1_divisor[11]), 
      .QN());
   DFF_X1 \div1_divisor_reg[10]  (.D(n_61), .CK(n_1_5), .Q(div1_divisor[10]), 
      .QN());
   DFF_X1 \div1_divisor_reg[9]  (.D(n_60), .CK(n_1_5), .Q(div1_divisor[9]), 
      .QN());
   DFF_X1 \div1_divisor_reg[8]  (.D(n_59), .CK(n_1_5), .Q(div1_divisor[8]), 
      .QN());
   DFF_X1 \div1_divisor_reg[7]  (.D(n_58), .CK(n_1_5), .Q(div1_divisor[7]), 
      .QN());
   DFF_X1 \div1_divisor_reg[6]  (.D(n_57), .CK(n_1_5), .Q(div1_divisor[6]), 
      .QN());
   DFF_X1 \div1_divisor_reg[5]  (.D(n_56), .CK(n_1_5), .Q(div1_divisor[5]), 
      .QN());
   DFF_X1 \div1_divisor_reg[4]  (.D(n_55), .CK(n_1_5), .Q(div1_divisor[4]), 
      .QN());
   DFF_X1 \div1_divisor_reg[3]  (.D(n_54), .CK(n_1_5), .Q(div1_divisor[3]), 
      .QN());
   DFF_X1 \div1_divisor_reg[2]  (.D(n_53), .CK(n_1_5), .Q(div1_divisor[2]), 
      .QN());
   DFF_X1 \div1_divisor_reg[1]  (.D(n_52), .CK(n_1_5), .Q(div1_divisor[1]), 
      .QN());
   DFF_X1 \div1_divisor_reg[0]  (.D(n_51), .CK(n_1_5), .Q(div1_divisor[0]), 
      .QN());
   DFF_X1 \div1_dividend_reg[15]  (.D(n_99), .CK(n_1_5), .Q(div1_dividend[15]), 
      .QN());
   DFF_X1 \div1_dividend_reg[14]  (.D(n_97), .CK(n_1_5), .Q(div1_dividend[14]), 
      .QN());
   DFF_X1 \div1_dividend_reg[13]  (.D(n_95), .CK(n_1_5), .Q(div1_dividend[13]), 
      .QN());
   DFF_X1 \div1_dividend_reg[12]  (.D(n_93), .CK(n_1_5), .Q(div1_dividend[12]), 
      .QN());
   DFF_X1 \div1_dividend_reg[11]  (.D(n_91), .CK(n_1_5), .Q(div1_dividend[11]), 
      .QN());
   DFF_X1 \div1_dividend_reg[10]  (.D(n_89), .CK(n_1_5), .Q(div1_dividend[10]), 
      .QN());
   DFF_X1 \div1_dividend_reg[9]  (.D(n_87), .CK(n_1_5), .Q(div1_dividend[9]), 
      .QN());
   DFF_X1 \div1_dividend_reg[8]  (.D(n_85), .CK(n_1_5), .Q(div1_dividend[8]), 
      .QN());
   DFF_X1 \div1_dividend_reg[7]  (.D(n_83), .CK(n_1_5), .Q(div1_dividend[7]), 
      .QN());
   DFF_X1 \div1_dividend_reg[6]  (.D(n_81), .CK(n_1_5), .Q(div1_dividend[6]), 
      .QN());
   DFF_X1 \div1_dividend_reg[5]  (.D(n_79), .CK(n_1_5), .Q(div1_dividend[5]), 
      .QN());
   DFF_X1 \div1_dividend_reg[4]  (.D(n_77), .CK(n_1_5), .Q(div1_dividend[4]), 
      .QN());
   DFF_X1 \div1_dividend_reg[3]  (.D(n_75), .CK(n_1_5), .Q(div1_dividend[3]), 
      .QN());
   DFF_X1 \div1_dividend_reg[2]  (.D(n_73), .CK(n_1_5), .Q(div1_dividend[2]), 
      .QN());
   DFF_X1 \div1_dividend_reg[1]  (.D(n_71), .CK(n_1_5), .Q(div1_dividend[1]), 
      .QN());
   DFF_X1 \div1_dividend_reg[0]  (.D(n_5), .CK(n_1_5), .Q(div1_dividend[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_Interpolation_RAM_WR_Data_reg (.CK(CLK), .E(n_100), 
      .SE(1'b0), .GCK(n_1_0));
   DFF_X1 \Interpolation_RAM_WR_Data_reg[15]  (.D(n_98), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[15]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[14]  (.D(n_96), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[14]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[13]  (.D(n_94), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[13]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[12]  (.D(n_92), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[12]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[11]  (.D(n_90), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[11]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[10]  (.D(n_88), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[10]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[9]  (.D(n_86), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[9]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[8]  (.D(n_84), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[8]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[7]  (.D(n_82), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[7]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[6]  (.D(n_80), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[6]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[5]  (.D(n_78), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[5]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[4]  (.D(n_76), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[4]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[3]  (.D(n_74), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[3]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[2]  (.D(n_72), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[2]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[1]  (.D(n_70), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[1]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Data_reg[0]  (.D(n_69), .CK(n_1_0), .Q(
      Interpolation_RAM_WR_Data[0]), .QN());
   DFF_X1 mult1_enable_reg (.D(n_1_8), .CK(CLK), .Q(mult1_enable), .QN());
   DFF_X1 \mult1_second_operand_reg[15]  (.D(n_47), .CK(n_1_6), .Q(
      mult1_second_operand[15]), .QN());
   DFF_X1 \mult1_second_operand_reg[14]  (.D(n_46), .CK(n_1_6), .Q(
      mult1_second_operand[14]), .QN());
   DFF_X1 \mult1_second_operand_reg[13]  (.D(n_45), .CK(n_1_6), .Q(
      mult1_second_operand[13]), .QN());
   DFF_X1 \mult1_second_operand_reg[12]  (.D(n_44), .CK(n_1_6), .Q(
      mult1_second_operand[12]), .QN());
   DFF_X1 \mult1_second_operand_reg[11]  (.D(n_43), .CK(n_1_6), .Q(
      mult1_second_operand[11]), .QN());
   DFF_X1 \mult1_second_operand_reg[10]  (.D(n_42), .CK(n_1_6), .Q(
      mult1_second_operand[10]), .QN());
   DFF_X1 \mult1_second_operand_reg[9]  (.D(n_41), .CK(n_1_6), .Q(
      mult1_second_operand[9]), .QN());
   DFF_X1 \mult1_second_operand_reg[8]  (.D(n_40), .CK(n_1_6), .Q(
      mult1_second_operand[8]), .QN());
   DFF_X1 \mult1_second_operand_reg[7]  (.D(n_39), .CK(n_1_6), .Q(
      mult1_second_operand[7]), .QN());
   DFF_X1 \mult1_second_operand_reg[6]  (.D(n_38), .CK(n_1_6), .Q(
      mult1_second_operand[6]), .QN());
   DFF_X1 \mult1_second_operand_reg[5]  (.D(n_37), .CK(n_1_6), .Q(
      mult1_second_operand[5]), .QN());
   DFF_X1 \mult1_second_operand_reg[4]  (.D(n_36), .CK(n_1_6), .Q(
      mult1_second_operand[4]), .QN());
   DFF_X1 \mult1_second_operand_reg[3]  (.D(n_35), .CK(n_1_6), .Q(
      mult1_second_operand[3]), .QN());
   DFF_X1 \mult1_second_operand_reg[2]  (.D(n_34), .CK(n_1_6), .Q(
      mult1_second_operand[2]), .QN());
   DFF_X1 \mult1_second_operand_reg[1]  (.D(n_33), .CK(n_1_6), .Q(
      mult1_second_operand[1]), .QN());
   DFF_X1 \mult1_second_operand_reg[0]  (.D(n_32), .CK(n_1_6), .Q(
      mult1_second_operand[0]), .QN());
   DFF_X1 \mult1_first_operand_reg[15]  (.D(n_31), .CK(n_1_6), .Q(
      mult1_first_operand[15]), .QN());
   DFF_X1 \mult1_first_operand_reg[14]  (.D(n_30), .CK(n_1_6), .Q(
      mult1_first_operand[14]), .QN());
   DFF_X1 \mult1_first_operand_reg[13]  (.D(n_29), .CK(n_1_6), .Q(
      mult1_first_operand[13]), .QN());
   DFF_X1 \mult1_first_operand_reg[12]  (.D(n_28), .CK(n_1_6), .Q(
      mult1_first_operand[12]), .QN());
   DFF_X1 \mult1_first_operand_reg[11]  (.D(n_27), .CK(n_1_6), .Q(
      mult1_first_operand[11]), .QN());
   DFF_X1 \mult1_first_operand_reg[10]  (.D(n_26), .CK(n_1_6), .Q(
      mult1_first_operand[10]), .QN());
   DFF_X1 \mult1_first_operand_reg[9]  (.D(n_25), .CK(n_1_6), .Q(
      mult1_first_operand[9]), .QN());
   DFF_X1 \mult1_first_operand_reg[8]  (.D(n_24), .CK(n_1_6), .Q(
      mult1_first_operand[8]), .QN());
   DFF_X1 \mult1_first_operand_reg[7]  (.D(n_23), .CK(n_1_6), .Q(
      mult1_first_operand[7]), .QN());
   DFF_X1 \mult1_first_operand_reg[6]  (.D(n_22), .CK(n_1_6), .Q(
      mult1_first_operand[6]), .QN());
   DFF_X1 \mult1_first_operand_reg[5]  (.D(n_21), .CK(n_1_6), .Q(
      mult1_first_operand[5]), .QN());
   DFF_X1 \mult1_first_operand_reg[4]  (.D(n_20), .CK(n_1_6), .Q(
      mult1_first_operand[4]), .QN());
   DFF_X1 \mult1_first_operand_reg[3]  (.D(n_19), .CK(n_1_6), .Q(
      mult1_first_operand[3]), .QN());
   DFF_X1 \mult1_first_operand_reg[2]  (.D(n_18), .CK(n_1_6), .Q(
      mult1_first_operand[2]), .QN());
   DFF_X1 \mult1_first_operand_reg[1]  (.D(n_17), .CK(n_1_6), .Q(
      mult1_first_operand[1]), .QN());
   DFF_X1 \mult1_first_operand_reg[0]  (.D(n_16), .CK(n_1_6), .Q(
      mult1_first_operand[0]), .QN());
   DFF_X1 div1_reset_reg (.D(n_1_9), .CK(CLK), .Q(div1_reset), .QN());
   DFF_X1 \adder_sub2_In1_reg[12]  (.D(n_127), .CK(n_1_7), .Q(adder_sub2_In1[12]), 
      .QN());
   DFF_X1 \adder_sub2_In1_reg[11]  (.D(n_126), .CK(n_1_7), .Q(adder_sub2_In1[11]), 
      .QN());
   DFF_X1 \adder_sub2_In1_reg[10]  (.D(n_125), .CK(n_1_7), .Q(adder_sub2_In1[10]), 
      .QN());
   DFF_X1 \adder_sub2_In1_reg[9]  (.D(n_124), .CK(n_1_7), .Q(adder_sub2_In1[9]), 
      .QN());
   DFF_X1 \adder_sub2_In1_reg[8]  (.D(n_123), .CK(n_1_7), .Q(adder_sub2_In1[8]), 
      .QN());
   DFF_X1 \adder_sub2_In1_reg[7]  (.D(n_122), .CK(n_1_7), .Q(adder_sub2_In1[7]), 
      .QN());
   DFF_X1 \adder_sub2_In1_reg[6]  (.D(n_121), .CK(n_1_7), .Q(adder_sub2_In1[6]), 
      .QN());
   DFF_X1 \adder_sub2_In1_reg[5]  (.D(n_120), .CK(n_1_7), .Q(adder_sub2_In1[5]), 
      .QN());
   DFF_X1 \adder_sub2_In1_reg[4]  (.D(n_119), .CK(n_1_7), .Q(adder_sub2_In1[4]), 
      .QN());
   DFF_X1 \adder_sub2_In1_reg[3]  (.D(n_118), .CK(n_1_7), .Q(adder_sub2_In1[3]), 
      .QN());
   DFF_X1 \adder_sub2_In1_reg[2]  (.D(n_117), .CK(n_1_7), .Q(adder_sub2_In1[2]), 
      .QN());
   DFF_X1 \adder_sub2_In1_reg[1]  (.D(n_116), .CK(n_1_7), .Q(adder_sub2_In1[1]), 
      .QN());
   DFF_X1 \adder_sub2_In1_reg[0]  (.D(n_115), .CK(n_1_7), .Q(adder_sub2_In1[0]), 
      .QN());
   DFF_X1 \adder_sub2_In2_reg[8]  (.D(n_134), .CK(n_1_7), .Q(adder_sub2_In2[8]), 
      .QN());
   DFF_X1 \adder_sub2_In2_reg[5]  (.D(n_133), .CK(n_1_7), .Q(adder_sub2_In2[5]), 
      .QN());
   DFF_X1 \adder_sub2_In2_reg[4]  (.D(n_132), .CK(n_1_7), .Q(adder_sub2_In2[4]), 
      .QN());
   DFF_X1 \adder_sub2_In2_reg[2]  (.D(n_131), .CK(n_1_7), .Q(adder_sub2_In2[2]), 
      .QN());
   DFF_X1 \adder_sub2_In2_reg[1]  (.D(n_130), .CK(n_1_7), .Q(adder_sub2_In2[1]), 
      .QN());
   DFF_X1 \adder_sub2_In2_reg[0]  (.D(n_129), .CK(n_1_7), .Q(adder_sub2_In2[0]), 
      .QN());
   DFF_X1 Start_Intialization_reg (.D(n_1), .CK(CLK), .Q(Start_Intialization), 
      .QN());
   DFF_X1 Start_Interpolation_reg (.D(n_0), .CK(CLK), .Q(Start_Interpolation), 
      .QN());
   CLKGATETST_X1 clk_gate_Interpolation_RAM_RD1_Address_reg (.CK(CLK), .E(n_135), 
      .SE(1'b0), .GCK(n_1_1));
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[12]  (.D(n_114), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[12]), .QN());
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[11]  (.D(n_113), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[11]), .QN());
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[10]  (.D(n_112), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[10]), .QN());
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[9]  (.D(n_111), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[9]), .QN());
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[8]  (.D(n_110), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[8]), .QN());
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[7]  (.D(n_109), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[7]), .QN());
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[6]  (.D(n_108), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[6]), .QN());
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[5]  (.D(n_107), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[5]), .QN());
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[4]  (.D(n_106), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[4]), .QN());
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[3]  (.D(n_105), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[3]), .QN());
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[2]  (.D(n_104), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[2]), .QN());
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[1]  (.D(n_103), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[1]), .QN());
   DFF_X1 \Interpolation_RAM_RD1_Address_reg[0]  (.D(n_102), .CK(n_1_1), 
      .Q(Interpolation_RAM_RD1_Address[0]), .QN());
   DFF_X1 \Count2_reg[2]  (.D(n_10), .CK(CLK), .Q(Count2[2]), .QN());
   DFF_X1 \Count2_reg[1]  (.D(n_8), .CK(CLK), .Q(Count2[1]), .QN());
   DFF_X1 \Count2_reg[0]  (.D(n_6), .CK(CLK), .Q(Count2[0]), .QN());
   CLKGATETST_X1 clk_gate_Interpolation_RAM_RD2_Address_reg (.CK(CLK), .E(n_149), 
      .SE(1'b0), .GCK(n_1_2));
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[12]  (.D(n_148), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[12]), .QN());
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[11]  (.D(n_147), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[11]), .QN());
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[10]  (.D(n_146), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[10]), .QN());
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[9]  (.D(n_145), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[9]), .QN());
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[8]  (.D(n_144), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[8]), .QN());
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[7]  (.D(n_143), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[7]), .QN());
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[6]  (.D(n_142), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[6]), .QN());
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[5]  (.D(n_141), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[5]), .QN());
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[4]  (.D(n_140), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[4]), .QN());
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[3]  (.D(n_139), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[3]), .QN());
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[2]  (.D(n_138), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[2]), .QN());
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[1]  (.D(n_137), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[1]), .QN());
   DFF_X1 \Interpolation_RAM_RD2_Address_reg[0]  (.D(n_136), .CK(n_1_2), 
      .Q(Interpolation_RAM_RD2_Address[0]), .QN());
   CLKGATETST_X1 clk_gate_Interpolation_RAM_WR_Address_reg (.CK(CLK), .E(n_163), 
      .SE(1'b0), .GCK(n_1_3));
   DFF_X1 \Interpolation_RAM_WR_Address_reg[12]  (.D(n_162), .CK(n_1_3), 
      .Q(Interpolation_RAM_WR_Address[12]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Address_reg[11]  (.D(n_161), .CK(n_1_3), 
      .Q(Interpolation_RAM_WR_Address[11]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Address_reg[10]  (.D(n_160), .CK(n_1_3), 
      .Q(Interpolation_RAM_WR_Address[10]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Address_reg[9]  (.D(n_159), .CK(n_1_3), .Q(
      Interpolation_RAM_WR_Address[9]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Address_reg[8]  (.D(n_158), .CK(n_1_3), .Q(
      Interpolation_RAM_WR_Address[8]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Address_reg[7]  (.D(n_157), .CK(n_1_3), .Q(
      Interpolation_RAM_WR_Address[7]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Address_reg[6]  (.D(n_156), .CK(n_1_3), .Q(
      Interpolation_RAM_WR_Address[6]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Address_reg[5]  (.D(n_155), .CK(n_1_3), .Q(
      Interpolation_RAM_WR_Address[5]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Address_reg[4]  (.D(n_154), .CK(n_1_3), .Q(
      Interpolation_RAM_WR_Address[4]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Address_reg[3]  (.D(n_153), .CK(n_1_3), .Q(
      Interpolation_RAM_WR_Address[3]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Address_reg[2]  (.D(n_152), .CK(n_1_3), .Q(
      Interpolation_RAM_WR_Address[2]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Address_reg[1]  (.D(n_151), .CK(n_1_3), .Q(
      Interpolation_RAM_WR_Address[1]), .QN());
   DFF_X1 \Interpolation_RAM_WR_Address_reg[0]  (.D(n_150), .CK(n_1_3), .Q(
      Interpolation_RAM_WR_Address[0]), .QN());
   DFF_X1 Div_Count_reg (.D(n_1_10), .CK(CLK), .Q(Div_Count), .QN());
   CLKGATETST_X1 clk_gate_USIZE_reg (.CK(CLK), .E(n_177), .SE(1'b0), .GCK(n_1_14));
   DFF_X1 \USIZE_reg[4]  (.D(n_176), .CK(n_1_14), .Q(USIZE[4]), .QN());
   DFF_X1 \USIZE_reg[3]  (.D(n_175), .CK(n_1_14), .Q(USIZE[3]), .QN());
   DFF_X1 \USIZE_reg[2]  (.D(n_174), .CK(n_1_14), .Q(USIZE[2]), .QN());
   DFF_X1 \USIZE_reg[1]  (.D(n_173), .CK(n_1_14), .Q(USIZE[1]), .QN());
   DFF_X1 \USIZE_reg[0]  (.D(n_172), .CK(n_1_14), .Q(USIZE[0]), .QN());
   DFF_X1 Error_reg (.D(n_1_11), .CK(CLK), .Q(Error), .QN());
   DFF_X1 \U_CURRENT_SIZE_reg[5]  (.D(n_1_15), .CK(CLK), .Q(U_CURRENT_SIZE[5]), 
      .QN());
   DFF_X1 \U_CURRENT_SIZE_reg[4]  (.D(n_1_13), .CK(CLK), .Q(U_CURRENT_SIZE[4]), 
      .QN());
   DFF_X1 \U_CURRENT_SIZE_reg[1]  (.D(n_1_12), .CK(CLK), .Q(U_CURRENT_SIZE[1]), 
      .QN());
   DFF_X1 \interpolation_state_reg[3]  (.D(n_171), .CK(CLK), .Q(
      interpolation_state[3]), .QN());
   DFF_X1 \interpolation_state_reg[2]  (.D(n_170), .CK(CLK), .Q(
      interpolation_state[2]), .QN());
   DFF_X1 \interpolation_state_reg[1]  (.D(n_169), .CK(CLK), .Q(
      interpolation_state[1]), .QN());
   DFF_X1 \interpolation_state_reg[0]  (.D(n_168), .CK(CLK), .Q(
      interpolation_state[0]), .QN());
   CLKGATETST_X1 clk_gate_adder_sub3_Cin_reg (.CK(CLK), .E(n_101), .SE(1'b0), 
      .GCK(n_1_4));
   CLKGATETST_X1 clk_gate_div1_divisor_reg (.CK(CLK), .E(n_164), .SE(1'b0), 
      .GCK(n_1_5));
   CLKGATETST_X1 clk_gate_mult1_second_operand_reg (.CK(CLK), .E(n_50), .SE(1'b0), 
      .GCK(n_1_6));
   CLKGATETST_X1 clk_gate_adder_sub2_Sub_reg (.CK(CLK), .E(n_128), .SE(1'b0), 
      .GCK(n_1_7));
   DFF_X1 adder_sub1_Sub_reg (.D(n_1_16), .CK(CLK), .Q(adder_sub1_Sub), .QN());
   MUX2_X1 mult1_enable_reg_enable_mux_0 (.A(mult1_enable), .B(n_48), .S(n_49), 
      .Z(n_1_8));
   MUX2_X1 div1_reset_reg_enable_mux_0 (.A(div1_reset), .B(n_165), .S(n_2), 
      .Z(n_1_9));
   MUX2_X1 Div_Count_reg_enable_mux_0 (.A(Div_Count), .B(n_67), .S(n_68), 
      .Z(n_1_10));
   MUX2_X1 Error_reg_enable_mux_0 (.A(Error), .B(n_166), .S(n_167), .Z(n_1_11));
   MUX2_X1 i_1_0_0 (.A(U_CURRENT_SIZE[5]), .B(n_14), .S(n_15), .Z(n_1_15));
   MUX2_X1 i_1_0_1 (.A(U_CURRENT_SIZE[4]), .B(n_13), .S(n_15), .Z(n_1_13));
   MUX2_X1 i_1_0_2 (.A(U_CURRENT_SIZE[1]), .B(n_12), .S(n_15), .Z(n_1_12));
   MUX2_X1 adder_sub1_Sub_reg_enable_mux_0 (.A(adder_sub1_Sub), .B(n_3), 
      .S(n_4), .Z(n_1_16));
   multiplier_16bit mult1 (.first_operand(mult1_first_operand), .second_operand(
      mult1_second_operand), .out(mult1_out), .enable(mult1_enable), .overflow());
   Division_CLHA div1 (.reset(div1_reset), .clk(CLK), .dividend(div1_dividend), 
      .divisor(div1_divisor), .Q({uc_0, div1_Q[14], uc_1, div1_Q[12], div1_Q[11], 
      div1_Q[10], div1_Q[9], div1_Q[8], div1_Q[7], div1_Q[6], div1_Q[5], 
      div1_Q[4], div1_Q[3], div1_Q[2], div1_Q[1], div1_Q[0]}), .ready(div1_ready), 
      .overFlow(div1_overFlow), .divideByZero(div1_divideByZero));
   OAI21_X1 adder_sub1_i_0_0 (.A(adder_sub1_i_0_n_59), .B1(adder_sub1_i_0_n_57), 
      .B2(adder_sub1_i_0_n_58), .ZN(adder_sub1_Out[0]));
   XNOR2_X1 adder_sub1_i_0_1 (.A(adder_sub1_i_0_n_60), .B(adder_sub1_i_0_n_73), 
      .ZN(adder_sub1_Out[1]));
   XNOR2_X1 adder_sub1_i_0_2 (.A(adder_sub1_i_0_n_78), .B(adder_sub1_i_0_n_113), 
      .ZN(adder_sub1_Out[2]));
   XNOR2_X1 adder_sub1_i_0_3 (.A(adder_sub1_i_0_n_123), .B(adder_sub1_i_0_n_158), 
      .ZN(adder_sub1_Out[3]));
   XNOR2_X1 adder_sub1_i_0_4 (.A(adder_sub1_i_0_n_159), .B(adder_sub1_i_0_n_182), 
      .ZN(adder_sub1_Out[4]));
   XNOR2_X1 adder_sub1_i_0_5 (.A(adder_sub1_i_0_n_13), .B(adder_sub1_i_0_n_12), 
      .ZN(adder_sub1_Out[6]));
   XNOR2_X1 adder_sub1_i_0_6 (.A(adder_sub1_i_0_n_11), .B(adder_sub1_i_0_n_10), 
      .ZN(adder_sub1_Out[7]));
   XNOR2_X1 adder_sub1_i_0_7 (.A(adder_sub1_i_0_n_9), .B(adder_sub1_i_0_n_0), 
      .ZN(adder_sub1_Out[8]));
   AOI21_X1 adder_sub1_i_0_8 (.A(adder_sub1_i_0_n_93), .B1(adder_sub1_i_0_n_100), 
      .B2(adder_sub1_i_0_n_94), .ZN(adder_sub1_i_0_n_0));
   XOR2_X1 adder_sub1_i_0_9 (.A(adder_sub1_i_0_n_105), .B(adder_sub1_i_0_n_8), 
      .Z(adder_sub1_Out[9]));
   XOR2_X1 adder_sub1_i_0_10 (.A(adder_sub1_i_0_n_7), .B(adder_sub1_i_0_n_6), 
      .Z(adder_sub1_Out[10]));
   XNOR2_X1 adder_sub1_i_0_11 (.A(adder_sub1_i_0_n_4), .B(adder_sub1_i_0_n_3), 
      .ZN(adder_sub1_Out[11]));
   XOR2_X1 adder_sub1_i_0_12 (.A(adder_sub1_i_0_n_161), .B(adder_sub1_i_0_n_1), 
      .Z(adder_sub1_Out[12]));
   XNOR2_X1 adder_sub1_i_0_13 (.A(adder_sub1_i_0_n_144), .B(adder_sub1_i_0_n_2), 
      .ZN(adder_sub1_i_0_n_1));
   AOI21_X1 adder_sub1_i_0_14 (.A(adder_sub1_i_0_n_131), .B1(adder_sub1_i_0_n_4), 
      .B2(adder_sub1_i_0_n_3), .ZN(adder_sub1_i_0_n_2));
   AOI21_X1 adder_sub1_i_0_15 (.A(adder_sub1_i_0_n_131), .B1(
      adder_sub1_i_0_n_139), .B2(adder_sub1_i_0_n_132), .ZN(adder_sub1_i_0_n_3));
   INV_X1 adder_sub1_i_0_16 (.A(adder_sub1_i_0_n_5), .ZN(adder_sub1_i_0_n_4));
   OAI22_X1 adder_sub1_i_0_17 (.A1(adder_sub1_i_0_n_124), .A2(
      adder_sub1_i_0_n_119), .B1(adder_sub1_i_0_n_7), .B2(adder_sub1_i_0_n_6), 
      .ZN(adder_sub1_i_0_n_5));
   XNOR2_X1 adder_sub1_i_0_18 (.A(adder_sub1_i_0_n_124), .B(adder_sub1_i_0_n_119), 
      .ZN(adder_sub1_i_0_n_6));
   AOI21_X1 adder_sub1_i_0_19 (.A(adder_sub1_i_0_n_106), .B1(
      adder_sub1_i_0_n_105), .B2(adder_sub1_i_0_n_8), .ZN(adder_sub1_i_0_n_7));
   AOI22_X1 adder_sub1_i_0_20 (.A1(adder_sub1_i_0_n_100), .A2(
      adder_sub1_i_0_n_94), .B1(adder_sub1_i_0_n_92), .B2(adder_sub1_i_0_n_9), 
      .ZN(adder_sub1_i_0_n_8));
   OAI22_X1 adder_sub1_i_0_21 (.A1(adder_sub1_i_0_n_86), .A2(adder_sub1_i_0_n_80), 
      .B1(adder_sub1_i_0_n_11), .B2(adder_sub1_i_0_n_10), .ZN(adder_sub1_i_0_n_9));
   XNOR2_X1 adder_sub1_i_0_22 (.A(adder_sub1_i_0_n_86), .B(adder_sub1_i_0_n_80), 
      .ZN(adder_sub1_i_0_n_10));
   AOI21_X1 adder_sub1_i_0_23 (.A(adder_sub1_i_0_n_67), .B1(adder_sub1_i_0_n_13), 
      .B2(adder_sub1_i_0_n_12), .ZN(adder_sub1_i_0_n_11));
   AOI21_X1 adder_sub1_i_0_24 (.A(adder_sub1_i_0_n_67), .B1(adder_sub1_i_0_n_74), 
      .B2(adder_sub1_i_0_n_68), .ZN(adder_sub1_i_0_n_12));
   INV_X1 adder_sub1_i_0_25 (.A(adder_sub1_i_0_n_14), .ZN(adder_sub1_i_0_n_13));
   OAI22_X1 adder_sub1_i_0_26 (.A1(adder_sub1_i_0_n_191), .A2(
      adder_sub1_i_0_n_197), .B1(adder_sub1_i_0_n_183), .B2(adder_sub1_i_0_n_199), 
      .ZN(adder_sub1_i_0_n_14));
   NOR2_X1 adder_sub1_i_0_27 (.A1(adder_sub1_i_0_n_74), .A2(adder_sub1_i_0_n_68), 
      .ZN(adder_sub1_i_0_n_67));
   OAI22_X1 adder_sub1_i_0_28 (.A1(adder_sub1_i_0_n_45), .A2(adder_sub1_i_0_n_69), 
      .B1(adder_sub1_i_0_n_198), .B2(adder_sub1_i_0_n_51), .ZN(
      adder_sub1_i_0_n_68));
   INV_X1 adder_sub1_i_0_29 (.A(adder_sub1_i_0_n_70), .ZN(adder_sub1_i_0_n_69));
   OAI22_X1 adder_sub1_i_0_30 (.A1(adder_sub1_i_0_n_34), .A2(adder_sub1_i_0_n_83), 
      .B1(adder_sub1_i_0_n_35), .B2(adder_sub1_i_0_n_195), .ZN(
      adder_sub1_i_0_n_70));
   XNOR2_X1 adder_sub1_i_0_31 (.A(adder_sub1_Sub), .B(adder_sub1_i_0_n_75), 
      .ZN(adder_sub1_i_0_n_74));
   OAI21_X1 adder_sub1_i_0_32 (.A(adder_sub1_i_0_n_76), .B1(adder_sub1_In2[6]), 
      .B2(adder_sub1_i_0_n_30), .ZN(adder_sub1_i_0_n_75));
   OAI221_X1 adder_sub1_i_0_33 (.A(adder_sub1_i_0_n_30), .B1(adder_sub1_i_0_n_34), 
      .B2(adder_sub1_i_0_n_89), .C1(adder_sub1_i_0_n_35), .C2(
      adder_sub1_i_0_n_187), .ZN(adder_sub1_i_0_n_76));
   INV_X1 adder_sub1_i_0_34 (.A(adder_sub1_i_0_n_81), .ZN(adder_sub1_i_0_n_80));
   OAI22_X1 adder_sub1_i_0_35 (.A1(adder_sub1_i_0_n_45), .A2(adder_sub1_i_0_n_82), 
      .B1(adder_sub1_In1[7]), .B2(adder_sub1_i_0_n_51), .ZN(adder_sub1_i_0_n_81));
   AOI22_X1 adder_sub1_i_0_36 (.A1(adder_sub1_i_0_n_35), .A2(
      adder_sub1_i_0_n_102), .B1(adder_sub1_i_0_n_34), .B2(adder_sub1_i_0_n_83), 
      .ZN(adder_sub1_i_0_n_82));
   AOI22_X1 adder_sub1_i_0_37 (.A1(adder_sub1_i_0_n_46), .A2(adder_sub1_i_0_n_55), 
      .B1(adder_sub1_i_0_n_53), .B2(adder_sub1_i_0_n_143), .ZN(
      adder_sub1_i_0_n_83));
   XNOR2_X1 adder_sub1_i_0_38 (.A(adder_sub1_Sub), .B(adder_sub1_i_0_n_87), 
      .ZN(adder_sub1_i_0_n_86));
   OAI21_X1 adder_sub1_i_0_39 (.A(adder_sub1_i_0_n_88), .B1(adder_sub1_In2[7]), 
      .B2(adder_sub1_i_0_n_30), .ZN(adder_sub1_i_0_n_87));
   OAI221_X1 adder_sub1_i_0_40 (.A(adder_sub1_i_0_n_30), .B1(adder_sub1_i_0_n_34), 
      .B2(adder_sub1_i_0_n_97), .C1(adder_sub1_i_0_n_35), .C2(
      adder_sub1_i_0_n_89), .ZN(adder_sub1_i_0_n_88));
   INV_X1 adder_sub1_i_0_41 (.A(adder_sub1_i_0_n_90), .ZN(adder_sub1_i_0_n_89));
   OAI22_X1 adder_sub1_i_0_42 (.A1(adder_sub1_i_0_n_42), .A2(
      adder_sub1_i_0_n_137), .B1(adder_sub1_i_0_n_38), .B2(adder_sub1_i_0_n_52), 
      .ZN(adder_sub1_i_0_n_90));
   INV_X1 adder_sub1_i_0_43 (.A(adder_sub1_i_0_n_93), .ZN(adder_sub1_i_0_n_92));
   NOR2_X1 adder_sub1_i_0_44 (.A1(adder_sub1_i_0_n_100), .A2(adder_sub1_i_0_n_94), 
      .ZN(adder_sub1_i_0_n_93));
   XOR2_X1 adder_sub1_i_0_45 (.A(adder_sub1_Sub), .B(adder_sub1_i_0_n_95), 
      .Z(adder_sub1_i_0_n_94));
   OAI21_X1 adder_sub1_i_0_46 (.A(adder_sub1_i_0_n_96), .B1(adder_sub1_In2[8]), 
      .B2(adder_sub1_i_0_n_30), .ZN(adder_sub1_i_0_n_95));
   OAI221_X1 adder_sub1_i_0_47 (.A(adder_sub1_i_0_n_30), .B1(adder_sub1_i_0_n_35), 
      .B2(adder_sub1_i_0_n_97), .C1(adder_sub1_i_0_n_34), .C2(
      adder_sub1_i_0_n_110), .ZN(adder_sub1_i_0_n_96));
   INV_X1 adder_sub1_i_0_48 (.A(adder_sub1_i_0_n_98), .ZN(adder_sub1_i_0_n_97));
   OAI22_X1 adder_sub1_i_0_49 (.A1(adder_sub1_i_0_n_42), .A2(
      adder_sub1_i_0_n_170), .B1(adder_sub1_i_0_n_38), .B2(adder_sub1_i_0_n_41), 
      .ZN(adder_sub1_i_0_n_98));
   OAI22_X1 adder_sub1_i_0_50 (.A1(adder_sub1_i_0_n_45), .A2(
      adder_sub1_i_0_n_101), .B1(adder_sub1_In1[8]), .B2(adder_sub1_i_0_n_51), 
      .ZN(adder_sub1_i_0_n_100));
   AOI22_X1 adder_sub1_i_0_51 (.A1(adder_sub1_i_0_n_35), .A2(
      adder_sub1_i_0_n_116), .B1(adder_sub1_i_0_n_34), .B2(adder_sub1_i_0_n_102), 
      .ZN(adder_sub1_i_0_n_101));
   INV_X1 adder_sub1_i_0_52 (.A(adder_sub1_i_0_n_103), .ZN(adder_sub1_i_0_n_102));
   OAI22_X1 adder_sub1_i_0_53 (.A1(adder_sub1_i_0_n_53), .A2(adder_sub1_i_0_n_49), 
      .B1(adder_sub1_i_0_n_46), .B2(adder_sub1_i_0_n_152), .ZN(
      adder_sub1_i_0_n_103));
   AOI21_X1 adder_sub1_i_0_54 (.A(adder_sub1_i_0_n_106), .B1(
      adder_sub1_i_0_n_114), .B2(adder_sub1_i_0_n_107), .ZN(adder_sub1_i_0_n_105));
   NOR2_X1 adder_sub1_i_0_55 (.A1(adder_sub1_i_0_n_114), .A2(
      adder_sub1_i_0_n_107), .ZN(adder_sub1_i_0_n_106));
   XOR2_X1 adder_sub1_i_0_56 (.A(adder_sub1_Sub), .B(adder_sub1_i_0_n_108), 
      .Z(adder_sub1_i_0_n_107));
   OAI21_X1 adder_sub1_i_0_57 (.A(adder_sub1_i_0_n_109), .B1(adder_sub1_In2[9]), 
      .B2(adder_sub1_i_0_n_30), .ZN(adder_sub1_i_0_n_108));
   OAI221_X1 adder_sub1_i_0_58 (.A(adder_sub1_i_0_n_30), .B1(adder_sub1_i_0_n_34), 
      .B2(adder_sub1_i_0_n_127), .C1(adder_sub1_i_0_n_35), .C2(
      adder_sub1_i_0_n_110), .ZN(adder_sub1_i_0_n_109));
   INV_X1 adder_sub1_i_0_59 (.A(adder_sub1_i_0_n_111), .ZN(adder_sub1_i_0_n_110));
   OAI22_X1 adder_sub1_i_0_60 (.A1(adder_sub1_i_0_n_42), .A2(
      adder_sub1_i_0_n_167), .B1(adder_sub1_i_0_n_38), .B2(adder_sub1_i_0_n_43), 
      .ZN(adder_sub1_i_0_n_111));
   OAI22_X1 adder_sub1_i_0_61 (.A1(adder_sub1_i_0_n_45), .A2(
      adder_sub1_i_0_n_115), .B1(adder_sub1_In1[9]), .B2(adder_sub1_i_0_n_51), 
      .ZN(adder_sub1_i_0_n_114));
   AOI22_X1 adder_sub1_i_0_62 (.A1(adder_sub1_i_0_n_35), .A2(
      adder_sub1_i_0_n_121), .B1(adder_sub1_i_0_n_34), .B2(adder_sub1_i_0_n_116), 
      .ZN(adder_sub1_i_0_n_115));
   INV_X1 adder_sub1_i_0_63 (.A(adder_sub1_i_0_n_117), .ZN(adder_sub1_i_0_n_116));
   OAI22_X1 adder_sub1_i_0_64 (.A1(adder_sub1_i_0_n_53), .A2(adder_sub1_i_0_n_50), 
      .B1(adder_sub1_i_0_n_46), .B2(adder_sub1_i_0_n_149), .ZN(
      adder_sub1_i_0_n_117));
   OAI22_X1 adder_sub1_i_0_65 (.A1(adder_sub1_i_0_n_45), .A2(
      adder_sub1_i_0_n_120), .B1(adder_sub1_In1[10]), .B2(adder_sub1_i_0_n_51), 
      .ZN(adder_sub1_i_0_n_119));
   AOI22_X1 adder_sub1_i_0_66 (.A1(adder_sub1_i_0_n_34), .A2(
      adder_sub1_i_0_n_121), .B1(adder_sub1_i_0_n_35), .B2(adder_sub1_i_0_n_142), 
      .ZN(adder_sub1_i_0_n_120));
   OAI222_X1 adder_sub1_i_0_67 (.A1(adder_sub1_In1[9]), .A2(adder_sub1_i_0_n_56), 
      .B1(adder_sub1_i_0_n_53), .B2(adder_sub1_i_0_n_194), .C1(adder_sub1_In1[7]), 
      .C2(adder_sub1_i_0_n_153), .ZN(adder_sub1_i_0_n_121));
   XOR2_X1 adder_sub1_i_0_68 (.A(adder_sub1_Sub), .B(adder_sub1_i_0_n_125), 
      .Z(adder_sub1_i_0_n_124));
   OAI21_X1 adder_sub1_i_0_69 (.A(adder_sub1_i_0_n_126), .B1(adder_sub1_In2[10]), 
      .B2(adder_sub1_i_0_n_30), .ZN(adder_sub1_i_0_n_125));
   OAI221_X1 adder_sub1_i_0_70 (.A(adder_sub1_i_0_n_30), .B1(adder_sub1_i_0_n_35), 
      .B2(adder_sub1_i_0_n_127), .C1(adder_sub1_i_0_n_34), .C2(
      adder_sub1_i_0_n_135), .ZN(adder_sub1_i_0_n_126));
   INV_X1 adder_sub1_i_0_71 (.A(adder_sub1_i_0_n_128), .ZN(adder_sub1_i_0_n_127));
   OAI22_X1 adder_sub1_i_0_72 (.A1(adder_sub1_i_0_n_42), .A2(
      adder_sub1_i_0_n_130), .B1(adder_sub1_i_0_n_38), .B2(adder_sub1_i_0_n_184), 
      .ZN(adder_sub1_i_0_n_128));
   AOI22_X1 adder_sub1_i_0_73 (.A1(adder_sub1_In2[7]), .A2(adder_sub1_i_0_n_39), 
      .B1(adder_sub1_In2[9]), .B2(adder_sub1_i_0_n_40), .ZN(adder_sub1_i_0_n_130));
   NOR2_X1 adder_sub1_i_0_74 (.A1(adder_sub1_i_0_n_139), .A2(
      adder_sub1_i_0_n_132), .ZN(adder_sub1_i_0_n_131));
   XNOR2_X1 adder_sub1_i_0_75 (.A(adder_sub1_Sub), .B(adder_sub1_i_0_n_133), 
      .ZN(adder_sub1_i_0_n_132));
   OAI21_X1 adder_sub1_i_0_76 (.A(adder_sub1_i_0_n_134), .B1(adder_sub1_In2[11]), 
      .B2(adder_sub1_i_0_n_30), .ZN(adder_sub1_i_0_n_133));
   OAI221_X1 adder_sub1_i_0_77 (.A(adder_sub1_i_0_n_30), .B1(adder_sub1_i_0_n_35), 
      .B2(adder_sub1_i_0_n_135), .C1(adder_sub1_i_0_n_34), .C2(
      adder_sub1_i_0_n_168), .ZN(adder_sub1_i_0_n_134));
   INV_X1 adder_sub1_i_0_78 (.A(adder_sub1_i_0_n_136), .ZN(adder_sub1_i_0_n_135));
   OAI22_X1 adder_sub1_i_0_79 (.A1(adder_sub1_i_0_n_42), .A2(
      adder_sub1_i_0_n_138), .B1(adder_sub1_i_0_n_38), .B2(adder_sub1_i_0_n_137), 
      .ZN(adder_sub1_i_0_n_136));
   AOI22_X1 adder_sub1_i_0_80 (.A1(adder_sub1_In2[4]), .A2(adder_sub1_i_0_n_39), 
      .B1(adder_sub1_In2[6]), .B2(adder_sub1_i_0_n_40), .ZN(adder_sub1_i_0_n_137));
   AOI22_X1 adder_sub1_i_0_81 (.A1(adder_sub1_In2[8]), .A2(adder_sub1_i_0_n_39), 
      .B1(adder_sub1_In2[10]), .B2(adder_sub1_i_0_n_40), .ZN(
      adder_sub1_i_0_n_138));
   INV_X1 adder_sub1_i_0_82 (.A(adder_sub1_i_0_n_140), .ZN(adder_sub1_i_0_n_139));
   OAI22_X1 adder_sub1_i_0_83 (.A1(adder_sub1_i_0_n_45), .A2(
      adder_sub1_i_0_n_141), .B1(adder_sub1_In1[11]), .B2(adder_sub1_i_0_n_51), 
      .ZN(adder_sub1_i_0_n_140));
   AOI22_X1 adder_sub1_i_0_84 (.A1(adder_sub1_i_0_n_34), .A2(
      adder_sub1_i_0_n_142), .B1(adder_sub1_i_0_n_35), .B2(adder_sub1_i_0_n_150), 
      .ZN(adder_sub1_i_0_n_141));
   OAI222_X1 adder_sub1_i_0_85 (.A1(adder_sub1_In1[8]), .A2(adder_sub1_i_0_n_153), 
      .B1(adder_sub1_i_0_n_53), .B2(adder_sub1_i_0_n_143), .C1(
      adder_sub1_In1[10]), .C2(adder_sub1_i_0_n_56), .ZN(adder_sub1_i_0_n_142));
   OAI22_X1 adder_sub1_i_0_86 (.A1(adder_sub1_i_0_n_200), .A2(
      adder_sub1_i_0_n_48), .B1(adder_sub1_i_0_n_198), .B2(adder_sub1_i_0_n_47), 
      .ZN(adder_sub1_i_0_n_143));
   XNOR2_X1 adder_sub1_i_0_87 (.A(adder_sub1_Sub), .B(adder_sub1_i_0_n_145), 
      .ZN(adder_sub1_i_0_n_144));
   OAI21_X1 adder_sub1_i_0_88 (.A(adder_sub1_i_0_n_146), .B1(adder_sub1_In1[12]), 
      .B2(adder_sub1_i_0_n_51), .ZN(adder_sub1_i_0_n_145));
   OAI211_X1 adder_sub1_i_0_89 (.A(adder_sub1_i_0_n_51), .B(adder_sub1_i_0_n_147), 
      .C1(adder_sub1_i_0_n_35), .C2(adder_sub1_i_0_n_150), .ZN(
      adder_sub1_i_0_n_146));
   OAI221_X1 adder_sub1_i_0_90 (.A(adder_sub1_i_0_n_35), .B1(adder_sub1_i_0_n_53), 
      .B2(adder_sub1_i_0_n_148), .C1(adder_sub1_In1[10]), .C2(
      adder_sub1_i_0_n_153), .ZN(adder_sub1_i_0_n_147));
   INV_X1 adder_sub1_i_0_91 (.A(adder_sub1_i_0_n_149), .ZN(adder_sub1_i_0_n_148));
   AOI22_X1 adder_sub1_i_0_92 (.A1(adder_sub1_In1[6]), .A2(adder_sub1_i_0_n_47), 
      .B1(adder_sub1_In1[8]), .B2(adder_sub1_i_0_n_48), .ZN(adder_sub1_i_0_n_149));
   OAI222_X1 adder_sub1_i_0_93 (.A1(adder_sub1_In1[9]), .A2(adder_sub1_i_0_n_153), 
      .B1(adder_sub1_i_0_n_53), .B2(adder_sub1_i_0_n_151), .C1(
      adder_sub1_In1[11]), .C2(adder_sub1_i_0_n_56), .ZN(adder_sub1_i_0_n_150));
   INV_X1 adder_sub1_i_0_94 (.A(adder_sub1_i_0_n_152), .ZN(adder_sub1_i_0_n_151));
   AOI22_X1 adder_sub1_i_0_95 (.A1(adder_sub1_In1[5]), .A2(adder_sub1_i_0_n_47), 
      .B1(adder_sub1_In1[7]), .B2(adder_sub1_i_0_n_48), .ZN(adder_sub1_i_0_n_152));
   NAND2_X1 adder_sub1_i_0_96 (.A1(adder_sub1_i_0_n_53), .A2(adder_sub1_i_0_n_47), 
      .ZN(adder_sub1_i_0_n_153));
   OAI21_X1 adder_sub1_i_0_97 (.A(adder_sub1_i_0_n_162), .B1(adder_sub1_In2[12]), 
      .B2(adder_sub1_i_0_n_30), .ZN(adder_sub1_i_0_n_161));
   OAI21_X1 adder_sub1_i_0_98 (.A(adder_sub1_i_0_n_163), .B1(adder_sub1_i_0_n_35), 
      .B2(adder_sub1_i_0_n_168), .ZN(adder_sub1_i_0_n_162));
   NOR3_X1 adder_sub1_i_0_99 (.A1(adder_sub1_i_0_n_31), .A2(adder_sub1_i_0_n_164), 
      .A3(adder_sub1_i_0_n_166), .ZN(adder_sub1_i_0_n_163));
   NOR3_X1 adder_sub1_i_0_100 (.A1(adder_sub1_i_0_n_190), .A2(
      adder_sub1_i_0_n_40), .A3(adder_sub1_i_0_n_44), .ZN(adder_sub1_i_0_n_164));
   NOR3_X1 adder_sub1_i_0_101 (.A1(adder_sub1_i_0_n_34), .A2(adder_sub1_i_0_n_38), 
      .A3(adder_sub1_i_0_n_167), .ZN(adder_sub1_i_0_n_166));
   AOI22_X1 adder_sub1_i_0_102 (.A1(adder_sub1_In2[6]), .A2(adder_sub1_i_0_n_39), 
      .B1(adder_sub1_In2[8]), .B2(adder_sub1_i_0_n_40), .ZN(adder_sub1_i_0_n_167));
   INV_X1 adder_sub1_i_0_103 (.A(adder_sub1_i_0_n_169), .ZN(adder_sub1_i_0_n_168));
   OAI22_X1 adder_sub1_i_0_104 (.A1(adder_sub1_i_0_n_42), .A2(
      adder_sub1_i_0_n_171), .B1(adder_sub1_i_0_n_38), .B2(adder_sub1_i_0_n_170), 
      .ZN(adder_sub1_i_0_n_169));
   AOI22_X1 adder_sub1_i_0_105 (.A1(adder_sub1_In2[5]), .A2(adder_sub1_i_0_n_39), 
      .B1(adder_sub1_In2[7]), .B2(adder_sub1_i_0_n_40), .ZN(adder_sub1_i_0_n_170));
   AOI22_X1 adder_sub1_i_0_106 (.A1(adder_sub1_In2[9]), .A2(adder_sub1_i_0_n_39), 
      .B1(adder_sub1_In2[11]), .B2(adder_sub1_i_0_n_40), .ZN(
      adder_sub1_i_0_n_171));
   OAI22_X1 adder_sub1_i_0_193 (.A1(adder_sub1_i_0_n_17), .A2(
      adder_sub1_i_0_n_31), .B1(adder_sub1_i_0_n_32), .B2(adder_sub1_i_0_n_30), 
      .ZN(adder_sub1_Out[13]));
   OAI22_X1 adder_sub1_i_0_194 (.A1(adder_sub1_i_0_n_15), .A2(
      adder_sub1_i_0_n_31), .B1(adder_sub1_i_0_n_16), .B2(adder_sub1_i_0_n_30), 
      .ZN(adder_sub1_Out[14]));
   INV_X1 adder_sub1_i_0_107 (.A(adder_sub1_In2[10]), .ZN(adder_sub1_i_0_n_190));
   INV_X1 adder_sub1_i_0_108 (.A(adder_sub1_In1[6]), .ZN(adder_sub1_i_0_n_198));
   INV_X1 adder_sub1_i_0_109 (.A(adder_sub1_In1[14]), .ZN(adder_sub1_i_0_n_15));
   INV_X1 adder_sub1_i_0_110 (.A(adder_sub1_In2[14]), .ZN(adder_sub1_i_0_n_16));
   INV_X1 adder_sub1_i_0_111 (.A(adder_sub1_In1[13]), .ZN(adder_sub1_i_0_n_17));
   INV_X1 adder_sub1_i_0_112 (.A(adder_sub1_In2[15]), .ZN(adder_sub1_i_0_n_18));
   INV_X1 adder_sub1_i_0_113 (.A(adder_sub1_In1[15]), .ZN(adder_sub1_i_0_n_19));
   NAND2_X1 adder_sub1_i_0_114 (.A1(adder_sub1_i_0_n_18), .A2(
      adder_sub1_i_0_n_19), .ZN(adder_sub1_Out[15]));
   NAND2_X1 adder_sub1_i_0_115 (.A1(adder_sub1_i_0_n_16), .A2(adder_sub1_In1[14]), 
      .ZN(adder_sub1_i_0_n_20));
   NAND2_X1 adder_sub1_i_0_116 (.A1(adder_sub1_i_0_n_15), .A2(adder_sub1_In2[14]), 
      .ZN(adder_sub1_i_0_n_21));
   NAND2_X1 adder_sub1_i_0_117 (.A1(adder_sub1_i_0_n_20), .A2(
      adder_sub1_i_0_n_21), .ZN(adder_sub1_i_0_n_22));
   INV_X1 adder_sub1_i_0_118 (.A(adder_sub1_i_0_n_22), .ZN(adder_sub1_i_0_n_23));
   NOR2_X1 adder_sub1_i_0_119 (.A1(adder_sub1_i_0_n_17), .A2(adder_sub1_In2[13]), 
      .ZN(adder_sub1_i_0_n_24));
   NAND2_X1 adder_sub1_i_0_120 (.A1(adder_sub1_i_0_n_23), .A2(
      adder_sub1_i_0_n_24), .ZN(adder_sub1_i_0_n_25));
   NAND2_X1 adder_sub1_i_0_121 (.A1(adder_sub1_i_0_n_25), .A2(
      adder_sub1_i_0_n_20), .ZN(adder_sub1_i_0_n_26));
   OAI21_X1 adder_sub1_i_0_122 (.A(adder_sub1_Out[15]), .B1(adder_sub1_i_0_n_18), 
      .B2(adder_sub1_i_0_n_19), .ZN(adder_sub1_i_0_n_27));
   NAND2_X1 adder_sub1_i_0_123 (.A1(adder_sub1_i_0_n_26), .A2(
      adder_sub1_i_0_n_27), .ZN(adder_sub1_i_0_n_28));
   NAND2_X1 adder_sub1_i_0_124 (.A1(adder_sub1_i_0_n_18), .A2(adder_sub1_In1[15]), 
      .ZN(adder_sub1_i_0_n_29));
   NAND2_X1 adder_sub1_i_0_125 (.A1(adder_sub1_i_0_n_28), .A2(
      adder_sub1_i_0_n_29), .ZN(adder_sub1_i_0_n_30));
   INV_X1 adder_sub1_i_0_126 (.A(adder_sub1_i_0_n_30), .ZN(adder_sub1_i_0_n_31));
   INV_X1 adder_sub1_i_0_127 (.A(adder_sub1_In2[13]), .ZN(adder_sub1_i_0_n_32));
   NOR2_X1 adder_sub1_i_0_128 (.A1(adder_sub1_i_0_n_32), .A2(adder_sub1_In1[13]), 
      .ZN(adder_sub1_i_0_n_33));
   OR2_X1 adder_sub1_i_0_129 (.A1(adder_sub1_i_0_n_24), .A2(adder_sub1_i_0_n_33), 
      .ZN(adder_sub1_i_0_n_34));
   INV_X1 adder_sub1_i_0_130 (.A(adder_sub1_i_0_n_34), .ZN(adder_sub1_i_0_n_35));
   NAND2_X1 adder_sub1_i_0_131 (.A1(adder_sub1_i_0_n_23), .A2(
      adder_sub1_i_0_n_33), .ZN(adder_sub1_i_0_n_36));
   NAND2_X1 adder_sub1_i_0_132 (.A1(adder_sub1_i_0_n_36), .A2(
      adder_sub1_i_0_n_21), .ZN(adder_sub1_i_0_n_37));
   XOR2_X1 adder_sub1_i_0_133 (.A(adder_sub1_i_0_n_37), .B(adder_sub1_i_0_n_27), 
      .Z(adder_sub1_i_0_n_38));
   OAI21_X1 adder_sub1_i_0_134 (.A(adder_sub1_i_0_n_36), .B1(adder_sub1_i_0_n_23), 
      .B2(adder_sub1_i_0_n_33), .ZN(adder_sub1_i_0_n_39));
   INV_X1 adder_sub1_i_0_135 (.A(adder_sub1_i_0_n_39), .ZN(adder_sub1_i_0_n_40));
   OAI22_X1 adder_sub1_i_0_136 (.A1(adder_sub1_i_0_n_40), .A2(adder_sub1_In2[1]), 
      .B1(adder_sub1_i_0_n_39), .B2(adder_sub1_In2[3]), .ZN(adder_sub1_i_0_n_41));
   INV_X1 adder_sub1_i_0_137 (.A(adder_sub1_i_0_n_38), .ZN(adder_sub1_i_0_n_42));
   OAI22_X1 adder_sub1_i_0_138 (.A1(adder_sub1_i_0_n_40), .A2(adder_sub1_In2[2]), 
      .B1(adder_sub1_i_0_n_39), .B2(adder_sub1_In2[4]), .ZN(adder_sub1_i_0_n_43));
   NAND2_X1 adder_sub1_i_0_139 (.A1(adder_sub1_i_0_n_38), .A2(
      adder_sub1_i_0_n_35), .ZN(adder_sub1_i_0_n_44));
   OAI21_X1 adder_sub1_i_0_140 (.A(adder_sub1_i_0_n_31), .B1(adder_sub1_i_0_n_44), 
      .B2(adder_sub1_i_0_n_22), .ZN(adder_sub1_i_0_n_45));
   OAI21_X1 adder_sub1_i_0_141 (.A(adder_sub1_i_0_n_28), .B1(adder_sub1_i_0_n_26), 
      .B2(adder_sub1_i_0_n_27), .ZN(adder_sub1_i_0_n_46));
   OAI21_X1 adder_sub1_i_0_142 (.A(adder_sub1_i_0_n_25), .B1(adder_sub1_i_0_n_23), 
      .B2(adder_sub1_i_0_n_24), .ZN(adder_sub1_i_0_n_47));
   INV_X1 adder_sub1_i_0_143 (.A(adder_sub1_i_0_n_47), .ZN(adder_sub1_i_0_n_48));
   OAI22_X1 adder_sub1_i_0_144 (.A1(adder_sub1_i_0_n_48), .A2(adder_sub1_In1[1]), 
      .B1(adder_sub1_i_0_n_47), .B2(adder_sub1_In1[3]), .ZN(adder_sub1_i_0_n_49));
   OAI22_X1 adder_sub1_i_0_145 (.A1(adder_sub1_i_0_n_48), .A2(adder_sub1_In1[2]), 
      .B1(adder_sub1_i_0_n_47), .B2(adder_sub1_In1[4]), .ZN(adder_sub1_i_0_n_50));
   INV_X1 adder_sub1_i_0_146 (.A(adder_sub1_i_0_n_45), .ZN(adder_sub1_i_0_n_51));
   OAI22_X1 adder_sub1_i_0_147 (.A1(adder_sub1_i_0_n_40), .A2(adder_sub1_In2[0]), 
      .B1(adder_sub1_i_0_n_39), .B2(adder_sub1_In2[2]), .ZN(adder_sub1_i_0_n_52));
   INV_X1 adder_sub1_i_0_148 (.A(adder_sub1_i_0_n_46), .ZN(adder_sub1_i_0_n_53));
   OAI22_X1 adder_sub1_i_0_149 (.A1(adder_sub1_i_0_n_48), .A2(adder_sub1_In1[0]), 
      .B1(adder_sub1_i_0_n_47), .B2(adder_sub1_In1[2]), .ZN(adder_sub1_i_0_n_54));
   INV_X1 adder_sub1_i_0_150 (.A(adder_sub1_i_0_n_54), .ZN(adder_sub1_i_0_n_55));
   NAND2_X1 adder_sub1_i_0_151 (.A1(adder_sub1_i_0_n_53), .A2(
      adder_sub1_i_0_n_48), .ZN(adder_sub1_i_0_n_56));
   NAND2_X1 adder_sub1_i_0_152 (.A1(adder_sub1_i_0_n_45), .A2(adder_sub1_In1[0]), 
      .ZN(adder_sub1_i_0_n_57));
   AND2_X1 adder_sub1_i_0_153 (.A1(adder_sub1_i_0_n_31), .A2(adder_sub1_In2[0]), 
      .ZN(adder_sub1_i_0_n_58));
   NAND2_X1 adder_sub1_i_0_154 (.A1(adder_sub1_i_0_n_57), .A2(
      adder_sub1_i_0_n_58), .ZN(adder_sub1_i_0_n_59));
   OAI21_X1 adder_sub1_i_0_155 (.A(adder_sub1_i_0_n_59), .B1(adder_sub1_Sub), 
      .B2(adder_sub1_i_0_n_58), .ZN(adder_sub1_i_0_n_60));
   NAND2_X1 adder_sub1_i_0_156 (.A1(adder_sub1_i_0_n_38), .A2(
      adder_sub1_i_0_n_34), .ZN(adder_sub1_i_0_n_61));
   NAND2_X1 adder_sub1_i_0_157 (.A1(adder_sub1_i_0_n_40), .A2(adder_sub1_In2[0]), 
      .ZN(adder_sub1_i_0_n_62));
   NOR3_X1 adder_sub1_i_0_158 (.A1(adder_sub1_i_0_n_61), .A2(adder_sub1_i_0_n_31), 
      .A3(adder_sub1_i_0_n_62), .ZN(adder_sub1_i_0_n_63));
   AOI21_X1 adder_sub1_i_0_159 (.A(adder_sub1_i_0_n_63), .B1(adder_sub1_In2[1]), 
      .B2(adder_sub1_i_0_n_31), .ZN(adder_sub1_i_0_n_64));
   XOR2_X1 adder_sub1_i_0_160 (.A(adder_sub1_i_0_n_64), .B(adder_sub1_Sub), 
      .Z(adder_sub1_i_0_n_65));
   INV_X1 adder_sub1_i_0_161 (.A(adder_sub1_i_0_n_29), .ZN(adder_sub1_i_0_n_66));
   NOR3_X1 adder_sub1_i_0_162 (.A1(adder_sub1_i_0_n_56), .A2(adder_sub1_i_0_n_66), 
      .A3(adder_sub1_i_0_n_35), .ZN(adder_sub1_i_0_n_71));
   AOI22_X1 adder_sub1_i_0_163 (.A1(adder_sub1_i_0_n_71), .A2(adder_sub1_In1[0]), 
      .B1(adder_sub1_i_0_n_45), .B2(adder_sub1_In1[1]), .ZN(adder_sub1_i_0_n_72));
   XOR2_X1 adder_sub1_i_0_164 (.A(adder_sub1_i_0_n_65), .B(adder_sub1_i_0_n_72), 
      .Z(adder_sub1_i_0_n_73));
   AOI22_X1 adder_sub1_i_0_165 (.A1(adder_sub1_i_0_n_73), .A2(
      adder_sub1_i_0_n_60), .B1(adder_sub1_i_0_n_65), .B2(adder_sub1_i_0_n_72), 
      .ZN(adder_sub1_i_0_n_77));
   INV_X1 adder_sub1_i_0_166 (.A(adder_sub1_i_0_n_77), .ZN(adder_sub1_i_0_n_78));
   INV_X1 adder_sub1_i_0_167 (.A(adder_sub1_In2[1]), .ZN(adder_sub1_i_0_n_79));
   OAI33_X1 adder_sub1_i_0_168 (.A1(adder_sub1_i_0_n_61), .A2(
      adder_sub1_i_0_n_79), .A3(adder_sub1_i_0_n_39), .B1(adder_sub1_i_0_n_42), 
      .B2(adder_sub1_i_0_n_52), .B3(adder_sub1_i_0_n_34), .ZN(
      adder_sub1_i_0_n_84));
   AOI22_X1 adder_sub1_i_0_169 (.A1(adder_sub1_i_0_n_84), .A2(
      adder_sub1_i_0_n_30), .B1(adder_sub1_In2[2]), .B2(adder_sub1_i_0_n_31), 
      .ZN(adder_sub1_i_0_n_85));
   XNOR2_X1 adder_sub1_i_0_170 (.A(adder_sub1_i_0_n_85), .B(adder_sub1_Sub), 
      .ZN(adder_sub1_i_0_n_91));
   AOI21_X1 adder_sub1_i_0_171 (.A(adder_sub1_i_0_n_35), .B1(adder_sub1_i_0_n_48), 
      .B2(adder_sub1_In1[1]), .ZN(adder_sub1_i_0_n_99));
   AOI211_X1 adder_sub1_i_0_172 (.A(adder_sub1_i_0_n_99), .B(adder_sub1_i_0_n_46), 
      .C1(adder_sub1_i_0_n_54), .C2(adder_sub1_i_0_n_35), .ZN(
      adder_sub1_i_0_n_104));
   OAI22_X1 adder_sub1_i_0_173 (.A1(adder_sub1_i_0_n_104), .A2(
      adder_sub1_i_0_n_45), .B1(adder_sub1_i_0_n_51), .B2(adder_sub1_In1[2]), 
      .ZN(adder_sub1_i_0_n_112));
   XNOR2_X1 adder_sub1_i_0_174 (.A(adder_sub1_i_0_n_91), .B(adder_sub1_i_0_n_112), 
      .ZN(adder_sub1_i_0_n_113));
   INV_X1 adder_sub1_i_0_175 (.A(adder_sub1_i_0_n_113), .ZN(adder_sub1_i_0_n_118));
   INV_X1 adder_sub1_i_0_176 (.A(adder_sub1_i_0_n_112), .ZN(adder_sub1_i_0_n_122));
   OAI22_X1 adder_sub1_i_0_177 (.A1(adder_sub1_i_0_n_118), .A2(
      adder_sub1_i_0_n_77), .B1(adder_sub1_i_0_n_91), .B2(adder_sub1_i_0_n_122), 
      .ZN(adder_sub1_i_0_n_123));
   OAI22_X1 adder_sub1_i_0_178 (.A1(adder_sub1_i_0_n_61), .A2(
      adder_sub1_i_0_n_52), .B1(adder_sub1_i_0_n_44), .B2(adder_sub1_i_0_n_41), 
      .ZN(adder_sub1_i_0_n_129));
   AOI22_X1 adder_sub1_i_0_179 (.A1(adder_sub1_i_0_n_129), .A2(
      adder_sub1_i_0_n_30), .B1(adder_sub1_In2[3]), .B2(adder_sub1_i_0_n_31), 
      .ZN(adder_sub1_i_0_n_154));
   XOR2_X1 adder_sub1_i_0_180 (.A(adder_sub1_i_0_n_154), .B(adder_sub1_Sub), 
      .Z(adder_sub1_i_0_n_155));
   AOI221_X1 adder_sub1_i_0_181 (.A(adder_sub1_i_0_n_46), .B1(
      adder_sub1_i_0_n_49), .B2(adder_sub1_i_0_n_35), .C1(adder_sub1_i_0_n_34), 
      .C2(adder_sub1_i_0_n_54), .ZN(adder_sub1_i_0_n_156));
   OAI22_X1 adder_sub1_i_0_182 (.A1(adder_sub1_i_0_n_156), .A2(
      adder_sub1_i_0_n_45), .B1(adder_sub1_i_0_n_51), .B2(adder_sub1_In1[3]), 
      .ZN(adder_sub1_i_0_n_157));
   XOR2_X1 adder_sub1_i_0_183 (.A(adder_sub1_i_0_n_155), .B(adder_sub1_i_0_n_157), 
      .Z(adder_sub1_i_0_n_158));
   AOI22_X1 adder_sub1_i_0_184 (.A1(adder_sub1_i_0_n_123), .A2(
      adder_sub1_i_0_n_158), .B1(adder_sub1_i_0_n_155), .B2(adder_sub1_i_0_n_157), 
      .ZN(adder_sub1_i_0_n_159));
   NOR2_X1 adder_sub1_i_0_185 (.A1(adder_sub1_i_0_n_53), .A2(adder_sub1_i_0_n_47), 
      .ZN(adder_sub1_i_0_n_160));
   INV_X1 adder_sub1_i_0_186 (.A(adder_sub1_i_0_n_50), .ZN(adder_sub1_i_0_n_165));
   AOI22_X1 adder_sub1_i_0_187 (.A1(adder_sub1_i_0_n_160), .A2(adder_sub1_In1[0]), 
      .B1(adder_sub1_i_0_n_53), .B2(adder_sub1_i_0_n_165), .ZN(
      adder_sub1_i_0_n_172));
   OAI33_X1 adder_sub1_i_0_188 (.A1(adder_sub1_i_0_n_172), .A2(
      adder_sub1_i_0_n_24), .A3(adder_sub1_i_0_n_33), .B1(adder_sub1_i_0_n_49), 
      .B2(adder_sub1_i_0_n_46), .B3(adder_sub1_i_0_n_35), .ZN(
      adder_sub1_i_0_n_173));
   OAI22_X1 adder_sub1_i_0_189 (.A1(adder_sub1_i_0_n_173), .A2(
      adder_sub1_i_0_n_45), .B1(adder_sub1_In1[4]), .B2(adder_sub1_i_0_n_51), 
      .ZN(adder_sub1_i_0_n_174));
   INV_X1 adder_sub1_i_0_190 (.A(adder_sub1_i_0_n_43), .ZN(adder_sub1_i_0_n_175));
   INV_X1 adder_sub1_i_0_191 (.A(adder_sub1_i_0_n_62), .ZN(adder_sub1_i_0_n_176));
   AOI22_X1 adder_sub1_i_0_192 (.A1(adder_sub1_i_0_n_38), .A2(
      adder_sub1_i_0_n_175), .B1(adder_sub1_i_0_n_42), .B2(adder_sub1_i_0_n_176), 
      .ZN(adder_sub1_i_0_n_177));
   OAI22_X1 adder_sub1_i_0_195 (.A1(adder_sub1_i_0_n_177), .A2(
      adder_sub1_i_0_n_34), .B1(adder_sub1_i_0_n_61), .B2(adder_sub1_i_0_n_41), 
      .ZN(adder_sub1_i_0_n_178));
   AOI22_X1 adder_sub1_i_0_196 (.A1(adder_sub1_i_0_n_178), .A2(
      adder_sub1_i_0_n_30), .B1(adder_sub1_In2[4]), .B2(adder_sub1_i_0_n_31), 
      .ZN(adder_sub1_i_0_n_179));
   XOR2_X1 adder_sub1_i_0_197 (.A(adder_sub1_i_0_n_179), .B(adder_sub1_Sub), 
      .Z(adder_sub1_i_0_n_180));
   NAND2_X1 adder_sub1_i_0_198 (.A1(adder_sub1_i_0_n_174), .A2(
      adder_sub1_i_0_n_180), .ZN(adder_sub1_i_0_n_181));
   OAI21_X1 adder_sub1_i_0_199 (.A(adder_sub1_i_0_n_181), .B1(
      adder_sub1_i_0_n_174), .B2(adder_sub1_i_0_n_180), .ZN(adder_sub1_i_0_n_182));
   OAI21_X1 adder_sub1_i_0_200 (.A(adder_sub1_i_0_n_181), .B1(
      adder_sub1_i_0_n_159), .B2(adder_sub1_i_0_n_182), .ZN(adder_sub1_i_0_n_183));
   OAI22_X1 adder_sub1_i_0_201 (.A1(adder_sub1_i_0_n_40), .A2(adder_sub1_In2[3]), 
      .B1(adder_sub1_i_0_n_39), .B2(adder_sub1_In2[5]), .ZN(adder_sub1_i_0_n_184));
   INV_X1 adder_sub1_i_0_202 (.A(adder_sub1_i_0_n_184), .ZN(adder_sub1_i_0_n_185));
   NOR2_X1 adder_sub1_i_0_203 (.A1(adder_sub1_i_0_n_39), .A2(adder_sub1_i_0_n_79), 
      .ZN(adder_sub1_i_0_n_186));
   OAI22_X1 adder_sub1_i_0_204 (.A1(adder_sub1_i_0_n_42), .A2(
      adder_sub1_i_0_n_185), .B1(adder_sub1_i_0_n_38), .B2(adder_sub1_i_0_n_186), 
      .ZN(adder_sub1_i_0_n_187));
   OAI22_X1 adder_sub1_i_0_205 (.A1(adder_sub1_i_0_n_177), .A2(
      adder_sub1_i_0_n_35), .B1(adder_sub1_i_0_n_187), .B2(adder_sub1_i_0_n_34), 
      .ZN(adder_sub1_i_0_n_188));
   AOI22_X1 adder_sub1_i_0_206 (.A1(adder_sub1_i_0_n_188), .A2(
      adder_sub1_i_0_n_30), .B1(adder_sub1_In2[5]), .B2(adder_sub1_i_0_n_31), 
      .ZN(adder_sub1_i_0_n_189));
   XOR2_X1 adder_sub1_i_0_207 (.A(adder_sub1_i_0_n_189), .B(adder_sub1_Sub), 
      .Z(adder_sub1_i_0_n_191));
   INV_X1 adder_sub1_i_0_208 (.A(adder_sub1_In1[5]), .ZN(adder_sub1_i_0_n_192));
   INV_X1 adder_sub1_i_0_209 (.A(adder_sub1_In1[3]), .ZN(adder_sub1_i_0_n_193));
   AOI22_X1 adder_sub1_i_0_210 (.A1(adder_sub1_i_0_n_48), .A2(
      adder_sub1_i_0_n_192), .B1(adder_sub1_i_0_n_47), .B2(adder_sub1_i_0_n_193), 
      .ZN(adder_sub1_i_0_n_194));
   AOI22_X1 adder_sub1_i_0_211 (.A1(adder_sub1_i_0_n_160), .A2(adder_sub1_In1[1]), 
      .B1(adder_sub1_i_0_n_53), .B2(adder_sub1_i_0_n_194), .ZN(
      adder_sub1_i_0_n_195));
   AOI22_X1 adder_sub1_i_0_212 (.A1(adder_sub1_i_0_n_195), .A2(
      adder_sub1_i_0_n_35), .B1(adder_sub1_i_0_n_172), .B2(adder_sub1_i_0_n_34), 
      .ZN(adder_sub1_i_0_n_196));
   OAI22_X1 adder_sub1_i_0_213 (.A1(adder_sub1_i_0_n_196), .A2(
      adder_sub1_i_0_n_45), .B1(adder_sub1_In1[5]), .B2(adder_sub1_i_0_n_51), 
      .ZN(adder_sub1_i_0_n_197));
   XNOR2_X1 adder_sub1_i_0_214 (.A(adder_sub1_i_0_n_191), .B(
      adder_sub1_i_0_n_197), .ZN(adder_sub1_i_0_n_199));
   XOR2_X1 adder_sub1_i_0_215 (.A(adder_sub1_i_0_n_183), .B(adder_sub1_i_0_n_199), 
      .Z(adder_sub1_Out[5]));
   INV_X1 adder_sub1_i_0_216 (.A(adder_sub1_In1[4]), .ZN(adder_sub1_i_0_n_200));
   XOR2_X1 adder_sub2_i_0_0 (.A(adder_sub2_In1[0]), .B(adder_sub2_In2[0]), 
      .Z(n_178));
   XNOR2_X1 adder_sub2_i_0_1 (.A(adder_sub2_i_0_n_3), .B(adder_sub2_i_0_n_15), 
      .ZN(n_179));
   XNOR2_X1 adder_sub2_i_0_2 (.A(adder_sub2_i_0_n_24), .B(adder_sub2_i_0_n_22), 
      .ZN(n_180));
   XNOR2_X1 adder_sub2_i_0_3 (.A(adder_sub2_In1[6]), .B(adder_sub2_i_0_n_12), 
      .ZN(n_181));
   XNOR2_X1 adder_sub2_i_0_4 (.A(adder_sub2_i_0_n_11), .B(adder_sub2_i_0_n_2), 
      .ZN(n_182));
   XOR2_X1 adder_sub2_i_0_5 (.A(adder_sub2_In1[7]), .B(adder_sub2_In2[8]), 
      .Z(adder_sub2_i_0_n_2));
   XNOR2_X1 adder_sub2_i_0_6 (.A(adder_sub2_i_0_n_9), .B(adder_sub2_i_0_n_25), 
      .ZN(n_183));
   XOR2_X1 adder_sub2_i_0_7 (.A(adder_sub2_In1[9]), .B(adder_sub2_i_0_n_8), 
      .Z(n_184));
   NOR2_X1 adder_sub2_i_0_8 (.A1(adder_sub2_i_0_n_5), .A2(adder_sub2_i_0_n_4), 
      .ZN(n_185));
   AOI21_X1 adder_sub2_i_0_9 (.A(adder_sub2_In1[10]), .B1(adder_sub2_i_0_n_8), 
      .B2(adder_sub2_In1[9]), .ZN(adder_sub2_i_0_n_4));
   XNOR2_X1 adder_sub2_i_0_10 (.A(adder_sub2_In1[11]), .B(adder_sub2_i_0_n_6), 
      .ZN(n_186));
   INV_X1 adder_sub2_i_0_11 (.A(adder_sub2_i_0_n_6), .ZN(adder_sub2_i_0_n_5));
   NAND3_X1 adder_sub2_i_0_12 (.A1(adder_sub2_i_0_n_8), .A2(adder_sub2_In1[9]), 
      .A3(adder_sub2_In1[10]), .ZN(adder_sub2_i_0_n_6));
   XNOR2_X1 adder_sub2_i_0_13 (.A(adder_sub2_In1[12]), .B(adder_sub2_i_0_n_7), 
      .ZN(n_187));
   NAND4_X1 adder_sub2_i_0_14 (.A1(adder_sub2_i_0_n_8), .A2(adder_sub2_In1[9]), 
      .A3(adder_sub2_In1[10]), .A4(adder_sub2_In1[11]), .ZN(adder_sub2_i_0_n_7));
   AOI21_X1 adder_sub2_i_0_15 (.A(adder_sub2_i_0_n_27), .B1(adder_sub2_i_0_n_9), 
      .B2(adder_sub2_i_0_n_28), .ZN(adder_sub2_i_0_n_8));
   OAI21_X1 adder_sub2_i_0_16 (.A(adder_sub2_i_0_n_10), .B1(adder_sub2_In2[8]), 
      .B2(adder_sub2_In1[7]), .ZN(adder_sub2_i_0_n_9));
   NAND2_X1 adder_sub2_i_0_17 (.A1(adder_sub2_i_0_n_26), .A2(adder_sub2_i_0_n_11), 
      .ZN(adder_sub2_i_0_n_10));
   OAI211_X1 adder_sub2_i_0_18 (.A(adder_sub2_i_0_n_13), .B(adder_sub2_In1[6]), 
      .C1(adder_sub2_In1[5]), .C2(adder_sub2_In2[5]), .ZN(adder_sub2_i_0_n_11));
   OAI21_X1 adder_sub2_i_0_19 (.A(adder_sub2_i_0_n_13), .B1(adder_sub2_In2[5]), 
      .B2(adder_sub2_In1[5]), .ZN(adder_sub2_i_0_n_12));
   INV_X1 adder_sub2_i_0_20 (.A(adder_sub2_i_0_n_14), .ZN(adder_sub2_i_0_n_13));
   AOI21_X1 adder_sub2_i_0_21 (.A(adder_sub2_i_0_n_21), .B1(adder_sub2_In2[5]), 
      .B2(adder_sub2_In1[5]), .ZN(adder_sub2_i_0_n_14));
   NAND2_X1 adder_sub2_i_0_22 (.A1(adder_sub2_In1[7]), .A2(adder_sub2_In2[8]), 
      .ZN(adder_sub2_i_0_n_26));
   XOR2_X1 adder_sub2_i_0_23 (.A(adder_sub2_i_0_n_1), .B(adder_sub2_i_0_n_0), 
      .Z(n_188));
   XOR2_X1 adder_sub2_i_0_24 (.A(adder_sub2_In1[2]), .B(adder_sub2_In2[2]), 
      .Z(adder_sub2_i_0_n_0));
   AOI21_X1 adder_sub2_i_0_25 (.A(adder_sub2_i_0_n_16), .B1(adder_sub2_i_0_n_15), 
      .B2(adder_sub2_i_0_n_3), .ZN(adder_sub2_i_0_n_1));
   NAND2_X1 adder_sub2_i_0_26 (.A1(adder_sub2_In1[0]), .A2(adder_sub2_In2[0]), 
      .ZN(adder_sub2_i_0_n_3));
   AOI21_X1 adder_sub2_i_0_27 (.A(adder_sub2_i_0_n_16), .B1(adder_sub2_In1[1]), 
      .B2(adder_sub2_In2[1]), .ZN(adder_sub2_i_0_n_15));
   NOR2_X1 adder_sub2_i_0_28 (.A1(adder_sub2_In1[1]), .A2(adder_sub2_In2[1]), 
      .ZN(adder_sub2_i_0_n_16));
   XNOR2_X1 adder_sub2_i_0_29 (.A(adder_sub2_In1[3]), .B(adder_sub2_i_0_n_17), 
      .ZN(n_189));
   OAI21_X1 adder_sub2_i_0_30 (.A(adder_sub2_i_0_n_18), .B1(adder_sub2_In1[2]), 
      .B2(adder_sub2_In2[2]), .ZN(adder_sub2_i_0_n_17));
   INV_X1 adder_sub2_i_0_31 (.A(adder_sub2_i_0_n_19), .ZN(adder_sub2_i_0_n_18));
   AOI21_X1 adder_sub2_i_0_32 (.A(adder_sub2_i_0_n_1), .B1(adder_sub2_In1[2]), 
      .B2(adder_sub2_In2[2]), .ZN(adder_sub2_i_0_n_19));
   XOR2_X1 adder_sub2_i_0_33 (.A(adder_sub2_i_0_n_21), .B(adder_sub2_i_0_n_20), 
      .Z(n_190));
   XOR2_X1 adder_sub2_i_0_34 (.A(adder_sub2_In1[5]), .B(adder_sub2_In2[5]), 
      .Z(adder_sub2_i_0_n_20));
   AOI21_X1 adder_sub2_i_0_35 (.A(adder_sub2_i_0_n_23), .B1(adder_sub2_i_0_n_24), 
      .B2(adder_sub2_i_0_n_22), .ZN(adder_sub2_i_0_n_21));
   AOI21_X1 adder_sub2_i_0_36 (.A(adder_sub2_i_0_n_23), .B1(adder_sub2_In1[4]), 
      .B2(adder_sub2_In2[4]), .ZN(adder_sub2_i_0_n_22));
   NOR2_X1 adder_sub2_i_0_37 (.A1(adder_sub2_In1[4]), .A2(adder_sub2_In2[4]), 
      .ZN(adder_sub2_i_0_n_23));
   OAI211_X1 adder_sub2_i_0_38 (.A(adder_sub2_In1[3]), .B(adder_sub2_i_0_n_18), 
      .C1(adder_sub2_In1[2]), .C2(adder_sub2_In2[2]), .ZN(adder_sub2_i_0_n_24));
   AOI21_X1 adder_sub2_i_0_39 (.A(adder_sub2_i_0_n_27), .B1(adder_sub2_In1[8]), 
      .B2(adder_sub2_In2[8]), .ZN(adder_sub2_i_0_n_25));
   NOR2_X1 adder_sub2_i_0_40 (.A1(adder_sub2_In1[8]), .A2(adder_sub2_In2[8]), 
      .ZN(adder_sub2_i_0_n_27));
   NAND2_X1 adder_sub2_i_0_41 (.A1(adder_sub2_In1[8]), .A2(adder_sub2_In2[8]), 
      .ZN(adder_sub2_i_0_n_28));
   XOR2_X1 i_2_0_0 (.A(adder_sub3_In1[0]), .B(adder_sub3_In2[0]), .Z(n_191));
   XNOR2_X1 i_2_0_1 (.A(adder_sub3_In1[1]), .B(n_2_0_1), .ZN(n_192));
   XNOR2_X1 i_2_0_2 (.A(adder_sub3_In1[2]), .B(n_2_0_0), .ZN(n_193));
   NAND3_X1 i_2_0_3 (.A1(adder_sub3_In1[1]), .A2(adder_sub3_In1[0]), .A3(
      adder_sub3_In2[0]), .ZN(n_2_0_0));
   NAND2_X1 i_2_0_4 (.A1(adder_sub3_In1[0]), .A2(adder_sub3_In2[0]), .ZN(n_2_0_1));
endmodule
