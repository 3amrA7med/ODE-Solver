/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Apr 24 04:09:15 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 230966499 */

module add_sub_cla__0_283__GU(enable, sub, in1, in2, cin, out, cout, invalid);
   input enable;
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   wire [19:0]tempIn11;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;

   DLH_X1 \tempIn11_reg[12]  (.D(n_12), .G(n_13), .Q(tempIn11[12]));
   DLH_X1 \tempIn11_reg[11]  (.D(n_11), .G(n_13), .Q(tempIn11[11]));
   DLH_X1 \tempIn11_reg[10]  (.D(n_10), .G(n_13), .Q(tempIn11[10]));
   DLH_X1 \tempIn11_reg[9]  (.D(n_9), .G(n_13), .Q(tempIn11[9]));
   DLH_X1 \tempIn11_reg[8]  (.D(n_8), .G(n_13), .Q(tempIn11[8]));
   DLH_X1 \tempIn11_reg[7]  (.D(n_7), .G(n_13), .Q(tempIn11[7]));
   DLH_X1 \tempIn11_reg[6]  (.D(n_6), .G(n_13), .Q(tempIn11[6]));
   DLH_X1 \tempIn11_reg[5]  (.D(n_5), .G(n_13), .Q(tempIn11[5]));
   DLH_X1 \tempIn11_reg[4]  (.D(n_4), .G(n_13), .Q(tempIn11[4]));
   DLH_X1 \tempIn11_reg[3]  (.D(n_3), .G(n_13), .Q(tempIn11[3]));
   DLH_X1 \tempIn11_reg[2]  (.D(n_2), .G(n_13), .Q(tempIn11[2]));
   DLH_X1 \tempIn11_reg[1]  (.D(n_1), .G(n_13), .Q(tempIn11[1]));
   DLH_X1 \tempIn11_reg[0]  (.D(n_0), .G(n_13), .Q(tempIn11[0]));
   AND2_X1 i_0_0 (.A1(in1[0]), .A2(n_13), .ZN(n_0));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(n_1));
   NAND4_X1 i_0_2 (.A1(in1[15]), .A2(in1[14]), .A3(in1[13]), .A4(in1[0]), 
      .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in1[1]), .A2(n_13), .ZN(n_0_1));
   OAI21_X1 i_0_4 (.A(n_0_2), .B1(n_0_4), .B2(in1[13]), .ZN(n_2));
   NAND4_X1 i_0_5 (.A1(in1[15]), .A2(in1[14]), .A3(in1[13]), .A4(in1[1]), 
      .ZN(n_0_2));
   OAI21_X1 i_0_6 (.A(n_0_3), .B1(n_0_4), .B2(n_0_36), .ZN(n_3));
   NAND3_X1 i_0_7 (.A1(n_0_14), .A2(n_0_33), .A3(n_0_36), .ZN(n_0_3));
   NAND2_X1 i_0_8 (.A1(n_0_12), .A2(n_0_33), .ZN(n_0_4));
   OAI21_X1 i_0_9 (.A(n_0_5), .B1(n_0_7), .B2(in1[13]), .ZN(n_4));
   NAND3_X1 i_0_10 (.A1(in1[15]), .A2(in1[13]), .A3(n_0_14), .ZN(n_0_5));
   OAI21_X1 i_0_11 (.A(n_0_6), .B1(n_0_7), .B2(n_0_36), .ZN(n_5));
   OR2_X1 i_0_12 (.A1(in1[13]), .A2(n_0_9), .ZN(n_0_6));
   AOI22_X1 i_0_13 (.A1(n_0_16), .A2(n_0_33), .B1(in1[0]), .B2(n_0_10), .ZN(
      n_0_7));
   OAI21_X1 i_0_14 (.A(n_0_8), .B1(n_0_9), .B2(n_0_36), .ZN(n_6));
   NAND2_X1 i_0_15 (.A1(n_0_11), .A2(n_0_36), .ZN(n_0_8));
   AOI22_X1 i_0_16 (.A1(n_0_18), .A2(n_0_33), .B1(in1[1]), .B2(n_0_10), .ZN(
      n_0_9));
   NOR2_X1 i_0_17 (.A1(n_0_33), .A2(n_0_31), .ZN(n_0_10));
   MUX2_X1 i_0_18 (.A(n_0_13), .B(n_0_11), .S(in1[13]), .Z(n_7));
   MUX2_X1 i_0_19 (.A(n_0_12), .B(n_0_21), .S(n_0_33), .Z(n_0_11));
   MUX2_X1 i_0_20 (.A(in1[0]), .B(in1[2]), .S(n_0_32), .Z(n_0_12));
   MUX2_X1 i_0_21 (.A(n_0_15), .B(n_0_13), .S(in1[13]), .Z(n_8));
   MUX2_X1 i_0_22 (.A(n_0_14), .B(n_0_25), .S(n_0_33), .Z(n_0_13));
   MUX2_X1 i_0_23 (.A(in1[1]), .B(in1[3]), .S(n_0_32), .Z(n_0_14));
   MUX2_X1 i_0_24 (.A(n_0_17), .B(n_0_15), .S(in1[13]), .Z(n_9));
   MUX2_X1 i_0_25 (.A(n_0_16), .B(n_0_30), .S(n_0_33), .Z(n_0_15));
   MUX2_X1 i_0_26 (.A(in1[2]), .B(in1[4]), .S(n_0_32), .Z(n_0_16));
   MUX2_X1 i_0_27 (.A(n_0_20), .B(n_0_17), .S(in1[13]), .Z(n_10));
   MUX2_X1 i_0_28 (.A(n_0_18), .B(n_0_19), .S(n_0_33), .Z(n_0_17));
   MUX2_X1 i_0_29 (.A(in1[3]), .B(in1[5]), .S(n_0_32), .Z(n_0_18));
   MUX2_X1 i_0_30 (.A(in1[7]), .B(in1[9]), .S(n_0_32), .Z(n_0_19));
   MUX2_X1 i_0_31 (.A(n_0_24), .B(n_0_20), .S(in1[13]), .Z(n_11));
   MUX2_X1 i_0_32 (.A(n_0_21), .B(n_0_22), .S(n_0_33), .Z(n_0_20));
   MUX2_X1 i_0_33 (.A(in1[4]), .B(in1[6]), .S(n_0_32), .Z(n_0_21));
   MUX2_X1 i_0_34 (.A(in1[8]), .B(in1[10]), .S(n_0_32), .Z(n_0_22));
   OAI21_X1 i_0_35 (.A(n_0_23), .B1(n_0_27), .B2(in1[13]), .ZN(n_12));
   NAND2_X1 i_0_36 (.A1(in1[13]), .A2(n_0_24), .ZN(n_0_23));
   MUX2_X1 i_0_37 (.A(n_0_25), .B(n_0_26), .S(n_0_33), .Z(n_0_24));
   MUX2_X1 i_0_38 (.A(in1[5]), .B(in1[7]), .S(n_0_32), .Z(n_0_25));
   MUX2_X1 i_0_39 (.A(in1[9]), .B(in1[11]), .S(n_0_32), .Z(n_0_26));
   OAI21_X1 i_0_40 (.A(n_0_28), .B1(n_0_30), .B2(n_0_33), .ZN(n_0_27));
   OAI211_X1 i_0_41 (.A(n_0_33), .B(n_0_29), .C1(in1[14]), .C2(n_0_35), .ZN(
      n_0_28));
   NAND2_X1 i_0_42 (.A1(in1[10]), .A2(n_0_31), .ZN(n_0_29));
   MUX2_X1 i_0_43 (.A(in1[6]), .B(in1[8]), .S(n_0_32), .Z(n_0_30));
   INV_X1 i_0_44 (.A(n_0_32), .ZN(n_0_31));
   XNOR2_X1 i_0_45 (.A(in1[14]), .B(in1[13]), .ZN(n_0_32));
   XOR2_X1 i_0_46 (.A(in1[15]), .B(n_0_34), .Z(n_0_33));
   NOR3_X1 i_0_47 (.A1(in1[15]), .A2(in1[14]), .A3(in1[13]), .ZN(n_13));
   NOR2_X1 i_0_48 (.A1(in1[14]), .A2(in1[13]), .ZN(n_0_34));
   INV_X1 i_0_49 (.A(in1[12]), .ZN(n_0_35));
   INV_X1 i_0_50 (.A(in1[13]), .ZN(n_0_36));
   XNOR2_X1 i_1_0 (.A(tempIn11[1]), .B(out[0]), .ZN(out[1]));
   NOR2_X1 i_1_1 (.A1(n_1_10), .A2(n_1_0), .ZN(out[2]));
   AOI21_X1 i_1_2 (.A(tempIn11[2]), .B1(tempIn11[1]), .B2(tempIn11[0]), .ZN(
      n_1_0));
   XNOR2_X1 i_1_3 (.A(tempIn11[3]), .B(n_1_11), .ZN(out[3]));
   XOR2_X1 i_1_4 (.A(tempIn11[4]), .B(n_1_9), .Z(out[4]));
   NOR2_X1 i_1_5 (.A1(n_1_8), .A2(n_1_1), .ZN(out[5]));
   AOI21_X1 i_1_6 (.A(tempIn11[5]), .B1(tempIn11[4]), .B2(n_1_9), .ZN(n_1_1));
   XOR2_X1 i_1_7 (.A(tempIn11[6]), .B(n_1_8), .Z(out[6]));
   XNOR2_X1 i_1_8 (.A(tempIn11[7]), .B(n_1_2), .ZN(out[7]));
   NAND2_X1 i_1_9 (.A1(tempIn11[6]), .A2(n_1_8), .ZN(n_1_2));
   XOR2_X1 i_1_10 (.A(tempIn11[8]), .B(n_1_7), .Z(out[8]));
   XNOR2_X1 i_1_11 (.A(tempIn11[9]), .B(n_1_3), .ZN(out[9]));
   NAND2_X1 i_1_12 (.A1(tempIn11[8]), .A2(n_1_7), .ZN(n_1_3));
   XOR2_X1 i_1_13 (.A(tempIn11[10]), .B(n_1_6), .Z(out[10]));
   XNOR2_X1 i_1_14 (.A(tempIn11[11]), .B(n_1_4), .ZN(out[11]));
   NAND2_X1 i_1_15 (.A1(tempIn11[10]), .A2(n_1_6), .ZN(n_1_4));
   XNOR2_X1 i_1_16 (.A(tempIn11[12]), .B(n_1_5), .ZN(out[12]));
   NAND3_X1 i_1_17 (.A1(tempIn11[11]), .A2(tempIn11[10]), .A3(n_1_6), .ZN(n_1_5));
   AND3_X1 i_1_18 (.A1(tempIn11[9]), .A2(tempIn11[8]), .A3(n_1_7), .ZN(n_1_6));
   AND3_X1 i_1_19 (.A1(tempIn11[7]), .A2(tempIn11[6]), .A3(n_1_8), .ZN(n_1_7));
   AND3_X1 i_1_20 (.A1(tempIn11[5]), .A2(tempIn11[4]), .A3(n_1_9), .ZN(n_1_8));
   AND2_X1 i_1_21 (.A1(tempIn11[3]), .A2(n_1_10), .ZN(n_1_9));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_1_10));
   NAND3_X1 i_1_23 (.A1(tempIn11[2]), .A2(tempIn11[1]), .A3(tempIn11[0]), 
      .ZN(n_1_11));
   INV_X1 i_1_24 (.A(tempIn11[0]), .ZN(out[0]));
endmodule

module add_sub_cla__0_254__GU(enable, sub, in1, in2, cin, out, cout, invalid);
   input enable;
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   wire [19:0]tempIn11;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;

   DLH_X1 \tempIn11_reg[12]  (.D(n_12), .G(n_13), .Q(tempIn11[12]));
   DLH_X1 \tempIn11_reg[11]  (.D(n_11), .G(n_13), .Q(tempIn11[11]));
   DLH_X1 \tempIn11_reg[10]  (.D(n_10), .G(n_13), .Q(tempIn11[10]));
   DLH_X1 \tempIn11_reg[9]  (.D(n_9), .G(n_13), .Q(tempIn11[9]));
   DLH_X1 \tempIn11_reg[8]  (.D(n_8), .G(n_13), .Q(tempIn11[8]));
   DLH_X1 \tempIn11_reg[7]  (.D(n_7), .G(n_13), .Q(tempIn11[7]));
   DLH_X1 \tempIn11_reg[6]  (.D(n_6), .G(n_13), .Q(tempIn11[6]));
   DLH_X1 \tempIn11_reg[5]  (.D(n_5), .G(n_13), .Q(tempIn11[5]));
   DLH_X1 \tempIn11_reg[4]  (.D(n_4), .G(n_13), .Q(tempIn11[4]));
   DLH_X1 \tempIn11_reg[3]  (.D(n_3), .G(n_13), .Q(tempIn11[3]));
   DLH_X1 \tempIn11_reg[2]  (.D(n_2), .G(n_13), .Q(tempIn11[2]));
   DLH_X1 \tempIn11_reg[1]  (.D(n_1), .G(n_13), .Q(tempIn11[1]));
   DLH_X1 \tempIn11_reg[0]  (.D(n_0), .G(n_13), .Q(tempIn11[0]));
   AND2_X1 i_0_0 (.A1(in1[0]), .A2(n_13), .ZN(n_0));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(n_1));
   NAND4_X1 i_0_2 (.A1(in1[15]), .A2(in1[14]), .A3(in1[13]), .A4(in1[0]), 
      .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in1[1]), .A2(n_13), .ZN(n_0_1));
   OAI21_X1 i_0_4 (.A(n_0_2), .B1(n_0_4), .B2(in1[13]), .ZN(n_2));
   NAND4_X1 i_0_5 (.A1(in1[15]), .A2(in1[14]), .A3(in1[13]), .A4(in1[1]), 
      .ZN(n_0_2));
   OAI21_X1 i_0_6 (.A(n_0_3), .B1(n_0_4), .B2(n_0_36), .ZN(n_3));
   NAND3_X1 i_0_7 (.A1(n_0_14), .A2(n_0_33), .A3(n_0_36), .ZN(n_0_3));
   NAND2_X1 i_0_8 (.A1(n_0_12), .A2(n_0_33), .ZN(n_0_4));
   OAI21_X1 i_0_9 (.A(n_0_5), .B1(n_0_7), .B2(in1[13]), .ZN(n_4));
   NAND3_X1 i_0_10 (.A1(in1[15]), .A2(in1[13]), .A3(n_0_14), .ZN(n_0_5));
   OAI21_X1 i_0_11 (.A(n_0_6), .B1(n_0_7), .B2(n_0_36), .ZN(n_5));
   OR2_X1 i_0_12 (.A1(in1[13]), .A2(n_0_9), .ZN(n_0_6));
   AOI22_X1 i_0_13 (.A1(n_0_16), .A2(n_0_33), .B1(in1[0]), .B2(n_0_10), .ZN(
      n_0_7));
   OAI21_X1 i_0_14 (.A(n_0_8), .B1(n_0_9), .B2(n_0_36), .ZN(n_6));
   NAND2_X1 i_0_15 (.A1(n_0_11), .A2(n_0_36), .ZN(n_0_8));
   AOI22_X1 i_0_16 (.A1(n_0_18), .A2(n_0_33), .B1(in1[1]), .B2(n_0_10), .ZN(
      n_0_9));
   NOR2_X1 i_0_17 (.A1(n_0_33), .A2(n_0_31), .ZN(n_0_10));
   MUX2_X1 i_0_18 (.A(n_0_13), .B(n_0_11), .S(in1[13]), .Z(n_7));
   MUX2_X1 i_0_19 (.A(n_0_12), .B(n_0_21), .S(n_0_33), .Z(n_0_11));
   MUX2_X1 i_0_20 (.A(in1[0]), .B(in1[2]), .S(n_0_32), .Z(n_0_12));
   MUX2_X1 i_0_21 (.A(n_0_15), .B(n_0_13), .S(in1[13]), .Z(n_8));
   MUX2_X1 i_0_22 (.A(n_0_14), .B(n_0_25), .S(n_0_33), .Z(n_0_13));
   MUX2_X1 i_0_23 (.A(in1[1]), .B(in1[3]), .S(n_0_32), .Z(n_0_14));
   MUX2_X1 i_0_24 (.A(n_0_17), .B(n_0_15), .S(in1[13]), .Z(n_9));
   MUX2_X1 i_0_25 (.A(n_0_16), .B(n_0_30), .S(n_0_33), .Z(n_0_15));
   MUX2_X1 i_0_26 (.A(in1[2]), .B(in1[4]), .S(n_0_32), .Z(n_0_16));
   MUX2_X1 i_0_27 (.A(n_0_20), .B(n_0_17), .S(in1[13]), .Z(n_10));
   MUX2_X1 i_0_28 (.A(n_0_18), .B(n_0_19), .S(n_0_33), .Z(n_0_17));
   MUX2_X1 i_0_29 (.A(in1[3]), .B(in1[5]), .S(n_0_32), .Z(n_0_18));
   MUX2_X1 i_0_30 (.A(in1[7]), .B(in1[9]), .S(n_0_32), .Z(n_0_19));
   MUX2_X1 i_0_31 (.A(n_0_24), .B(n_0_20), .S(in1[13]), .Z(n_11));
   MUX2_X1 i_0_32 (.A(n_0_21), .B(n_0_22), .S(n_0_33), .Z(n_0_20));
   MUX2_X1 i_0_33 (.A(in1[4]), .B(in1[6]), .S(n_0_32), .Z(n_0_21));
   MUX2_X1 i_0_34 (.A(in1[8]), .B(in1[10]), .S(n_0_32), .Z(n_0_22));
   OAI21_X1 i_0_35 (.A(n_0_23), .B1(n_0_27), .B2(in1[13]), .ZN(n_12));
   NAND2_X1 i_0_36 (.A1(in1[13]), .A2(n_0_24), .ZN(n_0_23));
   MUX2_X1 i_0_37 (.A(n_0_25), .B(n_0_26), .S(n_0_33), .Z(n_0_24));
   MUX2_X1 i_0_38 (.A(in1[5]), .B(in1[7]), .S(n_0_32), .Z(n_0_25));
   MUX2_X1 i_0_39 (.A(in1[9]), .B(in1[11]), .S(n_0_32), .Z(n_0_26));
   OAI21_X1 i_0_40 (.A(n_0_28), .B1(n_0_30), .B2(n_0_33), .ZN(n_0_27));
   OAI211_X1 i_0_41 (.A(n_0_33), .B(n_0_29), .C1(in1[14]), .C2(n_0_35), .ZN(
      n_0_28));
   NAND2_X1 i_0_42 (.A1(in1[10]), .A2(n_0_31), .ZN(n_0_29));
   MUX2_X1 i_0_43 (.A(in1[6]), .B(in1[8]), .S(n_0_32), .Z(n_0_30));
   INV_X1 i_0_44 (.A(n_0_32), .ZN(n_0_31));
   XNOR2_X1 i_0_45 (.A(in1[14]), .B(in1[13]), .ZN(n_0_32));
   XOR2_X1 i_0_46 (.A(in1[15]), .B(n_0_34), .Z(n_0_33));
   NOR3_X1 i_0_47 (.A1(in1[15]), .A2(in1[14]), .A3(in1[13]), .ZN(n_13));
   NOR2_X1 i_0_48 (.A1(in1[14]), .A2(in1[13]), .ZN(n_0_34));
   INV_X1 i_0_49 (.A(in1[12]), .ZN(n_0_35));
   INV_X1 i_0_50 (.A(in1[13]), .ZN(n_0_36));
   XNOR2_X1 i_1_0 (.A(tempIn11[1]), .B(out[0]), .ZN(out[1]));
   NOR2_X1 i_1_1 (.A1(n_1_10), .A2(n_1_0), .ZN(out[2]));
   AOI21_X1 i_1_2 (.A(tempIn11[2]), .B1(tempIn11[1]), .B2(tempIn11[0]), .ZN(
      n_1_0));
   XNOR2_X1 i_1_3 (.A(tempIn11[3]), .B(n_1_11), .ZN(out[3]));
   XOR2_X1 i_1_4 (.A(tempIn11[4]), .B(n_1_9), .Z(out[4]));
   NOR2_X1 i_1_5 (.A1(n_1_8), .A2(n_1_1), .ZN(out[5]));
   AOI21_X1 i_1_6 (.A(tempIn11[5]), .B1(tempIn11[4]), .B2(n_1_9), .ZN(n_1_1));
   XOR2_X1 i_1_7 (.A(tempIn11[6]), .B(n_1_8), .Z(out[6]));
   XNOR2_X1 i_1_8 (.A(tempIn11[7]), .B(n_1_2), .ZN(out[7]));
   NAND2_X1 i_1_9 (.A1(tempIn11[6]), .A2(n_1_8), .ZN(n_1_2));
   XOR2_X1 i_1_10 (.A(tempIn11[8]), .B(n_1_7), .Z(out[8]));
   XNOR2_X1 i_1_11 (.A(tempIn11[9]), .B(n_1_3), .ZN(out[9]));
   NAND2_X1 i_1_12 (.A1(tempIn11[8]), .A2(n_1_7), .ZN(n_1_3));
   XOR2_X1 i_1_13 (.A(tempIn11[10]), .B(n_1_6), .Z(out[10]));
   XNOR2_X1 i_1_14 (.A(tempIn11[11]), .B(n_1_4), .ZN(out[11]));
   NAND2_X1 i_1_15 (.A1(tempIn11[10]), .A2(n_1_6), .ZN(n_1_4));
   XNOR2_X1 i_1_16 (.A(tempIn11[12]), .B(n_1_5), .ZN(out[12]));
   NAND3_X1 i_1_17 (.A1(tempIn11[11]), .A2(tempIn11[10]), .A3(n_1_6), .ZN(n_1_5));
   AND3_X1 i_1_18 (.A1(tempIn11[9]), .A2(tempIn11[8]), .A3(n_1_7), .ZN(n_1_6));
   AND3_X1 i_1_19 (.A1(tempIn11[7]), .A2(tempIn11[6]), .A3(n_1_8), .ZN(n_1_7));
   AND3_X1 i_1_20 (.A1(tempIn11[5]), .A2(tempIn11[4]), .A3(n_1_9), .ZN(n_1_8));
   AND2_X1 i_1_21 (.A1(tempIn11[3]), .A2(n_1_10), .ZN(n_1_9));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_1_10));
   NAND3_X1 i_1_23 (.A1(tempIn11[2]), .A2(tempIn11[1]), .A3(tempIn11[0]), 
      .ZN(n_1_11));
   INV_X1 i_1_24 (.A(tempIn11[0]), .ZN(out[0]));
endmodule

module add_sub_cla__GU(enable, sub, in1, in2, cin, out, cout, invalid);
   input enable;
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   wire [19:0]tempIn11;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;

   DLH_X1 \tempIn11_reg[12]  (.D(n_12), .G(n_13), .Q(tempIn11[12]));
   DLH_X1 \tempIn11_reg[11]  (.D(n_11), .G(n_13), .Q(tempIn11[11]));
   DLH_X1 \tempIn11_reg[10]  (.D(n_10), .G(n_13), .Q(tempIn11[10]));
   DLH_X1 \tempIn11_reg[9]  (.D(n_9), .G(n_13), .Q(tempIn11[9]));
   DLH_X1 \tempIn11_reg[8]  (.D(n_8), .G(n_13), .Q(tempIn11[8]));
   DLH_X1 \tempIn11_reg[7]  (.D(n_7), .G(n_13), .Q(tempIn11[7]));
   DLH_X1 \tempIn11_reg[6]  (.D(n_6), .G(n_13), .Q(tempIn11[6]));
   DLH_X1 \tempIn11_reg[5]  (.D(n_5), .G(n_13), .Q(tempIn11[5]));
   DLH_X1 \tempIn11_reg[4]  (.D(n_4), .G(n_13), .Q(tempIn11[4]));
   DLH_X1 \tempIn11_reg[3]  (.D(n_3), .G(n_13), .Q(tempIn11[3]));
   DLH_X1 \tempIn11_reg[2]  (.D(n_2), .G(n_13), .Q(tempIn11[2]));
   DLH_X1 \tempIn11_reg[1]  (.D(n_1), .G(n_13), .Q(tempIn11[1]));
   DLH_X1 \tempIn11_reg[0]  (.D(n_0), .G(n_13), .Q(tempIn11[0]));
   AND2_X1 i_0_0 (.A1(in1[0]), .A2(n_13), .ZN(n_0));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(n_1));
   NAND4_X1 i_0_2 (.A1(in1[15]), .A2(in1[14]), .A3(in1[13]), .A4(in1[0]), 
      .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in1[1]), .A2(n_13), .ZN(n_0_1));
   OAI21_X1 i_0_4 (.A(n_0_2), .B1(n_0_4), .B2(in1[13]), .ZN(n_2));
   NAND4_X1 i_0_5 (.A1(in1[15]), .A2(in1[14]), .A3(in1[13]), .A4(in1[1]), 
      .ZN(n_0_2));
   OAI21_X1 i_0_6 (.A(n_0_3), .B1(n_0_4), .B2(n_0_36), .ZN(n_3));
   NAND3_X1 i_0_7 (.A1(n_0_14), .A2(n_0_33), .A3(n_0_36), .ZN(n_0_3));
   NAND2_X1 i_0_8 (.A1(n_0_12), .A2(n_0_33), .ZN(n_0_4));
   OAI21_X1 i_0_9 (.A(n_0_5), .B1(n_0_7), .B2(in1[13]), .ZN(n_4));
   NAND3_X1 i_0_10 (.A1(in1[15]), .A2(in1[13]), .A3(n_0_14), .ZN(n_0_5));
   OAI21_X1 i_0_11 (.A(n_0_6), .B1(n_0_7), .B2(n_0_36), .ZN(n_5));
   OR2_X1 i_0_12 (.A1(in1[13]), .A2(n_0_9), .ZN(n_0_6));
   AOI22_X1 i_0_13 (.A1(n_0_16), .A2(n_0_33), .B1(in1[0]), .B2(n_0_10), .ZN(
      n_0_7));
   OAI21_X1 i_0_14 (.A(n_0_8), .B1(n_0_9), .B2(n_0_36), .ZN(n_6));
   NAND2_X1 i_0_15 (.A1(n_0_11), .A2(n_0_36), .ZN(n_0_8));
   AOI22_X1 i_0_16 (.A1(n_0_18), .A2(n_0_33), .B1(in1[1]), .B2(n_0_10), .ZN(
      n_0_9));
   NOR2_X1 i_0_17 (.A1(n_0_33), .A2(n_0_31), .ZN(n_0_10));
   MUX2_X1 i_0_18 (.A(n_0_13), .B(n_0_11), .S(in1[13]), .Z(n_7));
   MUX2_X1 i_0_19 (.A(n_0_12), .B(n_0_21), .S(n_0_33), .Z(n_0_11));
   MUX2_X1 i_0_20 (.A(in1[0]), .B(in1[2]), .S(n_0_32), .Z(n_0_12));
   MUX2_X1 i_0_21 (.A(n_0_15), .B(n_0_13), .S(in1[13]), .Z(n_8));
   MUX2_X1 i_0_22 (.A(n_0_14), .B(n_0_25), .S(n_0_33), .Z(n_0_13));
   MUX2_X1 i_0_23 (.A(in1[1]), .B(in1[3]), .S(n_0_32), .Z(n_0_14));
   MUX2_X1 i_0_24 (.A(n_0_17), .B(n_0_15), .S(in1[13]), .Z(n_9));
   MUX2_X1 i_0_25 (.A(n_0_16), .B(n_0_30), .S(n_0_33), .Z(n_0_15));
   MUX2_X1 i_0_26 (.A(in1[2]), .B(in1[4]), .S(n_0_32), .Z(n_0_16));
   MUX2_X1 i_0_27 (.A(n_0_20), .B(n_0_17), .S(in1[13]), .Z(n_10));
   MUX2_X1 i_0_28 (.A(n_0_18), .B(n_0_19), .S(n_0_33), .Z(n_0_17));
   MUX2_X1 i_0_29 (.A(in1[3]), .B(in1[5]), .S(n_0_32), .Z(n_0_18));
   MUX2_X1 i_0_30 (.A(in1[7]), .B(in1[9]), .S(n_0_32), .Z(n_0_19));
   MUX2_X1 i_0_31 (.A(n_0_24), .B(n_0_20), .S(in1[13]), .Z(n_11));
   MUX2_X1 i_0_32 (.A(n_0_21), .B(n_0_22), .S(n_0_33), .Z(n_0_20));
   MUX2_X1 i_0_33 (.A(in1[4]), .B(in1[6]), .S(n_0_32), .Z(n_0_21));
   MUX2_X1 i_0_34 (.A(in1[8]), .B(in1[10]), .S(n_0_32), .Z(n_0_22));
   OAI21_X1 i_0_35 (.A(n_0_23), .B1(n_0_27), .B2(in1[13]), .ZN(n_12));
   NAND2_X1 i_0_36 (.A1(in1[13]), .A2(n_0_24), .ZN(n_0_23));
   MUX2_X1 i_0_37 (.A(n_0_25), .B(n_0_26), .S(n_0_33), .Z(n_0_24));
   MUX2_X1 i_0_38 (.A(in1[5]), .B(in1[7]), .S(n_0_32), .Z(n_0_25));
   MUX2_X1 i_0_39 (.A(in1[9]), .B(in1[11]), .S(n_0_32), .Z(n_0_26));
   OAI21_X1 i_0_40 (.A(n_0_28), .B1(n_0_30), .B2(n_0_33), .ZN(n_0_27));
   OAI211_X1 i_0_41 (.A(n_0_33), .B(n_0_29), .C1(in1[14]), .C2(n_0_35), .ZN(
      n_0_28));
   NAND2_X1 i_0_42 (.A1(in1[10]), .A2(n_0_31), .ZN(n_0_29));
   MUX2_X1 i_0_43 (.A(in1[6]), .B(in1[8]), .S(n_0_32), .Z(n_0_30));
   INV_X1 i_0_44 (.A(n_0_32), .ZN(n_0_31));
   XNOR2_X1 i_0_45 (.A(in1[14]), .B(in1[13]), .ZN(n_0_32));
   XOR2_X1 i_0_46 (.A(in1[15]), .B(n_0_34), .Z(n_0_33));
   NOR3_X1 i_0_47 (.A1(in1[15]), .A2(in1[14]), .A3(in1[13]), .ZN(n_13));
   NOR2_X1 i_0_48 (.A1(in1[14]), .A2(in1[13]), .ZN(n_0_34));
   INV_X1 i_0_49 (.A(in1[12]), .ZN(n_0_35));
   INV_X1 i_0_50 (.A(in1[13]), .ZN(n_0_36));
   XNOR2_X1 i_1_0 (.A(tempIn11[1]), .B(out[0]), .ZN(out[1]));
   NOR2_X1 i_1_1 (.A1(n_1_10), .A2(n_1_0), .ZN(out[2]));
   AOI21_X1 i_1_2 (.A(tempIn11[2]), .B1(tempIn11[1]), .B2(tempIn11[0]), .ZN(
      n_1_0));
   XNOR2_X1 i_1_3 (.A(tempIn11[3]), .B(n_1_11), .ZN(out[3]));
   XOR2_X1 i_1_4 (.A(tempIn11[4]), .B(n_1_9), .Z(out[4]));
   NOR2_X1 i_1_5 (.A1(n_1_8), .A2(n_1_1), .ZN(out[5]));
   AOI21_X1 i_1_6 (.A(tempIn11[5]), .B1(tempIn11[4]), .B2(n_1_9), .ZN(n_1_1));
   XOR2_X1 i_1_7 (.A(tempIn11[6]), .B(n_1_8), .Z(out[6]));
   XNOR2_X1 i_1_8 (.A(tempIn11[7]), .B(n_1_2), .ZN(out[7]));
   NAND2_X1 i_1_9 (.A1(tempIn11[6]), .A2(n_1_8), .ZN(n_1_2));
   XOR2_X1 i_1_10 (.A(tempIn11[8]), .B(n_1_7), .Z(out[8]));
   XNOR2_X1 i_1_11 (.A(tempIn11[9]), .B(n_1_3), .ZN(out[9]));
   NAND2_X1 i_1_12 (.A1(tempIn11[8]), .A2(n_1_7), .ZN(n_1_3));
   XOR2_X1 i_1_13 (.A(tempIn11[10]), .B(n_1_6), .Z(out[10]));
   XNOR2_X1 i_1_14 (.A(tempIn11[11]), .B(n_1_4), .ZN(out[11]));
   NAND2_X1 i_1_15 (.A1(tempIn11[10]), .A2(n_1_6), .ZN(n_1_4));
   XNOR2_X1 i_1_16 (.A(tempIn11[12]), .B(n_1_5), .ZN(out[12]));
   NAND3_X1 i_1_17 (.A1(tempIn11[11]), .A2(tempIn11[10]), .A3(n_1_6), .ZN(n_1_5));
   AND3_X1 i_1_18 (.A1(tempIn11[9]), .A2(tempIn11[8]), .A3(n_1_7), .ZN(n_1_6));
   AND3_X1 i_1_19 (.A1(tempIn11[7]), .A2(tempIn11[6]), .A3(n_1_8), .ZN(n_1_7));
   AND3_X1 i_1_20 (.A1(tempIn11[5]), .A2(tempIn11[4]), .A3(n_1_9), .ZN(n_1_8));
   AND2_X1 i_1_21 (.A1(tempIn11[3]), .A2(n_1_10), .ZN(n_1_9));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_1_10));
   NAND3_X1 i_1_23 (.A1(tempIn11[2]), .A2(tempIn11[1]), .A3(tempIn11[0]), 
      .ZN(n_1_11));
   INV_X1 i_1_24 (.A(tempIn11[0]), .ZN(out[0]));
endmodule

module add_sub_cla__0_312__GU(enable, sub, in1, in2, cin, out, cout, invalid);
   input enable;
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   wire [19:0]tempIn11;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;

   DLH_X1 \tempIn11_reg[12]  (.D(n_12), .G(n_13), .Q(tempIn11[12]));
   DLH_X1 \tempIn11_reg[11]  (.D(n_11), .G(n_13), .Q(tempIn11[11]));
   DLH_X1 \tempIn11_reg[10]  (.D(n_10), .G(n_13), .Q(tempIn11[10]));
   DLH_X1 \tempIn11_reg[9]  (.D(n_9), .G(n_13), .Q(tempIn11[9]));
   DLH_X1 \tempIn11_reg[8]  (.D(n_8), .G(n_13), .Q(tempIn11[8]));
   DLH_X1 \tempIn11_reg[7]  (.D(n_7), .G(n_13), .Q(tempIn11[7]));
   DLH_X1 \tempIn11_reg[6]  (.D(n_6), .G(n_13), .Q(tempIn11[6]));
   DLH_X1 \tempIn11_reg[5]  (.D(n_5), .G(n_13), .Q(tempIn11[5]));
   DLH_X1 \tempIn11_reg[4]  (.D(n_4), .G(n_13), .Q(tempIn11[4]));
   DLH_X1 \tempIn11_reg[3]  (.D(n_3), .G(n_13), .Q(tempIn11[3]));
   DLH_X1 \tempIn11_reg[2]  (.D(n_2), .G(n_13), .Q(tempIn11[2]));
   DLH_X1 \tempIn11_reg[1]  (.D(n_1), .G(n_13), .Q(tempIn11[1]));
   DLH_X1 \tempIn11_reg[0]  (.D(n_0), .G(n_13), .Q(tempIn11[0]));
   AND2_X1 i_0_0 (.A1(in1[0]), .A2(n_13), .ZN(n_0));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(n_1));
   NAND4_X1 i_0_2 (.A1(in1[15]), .A2(in1[14]), .A3(in1[13]), .A4(in1[0]), 
      .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(in1[1]), .A2(n_13), .ZN(n_0_1));
   OAI21_X1 i_0_4 (.A(n_0_2), .B1(n_0_4), .B2(in1[13]), .ZN(n_2));
   NAND4_X1 i_0_5 (.A1(in1[15]), .A2(in1[14]), .A3(in1[13]), .A4(in1[1]), 
      .ZN(n_0_2));
   OAI21_X1 i_0_6 (.A(n_0_3), .B1(n_0_4), .B2(n_0_36), .ZN(n_3));
   NAND3_X1 i_0_7 (.A1(n_0_14), .A2(n_0_33), .A3(n_0_36), .ZN(n_0_3));
   NAND2_X1 i_0_8 (.A1(n_0_12), .A2(n_0_33), .ZN(n_0_4));
   OAI21_X1 i_0_9 (.A(n_0_5), .B1(n_0_7), .B2(in1[13]), .ZN(n_4));
   NAND3_X1 i_0_10 (.A1(in1[15]), .A2(in1[13]), .A3(n_0_14), .ZN(n_0_5));
   OAI21_X1 i_0_11 (.A(n_0_6), .B1(n_0_7), .B2(n_0_36), .ZN(n_5));
   OR2_X1 i_0_12 (.A1(in1[13]), .A2(n_0_9), .ZN(n_0_6));
   AOI22_X1 i_0_13 (.A1(n_0_16), .A2(n_0_33), .B1(in1[0]), .B2(n_0_10), .ZN(
      n_0_7));
   OAI21_X1 i_0_14 (.A(n_0_8), .B1(n_0_9), .B2(n_0_36), .ZN(n_6));
   NAND2_X1 i_0_15 (.A1(n_0_11), .A2(n_0_36), .ZN(n_0_8));
   AOI22_X1 i_0_16 (.A1(n_0_18), .A2(n_0_33), .B1(in1[1]), .B2(n_0_10), .ZN(
      n_0_9));
   NOR2_X1 i_0_17 (.A1(n_0_33), .A2(n_0_31), .ZN(n_0_10));
   MUX2_X1 i_0_18 (.A(n_0_13), .B(n_0_11), .S(in1[13]), .Z(n_7));
   MUX2_X1 i_0_19 (.A(n_0_12), .B(n_0_21), .S(n_0_33), .Z(n_0_11));
   MUX2_X1 i_0_20 (.A(in1[0]), .B(in1[2]), .S(n_0_32), .Z(n_0_12));
   MUX2_X1 i_0_21 (.A(n_0_15), .B(n_0_13), .S(in1[13]), .Z(n_8));
   MUX2_X1 i_0_22 (.A(n_0_14), .B(n_0_25), .S(n_0_33), .Z(n_0_13));
   MUX2_X1 i_0_23 (.A(in1[1]), .B(in1[3]), .S(n_0_32), .Z(n_0_14));
   MUX2_X1 i_0_24 (.A(n_0_17), .B(n_0_15), .S(in1[13]), .Z(n_9));
   MUX2_X1 i_0_25 (.A(n_0_16), .B(n_0_30), .S(n_0_33), .Z(n_0_15));
   MUX2_X1 i_0_26 (.A(in1[2]), .B(in1[4]), .S(n_0_32), .Z(n_0_16));
   MUX2_X1 i_0_27 (.A(n_0_20), .B(n_0_17), .S(in1[13]), .Z(n_10));
   MUX2_X1 i_0_28 (.A(n_0_18), .B(n_0_19), .S(n_0_33), .Z(n_0_17));
   MUX2_X1 i_0_29 (.A(in1[3]), .B(in1[5]), .S(n_0_32), .Z(n_0_18));
   MUX2_X1 i_0_30 (.A(in1[7]), .B(in1[9]), .S(n_0_32), .Z(n_0_19));
   MUX2_X1 i_0_31 (.A(n_0_24), .B(n_0_20), .S(in1[13]), .Z(n_11));
   MUX2_X1 i_0_32 (.A(n_0_21), .B(n_0_22), .S(n_0_33), .Z(n_0_20));
   MUX2_X1 i_0_33 (.A(in1[4]), .B(in1[6]), .S(n_0_32), .Z(n_0_21));
   MUX2_X1 i_0_34 (.A(in1[8]), .B(in1[10]), .S(n_0_32), .Z(n_0_22));
   OAI21_X1 i_0_35 (.A(n_0_23), .B1(n_0_27), .B2(in1[13]), .ZN(n_12));
   NAND2_X1 i_0_36 (.A1(in1[13]), .A2(n_0_24), .ZN(n_0_23));
   MUX2_X1 i_0_37 (.A(n_0_25), .B(n_0_26), .S(n_0_33), .Z(n_0_24));
   MUX2_X1 i_0_38 (.A(in1[5]), .B(in1[7]), .S(n_0_32), .Z(n_0_25));
   MUX2_X1 i_0_39 (.A(in1[9]), .B(in1[11]), .S(n_0_32), .Z(n_0_26));
   OAI21_X1 i_0_40 (.A(n_0_28), .B1(n_0_30), .B2(n_0_33), .ZN(n_0_27));
   OAI211_X1 i_0_41 (.A(n_0_33), .B(n_0_29), .C1(in1[14]), .C2(n_0_35), .ZN(
      n_0_28));
   NAND2_X1 i_0_42 (.A1(in1[10]), .A2(n_0_31), .ZN(n_0_29));
   MUX2_X1 i_0_43 (.A(in1[6]), .B(in1[8]), .S(n_0_32), .Z(n_0_30));
   INV_X1 i_0_44 (.A(n_0_32), .ZN(n_0_31));
   XNOR2_X1 i_0_45 (.A(in1[14]), .B(in1[13]), .ZN(n_0_32));
   XOR2_X1 i_0_46 (.A(in1[15]), .B(n_0_34), .Z(n_0_33));
   NOR3_X1 i_0_47 (.A1(in1[15]), .A2(in1[14]), .A3(in1[13]), .ZN(n_13));
   NOR2_X1 i_0_48 (.A1(in1[14]), .A2(in1[13]), .ZN(n_0_34));
   INV_X1 i_0_49 (.A(in1[12]), .ZN(n_0_35));
   INV_X1 i_0_50 (.A(in1[13]), .ZN(n_0_36));
   XNOR2_X1 i_1_0 (.A(tempIn11[1]), .B(out[0]), .ZN(out[1]));
   NOR2_X1 i_1_1 (.A1(n_1_10), .A2(n_1_0), .ZN(out[2]));
   AOI21_X1 i_1_2 (.A(tempIn11[2]), .B1(tempIn11[1]), .B2(tempIn11[0]), .ZN(
      n_1_0));
   XNOR2_X1 i_1_3 (.A(tempIn11[3]), .B(n_1_11), .ZN(out[3]));
   XOR2_X1 i_1_4 (.A(tempIn11[4]), .B(n_1_9), .Z(out[4]));
   NOR2_X1 i_1_5 (.A1(n_1_8), .A2(n_1_1), .ZN(out[5]));
   AOI21_X1 i_1_6 (.A(tempIn11[5]), .B1(tempIn11[4]), .B2(n_1_9), .ZN(n_1_1));
   XOR2_X1 i_1_7 (.A(tempIn11[6]), .B(n_1_8), .Z(out[6]));
   XNOR2_X1 i_1_8 (.A(tempIn11[7]), .B(n_1_2), .ZN(out[7]));
   NAND2_X1 i_1_9 (.A1(tempIn11[6]), .A2(n_1_8), .ZN(n_1_2));
   XOR2_X1 i_1_10 (.A(tempIn11[8]), .B(n_1_7), .Z(out[8]));
   XNOR2_X1 i_1_11 (.A(tempIn11[9]), .B(n_1_3), .ZN(out[9]));
   NAND2_X1 i_1_12 (.A1(tempIn11[8]), .A2(n_1_7), .ZN(n_1_3));
   XOR2_X1 i_1_13 (.A(tempIn11[10]), .B(n_1_6), .Z(out[10]));
   XNOR2_X1 i_1_14 (.A(tempIn11[11]), .B(n_1_4), .ZN(out[11]));
   NAND2_X1 i_1_15 (.A1(tempIn11[10]), .A2(n_1_6), .ZN(n_1_4));
   XNOR2_X1 i_1_16 (.A(tempIn11[12]), .B(n_1_5), .ZN(out[12]));
   NAND3_X1 i_1_17 (.A1(tempIn11[11]), .A2(tempIn11[10]), .A3(n_1_6), .ZN(n_1_5));
   AND3_X1 i_1_18 (.A1(tempIn11[9]), .A2(tempIn11[8]), .A3(n_1_7), .ZN(n_1_6));
   AND3_X1 i_1_19 (.A1(tempIn11[7]), .A2(tempIn11[6]), .A3(n_1_8), .ZN(n_1_7));
   AND3_X1 i_1_20 (.A1(tempIn11[5]), .A2(tempIn11[4]), .A3(n_1_9), .ZN(n_1_8));
   AND2_X1 i_1_21 (.A1(tempIn11[3]), .A2(n_1_10), .ZN(n_1_9));
   INV_X1 i_1_22 (.A(n_1_11), .ZN(n_1_10));
   NAND3_X1 i_1_23 (.A1(tempIn11[2]), .A2(tempIn11[1]), .A3(tempIn11[0]), 
      .ZN(n_1_11));
   INV_X1 i_1_24 (.A(tempIn11[0]), .ZN(out[0]));
endmodule

module datapath__0_1(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_0 (.A(B[0]), .B(p_0[0]), .CO(n_0), .S(p_1[0]));
   FA_X1 i_1 (.A(B[1]), .B(p_0[1]), .CI(n_0), .CO(n_1), .S(p_1[1]));
   FA_X1 i_2 (.A(B[2]), .B(p_0[2]), .CI(n_1), .CO(n_2), .S(p_1[2]));
   FA_X1 i_3 (.A(B[3]), .B(p_0[3]), .CI(n_2), .CO(n_3), .S(p_1[3]));
   FA_X1 i_4 (.A(B[4]), .B(p_0[4]), .CI(n_3), .CO(n_4), .S(p_1[4]));
   FA_X1 i_5 (.A(B[5]), .B(p_0[5]), .CI(n_4), .CO(n_5), .S(p_1[5]));
   FA_X1 i_6 (.A(B[6]), .B(p_0[6]), .CI(n_5), .CO(n_6), .S(p_1[6]));
   FA_X1 i_7 (.A(B[7]), .B(p_0[7]), .CI(n_6), .CO(n_7), .S(p_1[7]));
   FA_X1 i_8 (.A(B[8]), .B(p_0[8]), .CI(n_7), .CO(n_8), .S(p_1[8]));
   FA_X1 i_9 (.A(B[9]), .B(p_0[9]), .CI(n_8), .CO(n_9), .S(p_1[9]));
   FA_X1 i_10 (.A(B[10]), .B(p_0[10]), .CI(n_9), .CO(n_10), .S(p_1[10]));
   FA_X1 i_11 (.A(B[11]), .B(p_0[11]), .CI(n_10), .CO(n_11), .S(p_1[11]));
   FA_X1 i_12 (.A(B[15]), .B(p_0[12]), .CI(n_11), .CO(n_12), .S(p_1[12]));
   FA_X1 i_13 (.A(B[15]), .B(p_0[13]), .CI(n_12), .CO(n_13), .S(p_1[13]));
   FA_X1 i_14 (.A(B[15]), .B(p_0[14]), .CI(n_13), .CO(n_14), .S(p_1[14]));
   XNOR2_X1 i_15 (.A(B[15]), .B(p_0[15]), .ZN(n_15));
   XNOR2_X1 i_16 (.A(n_15), .B(n_14), .ZN(p_1[15]));
endmodule

module datapath__0_6(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[15]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[15]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[15]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[15]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_7(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[14]), .B1(p_0[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[15]), .B(n_15), .Z(p_2[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[14]), .A3(n_16), .B1(p_0[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[14]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[14]), .ZN(n_18));
endmodule

module datapath__0_12(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[15]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[15]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[15]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[15]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_13(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[14]), .B1(p_0[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[15]), .B(n_15), .Z(p_2[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[14]), .A3(n_16), .B1(p_0[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[14]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[14]), .ZN(n_18));
endmodule

module datapath__0_18(B, p_0, p_1);
   input [15:0]B;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(B[0]), .B(p_0[0]), .CO(n_1), .S(p_1[0]));
   FA_X1 i_2 (.A(B[1]), .B(p_0[1]), .CI(n_1), .CO(n_2), .S(p_1[1]));
   FA_X1 i_3 (.A(B[2]), .B(p_0[2]), .CI(n_2), .CO(n_3), .S(p_1[2]));
   FA_X1 i_4 (.A(B[3]), .B(p_0[3]), .CI(n_3), .CO(n_4), .S(p_1[3]));
   FA_X1 i_5 (.A(B[4]), .B(p_0[4]), .CI(n_4), .CO(n_5), .S(p_1[4]));
   FA_X1 i_6 (.A(B[5]), .B(p_0[5]), .CI(n_5), .CO(n_6), .S(p_1[5]));
   FA_X1 i_7 (.A(B[6]), .B(p_0[6]), .CI(n_6), .CO(n_7), .S(p_1[6]));
   FA_X1 i_8 (.A(B[7]), .B(p_0[7]), .CI(n_7), .CO(n_8), .S(p_1[7]));
   FA_X1 i_9 (.A(B[8]), .B(p_0[8]), .CI(n_8), .CO(n_9), .S(p_1[8]));
   FA_X1 i_10 (.A(B[9]), .B(p_0[9]), .CI(n_9), .CO(n_10), .S(p_1[9]));
   FA_X1 i_11 (.A(B[10]), .B(p_0[10]), .CI(n_10), .CO(n_11), .S(p_1[10]));
   FA_X1 i_12 (.A(B[11]), .B(p_0[11]), .CI(n_11), .CO(n_12), .S(p_1[11]));
   FA_X1 i_13 (.A(B[15]), .B(p_0[12]), .CI(n_12), .CO(n_13), .S(p_1[12]));
   FA_X1 i_14 (.A(B[15]), .B(p_0[13]), .CI(n_13), .CO(n_14), .S(p_1[13]));
   OAI21_X1 i_0 (.A(n_0), .B1(B[15]), .B2(n_15), .ZN(p_1[14]));
   OAI21_X1 i_15 (.A(n_0), .B1(n_16), .B2(n_14), .ZN(p_1[15]));
   NAND2_X1 i_16 (.A1(B[15]), .A2(n_15), .ZN(n_0));
   XNOR2_X1 i_17 (.A(p_0[14]), .B(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(p_0[14]), .ZN(n_16));
endmodule

module datapath__0_19(p_0, p_1, p_2);
   input [15:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   HA_X1 i_1 (.A(p_0[0]), .B(p_1[0]), .CO(n_1), .S(p_2[0]));
   FA_X1 i_2 (.A(p_0[1]), .B(p_1[1]), .CI(n_1), .CO(n_2), .S(p_2[1]));
   FA_X1 i_3 (.A(p_0[2]), .B(p_1[2]), .CI(n_2), .CO(n_3), .S(p_2[2]));
   FA_X1 i_4 (.A(p_0[3]), .B(p_1[3]), .CI(n_3), .CO(n_4), .S(p_2[3]));
   FA_X1 i_5 (.A(p_0[4]), .B(p_1[4]), .CI(n_4), .CO(n_5), .S(p_2[4]));
   FA_X1 i_6 (.A(p_0[5]), .B(p_1[5]), .CI(n_5), .CO(n_6), .S(p_2[5]));
   FA_X1 i_7 (.A(p_0[6]), .B(p_1[6]), .CI(n_6), .CO(n_7), .S(p_2[6]));
   FA_X1 i_8 (.A(p_0[7]), .B(p_1[7]), .CI(n_7), .CO(n_8), .S(p_2[7]));
   FA_X1 i_9 (.A(p_0[8]), .B(p_1[8]), .CI(n_8), .CO(n_9), .S(p_2[8]));
   FA_X1 i_10 (.A(p_0[9]), .B(p_1[9]), .CI(n_9), .CO(n_10), .S(p_2[9]));
   FA_X1 i_11 (.A(p_0[10]), .B(p_1[10]), .CI(n_10), .CO(n_11), .S(p_2[10]));
   FA_X1 i_12 (.A(p_0[11]), .B(p_1[11]), .CI(n_11), .CO(n_12), .S(p_2[11]));
   FA_X1 i_13 (.A(p_0[12]), .B(p_1[12]), .CI(n_12), .CO(n_13), .S(p_2[12]));
   FA_X1 i_14 (.A(p_0[13]), .B(p_1[13]), .CI(n_13), .CO(n_14), .S(p_2[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[14]), .B1(p_0[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[15]), .B(n_15), .Z(p_2[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[14]), .A3(n_16), .B1(p_0[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[14]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[14]), .ZN(n_18));
endmodule

module booth_16bit_multiplier__1(A, B, product);
   input [15:0]A;
   input [15:0]B;
   output [31:0]product;

   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_215;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_0;
   wire n_1_1;
   wire n_1_15;
   wire n_1_16;
   wire n_1_17;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;
   wire n_1_28;
   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire n_1_60;
   wire n_1_61;
   wire n_1_62;
   wire n_1_63;
   wire n_1_64;
   wire n_1_65;
   wire n_1_66;
   wire n_1_67;
   wire n_1_68;
   wire n_1_69;
   wire n_1_70;
   wire n_1_71;
   wire n_1_72;
   wire n_1_73;
   wire n_1_74;
   wire n_1_75;
   wire n_1_76;
   wire n_1_77;
   wire n_1_78;
   wire n_1_79;
   wire n_1_80;
   wire n_1_81;
   wire n_1_82;
   wire n_1_83;
   wire n_1_84;
   wire n_1_85;
   wire n_1_86;
   wire n_1_87;
   wire n_1_88;
   wire n_1_89;
   wire n_1_90;
   wire n_1_91;
   wire n_1_92;
   wire n_1_93;
   wire n_1_94;
   wire n_1_95;
   wire n_1_96;
   wire n_1_97;
   wire n_1_98;
   wire n_1_99;
   wire n_1_100;
   wire n_1_101;
   wire n_1_102;
   wire n_1_103;
   wire n_1_104;
   wire n_1_105;
   wire n_1_106;
   wire n_1_107;
   wire n_1_108;
   wire n_1_109;
   wire n_1_110;
   wire n_1_111;
   wire n_1_112;
   wire n_1_113;
   wire n_1_114;
   wire n_1_115;
   wire n_1_116;
   wire n_1_117;
   wire n_1_118;
   wire n_1_119;
   wire n_1_120;
   wire n_1_121;
   wire n_1_122;
   wire n_1_123;
   wire n_1_124;
   wire n_1_125;
   wire n_1_126;
   wire n_1_127;
   wire n_1_128;
   wire n_1_129;
   wire n_1_130;
   wire n_1_131;
   wire n_1_132;
   wire n_1_133;
   wire n_1_134;
   wire n_1_135;
   wire n_1_136;
   wire n_1_137;
   wire n_1_138;
   wire n_1_139;
   wire n_1_140;
   wire n_1_141;
   wire n_1_142;
   wire n_1_143;
   wire n_1_144;
   wire n_1_145;
   wire n_1_146;
   wire n_1_147;
   wire n_1_148;
   wire n_1_149;
   wire n_1_150;
   wire n_1_151;
   wire n_1_152;
   wire n_1_153;
   wire n_1_154;
   wire n_1_155;
   wire n_1_156;
   wire n_1_157;
   wire n_1_158;
   wire n_1_159;
   wire n_1_160;
   wire n_1_161;
   wire n_1_162;
   wire n_1_163;
   wire n_1_164;
   wire n_1_165;
   wire n_1_166;
   wire n_1_167;
   wire n_1_168;
   wire n_1_169;
   wire n_1_170;
   wire n_1_171;
   wire n_1_172;
   wire n_1_173;
   wire n_1_174;
   wire n_1_175;

   datapath__0_1 i_2 (.B({B[15], uc_0, uc_1, uc_2, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({n_249, n_264, 
      n_263, n_262, n_261, n_260, n_259, n_258, n_257, n_256, n_255, n_254, 
      n_253, n_252, n_251, n_250}), .p_1({n_15, n_14, n_13, n_12, n_11, n_10, 
      n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0}));
   datapath__0_6 i_5 (.B({B[15], uc_3, uc_4, uc_5, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_6, n_248, n_247, 
      n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, n_238, n_237, 
      n_236, n_235, n_234}), .p_1({n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
      n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16}));
   datapath__0_7 i_6 (.p_0({n_264, n_263, n_262, n_261, n_260, n_259, n_258, 
      n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, B[0]}), .p_1({uc_7, 
      n_248, n_247, n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, 
      n_238, n_237, n_236, n_235, n_234}), .p_2({n_47, n_46, n_45, n_44, n_43, 
      n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32}));
   datapath__0_12 i_9 (.B({B[15], uc_8, uc_9, uc_10, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_11, n_233, 
      n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, 
      n_222, n_221, n_220, n_219}), .p_1({n_63, n_62, n_61, n_60, n_59, n_58, 
      n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48}));
   datapath__0_13 i_10 (.p_0({n_264, n_263, n_262, n_261, n_260, n_259, n_258, 
      n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, B[0]}), .p_1({
      uc_12, n_233, n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, 
      n_224, n_223, n_222, n_221, n_220, n_219}), .p_2({n_79, n_78, n_77, n_76, 
      n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64}));
   datapath__0_18 i_13 (.B({B[15], uc_13, uc_14, uc_15, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_16, n_218, 
      n_217, n_216, n_215, n_214, n_213, n_212, n_211, n_210, n_209, n_208, 
      n_207, n_206, n_205, n_204}), .p_1({n_95, n_94, n_93, n_92, n_91, n_90, 
      n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80}));
   datapath__0_19 i_14 (.p_0({n_264, n_263, n_262, n_261, n_260, n_259, n_258, 
      n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, B[0]}), .p_1({
      uc_17, n_218, n_217, n_216, n_215, n_214, n_213, n_212, n_211, n_210, 
      n_209, n_208, n_207, n_206, n_205, n_204}), .p_2({n_111, n_110, n_109, 
      n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
      n_97, n_96}));
   INV_X1 i_0_108 (.A(n_0_60), .ZN(product[12]));
   AOI222_X1 i_0_109 (.A1(n_438), .A2(n_0_79), .B1(n_438), .B2(n_0_78), .C1(
      n_112), .C2(n_0_77), .ZN(n_0_60));
   INV_X1 i_0_110 (.A(n_0_61), .ZN(product[13]));
   AOI222_X1 i_0_111 (.A1(n_424), .A2(n_0_79), .B1(n_417), .B2(n_0_78), .C1(
      n_113), .C2(n_0_77), .ZN(n_0_61));
   INV_X1 i_0_112 (.A(n_0_62), .ZN(product[14]));
   AOI222_X1 i_0_113 (.A1(n_425), .A2(n_0_79), .B1(n_418), .B2(n_0_78), .C1(
      n_114), .C2(n_0_77), .ZN(n_0_62));
   INV_X1 i_0_114 (.A(n_0_63), .ZN(product[15]));
   AOI222_X1 i_0_115 (.A1(n_426), .A2(n_0_79), .B1(n_419), .B2(n_0_78), .C1(
      n_115), .C2(n_0_77), .ZN(n_0_63));
   INV_X1 i_0_116 (.A(n_0_64), .ZN(product[16]));
   AOI222_X1 i_0_117 (.A1(n_427), .A2(n_0_79), .B1(n_420), .B2(n_0_78), .C1(
      n_116), .C2(n_0_77), .ZN(n_0_64));
   INV_X1 i_0_118 (.A(n_0_65), .ZN(product[17]));
   AOI222_X1 i_0_119 (.A1(n_428), .A2(n_0_79), .B1(n_421), .B2(n_0_78), .C1(
      n_117), .C2(n_0_77), .ZN(n_0_65));
   INV_X1 i_0_120 (.A(n_0_66), .ZN(product[18]));
   AOI222_X1 i_0_121 (.A1(n_429), .A2(n_0_79), .B1(n_422), .B2(n_0_78), .C1(
      n_118), .C2(n_0_77), .ZN(n_0_66));
   INV_X1 i_0_122 (.A(n_0_67), .ZN(product[19]));
   AOI222_X1 i_0_123 (.A1(n_430), .A2(n_0_79), .B1(n_423), .B2(n_0_78), .C1(
      n_119), .C2(n_0_77), .ZN(n_0_67));
   NOR2_X1 i_0_141 (.A1(n_0_79), .A2(n_0_78), .ZN(n_0_77));
   NOR2_X1 i_0_142 (.A1(A[15]), .A2(n_0_196), .ZN(n_0_78));
   NOR2_X1 i_0_143 (.A1(n_0_215), .A2(A[11]), .ZN(n_0_79));
   INV_X1 i_0_144 (.A(n_0_80), .ZN(product[11]));
   AOI222_X1 i_0_145 (.A1(n_437), .A2(n_0_98), .B1(n_437), .B2(n_0_99), .C1(
      n_120), .C2(n_0_97), .ZN(n_0_80));
   INV_X1 i_0_146 (.A(n_0_81), .ZN(n_112));
   AOI222_X1 i_0_147 (.A1(n_409), .A2(n_0_99), .B1(n_401), .B2(n_0_98), .C1(
      n_121), .C2(n_0_97), .ZN(n_0_81));
   INV_X1 i_0_148 (.A(n_0_82), .ZN(n_113));
   AOI222_X1 i_0_149 (.A1(n_410), .A2(n_0_99), .B1(n_402), .B2(n_0_98), .C1(
      n_122), .C2(n_0_97), .ZN(n_0_82));
   INV_X1 i_0_150 (.A(n_0_83), .ZN(n_114));
   AOI222_X1 i_0_151 (.A1(n_411), .A2(n_0_99), .B1(n_403), .B2(n_0_98), .C1(
      n_123), .C2(n_0_97), .ZN(n_0_83));
   INV_X1 i_0_152 (.A(n_0_84), .ZN(n_115));
   AOI222_X1 i_0_153 (.A1(n_412), .A2(n_0_99), .B1(n_404), .B2(n_0_98), .C1(
      n_124), .C2(n_0_97), .ZN(n_0_84));
   INV_X1 i_0_154 (.A(n_0_85), .ZN(n_116));
   AOI222_X1 i_0_155 (.A1(n_413), .A2(n_0_99), .B1(n_405), .B2(n_0_98), .C1(
      n_125), .C2(n_0_97), .ZN(n_0_85));
   INV_X1 i_0_156 (.A(n_0_86), .ZN(n_117));
   AOI222_X1 i_0_157 (.A1(n_414), .A2(n_0_99), .B1(n_406), .B2(n_0_98), .C1(
      n_126), .C2(n_0_97), .ZN(n_0_86));
   INV_X1 i_0_158 (.A(n_0_87), .ZN(n_118));
   AOI222_X1 i_0_159 (.A1(n_415), .A2(n_0_99), .B1(n_407), .B2(n_0_98), .C1(
      n_127), .C2(n_0_97), .ZN(n_0_87));
   INV_X1 i_0_160 (.A(n_0_88), .ZN(n_119));
   AOI222_X1 i_0_161 (.A1(n_416), .A2(n_0_99), .B1(n_408), .B2(n_0_98), .C1(
      n_128), .C2(n_0_97), .ZN(n_0_88));
   NOR2_X1 i_0_177 (.A1(n_0_99), .A2(n_0_98), .ZN(n_0_97));
   NOR2_X1 i_0_178 (.A1(A[11]), .A2(n_0_195), .ZN(n_0_98));
   NOR2_X1 i_0_179 (.A1(n_0_196), .A2(A[10]), .ZN(n_0_99));
   INV_X1 i_0_180 (.A(n_0_100), .ZN(product[10]));
   AOI222_X1 i_0_181 (.A1(n_436), .A2(n_0_118), .B1(n_436), .B2(n_0_119), 
      .C1(n_129), .C2(n_0_117), .ZN(n_0_100));
   INV_X1 i_0_182 (.A(n_0_101), .ZN(n_120));
   AOI222_X1 i_0_183 (.A1(n_383), .A2(n_0_118), .B1(n_392), .B2(n_0_119), 
      .C1(n_130), .C2(n_0_117), .ZN(n_0_101));
   INV_X1 i_0_184 (.A(n_0_102), .ZN(n_121));
   AOI222_X1 i_0_185 (.A1(n_384), .A2(n_0_118), .B1(n_393), .B2(n_0_119), 
      .C1(n_131), .C2(n_0_117), .ZN(n_0_102));
   INV_X1 i_0_186 (.A(n_0_103), .ZN(n_122));
   AOI222_X1 i_0_187 (.A1(n_394), .A2(n_0_119), .B1(n_385), .B2(n_0_118), 
      .C1(n_132), .C2(n_0_117), .ZN(n_0_103));
   INV_X1 i_0_188 (.A(n_0_104), .ZN(n_123));
   AOI222_X1 i_0_189 (.A1(n_395), .A2(n_0_119), .B1(n_386), .B2(n_0_118), 
      .C1(n_133), .C2(n_0_117), .ZN(n_0_104));
   INV_X1 i_0_190 (.A(n_0_105), .ZN(n_124));
   AOI222_X1 i_0_191 (.A1(n_396), .A2(n_0_119), .B1(n_387), .B2(n_0_118), 
      .C1(n_134), .C2(n_0_117), .ZN(n_0_105));
   INV_X1 i_0_192 (.A(n_0_106), .ZN(n_125));
   AOI222_X1 i_0_193 (.A1(n_397), .A2(n_0_119), .B1(n_388), .B2(n_0_118), 
      .C1(n_135), .C2(n_0_117), .ZN(n_0_106));
   INV_X1 i_0_194 (.A(n_0_107), .ZN(n_126));
   AOI222_X1 i_0_195 (.A1(n_398), .A2(n_0_119), .B1(n_389), .B2(n_0_118), 
      .C1(n_136), .C2(n_0_117), .ZN(n_0_107));
   INV_X1 i_0_196 (.A(n_0_108), .ZN(n_127));
   AOI222_X1 i_0_197 (.A1(n_399), .A2(n_0_119), .B1(n_390), .B2(n_0_118), 
      .C1(n_137), .C2(n_0_117), .ZN(n_0_108));
   INV_X1 i_0_198 (.A(n_0_109), .ZN(n_128));
   AOI222_X1 i_0_199 (.A1(n_400), .A2(n_0_119), .B1(n_391), .B2(n_0_118), 
      .C1(n_138), .C2(n_0_117), .ZN(n_0_109));
   NOR2_X1 i_0_213 (.A1(n_0_119), .A2(n_0_118), .ZN(n_0_117));
   NOR2_X1 i_0_214 (.A1(A[10]), .A2(n_0_194), .ZN(n_0_118));
   NOR2_X1 i_0_215 (.A1(n_0_195), .A2(A[9]), .ZN(n_0_119));
   INV_X1 i_0_216 (.A(n_0_120), .ZN(product[9]));
   AOI222_X1 i_0_217 (.A1(n_435), .A2(n_0_138), .B1(n_435), .B2(n_0_139), 
      .C1(n_139), .C2(n_0_137), .ZN(n_0_120));
   INV_X1 i_0_218 (.A(n_0_121), .ZN(n_129));
   AOI222_X1 i_0_219 (.A1(n_363), .A2(n_0_138), .B1(n_373), .B2(n_0_139), 
      .C1(n_140), .C2(n_0_137), .ZN(n_0_121));
   INV_X1 i_0_220 (.A(n_0_122), .ZN(n_130));
   AOI222_X1 i_0_221 (.A1(n_364), .A2(n_0_138), .B1(n_374), .B2(n_0_139), 
      .C1(n_141), .C2(n_0_137), .ZN(n_0_122));
   INV_X1 i_0_222 (.A(n_0_123), .ZN(n_131));
   AOI222_X1 i_0_223 (.A1(n_365), .A2(n_0_138), .B1(n_375), .B2(n_0_139), 
      .C1(n_142), .C2(n_0_137), .ZN(n_0_123));
   INV_X1 i_0_224 (.A(n_0_124), .ZN(n_132));
   AOI222_X1 i_0_225 (.A1(n_376), .A2(n_0_139), .B1(n_366), .B2(n_0_138), 
      .C1(n_143), .C2(n_0_137), .ZN(n_0_124));
   INV_X1 i_0_226 (.A(n_0_125), .ZN(n_133));
   AOI222_X1 i_0_227 (.A1(n_377), .A2(n_0_139), .B1(n_367), .B2(n_0_138), 
      .C1(n_144), .C2(n_0_137), .ZN(n_0_125));
   INV_X1 i_0_228 (.A(n_0_126), .ZN(n_134));
   AOI222_X1 i_0_229 (.A1(n_378), .A2(n_0_139), .B1(n_368), .B2(n_0_138), 
      .C1(n_145), .C2(n_0_137), .ZN(n_0_126));
   INV_X1 i_0_230 (.A(n_0_127), .ZN(n_135));
   AOI222_X1 i_0_231 (.A1(n_379), .A2(n_0_139), .B1(n_369), .B2(n_0_138), 
      .C1(n_146), .C2(n_0_137), .ZN(n_0_127));
   INV_X1 i_0_232 (.A(n_0_128), .ZN(n_136));
   AOI222_X1 i_0_233 (.A1(n_380), .A2(n_0_139), .B1(n_370), .B2(n_0_138), 
      .C1(n_147), .C2(n_0_137), .ZN(n_0_128));
   INV_X1 i_0_234 (.A(n_0_129), .ZN(n_137));
   AOI222_X1 i_0_235 (.A1(n_381), .A2(n_0_139), .B1(n_371), .B2(n_0_138), 
      .C1(n_148), .C2(n_0_137), .ZN(n_0_129));
   INV_X1 i_0_236 (.A(n_0_130), .ZN(n_138));
   AOI222_X1 i_0_237 (.A1(n_382), .A2(n_0_139), .B1(n_372), .B2(n_0_138), 
      .C1(n_149), .C2(n_0_137), .ZN(n_0_130));
   NOR2_X1 i_0_249 (.A1(n_0_139), .A2(n_0_138), .ZN(n_0_137));
   NOR2_X1 i_0_250 (.A1(A[9]), .A2(n_0_176), .ZN(n_0_138));
   NOR2_X1 i_0_251 (.A1(n_0_194), .A2(A[8]), .ZN(n_0_139));
   INV_X1 i_0_252 (.A(n_0_140), .ZN(product[8]));
   AOI222_X1 i_0_253 (.A1(n_434), .A2(n_0_158), .B1(n_434), .B2(n_0_159), 
      .C1(n_150), .C2(n_0_157), .ZN(n_0_140));
   INV_X1 i_0_254 (.A(n_0_141), .ZN(n_139));
   AOI222_X1 i_0_255 (.A1(n_341), .A2(n_0_158), .B1(n_352), .B2(n_0_159), 
      .C1(n_151), .C2(n_0_157), .ZN(n_0_141));
   INV_X1 i_0_256 (.A(n_0_142), .ZN(n_140));
   AOI222_X1 i_0_257 (.A1(n_342), .A2(n_0_158), .B1(n_353), .B2(n_0_159), 
      .C1(n_152), .C2(n_0_157), .ZN(n_0_142));
   INV_X1 i_0_258 (.A(n_0_143), .ZN(n_141));
   AOI222_X1 i_0_259 (.A1(n_343), .A2(n_0_158), .B1(n_354), .B2(n_0_159), 
      .C1(n_153), .C2(n_0_157), .ZN(n_0_143));
   INV_X1 i_0_260 (.A(n_0_144), .ZN(n_142));
   AOI222_X1 i_0_261 (.A1(n_344), .A2(n_0_158), .B1(n_355), .B2(n_0_159), 
      .C1(n_154), .C2(n_0_157), .ZN(n_0_144));
   INV_X1 i_0_262 (.A(n_0_145), .ZN(n_143));
   AOI222_X1 i_0_263 (.A1(n_356), .A2(n_0_159), .B1(n_345), .B2(n_0_158), 
      .C1(n_155), .C2(n_0_157), .ZN(n_0_145));
   INV_X1 i_0_264 (.A(n_0_146), .ZN(n_144));
   AOI222_X1 i_0_265 (.A1(n_357), .A2(n_0_159), .B1(n_346), .B2(n_0_158), 
      .C1(n_156), .C2(n_0_157), .ZN(n_0_146));
   INV_X1 i_0_266 (.A(n_0_147), .ZN(n_145));
   AOI222_X1 i_0_267 (.A1(n_358), .A2(n_0_159), .B1(n_347), .B2(n_0_158), 
      .C1(n_157), .C2(n_0_157), .ZN(n_0_147));
   INV_X1 i_0_268 (.A(n_0_148), .ZN(n_146));
   AOI222_X1 i_0_269 (.A1(n_359), .A2(n_0_159), .B1(n_348), .B2(n_0_158), 
      .C1(n_158), .C2(n_0_157), .ZN(n_0_148));
   INV_X1 i_0_270 (.A(n_0_149), .ZN(n_147));
   AOI222_X1 i_0_271 (.A1(n_360), .A2(n_0_159), .B1(n_349), .B2(n_0_158), 
      .C1(n_159), .C2(n_0_157), .ZN(n_0_149));
   INV_X1 i_0_272 (.A(n_0_150), .ZN(n_148));
   AOI222_X1 i_0_273 (.A1(n_361), .A2(n_0_159), .B1(n_350), .B2(n_0_158), 
      .C1(n_160), .C2(n_0_157), .ZN(n_0_150));
   INV_X1 i_0_274 (.A(n_0_151), .ZN(n_149));
   AOI222_X1 i_0_275 (.A1(n_362), .A2(n_0_159), .B1(n_351), .B2(n_0_158), 
      .C1(n_161), .C2(n_0_157), .ZN(n_0_151));
   NOR2_X1 i_0_285 (.A1(n_0_159), .A2(n_0_158), .ZN(n_0_157));
   NOR2_X1 i_0_286 (.A1(A[8]), .A2(n_0_175), .ZN(n_0_158));
   NOR2_X1 i_0_287 (.A1(n_0_176), .A2(A[7]), .ZN(n_0_159));
   INV_X1 i_0_288 (.A(n_0_160), .ZN(product[7]));
   AOI222_X1 i_0_289 (.A1(n_433), .A2(n_0_178), .B1(n_433), .B2(n_0_179), 
      .C1(n_162), .C2(n_0_177), .ZN(n_0_160));
   INV_X1 i_0_290 (.A(n_0_161), .ZN(n_150));
   AOI222_X1 i_0_291 (.A1(n_317), .A2(n_0_178), .B1(n_329), .B2(n_0_179), 
      .C1(n_163), .C2(n_0_177), .ZN(n_0_161));
   INV_X1 i_0_292 (.A(n_0_162), .ZN(n_151));
   AOI222_X1 i_0_293 (.A1(n_318), .A2(n_0_178), .B1(n_330), .B2(n_0_179), 
      .C1(n_164), .C2(n_0_177), .ZN(n_0_162));
   INV_X1 i_0_294 (.A(n_0_163), .ZN(n_152));
   AOI222_X1 i_0_295 (.A1(n_319), .A2(n_0_178), .B1(n_331), .B2(n_0_179), 
      .C1(n_165), .C2(n_0_177), .ZN(n_0_163));
   INV_X1 i_0_296 (.A(n_0_164), .ZN(n_153));
   AOI222_X1 i_0_297 (.A1(n_320), .A2(n_0_178), .B1(n_332), .B2(n_0_179), 
      .C1(n_166), .C2(n_0_177), .ZN(n_0_164));
   INV_X1 i_0_298 (.A(n_0_165), .ZN(n_154));
   AOI222_X1 i_0_299 (.A1(n_321), .A2(n_0_178), .B1(n_333), .B2(n_0_179), 
      .C1(n_167), .C2(n_0_177), .ZN(n_0_165));
   INV_X1 i_0_300 (.A(n_0_166), .ZN(n_155));
   AOI222_X1 i_0_301 (.A1(n_322), .A2(n_0_178), .B1(n_334), .B2(n_0_179), 
      .C1(n_168), .C2(n_0_177), .ZN(n_0_166));
   INV_X1 i_0_302 (.A(n_0_167), .ZN(n_156));
   AOI222_X1 i_0_303 (.A1(n_335), .A2(n_0_179), .B1(n_323), .B2(n_0_178), 
      .C1(n_169), .C2(n_0_177), .ZN(n_0_167));
   INV_X1 i_0_304 (.A(n_0_168), .ZN(n_157));
   AOI222_X1 i_0_305 (.A1(n_336), .A2(n_0_179), .B1(n_324), .B2(n_0_178), 
      .C1(n_170), .C2(n_0_177), .ZN(n_0_168));
   INV_X1 i_0_306 (.A(n_0_169), .ZN(n_158));
   AOI222_X1 i_0_307 (.A1(n_337), .A2(n_0_179), .B1(n_325), .B2(n_0_178), 
      .C1(n_171), .C2(n_0_177), .ZN(n_0_169));
   INV_X1 i_0_308 (.A(n_0_170), .ZN(n_159));
   AOI222_X1 i_0_309 (.A1(n_338), .A2(n_0_179), .B1(n_326), .B2(n_0_178), 
      .C1(n_172), .C2(n_0_177), .ZN(n_0_170));
   INV_X1 i_0_310 (.A(n_0_171), .ZN(n_160));
   AOI222_X1 i_0_311 (.A1(n_339), .A2(n_0_179), .B1(n_327), .B2(n_0_178), 
      .C1(n_173), .C2(n_0_177), .ZN(n_0_171));
   INV_X1 i_0_312 (.A(n_0_172), .ZN(n_161));
   AOI222_X1 i_0_313 (.A1(n_340), .A2(n_0_179), .B1(n_328), .B2(n_0_178), 
      .C1(n_174), .C2(n_0_177), .ZN(n_0_172));
   NOR2_X1 i_0_321 (.A1(n_0_179), .A2(n_0_178), .ZN(n_0_177));
   NOR2_X1 i_0_322 (.A1(A[7]), .A2(n_0_174), .ZN(n_0_178));
   NOR2_X1 i_0_323 (.A1(n_0_175), .A2(A[6]), .ZN(n_0_179));
   INV_X1 i_0_324 (.A(n_0_180), .ZN(product[6]));
   AOI222_X1 i_0_325 (.A1(n_432), .A2(n_0_198), .B1(n_432), .B2(n_0_199), 
      .C1(n_175), .C2(n_0_197), .ZN(n_0_180));
   INV_X1 i_0_326 (.A(n_0_181), .ZN(n_162));
   AOI222_X1 i_0_327 (.A1(n_291), .A2(n_0_198), .B1(n_304), .B2(n_0_199), 
      .C1(n_176), .C2(n_0_197), .ZN(n_0_181));
   INV_X1 i_0_328 (.A(n_0_182), .ZN(n_163));
   AOI222_X1 i_0_329 (.A1(n_292), .A2(n_0_198), .B1(n_305), .B2(n_0_199), 
      .C1(n_177), .C2(n_0_197), .ZN(n_0_182));
   INV_X1 i_0_330 (.A(n_0_183), .ZN(n_164));
   AOI222_X1 i_0_331 (.A1(n_293), .A2(n_0_198), .B1(n_306), .B2(n_0_199), 
      .C1(n_178), .C2(n_0_197), .ZN(n_0_183));
   INV_X1 i_0_332 (.A(n_0_184), .ZN(n_165));
   AOI222_X1 i_0_333 (.A1(n_294), .A2(n_0_198), .B1(n_307), .B2(n_0_199), 
      .C1(n_179), .C2(n_0_197), .ZN(n_0_184));
   INV_X1 i_0_334 (.A(n_0_185), .ZN(n_166));
   AOI222_X1 i_0_335 (.A1(n_295), .A2(n_0_198), .B1(n_308), .B2(n_0_199), 
      .C1(n_180), .C2(n_0_197), .ZN(n_0_185));
   INV_X1 i_0_336 (.A(n_0_186), .ZN(n_167));
   AOI222_X1 i_0_337 (.A1(n_296), .A2(n_0_198), .B1(n_309), .B2(n_0_199), 
      .C1(n_181), .C2(n_0_197), .ZN(n_0_186));
   INV_X1 i_0_338 (.A(n_0_187), .ZN(n_168));
   AOI222_X1 i_0_339 (.A1(n_297), .A2(n_0_198), .B1(n_310), .B2(n_0_199), 
      .C1(n_182), .C2(n_0_197), .ZN(n_0_187));
   INV_X1 i_0_340 (.A(n_0_188), .ZN(n_169));
   AOI222_X1 i_0_341 (.A1(n_311), .A2(n_0_199), .B1(n_298), .B2(n_0_198), 
      .C1(n_183), .C2(n_0_197), .ZN(n_0_188));
   INV_X1 i_0_342 (.A(n_0_189), .ZN(n_170));
   AOI222_X1 i_0_343 (.A1(n_312), .A2(n_0_199), .B1(n_299), .B2(n_0_198), 
      .C1(n_184), .C2(n_0_197), .ZN(n_0_189));
   INV_X1 i_0_344 (.A(n_0_190), .ZN(n_171));
   AOI222_X1 i_0_345 (.A1(n_313), .A2(n_0_199), .B1(n_300), .B2(n_0_198), 
      .C1(n_185), .C2(n_0_197), .ZN(n_0_190));
   INV_X1 i_0_346 (.A(n_0_191), .ZN(n_172));
   AOI222_X1 i_0_347 (.A1(n_314), .A2(n_0_199), .B1(n_301), .B2(n_0_198), 
      .C1(n_186), .C2(n_0_197), .ZN(n_0_191));
   INV_X1 i_0_348 (.A(n_0_192), .ZN(n_173));
   AOI222_X1 i_0_349 (.A1(n_315), .A2(n_0_199), .B1(n_302), .B2(n_0_198), 
      .C1(n_187), .C2(n_0_197), .ZN(n_0_192));
   INV_X1 i_0_350 (.A(n_0_193), .ZN(n_174));
   AOI222_X1 i_0_351 (.A1(n_316), .A2(n_0_199), .B1(n_303), .B2(n_0_198), 
      .C1(n_188), .C2(n_0_197), .ZN(n_0_193));
   NOR2_X1 i_0_357 (.A1(n_0_199), .A2(n_0_198), .ZN(n_0_197));
   NOR2_X1 i_0_358 (.A1(A[6]), .A2(n_0_173), .ZN(n_0_198));
   NOR2_X1 i_0_359 (.A1(n_0_174), .A2(A[5]), .ZN(n_0_199));
   INV_X1 i_0_360 (.A(n_0_200), .ZN(product[5]));
   AOI222_X1 i_0_361 (.A1(n_431), .A2(n_0_218), .B1(n_431), .B2(n_0_219), 
      .C1(n_189), .C2(n_0_217), .ZN(n_0_200));
   INV_X1 i_0_362 (.A(n_0_201), .ZN(n_175));
   AOI222_X1 i_0_363 (.A1(n_265), .A2(n_0_218), .B1(n_278), .B2(n_0_219), 
      .C1(n_190), .C2(n_0_217), .ZN(n_0_201));
   INV_X1 i_0_364 (.A(n_0_202), .ZN(n_176));
   AOI222_X1 i_0_365 (.A1(n_266), .A2(n_0_218), .B1(n_279), .B2(n_0_219), 
      .C1(n_191), .C2(n_0_217), .ZN(n_0_202));
   INV_X1 i_0_366 (.A(n_0_203), .ZN(n_177));
   AOI222_X1 i_0_367 (.A1(n_267), .A2(n_0_218), .B1(n_280), .B2(n_0_219), 
      .C1(n_192), .C2(n_0_217), .ZN(n_0_203));
   INV_X1 i_0_368 (.A(n_0_204), .ZN(n_178));
   AOI222_X1 i_0_369 (.A1(n_268), .A2(n_0_218), .B1(n_281), .B2(n_0_219), 
      .C1(n_193), .C2(n_0_217), .ZN(n_0_204));
   INV_X1 i_0_370 (.A(n_0_205), .ZN(n_179));
   AOI222_X1 i_0_371 (.A1(n_269), .A2(n_0_218), .B1(n_282), .B2(n_0_219), 
      .C1(n_194), .C2(n_0_217), .ZN(n_0_205));
   INV_X1 i_0_372 (.A(n_0_206), .ZN(n_180));
   AOI222_X1 i_0_373 (.A1(n_270), .A2(n_0_218), .B1(n_283), .B2(n_0_219), 
      .C1(n_195), .C2(n_0_217), .ZN(n_0_206));
   INV_X1 i_0_374 (.A(n_0_207), .ZN(n_181));
   AOI222_X1 i_0_375 (.A1(n_271), .A2(n_0_218), .B1(n_284), .B2(n_0_219), 
      .C1(n_196), .C2(n_0_217), .ZN(n_0_207));
   INV_X1 i_0_376 (.A(n_0_208), .ZN(n_182));
   AOI222_X1 i_0_377 (.A1(n_272), .A2(n_0_218), .B1(n_285), .B2(n_0_219), 
      .C1(n_197), .C2(n_0_217), .ZN(n_0_208));
   INV_X1 i_0_378 (.A(n_0_209), .ZN(n_183));
   AOI222_X1 i_0_379 (.A1(n_286), .A2(n_0_219), .B1(n_273), .B2(n_0_218), 
      .C1(n_198), .C2(n_0_217), .ZN(n_0_209));
   INV_X1 i_0_380 (.A(n_0_210), .ZN(n_184));
   AOI222_X1 i_0_381 (.A1(n_287), .A2(n_0_219), .B1(n_274), .B2(n_0_218), 
      .C1(n_199), .C2(n_0_217), .ZN(n_0_210));
   INV_X1 i_0_382 (.A(n_0_211), .ZN(n_185));
   AOI222_X1 i_0_383 (.A1(n_288), .A2(n_0_219), .B1(n_275), .B2(n_0_218), 
      .C1(n_200), .C2(n_0_217), .ZN(n_0_211));
   INV_X1 i_0_384 (.A(n_0_212), .ZN(n_186));
   AOI222_X1 i_0_385 (.A1(n_289), .A2(n_0_219), .B1(n_276), .B2(n_0_218), 
      .C1(n_201), .C2(n_0_217), .ZN(n_0_212));
   INV_X1 i_0_386 (.A(n_0_213), .ZN(n_187));
   AOI222_X1 i_0_387 (.A1(n_290), .A2(n_0_219), .B1(n_277), .B2(n_0_218), 
      .C1(n_202), .C2(n_0_217), .ZN(n_0_213));
   INV_X1 i_0_388 (.A(n_0_214), .ZN(n_188));
   AOI221_X1 i_0_389 (.A(n_0_216), .B1(n_440), .B2(n_0_218), .C1(n_439), 
      .C2(n_0_219), .ZN(n_0_214));
   AND2_X1 i_0_392 (.A1(n_203), .A2(n_0_217), .ZN(n_0_216));
   NOR2_X1 i_0_393 (.A1(n_0_219), .A2(n_0_218), .ZN(n_0_217));
   NOR2_X1 i_0_394 (.A1(A[5]), .A2(n_0_156), .ZN(n_0_218));
   NOR2_X1 i_0_395 (.A1(n_0_173), .A2(A[4]), .ZN(n_0_219));
   INV_X1 i_0_396 (.A(n_0_220), .ZN(product[4]));
   AOI222_X1 i_0_397 (.A1(n_80), .A2(n_0_2), .B1(n_96), .B2(n_0_3), .C1(n_204), 
      .C2(n_0_1), .ZN(n_0_220));
   INV_X1 i_0_398 (.A(n_0_221), .ZN(n_189));
   AOI222_X1 i_0_399 (.A1(n_81), .A2(n_0_2), .B1(n_97), .B2(n_0_3), .C1(n_205), 
      .C2(n_0_1), .ZN(n_0_221));
   INV_X1 i_0_400 (.A(n_0_222), .ZN(n_190));
   AOI222_X1 i_0_401 (.A1(n_82), .A2(n_0_2), .B1(n_98), .B2(n_0_3), .C1(n_206), 
      .C2(n_0_1), .ZN(n_0_222));
   INV_X1 i_0_402 (.A(n_0_223), .ZN(n_191));
   AOI222_X1 i_0_403 (.A1(n_83), .A2(n_0_2), .B1(n_99), .B2(n_0_3), .C1(n_207), 
      .C2(n_0_1), .ZN(n_0_223));
   INV_X1 i_0_404 (.A(n_0_224), .ZN(n_192));
   AOI222_X1 i_0_405 (.A1(n_84), .A2(n_0_2), .B1(n_100), .B2(n_0_3), .C1(n_208), 
      .C2(n_0_1), .ZN(n_0_224));
   INV_X1 i_0_406 (.A(n_0_225), .ZN(n_193));
   AOI222_X1 i_0_407 (.A1(n_85), .A2(n_0_2), .B1(n_101), .B2(n_0_3), .C1(n_209), 
      .C2(n_0_1), .ZN(n_0_225));
   INV_X1 i_0_408 (.A(n_0_226), .ZN(n_194));
   AOI222_X1 i_0_409 (.A1(n_86), .A2(n_0_2), .B1(n_102), .B2(n_0_3), .C1(n_210), 
      .C2(n_0_1), .ZN(n_0_226));
   INV_X1 i_0_410 (.A(n_0_227), .ZN(n_195));
   AOI222_X1 i_0_411 (.A1(n_87), .A2(n_0_2), .B1(n_103), .B2(n_0_3), .C1(n_211), 
      .C2(n_0_1), .ZN(n_0_227));
   INV_X1 i_0_412 (.A(n_0_228), .ZN(n_196));
   AOI222_X1 i_0_413 (.A1(n_88), .A2(n_0_2), .B1(n_104), .B2(n_0_3), .C1(n_212), 
      .C2(n_0_1), .ZN(n_0_228));
   INV_X1 i_0_414 (.A(n_0_229), .ZN(n_197));
   AOI222_X1 i_0_415 (.A1(n_89), .A2(n_0_2), .B1(n_105), .B2(n_0_3), .C1(n_213), 
      .C2(n_0_1), .ZN(n_0_229));
   INV_X1 i_0_416 (.A(n_0_230), .ZN(n_198));
   AOI222_X1 i_0_417 (.A1(n_90), .A2(n_0_2), .B1(n_106), .B2(n_0_3), .C1(n_214), 
      .C2(n_0_1), .ZN(n_0_230));
   INV_X1 i_0_418 (.A(n_0_231), .ZN(n_199));
   AOI222_X1 i_0_419 (.A1(n_107), .A2(n_0_3), .B1(n_91), .B2(n_0_2), .C1(n_215), 
      .C2(n_0_1), .ZN(n_0_231));
   INV_X1 i_0_420 (.A(n_0_232), .ZN(n_200));
   AOI222_X1 i_0_421 (.A1(n_108), .A2(n_0_3), .B1(n_92), .B2(n_0_2), .C1(n_216), 
      .C2(n_0_1), .ZN(n_0_232));
   INV_X1 i_0_422 (.A(n_0_233), .ZN(n_201));
   AOI222_X1 i_0_423 (.A1(n_109), .A2(n_0_3), .B1(n_93), .B2(n_0_2), .C1(n_217), 
      .C2(n_0_1), .ZN(n_0_233));
   INV_X1 i_0_424 (.A(n_0_234), .ZN(n_202));
   AOI221_X1 i_0_425 (.A(n_0_0), .B1(n_94), .B2(n_0_2), .C1(n_110), .C2(n_0_3), 
      .ZN(n_0_234));
   INV_X1 i_0_426 (.A(n_0_235), .ZN(n_203));
   AOI221_X1 i_0_427 (.A(n_0_0), .B1(n_95), .B2(n_0_2), .C1(n_111), .C2(n_0_3), 
      .ZN(n_0_235));
   AND2_X1 i_0_428 (.A1(n_218), .A2(n_0_1), .ZN(n_0_0));
   NOR2_X1 i_0_429 (.A1(n_0_3), .A2(n_0_2), .ZN(n_0_1));
   NOR2_X1 i_0_430 (.A1(A[4]), .A2(n_0_155), .ZN(n_0_2));
   NOR2_X1 i_0_431 (.A1(n_0_156), .A2(A[3]), .ZN(n_0_3));
   INV_X1 i_0_432 (.A(n_0_4), .ZN(product[3]));
   AOI222_X1 i_0_433 (.A1(n_48), .A2(n_0_22), .B1(n_64), .B2(n_0_23), .C1(n_219), 
      .C2(n_0_21), .ZN(n_0_4));
   INV_X1 i_0_434 (.A(n_0_5), .ZN(n_204));
   AOI222_X1 i_0_435 (.A1(n_49), .A2(n_0_22), .B1(n_65), .B2(n_0_23), .C1(n_220), 
      .C2(n_0_21), .ZN(n_0_5));
   INV_X1 i_0_436 (.A(n_0_6), .ZN(n_205));
   AOI222_X1 i_0_437 (.A1(n_50), .A2(n_0_22), .B1(n_66), .B2(n_0_23), .C1(n_221), 
      .C2(n_0_21), .ZN(n_0_6));
   INV_X1 i_0_438 (.A(n_0_7), .ZN(n_206));
   AOI222_X1 i_0_439 (.A1(n_51), .A2(n_0_22), .B1(n_67), .B2(n_0_23), .C1(n_222), 
      .C2(n_0_21), .ZN(n_0_7));
   INV_X1 i_0_440 (.A(n_0_8), .ZN(n_207));
   AOI222_X1 i_0_441 (.A1(n_52), .A2(n_0_22), .B1(n_68), .B2(n_0_23), .C1(n_223), 
      .C2(n_0_21), .ZN(n_0_8));
   INV_X1 i_0_442 (.A(n_0_9), .ZN(n_208));
   AOI222_X1 i_0_443 (.A1(n_53), .A2(n_0_22), .B1(n_69), .B2(n_0_23), .C1(n_224), 
      .C2(n_0_21), .ZN(n_0_9));
   INV_X1 i_0_444 (.A(n_0_10), .ZN(n_209));
   AOI222_X1 i_0_445 (.A1(n_54), .A2(n_0_22), .B1(n_70), .B2(n_0_23), .C1(n_225), 
      .C2(n_0_21), .ZN(n_0_10));
   INV_X1 i_0_446 (.A(n_0_11), .ZN(n_210));
   AOI222_X1 i_0_447 (.A1(n_55), .A2(n_0_22), .B1(n_71), .B2(n_0_23), .C1(n_226), 
      .C2(n_0_21), .ZN(n_0_11));
   INV_X1 i_0_448 (.A(n_0_12), .ZN(n_211));
   AOI222_X1 i_0_449 (.A1(n_56), .A2(n_0_22), .B1(n_72), .B2(n_0_23), .C1(n_227), 
      .C2(n_0_21), .ZN(n_0_12));
   INV_X1 i_0_450 (.A(n_0_13), .ZN(n_212));
   AOI222_X1 i_0_451 (.A1(n_57), .A2(n_0_22), .B1(n_73), .B2(n_0_23), .C1(n_228), 
      .C2(n_0_21), .ZN(n_0_13));
   INV_X1 i_0_452 (.A(n_0_14), .ZN(n_213));
   AOI222_X1 i_0_453 (.A1(n_58), .A2(n_0_22), .B1(n_74), .B2(n_0_23), .C1(n_229), 
      .C2(n_0_21), .ZN(n_0_14));
   INV_X1 i_0_454 (.A(n_0_15), .ZN(n_214));
   AOI222_X1 i_0_455 (.A1(n_59), .A2(n_0_22), .B1(n_75), .B2(n_0_23), .C1(n_230), 
      .C2(n_0_21), .ZN(n_0_15));
   INV_X1 i_0_456 (.A(n_0_16), .ZN(n_215));
   AOI222_X1 i_0_457 (.A1(n_76), .A2(n_0_23), .B1(n_60), .B2(n_0_22), .C1(n_231), 
      .C2(n_0_21), .ZN(n_0_16));
   INV_X1 i_0_458 (.A(n_0_17), .ZN(n_216));
   AOI222_X1 i_0_459 (.A1(n_77), .A2(n_0_23), .B1(n_61), .B2(n_0_22), .C1(n_232), 
      .C2(n_0_21), .ZN(n_0_17));
   INV_X1 i_0_460 (.A(n_0_18), .ZN(n_217));
   AOI221_X1 i_0_461 (.A(n_0_20), .B1(n_62), .B2(n_0_22), .C1(n_78), .C2(n_0_23), 
      .ZN(n_0_18));
   INV_X1 i_0_462 (.A(n_0_19), .ZN(n_218));
   AOI221_X1 i_0_463 (.A(n_0_20), .B1(n_63), .B2(n_0_22), .C1(n_79), .C2(n_0_23), 
      .ZN(n_0_19));
   AND2_X1 i_0_464 (.A1(n_233), .A2(n_0_21), .ZN(n_0_20));
   NOR2_X1 i_0_465 (.A1(n_0_23), .A2(n_0_22), .ZN(n_0_21));
   NOR2_X1 i_0_466 (.A1(A[3]), .A2(n_0_154), .ZN(n_0_22));
   NOR2_X1 i_0_467 (.A1(n_0_155), .A2(A[2]), .ZN(n_0_23));
   INV_X1 i_0_468 (.A(n_0_24), .ZN(product[2]));
   AOI222_X1 i_0_469 (.A1(n_16), .A2(n_0_42), .B1(n_32), .B2(n_0_43), .C1(n_234), 
      .C2(n_0_41), .ZN(n_0_24));
   INV_X1 i_0_470 (.A(n_0_25), .ZN(n_219));
   AOI222_X1 i_0_471 (.A1(n_17), .A2(n_0_42), .B1(n_33), .B2(n_0_43), .C1(n_235), 
      .C2(n_0_41), .ZN(n_0_25));
   INV_X1 i_0_472 (.A(n_0_26), .ZN(n_220));
   AOI222_X1 i_0_473 (.A1(n_18), .A2(n_0_42), .B1(n_34), .B2(n_0_43), .C1(n_236), 
      .C2(n_0_41), .ZN(n_0_26));
   INV_X1 i_0_474 (.A(n_0_27), .ZN(n_221));
   AOI222_X1 i_0_475 (.A1(n_19), .A2(n_0_42), .B1(n_35), .B2(n_0_43), .C1(n_237), 
      .C2(n_0_41), .ZN(n_0_27));
   INV_X1 i_0_476 (.A(n_0_28), .ZN(n_222));
   AOI222_X1 i_0_477 (.A1(n_20), .A2(n_0_42), .B1(n_36), .B2(n_0_43), .C1(n_238), 
      .C2(n_0_41), .ZN(n_0_28));
   INV_X1 i_0_478 (.A(n_0_29), .ZN(n_223));
   AOI222_X1 i_0_479 (.A1(n_21), .A2(n_0_42), .B1(n_37), .B2(n_0_43), .C1(n_239), 
      .C2(n_0_41), .ZN(n_0_29));
   INV_X1 i_0_480 (.A(n_0_30), .ZN(n_224));
   AOI222_X1 i_0_481 (.A1(n_22), .A2(n_0_42), .B1(n_38), .B2(n_0_43), .C1(n_240), 
      .C2(n_0_41), .ZN(n_0_30));
   INV_X1 i_0_482 (.A(n_0_31), .ZN(n_225));
   AOI222_X1 i_0_483 (.A1(n_23), .A2(n_0_42), .B1(n_39), .B2(n_0_43), .C1(n_241), 
      .C2(n_0_41), .ZN(n_0_31));
   INV_X1 i_0_484 (.A(n_0_32), .ZN(n_226));
   AOI222_X1 i_0_485 (.A1(n_24), .A2(n_0_42), .B1(n_40), .B2(n_0_43), .C1(n_242), 
      .C2(n_0_41), .ZN(n_0_32));
   INV_X1 i_0_486 (.A(n_0_33), .ZN(n_227));
   AOI222_X1 i_0_487 (.A1(n_25), .A2(n_0_42), .B1(n_41), .B2(n_0_43), .C1(n_243), 
      .C2(n_0_41), .ZN(n_0_33));
   INV_X1 i_0_488 (.A(n_0_34), .ZN(n_228));
   AOI222_X1 i_0_489 (.A1(n_26), .A2(n_0_42), .B1(n_42), .B2(n_0_43), .C1(n_244), 
      .C2(n_0_41), .ZN(n_0_34));
   INV_X1 i_0_490 (.A(n_0_35), .ZN(n_229));
   AOI222_X1 i_0_491 (.A1(n_27), .A2(n_0_42), .B1(n_43), .B2(n_0_43), .C1(n_245), 
      .C2(n_0_41), .ZN(n_0_35));
   INV_X1 i_0_492 (.A(n_0_36), .ZN(n_230));
   AOI222_X1 i_0_493 (.A1(n_28), .A2(n_0_42), .B1(n_44), .B2(n_0_43), .C1(n_246), 
      .C2(n_0_41), .ZN(n_0_36));
   INV_X1 i_0_494 (.A(n_0_37), .ZN(n_231));
   AOI222_X1 i_0_495 (.A1(n_45), .A2(n_0_43), .B1(n_29), .B2(n_0_42), .C1(n_247), 
      .C2(n_0_41), .ZN(n_0_37));
   INV_X1 i_0_496 (.A(n_0_38), .ZN(n_232));
   AOI221_X1 i_0_497 (.A(n_0_40), .B1(n_30), .B2(n_0_42), .C1(n_46), .C2(n_0_43), 
      .ZN(n_0_38));
   INV_X1 i_0_498 (.A(n_0_39), .ZN(n_233));
   AOI221_X1 i_0_499 (.A(n_0_40), .B1(n_31), .B2(n_0_42), .C1(n_47), .C2(n_0_43), 
      .ZN(n_0_39));
   AND2_X1 i_0_500 (.A1(n_248), .A2(n_0_41), .ZN(n_0_40));
   NOR2_X1 i_0_501 (.A1(n_0_43), .A2(n_0_42), .ZN(n_0_41));
   NOR2_X1 i_0_502 (.A1(A[2]), .A2(n_0_153), .ZN(n_0_42));
   NOR2_X1 i_0_503 (.A1(n_0_154), .A2(A[1]), .ZN(n_0_43));
   INV_X1 i_0_504 (.A(n_0_44), .ZN(product[1]));
   AOI222_X1 i_0_505 (.A1(n_0), .A2(n_0_70), .B1(B[0]), .B2(n_0_59), .C1(n_250), 
      .C2(n_0_68), .ZN(n_0_44));
   INV_X1 i_0_506 (.A(n_0_45), .ZN(n_234));
   AOI222_X1 i_0_507 (.A1(n_1), .A2(n_0_70), .B1(n_250), .B2(n_0_59), .C1(n_251), 
      .C2(n_0_68), .ZN(n_0_45));
   INV_X1 i_0_508 (.A(n_0_46), .ZN(n_235));
   AOI222_X1 i_0_509 (.A1(n_2), .A2(n_0_70), .B1(n_251), .B2(n_0_59), .C1(n_252), 
      .C2(n_0_68), .ZN(n_0_46));
   INV_X1 i_0_510 (.A(n_0_47), .ZN(n_236));
   AOI222_X1 i_0_511 (.A1(n_252), .A2(n_0_59), .B1(n_3), .B2(n_0_70), .C1(n_253), 
      .C2(n_0_68), .ZN(n_0_47));
   INV_X1 i_0_512 (.A(n_0_48), .ZN(n_237));
   AOI222_X1 i_0_513 (.A1(n_253), .A2(n_0_59), .B1(n_4), .B2(n_0_70), .C1(n_254), 
      .C2(n_0_68), .ZN(n_0_48));
   INV_X1 i_0_514 (.A(n_0_49), .ZN(n_238));
   AOI222_X1 i_0_515 (.A1(n_5), .A2(n_0_70), .B1(n_254), .B2(n_0_59), .C1(n_255), 
      .C2(n_0_68), .ZN(n_0_49));
   INV_X1 i_0_516 (.A(n_0_50), .ZN(n_239));
   AOI222_X1 i_0_517 (.A1(n_6), .A2(n_0_70), .B1(n_255), .B2(n_0_59), .C1(n_256), 
      .C2(n_0_68), .ZN(n_0_50));
   INV_X1 i_0_518 (.A(n_0_51), .ZN(n_240));
   AOI222_X1 i_0_519 (.A1(n_7), .A2(n_0_70), .B1(n_256), .B2(n_0_59), .C1(n_257), 
      .C2(n_0_68), .ZN(n_0_51));
   INV_X1 i_0_520 (.A(n_0_52), .ZN(n_241));
   AOI222_X1 i_0_521 (.A1(n_8), .A2(n_0_70), .B1(n_257), .B2(n_0_59), .C1(n_258), 
      .C2(n_0_68), .ZN(n_0_52));
   INV_X1 i_0_522 (.A(n_0_53), .ZN(n_242));
   AOI222_X1 i_0_523 (.A1(n_9), .A2(n_0_70), .B1(n_258), .B2(n_0_59), .C1(n_259), 
      .C2(n_0_68), .ZN(n_0_53));
   INV_X1 i_0_524 (.A(n_0_54), .ZN(n_243));
   AOI222_X1 i_0_525 (.A1(n_259), .A2(n_0_59), .B1(n_10), .B2(n_0_70), .C1(n_260), 
      .C2(n_0_68), .ZN(n_0_54));
   INV_X1 i_0_526 (.A(n_0_55), .ZN(n_244));
   AOI222_X1 i_0_527 (.A1(n_260), .A2(n_0_59), .B1(n_11), .B2(n_0_70), .C1(n_261), 
      .C2(n_0_68), .ZN(n_0_55));
   INV_X1 i_0_528 (.A(n_0_56), .ZN(n_245));
   AOI222_X1 i_0_529 (.A1(n_12), .A2(n_0_70), .B1(n_261), .B2(n_0_59), .C1(n_262), 
      .C2(n_0_68), .ZN(n_0_56));
   INV_X1 i_0_530 (.A(n_0_57), .ZN(n_246));
   AOI222_X1 i_0_531 (.A1(n_13), .A2(n_0_70), .B1(n_262), .B2(n_0_59), .C1(n_263), 
      .C2(n_0_68), .ZN(n_0_57));
   INV_X1 i_0_532 (.A(n_0_58), .ZN(n_247));
   AOI222_X1 i_0_533 (.A1(n_263), .A2(n_0_59), .B1(n_14), .B2(n_0_70), .C1(n_264), 
      .C2(n_0_68), .ZN(n_0_58));
   NOR2_X1 i_0_534 (.A1(n_0_153), .A2(A[0]), .ZN(n_0_59));
   NOR2_X1 i_0_535 (.A1(n_0_152), .A2(n_0_70), .ZN(n_0_68));
   INV_X1 i_0_536 (.A(n_0_69), .ZN(n_248));
   AOI22_X1 i_0_537 (.A1(n_15), .A2(n_0_70), .B1(A[1]), .B2(n_264), .ZN(n_0_69));
   NOR2_X1 i_0_538 (.A1(A[1]), .A2(n_0_152), .ZN(n_0_70));
   AND2_X1 i_0_539 (.A1(B[0]), .A2(A[0]), .ZN(product[0]));
   AND2_X1 i_0_540 (.A1(A[0]), .A2(n_264), .ZN(n_249));
   AOI21_X1 i_0_541 (.A(n_0_136), .B1(B[1]), .B2(B[0]), .ZN(n_250));
   AOI21_X1 i_0_542 (.A(n_0_134), .B1(B[2]), .B2(n_0_135), .ZN(n_251));
   AOI21_X1 i_0_543 (.A(n_0_132), .B1(B[3]), .B2(n_0_133), .ZN(n_252));
   AOI21_X1 i_0_544 (.A(n_0_116), .B1(B[4]), .B2(n_0_131), .ZN(n_253));
   AOI21_X1 i_0_545 (.A(n_0_114), .B1(B[5]), .B2(n_0_115), .ZN(n_254));
   AOI21_X1 i_0_546 (.A(n_0_112), .B1(B[6]), .B2(n_0_113), .ZN(n_255));
   AOI21_X1 i_0_547 (.A(n_0_110), .B1(B[7]), .B2(n_0_111), .ZN(n_256));
   AOI21_X1 i_0_548 (.A(n_0_95), .B1(B[8]), .B2(n_0_96), .ZN(n_257));
   AOI21_X1 i_0_549 (.A(n_0_93), .B1(B[9]), .B2(n_0_94), .ZN(n_258));
   AOI21_X1 i_0_550 (.A(n_0_91), .B1(B[10]), .B2(n_0_92), .ZN(n_259));
   AOI21_X1 i_0_551 (.A(n_0_89), .B1(B[11]), .B2(n_0_90), .ZN(n_260));
   AOI21_X1 i_0_552 (.A(n_0_75), .B1(B[15]), .B2(n_0_76), .ZN(n_261));
   AOI21_X1 i_0_553 (.A(n_0_73), .B1(B[15]), .B2(n_0_74), .ZN(n_262));
   AOI21_X1 i_0_554 (.A(n_0_71), .B1(B[15]), .B2(n_0_72), .ZN(n_263));
   XNOR2_X1 i_0_555 (.A(B[15]), .B(n_0_71), .ZN(n_264));
   NOR2_X1 i_0_556 (.A1(B[15]), .A2(n_0_72), .ZN(n_0_71));
   INV_X1 i_0_557 (.A(n_0_73), .ZN(n_0_72));
   NOR2_X1 i_0_558 (.A1(B[15]), .A2(n_0_74), .ZN(n_0_73));
   INV_X1 i_0_559 (.A(n_0_75), .ZN(n_0_74));
   NOR2_X1 i_0_560 (.A1(B[15]), .A2(n_0_76), .ZN(n_0_75));
   INV_X1 i_0_561 (.A(n_0_89), .ZN(n_0_76));
   NOR2_X1 i_0_562 (.A1(B[11]), .A2(n_0_90), .ZN(n_0_89));
   INV_X1 i_0_563 (.A(n_0_91), .ZN(n_0_90));
   NOR2_X1 i_0_564 (.A1(B[10]), .A2(n_0_92), .ZN(n_0_91));
   INV_X1 i_0_565 (.A(n_0_93), .ZN(n_0_92));
   NOR2_X1 i_0_566 (.A1(B[9]), .A2(n_0_94), .ZN(n_0_93));
   INV_X1 i_0_567 (.A(n_0_95), .ZN(n_0_94));
   NOR2_X1 i_0_568 (.A1(B[8]), .A2(n_0_96), .ZN(n_0_95));
   INV_X1 i_0_569 (.A(n_0_110), .ZN(n_0_96));
   NOR2_X1 i_0_570 (.A1(B[7]), .A2(n_0_111), .ZN(n_0_110));
   INV_X1 i_0_571 (.A(n_0_112), .ZN(n_0_111));
   NOR2_X1 i_0_572 (.A1(B[6]), .A2(n_0_113), .ZN(n_0_112));
   INV_X1 i_0_573 (.A(n_0_114), .ZN(n_0_113));
   NOR2_X1 i_0_574 (.A1(B[5]), .A2(n_0_115), .ZN(n_0_114));
   INV_X1 i_0_575 (.A(n_0_116), .ZN(n_0_115));
   NOR2_X1 i_0_576 (.A1(B[4]), .A2(n_0_131), .ZN(n_0_116));
   INV_X1 i_0_577 (.A(n_0_132), .ZN(n_0_131));
   NOR2_X1 i_0_578 (.A1(B[3]), .A2(n_0_133), .ZN(n_0_132));
   INV_X1 i_0_579 (.A(n_0_134), .ZN(n_0_133));
   NOR2_X1 i_0_580 (.A1(B[2]), .A2(n_0_135), .ZN(n_0_134));
   INV_X1 i_0_581 (.A(n_0_136), .ZN(n_0_135));
   NOR2_X1 i_0_582 (.A1(B[1]), .A2(B[0]), .ZN(n_0_136));
   INV_X1 i_0_583 (.A(A[0]), .ZN(n_0_152));
   INV_X1 i_0_584 (.A(A[1]), .ZN(n_0_153));
   INV_X1 i_0_585 (.A(A[2]), .ZN(n_0_154));
   INV_X1 i_0_586 (.A(A[3]), .ZN(n_0_155));
   INV_X1 i_0_587 (.A(A[4]), .ZN(n_0_156));
   INV_X1 i_0_588 (.A(A[5]), .ZN(n_0_173));
   INV_X1 i_0_589 (.A(A[6]), .ZN(n_0_174));
   INV_X1 i_0_590 (.A(A[7]), .ZN(n_0_175));
   INV_X1 i_0_591 (.A(A[8]), .ZN(n_0_176));
   INV_X1 i_0_592 (.A(A[9]), .ZN(n_0_194));
   INV_X1 i_0_593 (.A(A[10]), .ZN(n_0_195));
   INV_X1 i_0_594 (.A(A[11]), .ZN(n_0_196));
   INV_X1 i_0_595 (.A(A[15]), .ZN(n_0_215));
   FA_X1 i_1_0 (.A(B[1]), .B(n_190), .CI(n_1_166), .CO(n_1_2), .S(n_265));
   FA_X1 i_1_1 (.A(B[2]), .B(n_191), .CI(n_1_2), .CO(n_1_3), .S(n_266));
   FA_X1 i_1_2 (.A(B[3]), .B(n_192), .CI(n_1_3), .CO(n_1_4), .S(n_267));
   FA_X1 i_1_3 (.A(B[4]), .B(n_193), .CI(n_1_4), .CO(n_1_5), .S(n_268));
   FA_X1 i_1_4 (.A(B[5]), .B(n_194), .CI(n_1_5), .CO(n_1_6), .S(n_269));
   FA_X1 i_1_5 (.A(B[6]), .B(n_195), .CI(n_1_6), .CO(n_1_7), .S(n_270));
   FA_X1 i_1_6 (.A(B[7]), .B(n_196), .CI(n_1_7), .CO(n_1_8), .S(n_271));
   FA_X1 i_1_7 (.A(B[8]), .B(n_197), .CI(n_1_8), .CO(n_1_9), .S(n_272));
   FA_X1 i_1_8 (.A(B[9]), .B(n_198), .CI(n_1_9), .CO(n_1_10), .S(n_273));
   FA_X1 i_1_9 (.A(B[10]), .B(n_199), .CI(n_1_10), .CO(n_1_11), .S(n_274));
   FA_X1 i_1_10 (.A(B[11]), .B(n_200), .CI(n_1_11), .CO(n_1_12), .S(n_275));
   FA_X1 i_1_11 (.A(B[15]), .B(n_201), .CI(n_1_12), .CO(n_1_13), .S(n_276));
   FA_X1 i_1_12 (.A(B[15]), .B(n_202), .CI(n_1_13), .CO(n_1_14), .S(n_277));
   FA_X1 i_1_13 (.A(n_250), .B(n_190), .CI(n_1_166), .CO(n_1_0), .S(n_278));
   FA_X1 i_1_14 (.A(n_251), .B(n_191), .CI(n_1_0), .CO(n_1_1), .S(n_279));
   FA_X1 i_1_15 (.A(n_252), .B(n_192), .CI(n_1_1), .CO(n_1_15), .S(n_280));
   FA_X1 i_1_16 (.A(n_253), .B(n_193), .CI(n_1_15), .CO(n_1_16), .S(n_281));
   FA_X1 i_1_17 (.A(n_254), .B(n_194), .CI(n_1_16), .CO(n_1_17), .S(n_282));
   FA_X1 i_1_18 (.A(n_255), .B(n_195), .CI(n_1_17), .CO(n_1_18), .S(n_283));
   FA_X1 i_1_19 (.A(n_256), .B(n_196), .CI(n_1_18), .CO(n_1_19), .S(n_284));
   FA_X1 i_1_20 (.A(n_257), .B(n_197), .CI(n_1_19), .CO(n_1_20), .S(n_285));
   FA_X1 i_1_21 (.A(n_258), .B(n_198), .CI(n_1_20), .CO(n_1_21), .S(n_286));
   FA_X1 i_1_22 (.A(n_259), .B(n_199), .CI(n_1_21), .CO(n_1_22), .S(n_287));
   FA_X1 i_1_23 (.A(n_260), .B(n_200), .CI(n_1_22), .CO(n_1_23), .S(n_288));
   FA_X1 i_1_24 (.A(n_261), .B(n_201), .CI(n_1_23), .CO(n_1_24), .S(n_289));
   FA_X1 i_1_25 (.A(n_262), .B(n_202), .CI(n_1_24), .CO(n_1_25), .S(n_290));
   FA_X1 i_1_26 (.A(B[1]), .B(n_176), .CI(n_1_167), .CO(n_1_26), .S(n_291));
   FA_X1 i_1_27 (.A(B[2]), .B(n_177), .CI(n_1_26), .CO(n_1_27), .S(n_292));
   FA_X1 i_1_28 (.A(B[3]), .B(n_178), .CI(n_1_27), .CO(n_1_28), .S(n_293));
   FA_X1 i_1_29 (.A(B[4]), .B(n_179), .CI(n_1_28), .CO(n_1_29), .S(n_294));
   FA_X1 i_1_30 (.A(B[5]), .B(n_180), .CI(n_1_29), .CO(n_1_30), .S(n_295));
   FA_X1 i_1_31 (.A(B[6]), .B(n_181), .CI(n_1_30), .CO(n_1_31), .S(n_296));
   FA_X1 i_1_32 (.A(B[7]), .B(n_182), .CI(n_1_31), .CO(n_1_32), .S(n_297));
   FA_X1 i_1_33 (.A(B[8]), .B(n_183), .CI(n_1_32), .CO(n_1_33), .S(n_298));
   FA_X1 i_1_34 (.A(B[9]), .B(n_184), .CI(n_1_33), .CO(n_1_34), .S(n_299));
   FA_X1 i_1_35 (.A(B[10]), .B(n_185), .CI(n_1_34), .CO(n_1_35), .S(n_300));
   FA_X1 i_1_36 (.A(B[11]), .B(n_186), .CI(n_1_35), .CO(n_1_36), .S(n_301));
   FA_X1 i_1_37 (.A(B[15]), .B(n_187), .CI(n_1_36), .CO(n_1_37), .S(n_302));
   FA_X1 i_1_38 (.A(B[15]), .B(n_188), .CI(n_1_37), .CO(n_1_38), .S(n_303));
   FA_X1 i_1_39 (.A(n_250), .B(n_176), .CI(n_1_167), .CO(n_1_39), .S(n_304));
   FA_X1 i_1_40 (.A(n_251), .B(n_177), .CI(n_1_39), .CO(n_1_40), .S(n_305));
   FA_X1 i_1_41 (.A(n_252), .B(n_178), .CI(n_1_40), .CO(n_1_41), .S(n_306));
   FA_X1 i_1_42 (.A(n_253), .B(n_179), .CI(n_1_41), .CO(n_1_42), .S(n_307));
   FA_X1 i_1_43 (.A(n_254), .B(n_180), .CI(n_1_42), .CO(n_1_43), .S(n_308));
   FA_X1 i_1_44 (.A(n_255), .B(n_181), .CI(n_1_43), .CO(n_1_44), .S(n_309));
   FA_X1 i_1_45 (.A(n_256), .B(n_182), .CI(n_1_44), .CO(n_1_45), .S(n_310));
   FA_X1 i_1_46 (.A(n_257), .B(n_183), .CI(n_1_45), .CO(n_1_46), .S(n_311));
   FA_X1 i_1_47 (.A(n_258), .B(n_184), .CI(n_1_46), .CO(n_1_47), .S(n_312));
   FA_X1 i_1_48 (.A(n_259), .B(n_185), .CI(n_1_47), .CO(n_1_48), .S(n_313));
   FA_X1 i_1_49 (.A(n_260), .B(n_186), .CI(n_1_48), .CO(n_1_49), .S(n_314));
   FA_X1 i_1_50 (.A(n_261), .B(n_187), .CI(n_1_49), .CO(n_1_50), .S(n_315));
   FA_X1 i_1_51 (.A(n_262), .B(n_188), .CI(n_1_50), .CO(n_1_51), .S(n_316));
   FA_X1 i_1_52 (.A(B[1]), .B(n_163), .CI(n_1_168), .CO(n_1_52), .S(n_317));
   FA_X1 i_1_53 (.A(B[2]), .B(n_164), .CI(n_1_52), .CO(n_1_53), .S(n_318));
   FA_X1 i_1_54 (.A(B[3]), .B(n_165), .CI(n_1_53), .CO(n_1_54), .S(n_319));
   FA_X1 i_1_55 (.A(B[4]), .B(n_166), .CI(n_1_54), .CO(n_1_55), .S(n_320));
   FA_X1 i_1_56 (.A(B[5]), .B(n_167), .CI(n_1_55), .CO(n_1_56), .S(n_321));
   FA_X1 i_1_57 (.A(B[6]), .B(n_168), .CI(n_1_56), .CO(n_1_57), .S(n_322));
   FA_X1 i_1_58 (.A(B[7]), .B(n_169), .CI(n_1_57), .CO(n_1_58), .S(n_323));
   FA_X1 i_1_59 (.A(B[8]), .B(n_170), .CI(n_1_58), .CO(n_1_59), .S(n_324));
   FA_X1 i_1_60 (.A(B[9]), .B(n_171), .CI(n_1_59), .CO(n_1_60), .S(n_325));
   FA_X1 i_1_61 (.A(B[10]), .B(n_172), .CI(n_1_60), .CO(n_1_61), .S(n_326));
   FA_X1 i_1_62 (.A(B[11]), .B(n_173), .CI(n_1_61), .CO(n_1_62), .S(n_327));
   FA_X1 i_1_63 (.A(B[15]), .B(n_174), .CI(n_1_62), .CO(n_1_63), .S(n_328));
   FA_X1 i_1_64 (.A(n_250), .B(n_163), .CI(n_1_168), .CO(n_1_64), .S(n_329));
   FA_X1 i_1_65 (.A(n_251), .B(n_164), .CI(n_1_64), .CO(n_1_65), .S(n_330));
   FA_X1 i_1_66 (.A(n_252), .B(n_165), .CI(n_1_65), .CO(n_1_66), .S(n_331));
   FA_X1 i_1_67 (.A(n_253), .B(n_166), .CI(n_1_66), .CO(n_1_67), .S(n_332));
   FA_X1 i_1_68 (.A(n_254), .B(n_167), .CI(n_1_67), .CO(n_1_68), .S(n_333));
   FA_X1 i_1_69 (.A(n_255), .B(n_168), .CI(n_1_68), .CO(n_1_69), .S(n_334));
   FA_X1 i_1_70 (.A(n_256), .B(n_169), .CI(n_1_69), .CO(n_1_70), .S(n_335));
   FA_X1 i_1_71 (.A(n_257), .B(n_170), .CI(n_1_70), .CO(n_1_71), .S(n_336));
   FA_X1 i_1_72 (.A(n_258), .B(n_171), .CI(n_1_71), .CO(n_1_72), .S(n_337));
   FA_X1 i_1_73 (.A(n_259), .B(n_172), .CI(n_1_72), .CO(n_1_73), .S(n_338));
   FA_X1 i_1_74 (.A(n_260), .B(n_173), .CI(n_1_73), .CO(n_1_74), .S(n_339));
   FA_X1 i_1_75 (.A(n_261), .B(n_174), .CI(n_1_74), .CO(n_1_75), .S(n_340));
   FA_X1 i_1_76 (.A(B[1]), .B(n_151), .CI(n_1_169), .CO(n_1_76), .S(n_341));
   FA_X1 i_1_77 (.A(B[2]), .B(n_152), .CI(n_1_76), .CO(n_1_77), .S(n_342));
   FA_X1 i_1_78 (.A(B[3]), .B(n_153), .CI(n_1_77), .CO(n_1_78), .S(n_343));
   FA_X1 i_1_79 (.A(B[4]), .B(n_154), .CI(n_1_78), .CO(n_1_79), .S(n_344));
   FA_X1 i_1_80 (.A(B[5]), .B(n_155), .CI(n_1_79), .CO(n_1_80), .S(n_345));
   FA_X1 i_1_81 (.A(B[6]), .B(n_156), .CI(n_1_80), .CO(n_1_81), .S(n_346));
   FA_X1 i_1_82 (.A(B[7]), .B(n_157), .CI(n_1_81), .CO(n_1_82), .S(n_347));
   FA_X1 i_1_83 (.A(B[8]), .B(n_158), .CI(n_1_82), .CO(n_1_83), .S(n_348));
   FA_X1 i_1_84 (.A(B[9]), .B(n_159), .CI(n_1_83), .CO(n_1_84), .S(n_349));
   FA_X1 i_1_85 (.A(B[10]), .B(n_160), .CI(n_1_84), .CO(n_1_85), .S(n_350));
   FA_X1 i_1_86 (.A(B[11]), .B(n_161), .CI(n_1_85), .CO(n_1_86), .S(n_351));
   FA_X1 i_1_87 (.A(n_250), .B(n_151), .CI(n_1_169), .CO(n_1_87), .S(n_352));
   FA_X1 i_1_88 (.A(n_251), .B(n_152), .CI(n_1_87), .CO(n_1_88), .S(n_353));
   FA_X1 i_1_89 (.A(n_252), .B(n_153), .CI(n_1_88), .CO(n_1_89), .S(n_354));
   FA_X1 i_1_90 (.A(n_253), .B(n_154), .CI(n_1_89), .CO(n_1_90), .S(n_355));
   FA_X1 i_1_91 (.A(n_254), .B(n_155), .CI(n_1_90), .CO(n_1_91), .S(n_356));
   FA_X1 i_1_92 (.A(n_255), .B(n_156), .CI(n_1_91), .CO(n_1_92), .S(n_357));
   FA_X1 i_1_93 (.A(n_256), .B(n_157), .CI(n_1_92), .CO(n_1_93), .S(n_358));
   FA_X1 i_1_94 (.A(n_257), .B(n_158), .CI(n_1_93), .CO(n_1_94), .S(n_359));
   FA_X1 i_1_95 (.A(n_258), .B(n_159), .CI(n_1_94), .CO(n_1_95), .S(n_360));
   FA_X1 i_1_96 (.A(n_259), .B(n_160), .CI(n_1_95), .CO(n_1_96), .S(n_361));
   FA_X1 i_1_97 (.A(n_260), .B(n_161), .CI(n_1_96), .CO(n_1_97), .S(n_362));
   FA_X1 i_1_98 (.A(B[1]), .B(n_140), .CI(n_1_170), .CO(n_1_98), .S(n_363));
   FA_X1 i_1_99 (.A(B[2]), .B(n_141), .CI(n_1_98), .CO(n_1_99), .S(n_364));
   FA_X1 i_1_100 (.A(B[3]), .B(n_142), .CI(n_1_99), .CO(n_1_100), .S(n_365));
   FA_X1 i_1_101 (.A(B[4]), .B(n_143), .CI(n_1_100), .CO(n_1_101), .S(n_366));
   FA_X1 i_1_102 (.A(B[5]), .B(n_144), .CI(n_1_101), .CO(n_1_102), .S(n_367));
   FA_X1 i_1_103 (.A(B[6]), .B(n_145), .CI(n_1_102), .CO(n_1_103), .S(n_368));
   FA_X1 i_1_104 (.A(B[7]), .B(n_146), .CI(n_1_103), .CO(n_1_104), .S(n_369));
   FA_X1 i_1_105 (.A(B[8]), .B(n_147), .CI(n_1_104), .CO(n_1_105), .S(n_370));
   FA_X1 i_1_106 (.A(B[9]), .B(n_148), .CI(n_1_105), .CO(n_1_106), .S(n_371));
   FA_X1 i_1_107 (.A(B[10]), .B(n_149), .CI(n_1_106), .CO(n_1_107), .S(n_372));
   FA_X1 i_1_108 (.A(n_250), .B(n_140), .CI(n_1_170), .CO(n_1_108), .S(n_373));
   FA_X1 i_1_109 (.A(n_251), .B(n_141), .CI(n_1_108), .CO(n_1_109), .S(n_374));
   FA_X1 i_1_110 (.A(n_252), .B(n_142), .CI(n_1_109), .CO(n_1_110), .S(n_375));
   FA_X1 i_1_111 (.A(n_253), .B(n_143), .CI(n_1_110), .CO(n_1_111), .S(n_376));
   FA_X1 i_1_112 (.A(n_254), .B(n_144), .CI(n_1_111), .CO(n_1_112), .S(n_377));
   FA_X1 i_1_113 (.A(n_255), .B(n_145), .CI(n_1_112), .CO(n_1_113), .S(n_378));
   FA_X1 i_1_114 (.A(n_256), .B(n_146), .CI(n_1_113), .CO(n_1_114), .S(n_379));
   FA_X1 i_1_115 (.A(n_257), .B(n_147), .CI(n_1_114), .CO(n_1_115), .S(n_380));
   FA_X1 i_1_116 (.A(n_258), .B(n_148), .CI(n_1_115), .CO(n_1_116), .S(n_381));
   FA_X1 i_1_117 (.A(n_259), .B(n_149), .CI(n_1_116), .CO(n_1_117), .S(n_382));
   FA_X1 i_1_118 (.A(B[1]), .B(n_130), .CI(n_1_171), .CO(n_1_118), .S(n_383));
   FA_X1 i_1_119 (.A(B[2]), .B(n_131), .CI(n_1_118), .CO(n_1_119), .S(n_384));
   FA_X1 i_1_120 (.A(B[3]), .B(n_132), .CI(n_1_119), .CO(n_1_120), .S(n_385));
   FA_X1 i_1_121 (.A(B[4]), .B(n_133), .CI(n_1_120), .CO(n_1_121), .S(n_386));
   FA_X1 i_1_122 (.A(B[5]), .B(n_134), .CI(n_1_121), .CO(n_1_122), .S(n_387));
   FA_X1 i_1_123 (.A(B[6]), .B(n_135), .CI(n_1_122), .CO(n_1_123), .S(n_388));
   FA_X1 i_1_124 (.A(B[7]), .B(n_136), .CI(n_1_123), .CO(n_1_124), .S(n_389));
   FA_X1 i_1_125 (.A(B[8]), .B(n_137), .CI(n_1_124), .CO(n_1_125), .S(n_390));
   FA_X1 i_1_126 (.A(B[9]), .B(n_138), .CI(n_1_125), .CO(n_1_126), .S(n_391));
   FA_X1 i_1_127 (.A(n_250), .B(n_130), .CI(n_1_171), .CO(n_1_127), .S(n_392));
   FA_X1 i_1_128 (.A(n_251), .B(n_131), .CI(n_1_127), .CO(n_1_128), .S(n_393));
   FA_X1 i_1_129 (.A(n_252), .B(n_132), .CI(n_1_128), .CO(n_1_129), .S(n_394));
   FA_X1 i_1_130 (.A(n_253), .B(n_133), .CI(n_1_129), .CO(n_1_130), .S(n_395));
   FA_X1 i_1_131 (.A(n_254), .B(n_134), .CI(n_1_130), .CO(n_1_131), .S(n_396));
   FA_X1 i_1_132 (.A(n_255), .B(n_135), .CI(n_1_131), .CO(n_1_132), .S(n_397));
   FA_X1 i_1_133 (.A(n_256), .B(n_136), .CI(n_1_132), .CO(n_1_133), .S(n_398));
   FA_X1 i_1_134 (.A(n_257), .B(n_137), .CI(n_1_133), .CO(n_1_134), .S(n_399));
   FA_X1 i_1_135 (.A(n_258), .B(n_138), .CI(n_1_134), .CO(n_1_135), .S(n_400));
   FA_X1 i_1_136 (.A(B[1]), .B(n_121), .CI(n_1_172), .CO(n_1_136), .S(n_401));
   FA_X1 i_1_137 (.A(B[2]), .B(n_122), .CI(n_1_136), .CO(n_1_137), .S(n_402));
   FA_X1 i_1_138 (.A(B[3]), .B(n_123), .CI(n_1_137), .CO(n_1_138), .S(n_403));
   FA_X1 i_1_139 (.A(B[4]), .B(n_124), .CI(n_1_138), .CO(n_1_139), .S(n_404));
   FA_X1 i_1_140 (.A(B[5]), .B(n_125), .CI(n_1_139), .CO(n_1_140), .S(n_405));
   FA_X1 i_1_141 (.A(B[6]), .B(n_126), .CI(n_1_140), .CO(n_1_141), .S(n_406));
   FA_X1 i_1_142 (.A(B[7]), .B(n_127), .CI(n_1_141), .CO(n_1_142), .S(n_407));
   FA_X1 i_1_143 (.A(B[8]), .B(n_128), .CI(n_1_142), .CO(n_1_143), .S(n_408));
   FA_X1 i_1_144 (.A(n_250), .B(n_121), .CI(n_1_172), .CO(n_1_144), .S(n_409));
   FA_X1 i_1_145 (.A(n_251), .B(n_122), .CI(n_1_144), .CO(n_1_145), .S(n_410));
   FA_X1 i_1_146 (.A(n_252), .B(n_123), .CI(n_1_145), .CO(n_1_146), .S(n_411));
   FA_X1 i_1_147 (.A(n_253), .B(n_124), .CI(n_1_146), .CO(n_1_147), .S(n_412));
   FA_X1 i_1_148 (.A(n_254), .B(n_125), .CI(n_1_147), .CO(n_1_148), .S(n_413));
   FA_X1 i_1_149 (.A(n_255), .B(n_126), .CI(n_1_148), .CO(n_1_149), .S(n_414));
   FA_X1 i_1_150 (.A(n_256), .B(n_127), .CI(n_1_149), .CO(n_1_150), .S(n_415));
   FA_X1 i_1_151 (.A(n_257), .B(n_128), .CI(n_1_150), .CO(n_1_151), .S(n_416));
   FA_X1 i_1_152 (.A(B[1]), .B(n_113), .CI(n_1_173), .CO(n_1_152), .S(n_417));
   FA_X1 i_1_153 (.A(B[2]), .B(n_114), .CI(n_1_152), .CO(n_1_153), .S(n_418));
   FA_X1 i_1_154 (.A(B[3]), .B(n_115), .CI(n_1_153), .CO(n_1_154), .S(n_419));
   FA_X1 i_1_155 (.A(B[4]), .B(n_116), .CI(n_1_154), .CO(n_1_155), .S(n_420));
   FA_X1 i_1_156 (.A(B[5]), .B(n_117), .CI(n_1_155), .CO(n_1_156), .S(n_421));
   FA_X1 i_1_157 (.A(B[6]), .B(n_118), .CI(n_1_156), .CO(n_1_157), .S(n_422));
   FA_X1 i_1_158 (.A(B[7]), .B(n_119), .CI(n_1_157), .CO(n_1_158), .S(n_423));
   FA_X1 i_1_159 (.A(n_250), .B(n_113), .CI(n_1_173), .CO(n_1_159), .S(n_424));
   FA_X1 i_1_160 (.A(n_251), .B(n_114), .CI(n_1_159), .CO(n_1_160), .S(n_425));
   FA_X1 i_1_161 (.A(n_252), .B(n_115), .CI(n_1_160), .CO(n_1_161), .S(n_426));
   FA_X1 i_1_162 (.A(n_253), .B(n_116), .CI(n_1_161), .CO(n_1_162), .S(n_427));
   FA_X1 i_1_163 (.A(n_254), .B(n_117), .CI(n_1_162), .CO(n_1_163), .S(n_428));
   FA_X1 i_1_164 (.A(n_255), .B(n_118), .CI(n_1_163), .CO(n_1_164), .S(n_429));
   FA_X1 i_1_165 (.A(n_256), .B(n_119), .CI(n_1_164), .CO(n_1_165), .S(n_430));
   HA_X1 i_1_166 (.A(B[0]), .B(n_189), .CO(n_1_166), .S(n_431));
   HA_X1 i_1_167 (.A(B[0]), .B(n_175), .CO(n_1_167), .S(n_432));
   HA_X1 i_1_168 (.A(B[0]), .B(n_162), .CO(n_1_168), .S(n_433));
   HA_X1 i_1_169 (.A(B[0]), .B(n_150), .CO(n_1_169), .S(n_434));
   HA_X1 i_1_170 (.A(B[0]), .B(n_139), .CO(n_1_170), .S(n_435));
   HA_X1 i_1_171 (.A(B[0]), .B(n_129), .CO(n_1_171), .S(n_436));
   HA_X1 i_1_172 (.A(B[0]), .B(n_120), .CO(n_1_172), .S(n_437));
   HA_X1 i_1_173 (.A(B[0]), .B(n_112), .CO(n_1_173), .S(n_438));
   XNOR2_X1 i_1_174 (.A(n_203), .B(n_1_174), .ZN(n_439));
   XNOR2_X1 i_1_175 (.A(n_263), .B(n_1_25), .ZN(n_1_174));
   XNOR2_X1 i_1_176 (.A(B[15]), .B(n_1_175), .ZN(n_440));
   XNOR2_X1 i_1_177 (.A(n_203), .B(n_1_14), .ZN(n_1_175));
endmodule

module multiplier_16bit__0_313(first_operand, second_operand, out, enable, 
      overflow);
   input [15:0]first_operand;
   input [15:0]second_operand;
   output [15:0]out;
   input enable;
   output overflow;

   wire [31:0]temp_result_wire;
   wire n_0_0_4;
   wire n_0_0_6;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_5;
   wire n_0_0_7;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;

   booth_16bit_multiplier__1 mult (.A({first_operand[12], uc_0, uc_1, uc_2, 
      first_operand[11], first_operand[10], first_operand[9], first_operand[8], 
      first_operand[7], first_operand[6], first_operand[5], first_operand[4], 
      first_operand[3], first_operand[2], first_operand[1], first_operand[0]}), 
      .B({second_operand[12], uc_3, uc_4, uc_5, second_operand[11], 
      second_operand[10], second_operand[9], second_operand[8], 
      second_operand[7], second_operand[6], second_operand[5], second_operand[4], 
      second_operand[3], second_operand[2], second_operand[1], second_operand[0]}), 
      .product({uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, 
      uc_16, uc_17, temp_result_wire[19], temp_result_wire[18], 
      temp_result_wire[17], temp_result_wire[16], temp_result_wire[15], 
      temp_result_wire[14], temp_result_wire[13], temp_result_wire[12], 
      temp_result_wire[11], temp_result_wire[10], temp_result_wire[9], 
      temp_result_wire[8], temp_result_wire[7], temp_result_wire[6], 
      temp_result_wire[5], temp_result_wire[4], temp_result_wire[3], 
      temp_result_wire[2], temp_result_wire[1], temp_result_wire[0]}));
   MUX2_X1 i_0_0_0 (.A(n_0_0_3), .B(n_0_0_4), .S(n_0_0_46), .Z(out[1]));
   MUX2_X1 i_0_0_1 (.A(n_0_0_4), .B(n_0_0_6), .S(n_0_0_46), .Z(out[2]));
   MUX2_X1 i_0_0_2 (.A(n_0_0_25), .B(n_0_0_9), .S(n_0_0_31), .Z(n_0_0_4));
   MUX2_X1 i_0_0_3 (.A(n_0_0_6), .B(n_0_0_8), .S(n_0_0_46), .Z(out[3]));
   MUX2_X1 i_0_0_4 (.A(n_0_0_7), .B(n_0_0_11), .S(n_0_0_31), .Z(n_0_0_6));
   MUX2_X1 i_0_0_5 (.A(n_0_0_8), .B(n_0_0_10), .S(n_0_0_46), .Z(out[4]));
   MUX2_X1 i_0_0_6 (.A(n_0_0_9), .B(n_0_0_13), .S(n_0_0_31), .Z(n_0_0_8));
   MUX2_X1 i_0_0_7 (.A(temp_result_wire[4]), .B(temp_result_wire[8]), .S(
      n_0_0_28), .Z(n_0_0_9));
   MUX2_X1 i_0_0_15 (.A(n_0_0_10), .B(n_0_0_12), .S(n_0_0_46), .Z(out[5]));
   MUX2_X1 i_0_0_8 (.A(n_0_0_11), .B(n_0_0_15), .S(n_0_0_31), .Z(n_0_0_10));
   MUX2_X1 i_0_0_9 (.A(temp_result_wire[5]), .B(temp_result_wire[9]), .S(
      n_0_0_28), .Z(n_0_0_11));
   MUX2_X1 i_0_0_18 (.A(n_0_0_12), .B(n_0_0_14), .S(n_0_0_46), .Z(out[6]));
   MUX2_X1 i_0_0_19 (.A(n_0_0_13), .B(n_0_0_17), .S(n_0_0_31), .Z(n_0_0_12));
   MUX2_X1 i_0_0_10 (.A(temp_result_wire[6]), .B(temp_result_wire[10]), .S(
      n_0_0_28), .Z(n_0_0_13));
   MUX2_X1 i_0_0_21 (.A(n_0_0_14), .B(n_0_0_16), .S(n_0_0_46), .Z(out[7]));
   MUX2_X1 i_0_0_22 (.A(n_0_0_15), .B(n_0_0_19), .S(n_0_0_31), .Z(n_0_0_14));
   MUX2_X1 i_0_0_11 (.A(temp_result_wire[7]), .B(temp_result_wire[11]), .S(
      n_0_0_28), .Z(n_0_0_15));
   MUX2_X1 i_0_0_24 (.A(n_0_0_16), .B(n_0_0_18), .S(n_0_0_46), .Z(out[8]));
   MUX2_X1 i_0_0_25 (.A(n_0_0_17), .B(n_0_0_21), .S(n_0_0_31), .Z(n_0_0_16));
   MUX2_X1 i_0_0_26 (.A(temp_result_wire[8]), .B(temp_result_wire[12]), .S(
      n_0_0_28), .Z(n_0_0_17));
   MUX2_X1 i_0_0_27 (.A(n_0_0_18), .B(n_0_0_20), .S(n_0_0_46), .Z(out[9]));
   MUX2_X1 i_0_0_28 (.A(n_0_0_19), .B(n_0_0_23), .S(n_0_0_31), .Z(n_0_0_18));
   MUX2_X1 i_0_0_29 (.A(temp_result_wire[9]), .B(temp_result_wire[13]), .S(
      n_0_0_28), .Z(n_0_0_19));
   MUX2_X1 i_0_0_30 (.A(n_0_0_20), .B(n_0_0_22), .S(n_0_0_46), .Z(out[10]));
   MUX2_X1 i_0_0_31 (.A(n_0_0_21), .B(n_0_0_63), .S(n_0_0_31), .Z(n_0_0_20));
   MUX2_X1 i_0_0_32 (.A(temp_result_wire[10]), .B(temp_result_wire[14]), 
      .S(n_0_0_28), .Z(n_0_0_21));
   MUX2_X1 i_0_0_12 (.A(n_0_0_22), .B(n_0_0_61), .S(n_0_0_46), .Z(out[11]));
   MUX2_X1 i_0_0_13 (.A(n_0_0_23), .B(n_0_0_58), .S(n_0_0_31), .Z(n_0_0_22));
   MUX2_X1 i_0_0_14 (.A(temp_result_wire[11]), .B(temp_result_wire[15]), 
      .S(n_0_0_28), .Z(n_0_0_23));
   AOI21_X1 i_0_0_16 (.A(n_0_0_40), .B1(n_0_0_37), .B2(n_0_0_52), .ZN(out[13]));
   NOR2_X1 i_0_0_17 (.A1(n_0_0_37), .A2(first_operand[13]), .ZN(n_0_0_40));
   AOI21_X1 i_0_0_55 (.A(n_0_0_41), .B1(n_0_0_37), .B2(n_0_0_53), .ZN(out[14]));
   NOR2_X1 i_0_0_56 (.A1(n_0_0_37), .A2(first_operand[14]), .ZN(n_0_0_41));
   OR2_X1 i_0_0_64 (.A1(second_operand[15]), .A2(first_operand[15]), .ZN(out[15]));
   INV_X1 i_0_0_20 (.A(n_0_0_0), .ZN(out[0]));
   AOI22_X1 i_0_0_23 (.A1(n_0_0_47), .A2(n_0_0_1), .B1(n_0_0_46), .B2(n_0_0_3), 
      .ZN(n_0_0_0));
   OAI22_X1 i_0_0_33 (.A1(n_0_0_31), .A2(n_0_0_2), .B1(n_0_0_30), .B2(n_0_0_26), 
      .ZN(n_0_0_1));
   AOI22_X1 i_0_0_34 (.A1(temp_result_wire[4]), .A2(n_0_0_28), .B1(
      temp_result_wire[0]), .B2(n_0_0_27), .ZN(n_0_0_2));
   AOI22_X1 i_0_0_35 (.A1(n_0_0_30), .A2(n_0_0_5), .B1(n_0_0_31), .B2(n_0_0_24), 
      .ZN(n_0_0_3));
   OAI22_X1 i_0_0_36 (.A1(temp_result_wire[5]), .A2(n_0_0_27), .B1(
      temp_result_wire[1]), .B2(n_0_0_28), .ZN(n_0_0_5));
   INV_X1 i_0_0_37 (.A(n_0_0_24), .ZN(n_0_0_7));
   OAI22_X1 i_0_0_38 (.A1(temp_result_wire[7]), .A2(n_0_0_27), .B1(
      temp_result_wire[3]), .B2(n_0_0_28), .ZN(n_0_0_24));
   INV_X1 i_0_0_39 (.A(n_0_0_26), .ZN(n_0_0_25));
   OAI22_X1 i_0_0_40 (.A1(temp_result_wire[6]), .A2(n_0_0_27), .B1(
      temp_result_wire[2]), .B2(n_0_0_28), .ZN(n_0_0_26));
   INV_X1 i_0_0_41 (.A(n_0_0_28), .ZN(n_0_0_27));
   OAI33_X1 i_0_0_42 (.A1(n_0_0_54), .A2(first_operand[15]), .A3(n_0_0_38), 
      .B1(n_0_0_45), .B2(n_0_0_39), .B3(n_0_0_29), .ZN(n_0_0_28));
   NOR2_X1 i_0_0_43 (.A1(n_0_0_48), .A2(n_0_0_42), .ZN(n_0_0_29));
   INV_X1 i_0_0_44 (.A(n_0_0_31), .ZN(n_0_0_30));
   OAI21_X1 i_0_0_45 (.A(n_0_0_32), .B1(n_0_0_36), .B2(n_0_0_33), .ZN(n_0_0_31));
   OAI221_X1 i_0_0_46 (.A(n_0_0_36), .B1(n_0_0_49), .B2(n_0_0_34), .C1(n_0_0_48), 
      .C2(n_0_0_35), .ZN(n_0_0_32));
   AOI22_X1 i_0_0_47 (.A1(n_0_0_51), .A2(n_0_0_34), .B1(n_0_0_50), .B2(n_0_0_35), 
      .ZN(n_0_0_33));
   INV_X1 i_0_0_48 (.A(n_0_0_35), .ZN(n_0_0_34));
   NOR2_X1 i_0_0_49 (.A1(n_0_0_42), .A2(n_0_0_39), .ZN(n_0_0_35));
   INV_X1 i_0_0_50 (.A(n_0_0_37), .ZN(n_0_0_36));
   OAI22_X1 i_0_0_51 (.A1(n_0_0_54), .A2(first_operand[15]), .B1(n_0_0_44), 
      .B2(n_0_0_38), .ZN(n_0_0_37));
   OAI21_X1 i_0_0_52 (.A(n_0_0_43), .B1(n_0_0_51), .B2(n_0_0_39), .ZN(n_0_0_38));
   NOR2_X1 i_0_0_53 (.A1(n_0_0_53), .A2(first_operand[14]), .ZN(n_0_0_39));
   INV_X1 i_0_0_54 (.A(n_0_0_43), .ZN(n_0_0_42));
   NAND2_X1 i_0_0_57 (.A1(n_0_0_53), .A2(first_operand[14]), .ZN(n_0_0_43));
   INV_X1 i_0_0_58 (.A(n_0_0_45), .ZN(n_0_0_44));
   NAND2_X1 i_0_0_59 (.A1(n_0_0_54), .A2(first_operand[15]), .ZN(n_0_0_45));
   INV_X1 i_0_0_60 (.A(n_0_0_47), .ZN(n_0_0_46));
   NOR2_X1 i_0_0_61 (.A1(n_0_0_50), .A2(n_0_0_49), .ZN(n_0_0_47));
   INV_X1 i_0_0_62 (.A(n_0_0_49), .ZN(n_0_0_48));
   NOR2_X1 i_0_0_63 (.A1(n_0_0_52), .A2(first_operand[13]), .ZN(n_0_0_49));
   INV_X1 i_0_0_65 (.A(n_0_0_51), .ZN(n_0_0_50));
   NAND2_X1 i_0_0_66 (.A1(n_0_0_52), .A2(first_operand[13]), .ZN(n_0_0_51));
   INV_X1 i_0_0_67 (.A(second_operand[13]), .ZN(n_0_0_52));
   INV_X1 i_0_0_68 (.A(second_operand[14]), .ZN(n_0_0_53));
   INV_X1 i_0_0_69 (.A(second_operand[15]), .ZN(n_0_0_54));
   OAI21_X1 i_0_0_70 (.A(n_0_0_55), .B1(n_0_0_46), .B2(n_0_0_60), .ZN(out[12]));
   NAND2_X1 i_0_0_71 (.A1(n_0_0_46), .A2(n_0_0_56), .ZN(n_0_0_55));
   OAI22_X1 i_0_0_72 (.A1(n_0_0_65), .A2(n_0_0_57), .B1(n_0_0_31), .B2(n_0_0_59), 
      .ZN(n_0_0_56));
   AOI22_X1 i_0_0_73 (.A1(n_0_0_66), .A2(temp_result_wire[15]), .B1(n_0_0_28), 
      .B2(temp_result_wire[19]), .ZN(n_0_0_57));
   INV_X1 i_0_0_74 (.A(n_0_0_59), .ZN(n_0_0_58));
   OAI22_X1 i_0_0_75 (.A1(n_0_0_28), .A2(temp_result_wire[13]), .B1(n_0_0_66), 
      .B2(temp_result_wire[17]), .ZN(n_0_0_59));
   INV_X1 i_0_0_76 (.A(n_0_0_61), .ZN(n_0_0_60));
   AOI22_X1 i_0_0_77 (.A1(n_0_0_31), .A2(n_0_0_62), .B1(n_0_0_65), .B2(n_0_0_64), 
      .ZN(n_0_0_61));
   OAI22_X1 i_0_0_78 (.A1(n_0_0_28), .A2(temp_result_wire[14]), .B1(n_0_0_66), 
      .B2(temp_result_wire[18]), .ZN(n_0_0_62));
   INV_X1 i_0_0_79 (.A(n_0_0_64), .ZN(n_0_0_63));
   OAI22_X1 i_0_0_80 (.A1(n_0_0_28), .A2(temp_result_wire[12]), .B1(n_0_0_66), 
      .B2(temp_result_wire[16]), .ZN(n_0_0_64));
   INV_X1 i_0_0_81 (.A(n_0_0_31), .ZN(n_0_0_65));
   INV_X1 i_0_0_82 (.A(n_0_0_28), .ZN(n_0_0_66));
endmodule

module booth_16bit_multiplier(A, B, product);
   input [15:0]A;
   input [15:0]B;
   output [31:0]product;

   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_215;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_14;
   wire n_1_0;
   wire n_1_1;
   wire n_1_15;
   wire n_1_16;
   wire n_1_17;
   wire n_1_18;
   wire n_1_19;
   wire n_1_20;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;
   wire n_1_28;
   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire n_1_60;
   wire n_1_61;
   wire n_1_62;
   wire n_1_63;
   wire n_1_64;
   wire n_1_65;
   wire n_1_66;
   wire n_1_67;
   wire n_1_68;
   wire n_1_69;
   wire n_1_70;
   wire n_1_71;
   wire n_1_72;
   wire n_1_73;
   wire n_1_74;
   wire n_1_75;
   wire n_1_76;
   wire n_1_77;
   wire n_1_78;
   wire n_1_79;
   wire n_1_80;
   wire n_1_81;
   wire n_1_82;
   wire n_1_83;
   wire n_1_84;
   wire n_1_85;
   wire n_1_86;
   wire n_1_87;
   wire n_1_88;
   wire n_1_89;
   wire n_1_90;
   wire n_1_91;
   wire n_1_92;
   wire n_1_93;
   wire n_1_94;
   wire n_1_95;
   wire n_1_96;
   wire n_1_97;
   wire n_1_98;
   wire n_1_99;
   wire n_1_100;
   wire n_1_101;
   wire n_1_102;
   wire n_1_103;
   wire n_1_104;
   wire n_1_105;
   wire n_1_106;
   wire n_1_107;
   wire n_1_108;
   wire n_1_109;
   wire n_1_110;
   wire n_1_111;
   wire n_1_112;
   wire n_1_113;
   wire n_1_114;
   wire n_1_115;
   wire n_1_116;
   wire n_1_117;
   wire n_1_118;
   wire n_1_119;
   wire n_1_120;
   wire n_1_121;
   wire n_1_122;
   wire n_1_123;
   wire n_1_124;
   wire n_1_125;
   wire n_1_126;
   wire n_1_127;
   wire n_1_128;
   wire n_1_129;
   wire n_1_130;
   wire n_1_131;
   wire n_1_132;
   wire n_1_133;
   wire n_1_134;
   wire n_1_135;
   wire n_1_136;
   wire n_1_137;
   wire n_1_138;
   wire n_1_139;
   wire n_1_140;
   wire n_1_141;
   wire n_1_142;
   wire n_1_143;
   wire n_1_144;
   wire n_1_145;
   wire n_1_146;
   wire n_1_147;
   wire n_1_148;
   wire n_1_149;
   wire n_1_150;
   wire n_1_151;
   wire n_1_152;
   wire n_1_153;
   wire n_1_154;
   wire n_1_155;
   wire n_1_156;
   wire n_1_157;
   wire n_1_158;
   wire n_1_159;
   wire n_1_160;
   wire n_1_161;
   wire n_1_162;
   wire n_1_163;
   wire n_1_164;
   wire n_1_165;
   wire n_1_166;
   wire n_1_167;
   wire n_1_168;
   wire n_1_169;
   wire n_1_170;
   wire n_1_171;
   wire n_1_172;
   wire n_1_173;
   wire n_1_174;
   wire n_1_175;

   datapath__0_1 i_2 (.B({B[15], uc_0, uc_1, uc_2, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({n_249, n_264, 
      n_263, n_262, n_261, n_260, n_259, n_258, n_257, n_256, n_255, n_254, 
      n_253, n_252, n_251, n_250}), .p_1({n_15, n_14, n_13, n_12, n_11, n_10, 
      n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0}));
   datapath__0_6 i_5 (.B({B[15], uc_3, uc_4, uc_5, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_6, n_248, n_247, 
      n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, n_238, n_237, 
      n_236, n_235, n_234}), .p_1({n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
      n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, n_16}));
   datapath__0_7 i_6 (.p_0({n_264, n_263, n_262, n_261, n_260, n_259, n_258, 
      n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, B[0]}), .p_1({uc_7, 
      n_248, n_247, n_246, n_245, n_244, n_243, n_242, n_241, n_240, n_239, 
      n_238, n_237, n_236, n_235, n_234}), .p_2({n_47, n_46, n_45, n_44, n_43, 
      n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32}));
   datapath__0_12 i_9 (.B({B[15], uc_8, uc_9, uc_10, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_11, n_233, 
      n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, n_224, n_223, 
      n_222, n_221, n_220, n_219}), .p_1({n_63, n_62, n_61, n_60, n_59, n_58, 
      n_57, n_56, n_55, n_54, n_53, n_52, n_51, n_50, n_49, n_48}));
   datapath__0_13 i_10 (.p_0({n_264, n_263, n_262, n_261, n_260, n_259, n_258, 
      n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, B[0]}), .p_1({
      uc_12, n_233, n_232, n_231, n_230, n_229, n_228, n_227, n_226, n_225, 
      n_224, n_223, n_222, n_221, n_220, n_219}), .p_2({n_79, n_78, n_77, n_76, 
      n_75, n_74, n_73, n_72, n_71, n_70, n_69, n_68, n_67, n_66, n_65, n_64}));
   datapath__0_18 i_13 (.B({B[15], uc_13, uc_14, uc_15, B[11], B[10], B[9], B[8], 
      B[7], B[6], B[5], B[4], B[3], B[2], B[1], B[0]}), .p_0({uc_16, n_218, 
      n_217, n_216, n_215, n_214, n_213, n_212, n_211, n_210, n_209, n_208, 
      n_207, n_206, n_205, n_204}), .p_1({n_95, n_94, n_93, n_92, n_91, n_90, 
      n_89, n_88, n_87, n_86, n_85, n_84, n_83, n_82, n_81, n_80}));
   datapath__0_19 i_14 (.p_0({n_264, n_263, n_262, n_261, n_260, n_259, n_258, 
      n_257, n_256, n_255, n_254, n_253, n_252, n_251, n_250, B[0]}), .p_1({
      uc_17, n_218, n_217, n_216, n_215, n_214, n_213, n_212, n_211, n_210, 
      n_209, n_208, n_207, n_206, n_205, n_204}), .p_2({n_111, n_110, n_109, 
      n_108, n_107, n_106, n_105, n_104, n_103, n_102, n_101, n_100, n_99, n_98, 
      n_97, n_96}));
   INV_X1 i_0_108 (.A(n_0_60), .ZN(product[12]));
   AOI222_X1 i_0_109 (.A1(n_438), .A2(n_0_79), .B1(n_438), .B2(n_0_78), .C1(
      n_112), .C2(n_0_77), .ZN(n_0_60));
   INV_X1 i_0_110 (.A(n_0_61), .ZN(product[13]));
   AOI222_X1 i_0_111 (.A1(n_424), .A2(n_0_79), .B1(n_417), .B2(n_0_78), .C1(
      n_113), .C2(n_0_77), .ZN(n_0_61));
   INV_X1 i_0_112 (.A(n_0_62), .ZN(product[14]));
   AOI222_X1 i_0_113 (.A1(n_425), .A2(n_0_79), .B1(n_418), .B2(n_0_78), .C1(
      n_114), .C2(n_0_77), .ZN(n_0_62));
   INV_X1 i_0_114 (.A(n_0_63), .ZN(product[15]));
   AOI222_X1 i_0_115 (.A1(n_426), .A2(n_0_79), .B1(n_419), .B2(n_0_78), .C1(
      n_115), .C2(n_0_77), .ZN(n_0_63));
   INV_X1 i_0_116 (.A(n_0_64), .ZN(product[16]));
   AOI222_X1 i_0_117 (.A1(n_427), .A2(n_0_79), .B1(n_420), .B2(n_0_78), .C1(
      n_116), .C2(n_0_77), .ZN(n_0_64));
   INV_X1 i_0_118 (.A(n_0_65), .ZN(product[17]));
   AOI222_X1 i_0_119 (.A1(n_428), .A2(n_0_79), .B1(n_421), .B2(n_0_78), .C1(
      n_117), .C2(n_0_77), .ZN(n_0_65));
   INV_X1 i_0_120 (.A(n_0_66), .ZN(product[18]));
   AOI222_X1 i_0_121 (.A1(n_429), .A2(n_0_79), .B1(n_422), .B2(n_0_78), .C1(
      n_118), .C2(n_0_77), .ZN(n_0_66));
   INV_X1 i_0_122 (.A(n_0_67), .ZN(product[19]));
   AOI222_X1 i_0_123 (.A1(n_430), .A2(n_0_79), .B1(n_423), .B2(n_0_78), .C1(
      n_119), .C2(n_0_77), .ZN(n_0_67));
   NOR2_X1 i_0_141 (.A1(n_0_79), .A2(n_0_78), .ZN(n_0_77));
   NOR2_X1 i_0_142 (.A1(A[15]), .A2(n_0_196), .ZN(n_0_78));
   NOR2_X1 i_0_143 (.A1(n_0_215), .A2(A[11]), .ZN(n_0_79));
   INV_X1 i_0_144 (.A(n_0_80), .ZN(product[11]));
   AOI222_X1 i_0_145 (.A1(n_437), .A2(n_0_98), .B1(n_437), .B2(n_0_99), .C1(
      n_120), .C2(n_0_97), .ZN(n_0_80));
   INV_X1 i_0_146 (.A(n_0_81), .ZN(n_112));
   AOI222_X1 i_0_147 (.A1(n_409), .A2(n_0_99), .B1(n_401), .B2(n_0_98), .C1(
      n_121), .C2(n_0_97), .ZN(n_0_81));
   INV_X1 i_0_148 (.A(n_0_82), .ZN(n_113));
   AOI222_X1 i_0_149 (.A1(n_410), .A2(n_0_99), .B1(n_402), .B2(n_0_98), .C1(
      n_122), .C2(n_0_97), .ZN(n_0_82));
   INV_X1 i_0_150 (.A(n_0_83), .ZN(n_114));
   AOI222_X1 i_0_151 (.A1(n_411), .A2(n_0_99), .B1(n_403), .B2(n_0_98), .C1(
      n_123), .C2(n_0_97), .ZN(n_0_83));
   INV_X1 i_0_152 (.A(n_0_84), .ZN(n_115));
   AOI222_X1 i_0_153 (.A1(n_412), .A2(n_0_99), .B1(n_404), .B2(n_0_98), .C1(
      n_124), .C2(n_0_97), .ZN(n_0_84));
   INV_X1 i_0_154 (.A(n_0_85), .ZN(n_116));
   AOI222_X1 i_0_155 (.A1(n_413), .A2(n_0_99), .B1(n_405), .B2(n_0_98), .C1(
      n_125), .C2(n_0_97), .ZN(n_0_85));
   INV_X1 i_0_156 (.A(n_0_86), .ZN(n_117));
   AOI222_X1 i_0_157 (.A1(n_414), .A2(n_0_99), .B1(n_406), .B2(n_0_98), .C1(
      n_126), .C2(n_0_97), .ZN(n_0_86));
   INV_X1 i_0_158 (.A(n_0_87), .ZN(n_118));
   AOI222_X1 i_0_159 (.A1(n_415), .A2(n_0_99), .B1(n_407), .B2(n_0_98), .C1(
      n_127), .C2(n_0_97), .ZN(n_0_87));
   INV_X1 i_0_160 (.A(n_0_88), .ZN(n_119));
   AOI222_X1 i_0_161 (.A1(n_416), .A2(n_0_99), .B1(n_408), .B2(n_0_98), .C1(
      n_128), .C2(n_0_97), .ZN(n_0_88));
   NOR2_X1 i_0_177 (.A1(n_0_99), .A2(n_0_98), .ZN(n_0_97));
   NOR2_X1 i_0_178 (.A1(A[11]), .A2(n_0_195), .ZN(n_0_98));
   NOR2_X1 i_0_179 (.A1(n_0_196), .A2(A[10]), .ZN(n_0_99));
   INV_X1 i_0_180 (.A(n_0_100), .ZN(product[10]));
   AOI222_X1 i_0_181 (.A1(n_436), .A2(n_0_118), .B1(n_436), .B2(n_0_119), 
      .C1(n_129), .C2(n_0_117), .ZN(n_0_100));
   INV_X1 i_0_182 (.A(n_0_101), .ZN(n_120));
   AOI222_X1 i_0_183 (.A1(n_383), .A2(n_0_118), .B1(n_392), .B2(n_0_119), 
      .C1(n_130), .C2(n_0_117), .ZN(n_0_101));
   INV_X1 i_0_184 (.A(n_0_102), .ZN(n_121));
   AOI222_X1 i_0_185 (.A1(n_384), .A2(n_0_118), .B1(n_393), .B2(n_0_119), 
      .C1(n_131), .C2(n_0_117), .ZN(n_0_102));
   INV_X1 i_0_186 (.A(n_0_103), .ZN(n_122));
   AOI222_X1 i_0_187 (.A1(n_394), .A2(n_0_119), .B1(n_385), .B2(n_0_118), 
      .C1(n_132), .C2(n_0_117), .ZN(n_0_103));
   INV_X1 i_0_188 (.A(n_0_104), .ZN(n_123));
   AOI222_X1 i_0_189 (.A1(n_395), .A2(n_0_119), .B1(n_386), .B2(n_0_118), 
      .C1(n_133), .C2(n_0_117), .ZN(n_0_104));
   INV_X1 i_0_190 (.A(n_0_105), .ZN(n_124));
   AOI222_X1 i_0_191 (.A1(n_396), .A2(n_0_119), .B1(n_387), .B2(n_0_118), 
      .C1(n_134), .C2(n_0_117), .ZN(n_0_105));
   INV_X1 i_0_192 (.A(n_0_106), .ZN(n_125));
   AOI222_X1 i_0_193 (.A1(n_397), .A2(n_0_119), .B1(n_388), .B2(n_0_118), 
      .C1(n_135), .C2(n_0_117), .ZN(n_0_106));
   INV_X1 i_0_194 (.A(n_0_107), .ZN(n_126));
   AOI222_X1 i_0_195 (.A1(n_398), .A2(n_0_119), .B1(n_389), .B2(n_0_118), 
      .C1(n_136), .C2(n_0_117), .ZN(n_0_107));
   INV_X1 i_0_196 (.A(n_0_108), .ZN(n_127));
   AOI222_X1 i_0_197 (.A1(n_399), .A2(n_0_119), .B1(n_390), .B2(n_0_118), 
      .C1(n_137), .C2(n_0_117), .ZN(n_0_108));
   INV_X1 i_0_198 (.A(n_0_109), .ZN(n_128));
   AOI222_X1 i_0_199 (.A1(n_400), .A2(n_0_119), .B1(n_391), .B2(n_0_118), 
      .C1(n_138), .C2(n_0_117), .ZN(n_0_109));
   NOR2_X1 i_0_213 (.A1(n_0_119), .A2(n_0_118), .ZN(n_0_117));
   NOR2_X1 i_0_214 (.A1(A[10]), .A2(n_0_194), .ZN(n_0_118));
   NOR2_X1 i_0_215 (.A1(n_0_195), .A2(A[9]), .ZN(n_0_119));
   INV_X1 i_0_216 (.A(n_0_120), .ZN(product[9]));
   AOI222_X1 i_0_217 (.A1(n_435), .A2(n_0_138), .B1(n_435), .B2(n_0_139), 
      .C1(n_139), .C2(n_0_137), .ZN(n_0_120));
   INV_X1 i_0_218 (.A(n_0_121), .ZN(n_129));
   AOI222_X1 i_0_219 (.A1(n_363), .A2(n_0_138), .B1(n_373), .B2(n_0_139), 
      .C1(n_140), .C2(n_0_137), .ZN(n_0_121));
   INV_X1 i_0_220 (.A(n_0_122), .ZN(n_130));
   AOI222_X1 i_0_221 (.A1(n_364), .A2(n_0_138), .B1(n_374), .B2(n_0_139), 
      .C1(n_141), .C2(n_0_137), .ZN(n_0_122));
   INV_X1 i_0_222 (.A(n_0_123), .ZN(n_131));
   AOI222_X1 i_0_223 (.A1(n_365), .A2(n_0_138), .B1(n_375), .B2(n_0_139), 
      .C1(n_142), .C2(n_0_137), .ZN(n_0_123));
   INV_X1 i_0_224 (.A(n_0_124), .ZN(n_132));
   AOI222_X1 i_0_225 (.A1(n_376), .A2(n_0_139), .B1(n_366), .B2(n_0_138), 
      .C1(n_143), .C2(n_0_137), .ZN(n_0_124));
   INV_X1 i_0_226 (.A(n_0_125), .ZN(n_133));
   AOI222_X1 i_0_227 (.A1(n_377), .A2(n_0_139), .B1(n_367), .B2(n_0_138), 
      .C1(n_144), .C2(n_0_137), .ZN(n_0_125));
   INV_X1 i_0_228 (.A(n_0_126), .ZN(n_134));
   AOI222_X1 i_0_229 (.A1(n_378), .A2(n_0_139), .B1(n_368), .B2(n_0_138), 
      .C1(n_145), .C2(n_0_137), .ZN(n_0_126));
   INV_X1 i_0_230 (.A(n_0_127), .ZN(n_135));
   AOI222_X1 i_0_231 (.A1(n_379), .A2(n_0_139), .B1(n_369), .B2(n_0_138), 
      .C1(n_146), .C2(n_0_137), .ZN(n_0_127));
   INV_X1 i_0_232 (.A(n_0_128), .ZN(n_136));
   AOI222_X1 i_0_233 (.A1(n_380), .A2(n_0_139), .B1(n_370), .B2(n_0_138), 
      .C1(n_147), .C2(n_0_137), .ZN(n_0_128));
   INV_X1 i_0_234 (.A(n_0_129), .ZN(n_137));
   AOI222_X1 i_0_235 (.A1(n_381), .A2(n_0_139), .B1(n_371), .B2(n_0_138), 
      .C1(n_148), .C2(n_0_137), .ZN(n_0_129));
   INV_X1 i_0_236 (.A(n_0_130), .ZN(n_138));
   AOI222_X1 i_0_237 (.A1(n_382), .A2(n_0_139), .B1(n_372), .B2(n_0_138), 
      .C1(n_149), .C2(n_0_137), .ZN(n_0_130));
   NOR2_X1 i_0_249 (.A1(n_0_139), .A2(n_0_138), .ZN(n_0_137));
   NOR2_X1 i_0_250 (.A1(A[9]), .A2(n_0_176), .ZN(n_0_138));
   NOR2_X1 i_0_251 (.A1(n_0_194), .A2(A[8]), .ZN(n_0_139));
   INV_X1 i_0_252 (.A(n_0_140), .ZN(product[8]));
   AOI222_X1 i_0_253 (.A1(n_434), .A2(n_0_158), .B1(n_434), .B2(n_0_159), 
      .C1(n_150), .C2(n_0_157), .ZN(n_0_140));
   INV_X1 i_0_254 (.A(n_0_141), .ZN(n_139));
   AOI222_X1 i_0_255 (.A1(n_341), .A2(n_0_158), .B1(n_352), .B2(n_0_159), 
      .C1(n_151), .C2(n_0_157), .ZN(n_0_141));
   INV_X1 i_0_256 (.A(n_0_142), .ZN(n_140));
   AOI222_X1 i_0_257 (.A1(n_342), .A2(n_0_158), .B1(n_353), .B2(n_0_159), 
      .C1(n_152), .C2(n_0_157), .ZN(n_0_142));
   INV_X1 i_0_258 (.A(n_0_143), .ZN(n_141));
   AOI222_X1 i_0_259 (.A1(n_343), .A2(n_0_158), .B1(n_354), .B2(n_0_159), 
      .C1(n_153), .C2(n_0_157), .ZN(n_0_143));
   INV_X1 i_0_260 (.A(n_0_144), .ZN(n_142));
   AOI222_X1 i_0_261 (.A1(n_344), .A2(n_0_158), .B1(n_355), .B2(n_0_159), 
      .C1(n_154), .C2(n_0_157), .ZN(n_0_144));
   INV_X1 i_0_262 (.A(n_0_145), .ZN(n_143));
   AOI222_X1 i_0_263 (.A1(n_356), .A2(n_0_159), .B1(n_345), .B2(n_0_158), 
      .C1(n_155), .C2(n_0_157), .ZN(n_0_145));
   INV_X1 i_0_264 (.A(n_0_146), .ZN(n_144));
   AOI222_X1 i_0_265 (.A1(n_357), .A2(n_0_159), .B1(n_346), .B2(n_0_158), 
      .C1(n_156), .C2(n_0_157), .ZN(n_0_146));
   INV_X1 i_0_266 (.A(n_0_147), .ZN(n_145));
   AOI222_X1 i_0_267 (.A1(n_358), .A2(n_0_159), .B1(n_347), .B2(n_0_158), 
      .C1(n_157), .C2(n_0_157), .ZN(n_0_147));
   INV_X1 i_0_268 (.A(n_0_148), .ZN(n_146));
   AOI222_X1 i_0_269 (.A1(n_359), .A2(n_0_159), .B1(n_348), .B2(n_0_158), 
      .C1(n_158), .C2(n_0_157), .ZN(n_0_148));
   INV_X1 i_0_270 (.A(n_0_149), .ZN(n_147));
   AOI222_X1 i_0_271 (.A1(n_360), .A2(n_0_159), .B1(n_349), .B2(n_0_158), 
      .C1(n_159), .C2(n_0_157), .ZN(n_0_149));
   INV_X1 i_0_272 (.A(n_0_150), .ZN(n_148));
   AOI222_X1 i_0_273 (.A1(n_361), .A2(n_0_159), .B1(n_350), .B2(n_0_158), 
      .C1(n_160), .C2(n_0_157), .ZN(n_0_150));
   INV_X1 i_0_274 (.A(n_0_151), .ZN(n_149));
   AOI222_X1 i_0_275 (.A1(n_362), .A2(n_0_159), .B1(n_351), .B2(n_0_158), 
      .C1(n_161), .C2(n_0_157), .ZN(n_0_151));
   NOR2_X1 i_0_285 (.A1(n_0_159), .A2(n_0_158), .ZN(n_0_157));
   NOR2_X1 i_0_286 (.A1(A[8]), .A2(n_0_175), .ZN(n_0_158));
   NOR2_X1 i_0_287 (.A1(n_0_176), .A2(A[7]), .ZN(n_0_159));
   INV_X1 i_0_288 (.A(n_0_160), .ZN(product[7]));
   AOI222_X1 i_0_289 (.A1(n_433), .A2(n_0_178), .B1(n_433), .B2(n_0_179), 
      .C1(n_162), .C2(n_0_177), .ZN(n_0_160));
   INV_X1 i_0_290 (.A(n_0_161), .ZN(n_150));
   AOI222_X1 i_0_291 (.A1(n_317), .A2(n_0_178), .B1(n_329), .B2(n_0_179), 
      .C1(n_163), .C2(n_0_177), .ZN(n_0_161));
   INV_X1 i_0_292 (.A(n_0_162), .ZN(n_151));
   AOI222_X1 i_0_293 (.A1(n_318), .A2(n_0_178), .B1(n_330), .B2(n_0_179), 
      .C1(n_164), .C2(n_0_177), .ZN(n_0_162));
   INV_X1 i_0_294 (.A(n_0_163), .ZN(n_152));
   AOI222_X1 i_0_295 (.A1(n_319), .A2(n_0_178), .B1(n_331), .B2(n_0_179), 
      .C1(n_165), .C2(n_0_177), .ZN(n_0_163));
   INV_X1 i_0_296 (.A(n_0_164), .ZN(n_153));
   AOI222_X1 i_0_297 (.A1(n_320), .A2(n_0_178), .B1(n_332), .B2(n_0_179), 
      .C1(n_166), .C2(n_0_177), .ZN(n_0_164));
   INV_X1 i_0_298 (.A(n_0_165), .ZN(n_154));
   AOI222_X1 i_0_299 (.A1(n_321), .A2(n_0_178), .B1(n_333), .B2(n_0_179), 
      .C1(n_167), .C2(n_0_177), .ZN(n_0_165));
   INV_X1 i_0_300 (.A(n_0_166), .ZN(n_155));
   AOI222_X1 i_0_301 (.A1(n_322), .A2(n_0_178), .B1(n_334), .B2(n_0_179), 
      .C1(n_168), .C2(n_0_177), .ZN(n_0_166));
   INV_X1 i_0_302 (.A(n_0_167), .ZN(n_156));
   AOI222_X1 i_0_303 (.A1(n_335), .A2(n_0_179), .B1(n_323), .B2(n_0_178), 
      .C1(n_169), .C2(n_0_177), .ZN(n_0_167));
   INV_X1 i_0_304 (.A(n_0_168), .ZN(n_157));
   AOI222_X1 i_0_305 (.A1(n_336), .A2(n_0_179), .B1(n_324), .B2(n_0_178), 
      .C1(n_170), .C2(n_0_177), .ZN(n_0_168));
   INV_X1 i_0_306 (.A(n_0_169), .ZN(n_158));
   AOI222_X1 i_0_307 (.A1(n_337), .A2(n_0_179), .B1(n_325), .B2(n_0_178), 
      .C1(n_171), .C2(n_0_177), .ZN(n_0_169));
   INV_X1 i_0_308 (.A(n_0_170), .ZN(n_159));
   AOI222_X1 i_0_309 (.A1(n_338), .A2(n_0_179), .B1(n_326), .B2(n_0_178), 
      .C1(n_172), .C2(n_0_177), .ZN(n_0_170));
   INV_X1 i_0_310 (.A(n_0_171), .ZN(n_160));
   AOI222_X1 i_0_311 (.A1(n_339), .A2(n_0_179), .B1(n_327), .B2(n_0_178), 
      .C1(n_173), .C2(n_0_177), .ZN(n_0_171));
   INV_X1 i_0_312 (.A(n_0_172), .ZN(n_161));
   AOI222_X1 i_0_313 (.A1(n_340), .A2(n_0_179), .B1(n_328), .B2(n_0_178), 
      .C1(n_174), .C2(n_0_177), .ZN(n_0_172));
   NOR2_X1 i_0_321 (.A1(n_0_179), .A2(n_0_178), .ZN(n_0_177));
   NOR2_X1 i_0_322 (.A1(A[7]), .A2(n_0_174), .ZN(n_0_178));
   NOR2_X1 i_0_323 (.A1(n_0_175), .A2(A[6]), .ZN(n_0_179));
   INV_X1 i_0_324 (.A(n_0_180), .ZN(product[6]));
   AOI222_X1 i_0_325 (.A1(n_432), .A2(n_0_198), .B1(n_432), .B2(n_0_199), 
      .C1(n_175), .C2(n_0_197), .ZN(n_0_180));
   INV_X1 i_0_326 (.A(n_0_181), .ZN(n_162));
   AOI222_X1 i_0_327 (.A1(n_291), .A2(n_0_198), .B1(n_304), .B2(n_0_199), 
      .C1(n_176), .C2(n_0_197), .ZN(n_0_181));
   INV_X1 i_0_328 (.A(n_0_182), .ZN(n_163));
   AOI222_X1 i_0_329 (.A1(n_292), .A2(n_0_198), .B1(n_305), .B2(n_0_199), 
      .C1(n_177), .C2(n_0_197), .ZN(n_0_182));
   INV_X1 i_0_330 (.A(n_0_183), .ZN(n_164));
   AOI222_X1 i_0_331 (.A1(n_293), .A2(n_0_198), .B1(n_306), .B2(n_0_199), 
      .C1(n_178), .C2(n_0_197), .ZN(n_0_183));
   INV_X1 i_0_332 (.A(n_0_184), .ZN(n_165));
   AOI222_X1 i_0_333 (.A1(n_294), .A2(n_0_198), .B1(n_307), .B2(n_0_199), 
      .C1(n_179), .C2(n_0_197), .ZN(n_0_184));
   INV_X1 i_0_334 (.A(n_0_185), .ZN(n_166));
   AOI222_X1 i_0_335 (.A1(n_295), .A2(n_0_198), .B1(n_308), .B2(n_0_199), 
      .C1(n_180), .C2(n_0_197), .ZN(n_0_185));
   INV_X1 i_0_336 (.A(n_0_186), .ZN(n_167));
   AOI222_X1 i_0_337 (.A1(n_296), .A2(n_0_198), .B1(n_309), .B2(n_0_199), 
      .C1(n_181), .C2(n_0_197), .ZN(n_0_186));
   INV_X1 i_0_338 (.A(n_0_187), .ZN(n_168));
   AOI222_X1 i_0_339 (.A1(n_297), .A2(n_0_198), .B1(n_310), .B2(n_0_199), 
      .C1(n_182), .C2(n_0_197), .ZN(n_0_187));
   INV_X1 i_0_340 (.A(n_0_188), .ZN(n_169));
   AOI222_X1 i_0_341 (.A1(n_311), .A2(n_0_199), .B1(n_298), .B2(n_0_198), 
      .C1(n_183), .C2(n_0_197), .ZN(n_0_188));
   INV_X1 i_0_342 (.A(n_0_189), .ZN(n_170));
   AOI222_X1 i_0_343 (.A1(n_312), .A2(n_0_199), .B1(n_299), .B2(n_0_198), 
      .C1(n_184), .C2(n_0_197), .ZN(n_0_189));
   INV_X1 i_0_344 (.A(n_0_190), .ZN(n_171));
   AOI222_X1 i_0_345 (.A1(n_313), .A2(n_0_199), .B1(n_300), .B2(n_0_198), 
      .C1(n_185), .C2(n_0_197), .ZN(n_0_190));
   INV_X1 i_0_346 (.A(n_0_191), .ZN(n_172));
   AOI222_X1 i_0_347 (.A1(n_314), .A2(n_0_199), .B1(n_301), .B2(n_0_198), 
      .C1(n_186), .C2(n_0_197), .ZN(n_0_191));
   INV_X1 i_0_348 (.A(n_0_192), .ZN(n_173));
   AOI222_X1 i_0_349 (.A1(n_315), .A2(n_0_199), .B1(n_302), .B2(n_0_198), 
      .C1(n_187), .C2(n_0_197), .ZN(n_0_192));
   INV_X1 i_0_350 (.A(n_0_193), .ZN(n_174));
   AOI222_X1 i_0_351 (.A1(n_316), .A2(n_0_199), .B1(n_303), .B2(n_0_198), 
      .C1(n_188), .C2(n_0_197), .ZN(n_0_193));
   NOR2_X1 i_0_357 (.A1(n_0_199), .A2(n_0_198), .ZN(n_0_197));
   NOR2_X1 i_0_358 (.A1(A[6]), .A2(n_0_173), .ZN(n_0_198));
   NOR2_X1 i_0_359 (.A1(n_0_174), .A2(A[5]), .ZN(n_0_199));
   INV_X1 i_0_360 (.A(n_0_200), .ZN(product[5]));
   AOI222_X1 i_0_361 (.A1(n_431), .A2(n_0_218), .B1(n_431), .B2(n_0_219), 
      .C1(n_189), .C2(n_0_217), .ZN(n_0_200));
   INV_X1 i_0_362 (.A(n_0_201), .ZN(n_175));
   AOI222_X1 i_0_363 (.A1(n_265), .A2(n_0_218), .B1(n_278), .B2(n_0_219), 
      .C1(n_190), .C2(n_0_217), .ZN(n_0_201));
   INV_X1 i_0_364 (.A(n_0_202), .ZN(n_176));
   AOI222_X1 i_0_365 (.A1(n_266), .A2(n_0_218), .B1(n_279), .B2(n_0_219), 
      .C1(n_191), .C2(n_0_217), .ZN(n_0_202));
   INV_X1 i_0_366 (.A(n_0_203), .ZN(n_177));
   AOI222_X1 i_0_367 (.A1(n_267), .A2(n_0_218), .B1(n_280), .B2(n_0_219), 
      .C1(n_192), .C2(n_0_217), .ZN(n_0_203));
   INV_X1 i_0_368 (.A(n_0_204), .ZN(n_178));
   AOI222_X1 i_0_369 (.A1(n_268), .A2(n_0_218), .B1(n_281), .B2(n_0_219), 
      .C1(n_193), .C2(n_0_217), .ZN(n_0_204));
   INV_X1 i_0_370 (.A(n_0_205), .ZN(n_179));
   AOI222_X1 i_0_371 (.A1(n_269), .A2(n_0_218), .B1(n_282), .B2(n_0_219), 
      .C1(n_194), .C2(n_0_217), .ZN(n_0_205));
   INV_X1 i_0_372 (.A(n_0_206), .ZN(n_180));
   AOI222_X1 i_0_373 (.A1(n_270), .A2(n_0_218), .B1(n_283), .B2(n_0_219), 
      .C1(n_195), .C2(n_0_217), .ZN(n_0_206));
   INV_X1 i_0_374 (.A(n_0_207), .ZN(n_181));
   AOI222_X1 i_0_375 (.A1(n_271), .A2(n_0_218), .B1(n_284), .B2(n_0_219), 
      .C1(n_196), .C2(n_0_217), .ZN(n_0_207));
   INV_X1 i_0_376 (.A(n_0_208), .ZN(n_182));
   AOI222_X1 i_0_377 (.A1(n_272), .A2(n_0_218), .B1(n_285), .B2(n_0_219), 
      .C1(n_197), .C2(n_0_217), .ZN(n_0_208));
   INV_X1 i_0_378 (.A(n_0_209), .ZN(n_183));
   AOI222_X1 i_0_379 (.A1(n_286), .A2(n_0_219), .B1(n_273), .B2(n_0_218), 
      .C1(n_198), .C2(n_0_217), .ZN(n_0_209));
   INV_X1 i_0_380 (.A(n_0_210), .ZN(n_184));
   AOI222_X1 i_0_381 (.A1(n_287), .A2(n_0_219), .B1(n_274), .B2(n_0_218), 
      .C1(n_199), .C2(n_0_217), .ZN(n_0_210));
   INV_X1 i_0_382 (.A(n_0_211), .ZN(n_185));
   AOI222_X1 i_0_383 (.A1(n_288), .A2(n_0_219), .B1(n_275), .B2(n_0_218), 
      .C1(n_200), .C2(n_0_217), .ZN(n_0_211));
   INV_X1 i_0_384 (.A(n_0_212), .ZN(n_186));
   AOI222_X1 i_0_385 (.A1(n_289), .A2(n_0_219), .B1(n_276), .B2(n_0_218), 
      .C1(n_201), .C2(n_0_217), .ZN(n_0_212));
   INV_X1 i_0_386 (.A(n_0_213), .ZN(n_187));
   AOI222_X1 i_0_387 (.A1(n_290), .A2(n_0_219), .B1(n_277), .B2(n_0_218), 
      .C1(n_202), .C2(n_0_217), .ZN(n_0_213));
   INV_X1 i_0_388 (.A(n_0_214), .ZN(n_188));
   AOI221_X1 i_0_389 (.A(n_0_216), .B1(n_440), .B2(n_0_218), .C1(n_439), 
      .C2(n_0_219), .ZN(n_0_214));
   AND2_X1 i_0_392 (.A1(n_203), .A2(n_0_217), .ZN(n_0_216));
   NOR2_X1 i_0_393 (.A1(n_0_219), .A2(n_0_218), .ZN(n_0_217));
   NOR2_X1 i_0_394 (.A1(A[5]), .A2(n_0_156), .ZN(n_0_218));
   NOR2_X1 i_0_395 (.A1(n_0_173), .A2(A[4]), .ZN(n_0_219));
   INV_X1 i_0_396 (.A(n_0_220), .ZN(product[4]));
   AOI222_X1 i_0_397 (.A1(n_80), .A2(n_0_2), .B1(n_96), .B2(n_0_3), .C1(n_204), 
      .C2(n_0_1), .ZN(n_0_220));
   INV_X1 i_0_398 (.A(n_0_221), .ZN(n_189));
   AOI222_X1 i_0_399 (.A1(n_81), .A2(n_0_2), .B1(n_97), .B2(n_0_3), .C1(n_205), 
      .C2(n_0_1), .ZN(n_0_221));
   INV_X1 i_0_400 (.A(n_0_222), .ZN(n_190));
   AOI222_X1 i_0_401 (.A1(n_82), .A2(n_0_2), .B1(n_98), .B2(n_0_3), .C1(n_206), 
      .C2(n_0_1), .ZN(n_0_222));
   INV_X1 i_0_402 (.A(n_0_223), .ZN(n_191));
   AOI222_X1 i_0_403 (.A1(n_83), .A2(n_0_2), .B1(n_99), .B2(n_0_3), .C1(n_207), 
      .C2(n_0_1), .ZN(n_0_223));
   INV_X1 i_0_404 (.A(n_0_224), .ZN(n_192));
   AOI222_X1 i_0_405 (.A1(n_84), .A2(n_0_2), .B1(n_100), .B2(n_0_3), .C1(n_208), 
      .C2(n_0_1), .ZN(n_0_224));
   INV_X1 i_0_406 (.A(n_0_225), .ZN(n_193));
   AOI222_X1 i_0_407 (.A1(n_85), .A2(n_0_2), .B1(n_101), .B2(n_0_3), .C1(n_209), 
      .C2(n_0_1), .ZN(n_0_225));
   INV_X1 i_0_408 (.A(n_0_226), .ZN(n_194));
   AOI222_X1 i_0_409 (.A1(n_86), .A2(n_0_2), .B1(n_102), .B2(n_0_3), .C1(n_210), 
      .C2(n_0_1), .ZN(n_0_226));
   INV_X1 i_0_410 (.A(n_0_227), .ZN(n_195));
   AOI222_X1 i_0_411 (.A1(n_87), .A2(n_0_2), .B1(n_103), .B2(n_0_3), .C1(n_211), 
      .C2(n_0_1), .ZN(n_0_227));
   INV_X1 i_0_412 (.A(n_0_228), .ZN(n_196));
   AOI222_X1 i_0_413 (.A1(n_88), .A2(n_0_2), .B1(n_104), .B2(n_0_3), .C1(n_212), 
      .C2(n_0_1), .ZN(n_0_228));
   INV_X1 i_0_414 (.A(n_0_229), .ZN(n_197));
   AOI222_X1 i_0_415 (.A1(n_89), .A2(n_0_2), .B1(n_105), .B2(n_0_3), .C1(n_213), 
      .C2(n_0_1), .ZN(n_0_229));
   INV_X1 i_0_416 (.A(n_0_230), .ZN(n_198));
   AOI222_X1 i_0_417 (.A1(n_90), .A2(n_0_2), .B1(n_106), .B2(n_0_3), .C1(n_214), 
      .C2(n_0_1), .ZN(n_0_230));
   INV_X1 i_0_418 (.A(n_0_231), .ZN(n_199));
   AOI222_X1 i_0_419 (.A1(n_107), .A2(n_0_3), .B1(n_91), .B2(n_0_2), .C1(n_215), 
      .C2(n_0_1), .ZN(n_0_231));
   INV_X1 i_0_420 (.A(n_0_232), .ZN(n_200));
   AOI222_X1 i_0_421 (.A1(n_108), .A2(n_0_3), .B1(n_92), .B2(n_0_2), .C1(n_216), 
      .C2(n_0_1), .ZN(n_0_232));
   INV_X1 i_0_422 (.A(n_0_233), .ZN(n_201));
   AOI222_X1 i_0_423 (.A1(n_109), .A2(n_0_3), .B1(n_93), .B2(n_0_2), .C1(n_217), 
      .C2(n_0_1), .ZN(n_0_233));
   INV_X1 i_0_424 (.A(n_0_234), .ZN(n_202));
   AOI221_X1 i_0_425 (.A(n_0_0), .B1(n_94), .B2(n_0_2), .C1(n_110), .C2(n_0_3), 
      .ZN(n_0_234));
   INV_X1 i_0_426 (.A(n_0_235), .ZN(n_203));
   AOI221_X1 i_0_427 (.A(n_0_0), .B1(n_95), .B2(n_0_2), .C1(n_111), .C2(n_0_3), 
      .ZN(n_0_235));
   AND2_X1 i_0_428 (.A1(n_218), .A2(n_0_1), .ZN(n_0_0));
   NOR2_X1 i_0_429 (.A1(n_0_3), .A2(n_0_2), .ZN(n_0_1));
   NOR2_X1 i_0_430 (.A1(A[4]), .A2(n_0_155), .ZN(n_0_2));
   NOR2_X1 i_0_431 (.A1(n_0_156), .A2(A[3]), .ZN(n_0_3));
   INV_X1 i_0_432 (.A(n_0_4), .ZN(product[3]));
   AOI222_X1 i_0_433 (.A1(n_48), .A2(n_0_22), .B1(n_64), .B2(n_0_23), .C1(n_219), 
      .C2(n_0_21), .ZN(n_0_4));
   INV_X1 i_0_434 (.A(n_0_5), .ZN(n_204));
   AOI222_X1 i_0_435 (.A1(n_49), .A2(n_0_22), .B1(n_65), .B2(n_0_23), .C1(n_220), 
      .C2(n_0_21), .ZN(n_0_5));
   INV_X1 i_0_436 (.A(n_0_6), .ZN(n_205));
   AOI222_X1 i_0_437 (.A1(n_50), .A2(n_0_22), .B1(n_66), .B2(n_0_23), .C1(n_221), 
      .C2(n_0_21), .ZN(n_0_6));
   INV_X1 i_0_438 (.A(n_0_7), .ZN(n_206));
   AOI222_X1 i_0_439 (.A1(n_51), .A2(n_0_22), .B1(n_67), .B2(n_0_23), .C1(n_222), 
      .C2(n_0_21), .ZN(n_0_7));
   INV_X1 i_0_440 (.A(n_0_8), .ZN(n_207));
   AOI222_X1 i_0_441 (.A1(n_52), .A2(n_0_22), .B1(n_68), .B2(n_0_23), .C1(n_223), 
      .C2(n_0_21), .ZN(n_0_8));
   INV_X1 i_0_442 (.A(n_0_9), .ZN(n_208));
   AOI222_X1 i_0_443 (.A1(n_53), .A2(n_0_22), .B1(n_69), .B2(n_0_23), .C1(n_224), 
      .C2(n_0_21), .ZN(n_0_9));
   INV_X1 i_0_444 (.A(n_0_10), .ZN(n_209));
   AOI222_X1 i_0_445 (.A1(n_54), .A2(n_0_22), .B1(n_70), .B2(n_0_23), .C1(n_225), 
      .C2(n_0_21), .ZN(n_0_10));
   INV_X1 i_0_446 (.A(n_0_11), .ZN(n_210));
   AOI222_X1 i_0_447 (.A1(n_55), .A2(n_0_22), .B1(n_71), .B2(n_0_23), .C1(n_226), 
      .C2(n_0_21), .ZN(n_0_11));
   INV_X1 i_0_448 (.A(n_0_12), .ZN(n_211));
   AOI222_X1 i_0_449 (.A1(n_56), .A2(n_0_22), .B1(n_72), .B2(n_0_23), .C1(n_227), 
      .C2(n_0_21), .ZN(n_0_12));
   INV_X1 i_0_450 (.A(n_0_13), .ZN(n_212));
   AOI222_X1 i_0_451 (.A1(n_57), .A2(n_0_22), .B1(n_73), .B2(n_0_23), .C1(n_228), 
      .C2(n_0_21), .ZN(n_0_13));
   INV_X1 i_0_452 (.A(n_0_14), .ZN(n_213));
   AOI222_X1 i_0_453 (.A1(n_58), .A2(n_0_22), .B1(n_74), .B2(n_0_23), .C1(n_229), 
      .C2(n_0_21), .ZN(n_0_14));
   INV_X1 i_0_454 (.A(n_0_15), .ZN(n_214));
   AOI222_X1 i_0_455 (.A1(n_59), .A2(n_0_22), .B1(n_75), .B2(n_0_23), .C1(n_230), 
      .C2(n_0_21), .ZN(n_0_15));
   INV_X1 i_0_456 (.A(n_0_16), .ZN(n_215));
   AOI222_X1 i_0_457 (.A1(n_76), .A2(n_0_23), .B1(n_60), .B2(n_0_22), .C1(n_231), 
      .C2(n_0_21), .ZN(n_0_16));
   INV_X1 i_0_458 (.A(n_0_17), .ZN(n_216));
   AOI222_X1 i_0_459 (.A1(n_77), .A2(n_0_23), .B1(n_61), .B2(n_0_22), .C1(n_232), 
      .C2(n_0_21), .ZN(n_0_17));
   INV_X1 i_0_460 (.A(n_0_18), .ZN(n_217));
   AOI221_X1 i_0_461 (.A(n_0_20), .B1(n_62), .B2(n_0_22), .C1(n_78), .C2(n_0_23), 
      .ZN(n_0_18));
   INV_X1 i_0_462 (.A(n_0_19), .ZN(n_218));
   AOI221_X1 i_0_463 (.A(n_0_20), .B1(n_63), .B2(n_0_22), .C1(n_79), .C2(n_0_23), 
      .ZN(n_0_19));
   AND2_X1 i_0_464 (.A1(n_233), .A2(n_0_21), .ZN(n_0_20));
   NOR2_X1 i_0_465 (.A1(n_0_23), .A2(n_0_22), .ZN(n_0_21));
   NOR2_X1 i_0_466 (.A1(A[3]), .A2(n_0_154), .ZN(n_0_22));
   NOR2_X1 i_0_467 (.A1(n_0_155), .A2(A[2]), .ZN(n_0_23));
   INV_X1 i_0_468 (.A(n_0_24), .ZN(product[2]));
   AOI222_X1 i_0_469 (.A1(n_16), .A2(n_0_42), .B1(n_32), .B2(n_0_43), .C1(n_234), 
      .C2(n_0_41), .ZN(n_0_24));
   INV_X1 i_0_470 (.A(n_0_25), .ZN(n_219));
   AOI222_X1 i_0_471 (.A1(n_17), .A2(n_0_42), .B1(n_33), .B2(n_0_43), .C1(n_235), 
      .C2(n_0_41), .ZN(n_0_25));
   INV_X1 i_0_472 (.A(n_0_26), .ZN(n_220));
   AOI222_X1 i_0_473 (.A1(n_18), .A2(n_0_42), .B1(n_34), .B2(n_0_43), .C1(n_236), 
      .C2(n_0_41), .ZN(n_0_26));
   INV_X1 i_0_474 (.A(n_0_27), .ZN(n_221));
   AOI222_X1 i_0_475 (.A1(n_19), .A2(n_0_42), .B1(n_35), .B2(n_0_43), .C1(n_237), 
      .C2(n_0_41), .ZN(n_0_27));
   INV_X1 i_0_476 (.A(n_0_28), .ZN(n_222));
   AOI222_X1 i_0_477 (.A1(n_20), .A2(n_0_42), .B1(n_36), .B2(n_0_43), .C1(n_238), 
      .C2(n_0_41), .ZN(n_0_28));
   INV_X1 i_0_478 (.A(n_0_29), .ZN(n_223));
   AOI222_X1 i_0_479 (.A1(n_21), .A2(n_0_42), .B1(n_37), .B2(n_0_43), .C1(n_239), 
      .C2(n_0_41), .ZN(n_0_29));
   INV_X1 i_0_480 (.A(n_0_30), .ZN(n_224));
   AOI222_X1 i_0_481 (.A1(n_22), .A2(n_0_42), .B1(n_38), .B2(n_0_43), .C1(n_240), 
      .C2(n_0_41), .ZN(n_0_30));
   INV_X1 i_0_482 (.A(n_0_31), .ZN(n_225));
   AOI222_X1 i_0_483 (.A1(n_23), .A2(n_0_42), .B1(n_39), .B2(n_0_43), .C1(n_241), 
      .C2(n_0_41), .ZN(n_0_31));
   INV_X1 i_0_484 (.A(n_0_32), .ZN(n_226));
   AOI222_X1 i_0_485 (.A1(n_24), .A2(n_0_42), .B1(n_40), .B2(n_0_43), .C1(n_242), 
      .C2(n_0_41), .ZN(n_0_32));
   INV_X1 i_0_486 (.A(n_0_33), .ZN(n_227));
   AOI222_X1 i_0_487 (.A1(n_25), .A2(n_0_42), .B1(n_41), .B2(n_0_43), .C1(n_243), 
      .C2(n_0_41), .ZN(n_0_33));
   INV_X1 i_0_488 (.A(n_0_34), .ZN(n_228));
   AOI222_X1 i_0_489 (.A1(n_26), .A2(n_0_42), .B1(n_42), .B2(n_0_43), .C1(n_244), 
      .C2(n_0_41), .ZN(n_0_34));
   INV_X1 i_0_490 (.A(n_0_35), .ZN(n_229));
   AOI222_X1 i_0_491 (.A1(n_27), .A2(n_0_42), .B1(n_43), .B2(n_0_43), .C1(n_245), 
      .C2(n_0_41), .ZN(n_0_35));
   INV_X1 i_0_492 (.A(n_0_36), .ZN(n_230));
   AOI222_X1 i_0_493 (.A1(n_28), .A2(n_0_42), .B1(n_44), .B2(n_0_43), .C1(n_246), 
      .C2(n_0_41), .ZN(n_0_36));
   INV_X1 i_0_494 (.A(n_0_37), .ZN(n_231));
   AOI222_X1 i_0_495 (.A1(n_45), .A2(n_0_43), .B1(n_29), .B2(n_0_42), .C1(n_247), 
      .C2(n_0_41), .ZN(n_0_37));
   INV_X1 i_0_496 (.A(n_0_38), .ZN(n_232));
   AOI221_X1 i_0_497 (.A(n_0_40), .B1(n_30), .B2(n_0_42), .C1(n_46), .C2(n_0_43), 
      .ZN(n_0_38));
   INV_X1 i_0_498 (.A(n_0_39), .ZN(n_233));
   AOI221_X1 i_0_499 (.A(n_0_40), .B1(n_31), .B2(n_0_42), .C1(n_47), .C2(n_0_43), 
      .ZN(n_0_39));
   AND2_X1 i_0_500 (.A1(n_248), .A2(n_0_41), .ZN(n_0_40));
   NOR2_X1 i_0_501 (.A1(n_0_43), .A2(n_0_42), .ZN(n_0_41));
   NOR2_X1 i_0_502 (.A1(A[2]), .A2(n_0_153), .ZN(n_0_42));
   NOR2_X1 i_0_503 (.A1(n_0_154), .A2(A[1]), .ZN(n_0_43));
   INV_X1 i_0_504 (.A(n_0_44), .ZN(product[1]));
   AOI222_X1 i_0_505 (.A1(n_0), .A2(n_0_70), .B1(B[0]), .B2(n_0_59), .C1(n_250), 
      .C2(n_0_68), .ZN(n_0_44));
   INV_X1 i_0_506 (.A(n_0_45), .ZN(n_234));
   AOI222_X1 i_0_507 (.A1(n_1), .A2(n_0_70), .B1(n_250), .B2(n_0_59), .C1(n_251), 
      .C2(n_0_68), .ZN(n_0_45));
   INV_X1 i_0_508 (.A(n_0_46), .ZN(n_235));
   AOI222_X1 i_0_509 (.A1(n_2), .A2(n_0_70), .B1(n_251), .B2(n_0_59), .C1(n_252), 
      .C2(n_0_68), .ZN(n_0_46));
   INV_X1 i_0_510 (.A(n_0_47), .ZN(n_236));
   AOI222_X1 i_0_511 (.A1(n_252), .A2(n_0_59), .B1(n_3), .B2(n_0_70), .C1(n_253), 
      .C2(n_0_68), .ZN(n_0_47));
   INV_X1 i_0_512 (.A(n_0_48), .ZN(n_237));
   AOI222_X1 i_0_513 (.A1(n_253), .A2(n_0_59), .B1(n_4), .B2(n_0_70), .C1(n_254), 
      .C2(n_0_68), .ZN(n_0_48));
   INV_X1 i_0_514 (.A(n_0_49), .ZN(n_238));
   AOI222_X1 i_0_515 (.A1(n_5), .A2(n_0_70), .B1(n_254), .B2(n_0_59), .C1(n_255), 
      .C2(n_0_68), .ZN(n_0_49));
   INV_X1 i_0_516 (.A(n_0_50), .ZN(n_239));
   AOI222_X1 i_0_517 (.A1(n_6), .A2(n_0_70), .B1(n_255), .B2(n_0_59), .C1(n_256), 
      .C2(n_0_68), .ZN(n_0_50));
   INV_X1 i_0_518 (.A(n_0_51), .ZN(n_240));
   AOI222_X1 i_0_519 (.A1(n_7), .A2(n_0_70), .B1(n_256), .B2(n_0_59), .C1(n_257), 
      .C2(n_0_68), .ZN(n_0_51));
   INV_X1 i_0_520 (.A(n_0_52), .ZN(n_241));
   AOI222_X1 i_0_521 (.A1(n_8), .A2(n_0_70), .B1(n_257), .B2(n_0_59), .C1(n_258), 
      .C2(n_0_68), .ZN(n_0_52));
   INV_X1 i_0_522 (.A(n_0_53), .ZN(n_242));
   AOI222_X1 i_0_523 (.A1(n_9), .A2(n_0_70), .B1(n_258), .B2(n_0_59), .C1(n_259), 
      .C2(n_0_68), .ZN(n_0_53));
   INV_X1 i_0_524 (.A(n_0_54), .ZN(n_243));
   AOI222_X1 i_0_525 (.A1(n_259), .A2(n_0_59), .B1(n_10), .B2(n_0_70), .C1(n_260), 
      .C2(n_0_68), .ZN(n_0_54));
   INV_X1 i_0_526 (.A(n_0_55), .ZN(n_244));
   AOI222_X1 i_0_527 (.A1(n_260), .A2(n_0_59), .B1(n_11), .B2(n_0_70), .C1(n_261), 
      .C2(n_0_68), .ZN(n_0_55));
   INV_X1 i_0_528 (.A(n_0_56), .ZN(n_245));
   AOI222_X1 i_0_529 (.A1(n_12), .A2(n_0_70), .B1(n_261), .B2(n_0_59), .C1(n_262), 
      .C2(n_0_68), .ZN(n_0_56));
   INV_X1 i_0_530 (.A(n_0_57), .ZN(n_246));
   AOI222_X1 i_0_531 (.A1(n_13), .A2(n_0_70), .B1(n_262), .B2(n_0_59), .C1(n_263), 
      .C2(n_0_68), .ZN(n_0_57));
   INV_X1 i_0_532 (.A(n_0_58), .ZN(n_247));
   AOI222_X1 i_0_533 (.A1(n_263), .A2(n_0_59), .B1(n_14), .B2(n_0_70), .C1(n_264), 
      .C2(n_0_68), .ZN(n_0_58));
   NOR2_X1 i_0_534 (.A1(n_0_153), .A2(A[0]), .ZN(n_0_59));
   NOR2_X1 i_0_535 (.A1(n_0_152), .A2(n_0_70), .ZN(n_0_68));
   INV_X1 i_0_536 (.A(n_0_69), .ZN(n_248));
   AOI22_X1 i_0_537 (.A1(n_15), .A2(n_0_70), .B1(A[1]), .B2(n_264), .ZN(n_0_69));
   NOR2_X1 i_0_538 (.A1(A[1]), .A2(n_0_152), .ZN(n_0_70));
   AND2_X1 i_0_539 (.A1(B[0]), .A2(A[0]), .ZN(product[0]));
   AND2_X1 i_0_540 (.A1(A[0]), .A2(n_264), .ZN(n_249));
   AOI21_X1 i_0_541 (.A(n_0_136), .B1(B[1]), .B2(B[0]), .ZN(n_250));
   AOI21_X1 i_0_542 (.A(n_0_134), .B1(B[2]), .B2(n_0_135), .ZN(n_251));
   AOI21_X1 i_0_543 (.A(n_0_132), .B1(B[3]), .B2(n_0_133), .ZN(n_252));
   AOI21_X1 i_0_544 (.A(n_0_116), .B1(B[4]), .B2(n_0_131), .ZN(n_253));
   AOI21_X1 i_0_545 (.A(n_0_114), .B1(B[5]), .B2(n_0_115), .ZN(n_254));
   AOI21_X1 i_0_546 (.A(n_0_112), .B1(B[6]), .B2(n_0_113), .ZN(n_255));
   AOI21_X1 i_0_547 (.A(n_0_110), .B1(B[7]), .B2(n_0_111), .ZN(n_256));
   AOI21_X1 i_0_548 (.A(n_0_95), .B1(B[8]), .B2(n_0_96), .ZN(n_257));
   AOI21_X1 i_0_549 (.A(n_0_93), .B1(B[9]), .B2(n_0_94), .ZN(n_258));
   AOI21_X1 i_0_550 (.A(n_0_91), .B1(B[10]), .B2(n_0_92), .ZN(n_259));
   AOI21_X1 i_0_551 (.A(n_0_89), .B1(B[11]), .B2(n_0_90), .ZN(n_260));
   AOI21_X1 i_0_552 (.A(n_0_75), .B1(B[15]), .B2(n_0_76), .ZN(n_261));
   AOI21_X1 i_0_553 (.A(n_0_73), .B1(B[15]), .B2(n_0_74), .ZN(n_262));
   AOI21_X1 i_0_554 (.A(n_0_71), .B1(B[15]), .B2(n_0_72), .ZN(n_263));
   XNOR2_X1 i_0_555 (.A(B[15]), .B(n_0_71), .ZN(n_264));
   NOR2_X1 i_0_556 (.A1(B[15]), .A2(n_0_72), .ZN(n_0_71));
   INV_X1 i_0_557 (.A(n_0_73), .ZN(n_0_72));
   NOR2_X1 i_0_558 (.A1(B[15]), .A2(n_0_74), .ZN(n_0_73));
   INV_X1 i_0_559 (.A(n_0_75), .ZN(n_0_74));
   NOR2_X1 i_0_560 (.A1(B[15]), .A2(n_0_76), .ZN(n_0_75));
   INV_X1 i_0_561 (.A(n_0_89), .ZN(n_0_76));
   NOR2_X1 i_0_562 (.A1(B[11]), .A2(n_0_90), .ZN(n_0_89));
   INV_X1 i_0_563 (.A(n_0_91), .ZN(n_0_90));
   NOR2_X1 i_0_564 (.A1(B[10]), .A2(n_0_92), .ZN(n_0_91));
   INV_X1 i_0_565 (.A(n_0_93), .ZN(n_0_92));
   NOR2_X1 i_0_566 (.A1(B[9]), .A2(n_0_94), .ZN(n_0_93));
   INV_X1 i_0_567 (.A(n_0_95), .ZN(n_0_94));
   NOR2_X1 i_0_568 (.A1(B[8]), .A2(n_0_96), .ZN(n_0_95));
   INV_X1 i_0_569 (.A(n_0_110), .ZN(n_0_96));
   NOR2_X1 i_0_570 (.A1(B[7]), .A2(n_0_111), .ZN(n_0_110));
   INV_X1 i_0_571 (.A(n_0_112), .ZN(n_0_111));
   NOR2_X1 i_0_572 (.A1(B[6]), .A2(n_0_113), .ZN(n_0_112));
   INV_X1 i_0_573 (.A(n_0_114), .ZN(n_0_113));
   NOR2_X1 i_0_574 (.A1(B[5]), .A2(n_0_115), .ZN(n_0_114));
   INV_X1 i_0_575 (.A(n_0_116), .ZN(n_0_115));
   NOR2_X1 i_0_576 (.A1(B[4]), .A2(n_0_131), .ZN(n_0_116));
   INV_X1 i_0_577 (.A(n_0_132), .ZN(n_0_131));
   NOR2_X1 i_0_578 (.A1(B[3]), .A2(n_0_133), .ZN(n_0_132));
   INV_X1 i_0_579 (.A(n_0_134), .ZN(n_0_133));
   NOR2_X1 i_0_580 (.A1(B[2]), .A2(n_0_135), .ZN(n_0_134));
   INV_X1 i_0_581 (.A(n_0_136), .ZN(n_0_135));
   NOR2_X1 i_0_582 (.A1(B[1]), .A2(B[0]), .ZN(n_0_136));
   INV_X1 i_0_583 (.A(A[0]), .ZN(n_0_152));
   INV_X1 i_0_584 (.A(A[1]), .ZN(n_0_153));
   INV_X1 i_0_585 (.A(A[2]), .ZN(n_0_154));
   INV_X1 i_0_586 (.A(A[3]), .ZN(n_0_155));
   INV_X1 i_0_587 (.A(A[4]), .ZN(n_0_156));
   INV_X1 i_0_588 (.A(A[5]), .ZN(n_0_173));
   INV_X1 i_0_589 (.A(A[6]), .ZN(n_0_174));
   INV_X1 i_0_590 (.A(A[7]), .ZN(n_0_175));
   INV_X1 i_0_591 (.A(A[8]), .ZN(n_0_176));
   INV_X1 i_0_592 (.A(A[9]), .ZN(n_0_194));
   INV_X1 i_0_593 (.A(A[10]), .ZN(n_0_195));
   INV_X1 i_0_594 (.A(A[11]), .ZN(n_0_196));
   INV_X1 i_0_595 (.A(A[15]), .ZN(n_0_215));
   FA_X1 i_1_0 (.A(B[1]), .B(n_190), .CI(n_1_166), .CO(n_1_2), .S(n_265));
   FA_X1 i_1_1 (.A(B[2]), .B(n_191), .CI(n_1_2), .CO(n_1_3), .S(n_266));
   FA_X1 i_1_2 (.A(B[3]), .B(n_192), .CI(n_1_3), .CO(n_1_4), .S(n_267));
   FA_X1 i_1_3 (.A(B[4]), .B(n_193), .CI(n_1_4), .CO(n_1_5), .S(n_268));
   FA_X1 i_1_4 (.A(B[5]), .B(n_194), .CI(n_1_5), .CO(n_1_6), .S(n_269));
   FA_X1 i_1_5 (.A(B[6]), .B(n_195), .CI(n_1_6), .CO(n_1_7), .S(n_270));
   FA_X1 i_1_6 (.A(B[7]), .B(n_196), .CI(n_1_7), .CO(n_1_8), .S(n_271));
   FA_X1 i_1_7 (.A(B[8]), .B(n_197), .CI(n_1_8), .CO(n_1_9), .S(n_272));
   FA_X1 i_1_8 (.A(B[9]), .B(n_198), .CI(n_1_9), .CO(n_1_10), .S(n_273));
   FA_X1 i_1_9 (.A(B[10]), .B(n_199), .CI(n_1_10), .CO(n_1_11), .S(n_274));
   FA_X1 i_1_10 (.A(B[11]), .B(n_200), .CI(n_1_11), .CO(n_1_12), .S(n_275));
   FA_X1 i_1_11 (.A(B[15]), .B(n_201), .CI(n_1_12), .CO(n_1_13), .S(n_276));
   FA_X1 i_1_12 (.A(B[15]), .B(n_202), .CI(n_1_13), .CO(n_1_14), .S(n_277));
   FA_X1 i_1_13 (.A(n_250), .B(n_190), .CI(n_1_166), .CO(n_1_0), .S(n_278));
   FA_X1 i_1_14 (.A(n_251), .B(n_191), .CI(n_1_0), .CO(n_1_1), .S(n_279));
   FA_X1 i_1_15 (.A(n_252), .B(n_192), .CI(n_1_1), .CO(n_1_15), .S(n_280));
   FA_X1 i_1_16 (.A(n_253), .B(n_193), .CI(n_1_15), .CO(n_1_16), .S(n_281));
   FA_X1 i_1_17 (.A(n_254), .B(n_194), .CI(n_1_16), .CO(n_1_17), .S(n_282));
   FA_X1 i_1_18 (.A(n_255), .B(n_195), .CI(n_1_17), .CO(n_1_18), .S(n_283));
   FA_X1 i_1_19 (.A(n_256), .B(n_196), .CI(n_1_18), .CO(n_1_19), .S(n_284));
   FA_X1 i_1_20 (.A(n_257), .B(n_197), .CI(n_1_19), .CO(n_1_20), .S(n_285));
   FA_X1 i_1_21 (.A(n_258), .B(n_198), .CI(n_1_20), .CO(n_1_21), .S(n_286));
   FA_X1 i_1_22 (.A(n_259), .B(n_199), .CI(n_1_21), .CO(n_1_22), .S(n_287));
   FA_X1 i_1_23 (.A(n_260), .B(n_200), .CI(n_1_22), .CO(n_1_23), .S(n_288));
   FA_X1 i_1_24 (.A(n_261), .B(n_201), .CI(n_1_23), .CO(n_1_24), .S(n_289));
   FA_X1 i_1_25 (.A(n_262), .B(n_202), .CI(n_1_24), .CO(n_1_25), .S(n_290));
   FA_X1 i_1_26 (.A(B[1]), .B(n_176), .CI(n_1_167), .CO(n_1_26), .S(n_291));
   FA_X1 i_1_27 (.A(B[2]), .B(n_177), .CI(n_1_26), .CO(n_1_27), .S(n_292));
   FA_X1 i_1_28 (.A(B[3]), .B(n_178), .CI(n_1_27), .CO(n_1_28), .S(n_293));
   FA_X1 i_1_29 (.A(B[4]), .B(n_179), .CI(n_1_28), .CO(n_1_29), .S(n_294));
   FA_X1 i_1_30 (.A(B[5]), .B(n_180), .CI(n_1_29), .CO(n_1_30), .S(n_295));
   FA_X1 i_1_31 (.A(B[6]), .B(n_181), .CI(n_1_30), .CO(n_1_31), .S(n_296));
   FA_X1 i_1_32 (.A(B[7]), .B(n_182), .CI(n_1_31), .CO(n_1_32), .S(n_297));
   FA_X1 i_1_33 (.A(B[8]), .B(n_183), .CI(n_1_32), .CO(n_1_33), .S(n_298));
   FA_X1 i_1_34 (.A(B[9]), .B(n_184), .CI(n_1_33), .CO(n_1_34), .S(n_299));
   FA_X1 i_1_35 (.A(B[10]), .B(n_185), .CI(n_1_34), .CO(n_1_35), .S(n_300));
   FA_X1 i_1_36 (.A(B[11]), .B(n_186), .CI(n_1_35), .CO(n_1_36), .S(n_301));
   FA_X1 i_1_37 (.A(B[15]), .B(n_187), .CI(n_1_36), .CO(n_1_37), .S(n_302));
   FA_X1 i_1_38 (.A(B[15]), .B(n_188), .CI(n_1_37), .CO(n_1_38), .S(n_303));
   FA_X1 i_1_39 (.A(n_250), .B(n_176), .CI(n_1_167), .CO(n_1_39), .S(n_304));
   FA_X1 i_1_40 (.A(n_251), .B(n_177), .CI(n_1_39), .CO(n_1_40), .S(n_305));
   FA_X1 i_1_41 (.A(n_252), .B(n_178), .CI(n_1_40), .CO(n_1_41), .S(n_306));
   FA_X1 i_1_42 (.A(n_253), .B(n_179), .CI(n_1_41), .CO(n_1_42), .S(n_307));
   FA_X1 i_1_43 (.A(n_254), .B(n_180), .CI(n_1_42), .CO(n_1_43), .S(n_308));
   FA_X1 i_1_44 (.A(n_255), .B(n_181), .CI(n_1_43), .CO(n_1_44), .S(n_309));
   FA_X1 i_1_45 (.A(n_256), .B(n_182), .CI(n_1_44), .CO(n_1_45), .S(n_310));
   FA_X1 i_1_46 (.A(n_257), .B(n_183), .CI(n_1_45), .CO(n_1_46), .S(n_311));
   FA_X1 i_1_47 (.A(n_258), .B(n_184), .CI(n_1_46), .CO(n_1_47), .S(n_312));
   FA_X1 i_1_48 (.A(n_259), .B(n_185), .CI(n_1_47), .CO(n_1_48), .S(n_313));
   FA_X1 i_1_49 (.A(n_260), .B(n_186), .CI(n_1_48), .CO(n_1_49), .S(n_314));
   FA_X1 i_1_50 (.A(n_261), .B(n_187), .CI(n_1_49), .CO(n_1_50), .S(n_315));
   FA_X1 i_1_51 (.A(n_262), .B(n_188), .CI(n_1_50), .CO(n_1_51), .S(n_316));
   FA_X1 i_1_52 (.A(B[1]), .B(n_163), .CI(n_1_168), .CO(n_1_52), .S(n_317));
   FA_X1 i_1_53 (.A(B[2]), .B(n_164), .CI(n_1_52), .CO(n_1_53), .S(n_318));
   FA_X1 i_1_54 (.A(B[3]), .B(n_165), .CI(n_1_53), .CO(n_1_54), .S(n_319));
   FA_X1 i_1_55 (.A(B[4]), .B(n_166), .CI(n_1_54), .CO(n_1_55), .S(n_320));
   FA_X1 i_1_56 (.A(B[5]), .B(n_167), .CI(n_1_55), .CO(n_1_56), .S(n_321));
   FA_X1 i_1_57 (.A(B[6]), .B(n_168), .CI(n_1_56), .CO(n_1_57), .S(n_322));
   FA_X1 i_1_58 (.A(B[7]), .B(n_169), .CI(n_1_57), .CO(n_1_58), .S(n_323));
   FA_X1 i_1_59 (.A(B[8]), .B(n_170), .CI(n_1_58), .CO(n_1_59), .S(n_324));
   FA_X1 i_1_60 (.A(B[9]), .B(n_171), .CI(n_1_59), .CO(n_1_60), .S(n_325));
   FA_X1 i_1_61 (.A(B[10]), .B(n_172), .CI(n_1_60), .CO(n_1_61), .S(n_326));
   FA_X1 i_1_62 (.A(B[11]), .B(n_173), .CI(n_1_61), .CO(n_1_62), .S(n_327));
   FA_X1 i_1_63 (.A(B[15]), .B(n_174), .CI(n_1_62), .CO(n_1_63), .S(n_328));
   FA_X1 i_1_64 (.A(n_250), .B(n_163), .CI(n_1_168), .CO(n_1_64), .S(n_329));
   FA_X1 i_1_65 (.A(n_251), .B(n_164), .CI(n_1_64), .CO(n_1_65), .S(n_330));
   FA_X1 i_1_66 (.A(n_252), .B(n_165), .CI(n_1_65), .CO(n_1_66), .S(n_331));
   FA_X1 i_1_67 (.A(n_253), .B(n_166), .CI(n_1_66), .CO(n_1_67), .S(n_332));
   FA_X1 i_1_68 (.A(n_254), .B(n_167), .CI(n_1_67), .CO(n_1_68), .S(n_333));
   FA_X1 i_1_69 (.A(n_255), .B(n_168), .CI(n_1_68), .CO(n_1_69), .S(n_334));
   FA_X1 i_1_70 (.A(n_256), .B(n_169), .CI(n_1_69), .CO(n_1_70), .S(n_335));
   FA_X1 i_1_71 (.A(n_257), .B(n_170), .CI(n_1_70), .CO(n_1_71), .S(n_336));
   FA_X1 i_1_72 (.A(n_258), .B(n_171), .CI(n_1_71), .CO(n_1_72), .S(n_337));
   FA_X1 i_1_73 (.A(n_259), .B(n_172), .CI(n_1_72), .CO(n_1_73), .S(n_338));
   FA_X1 i_1_74 (.A(n_260), .B(n_173), .CI(n_1_73), .CO(n_1_74), .S(n_339));
   FA_X1 i_1_75 (.A(n_261), .B(n_174), .CI(n_1_74), .CO(n_1_75), .S(n_340));
   FA_X1 i_1_76 (.A(B[1]), .B(n_151), .CI(n_1_169), .CO(n_1_76), .S(n_341));
   FA_X1 i_1_77 (.A(B[2]), .B(n_152), .CI(n_1_76), .CO(n_1_77), .S(n_342));
   FA_X1 i_1_78 (.A(B[3]), .B(n_153), .CI(n_1_77), .CO(n_1_78), .S(n_343));
   FA_X1 i_1_79 (.A(B[4]), .B(n_154), .CI(n_1_78), .CO(n_1_79), .S(n_344));
   FA_X1 i_1_80 (.A(B[5]), .B(n_155), .CI(n_1_79), .CO(n_1_80), .S(n_345));
   FA_X1 i_1_81 (.A(B[6]), .B(n_156), .CI(n_1_80), .CO(n_1_81), .S(n_346));
   FA_X1 i_1_82 (.A(B[7]), .B(n_157), .CI(n_1_81), .CO(n_1_82), .S(n_347));
   FA_X1 i_1_83 (.A(B[8]), .B(n_158), .CI(n_1_82), .CO(n_1_83), .S(n_348));
   FA_X1 i_1_84 (.A(B[9]), .B(n_159), .CI(n_1_83), .CO(n_1_84), .S(n_349));
   FA_X1 i_1_85 (.A(B[10]), .B(n_160), .CI(n_1_84), .CO(n_1_85), .S(n_350));
   FA_X1 i_1_86 (.A(B[11]), .B(n_161), .CI(n_1_85), .CO(n_1_86), .S(n_351));
   FA_X1 i_1_87 (.A(n_250), .B(n_151), .CI(n_1_169), .CO(n_1_87), .S(n_352));
   FA_X1 i_1_88 (.A(n_251), .B(n_152), .CI(n_1_87), .CO(n_1_88), .S(n_353));
   FA_X1 i_1_89 (.A(n_252), .B(n_153), .CI(n_1_88), .CO(n_1_89), .S(n_354));
   FA_X1 i_1_90 (.A(n_253), .B(n_154), .CI(n_1_89), .CO(n_1_90), .S(n_355));
   FA_X1 i_1_91 (.A(n_254), .B(n_155), .CI(n_1_90), .CO(n_1_91), .S(n_356));
   FA_X1 i_1_92 (.A(n_255), .B(n_156), .CI(n_1_91), .CO(n_1_92), .S(n_357));
   FA_X1 i_1_93 (.A(n_256), .B(n_157), .CI(n_1_92), .CO(n_1_93), .S(n_358));
   FA_X1 i_1_94 (.A(n_257), .B(n_158), .CI(n_1_93), .CO(n_1_94), .S(n_359));
   FA_X1 i_1_95 (.A(n_258), .B(n_159), .CI(n_1_94), .CO(n_1_95), .S(n_360));
   FA_X1 i_1_96 (.A(n_259), .B(n_160), .CI(n_1_95), .CO(n_1_96), .S(n_361));
   FA_X1 i_1_97 (.A(n_260), .B(n_161), .CI(n_1_96), .CO(n_1_97), .S(n_362));
   FA_X1 i_1_98 (.A(B[1]), .B(n_140), .CI(n_1_170), .CO(n_1_98), .S(n_363));
   FA_X1 i_1_99 (.A(B[2]), .B(n_141), .CI(n_1_98), .CO(n_1_99), .S(n_364));
   FA_X1 i_1_100 (.A(B[3]), .B(n_142), .CI(n_1_99), .CO(n_1_100), .S(n_365));
   FA_X1 i_1_101 (.A(B[4]), .B(n_143), .CI(n_1_100), .CO(n_1_101), .S(n_366));
   FA_X1 i_1_102 (.A(B[5]), .B(n_144), .CI(n_1_101), .CO(n_1_102), .S(n_367));
   FA_X1 i_1_103 (.A(B[6]), .B(n_145), .CI(n_1_102), .CO(n_1_103), .S(n_368));
   FA_X1 i_1_104 (.A(B[7]), .B(n_146), .CI(n_1_103), .CO(n_1_104), .S(n_369));
   FA_X1 i_1_105 (.A(B[8]), .B(n_147), .CI(n_1_104), .CO(n_1_105), .S(n_370));
   FA_X1 i_1_106 (.A(B[9]), .B(n_148), .CI(n_1_105), .CO(n_1_106), .S(n_371));
   FA_X1 i_1_107 (.A(B[10]), .B(n_149), .CI(n_1_106), .CO(n_1_107), .S(n_372));
   FA_X1 i_1_108 (.A(n_250), .B(n_140), .CI(n_1_170), .CO(n_1_108), .S(n_373));
   FA_X1 i_1_109 (.A(n_251), .B(n_141), .CI(n_1_108), .CO(n_1_109), .S(n_374));
   FA_X1 i_1_110 (.A(n_252), .B(n_142), .CI(n_1_109), .CO(n_1_110), .S(n_375));
   FA_X1 i_1_111 (.A(n_253), .B(n_143), .CI(n_1_110), .CO(n_1_111), .S(n_376));
   FA_X1 i_1_112 (.A(n_254), .B(n_144), .CI(n_1_111), .CO(n_1_112), .S(n_377));
   FA_X1 i_1_113 (.A(n_255), .B(n_145), .CI(n_1_112), .CO(n_1_113), .S(n_378));
   FA_X1 i_1_114 (.A(n_256), .B(n_146), .CI(n_1_113), .CO(n_1_114), .S(n_379));
   FA_X1 i_1_115 (.A(n_257), .B(n_147), .CI(n_1_114), .CO(n_1_115), .S(n_380));
   FA_X1 i_1_116 (.A(n_258), .B(n_148), .CI(n_1_115), .CO(n_1_116), .S(n_381));
   FA_X1 i_1_117 (.A(n_259), .B(n_149), .CI(n_1_116), .CO(n_1_117), .S(n_382));
   FA_X1 i_1_118 (.A(B[1]), .B(n_130), .CI(n_1_171), .CO(n_1_118), .S(n_383));
   FA_X1 i_1_119 (.A(B[2]), .B(n_131), .CI(n_1_118), .CO(n_1_119), .S(n_384));
   FA_X1 i_1_120 (.A(B[3]), .B(n_132), .CI(n_1_119), .CO(n_1_120), .S(n_385));
   FA_X1 i_1_121 (.A(B[4]), .B(n_133), .CI(n_1_120), .CO(n_1_121), .S(n_386));
   FA_X1 i_1_122 (.A(B[5]), .B(n_134), .CI(n_1_121), .CO(n_1_122), .S(n_387));
   FA_X1 i_1_123 (.A(B[6]), .B(n_135), .CI(n_1_122), .CO(n_1_123), .S(n_388));
   FA_X1 i_1_124 (.A(B[7]), .B(n_136), .CI(n_1_123), .CO(n_1_124), .S(n_389));
   FA_X1 i_1_125 (.A(B[8]), .B(n_137), .CI(n_1_124), .CO(n_1_125), .S(n_390));
   FA_X1 i_1_126 (.A(B[9]), .B(n_138), .CI(n_1_125), .CO(n_1_126), .S(n_391));
   FA_X1 i_1_127 (.A(n_250), .B(n_130), .CI(n_1_171), .CO(n_1_127), .S(n_392));
   FA_X1 i_1_128 (.A(n_251), .B(n_131), .CI(n_1_127), .CO(n_1_128), .S(n_393));
   FA_X1 i_1_129 (.A(n_252), .B(n_132), .CI(n_1_128), .CO(n_1_129), .S(n_394));
   FA_X1 i_1_130 (.A(n_253), .B(n_133), .CI(n_1_129), .CO(n_1_130), .S(n_395));
   FA_X1 i_1_131 (.A(n_254), .B(n_134), .CI(n_1_130), .CO(n_1_131), .S(n_396));
   FA_X1 i_1_132 (.A(n_255), .B(n_135), .CI(n_1_131), .CO(n_1_132), .S(n_397));
   FA_X1 i_1_133 (.A(n_256), .B(n_136), .CI(n_1_132), .CO(n_1_133), .S(n_398));
   FA_X1 i_1_134 (.A(n_257), .B(n_137), .CI(n_1_133), .CO(n_1_134), .S(n_399));
   FA_X1 i_1_135 (.A(n_258), .B(n_138), .CI(n_1_134), .CO(n_1_135), .S(n_400));
   FA_X1 i_1_136 (.A(B[1]), .B(n_121), .CI(n_1_172), .CO(n_1_136), .S(n_401));
   FA_X1 i_1_137 (.A(B[2]), .B(n_122), .CI(n_1_136), .CO(n_1_137), .S(n_402));
   FA_X1 i_1_138 (.A(B[3]), .B(n_123), .CI(n_1_137), .CO(n_1_138), .S(n_403));
   FA_X1 i_1_139 (.A(B[4]), .B(n_124), .CI(n_1_138), .CO(n_1_139), .S(n_404));
   FA_X1 i_1_140 (.A(B[5]), .B(n_125), .CI(n_1_139), .CO(n_1_140), .S(n_405));
   FA_X1 i_1_141 (.A(B[6]), .B(n_126), .CI(n_1_140), .CO(n_1_141), .S(n_406));
   FA_X1 i_1_142 (.A(B[7]), .B(n_127), .CI(n_1_141), .CO(n_1_142), .S(n_407));
   FA_X1 i_1_143 (.A(B[8]), .B(n_128), .CI(n_1_142), .CO(n_1_143), .S(n_408));
   FA_X1 i_1_144 (.A(n_250), .B(n_121), .CI(n_1_172), .CO(n_1_144), .S(n_409));
   FA_X1 i_1_145 (.A(n_251), .B(n_122), .CI(n_1_144), .CO(n_1_145), .S(n_410));
   FA_X1 i_1_146 (.A(n_252), .B(n_123), .CI(n_1_145), .CO(n_1_146), .S(n_411));
   FA_X1 i_1_147 (.A(n_253), .B(n_124), .CI(n_1_146), .CO(n_1_147), .S(n_412));
   FA_X1 i_1_148 (.A(n_254), .B(n_125), .CI(n_1_147), .CO(n_1_148), .S(n_413));
   FA_X1 i_1_149 (.A(n_255), .B(n_126), .CI(n_1_148), .CO(n_1_149), .S(n_414));
   FA_X1 i_1_150 (.A(n_256), .B(n_127), .CI(n_1_149), .CO(n_1_150), .S(n_415));
   FA_X1 i_1_151 (.A(n_257), .B(n_128), .CI(n_1_150), .CO(n_1_151), .S(n_416));
   FA_X1 i_1_152 (.A(B[1]), .B(n_113), .CI(n_1_173), .CO(n_1_152), .S(n_417));
   FA_X1 i_1_153 (.A(B[2]), .B(n_114), .CI(n_1_152), .CO(n_1_153), .S(n_418));
   FA_X1 i_1_154 (.A(B[3]), .B(n_115), .CI(n_1_153), .CO(n_1_154), .S(n_419));
   FA_X1 i_1_155 (.A(B[4]), .B(n_116), .CI(n_1_154), .CO(n_1_155), .S(n_420));
   FA_X1 i_1_156 (.A(B[5]), .B(n_117), .CI(n_1_155), .CO(n_1_156), .S(n_421));
   FA_X1 i_1_157 (.A(B[6]), .B(n_118), .CI(n_1_156), .CO(n_1_157), .S(n_422));
   FA_X1 i_1_158 (.A(B[7]), .B(n_119), .CI(n_1_157), .CO(n_1_158), .S(n_423));
   FA_X1 i_1_159 (.A(n_250), .B(n_113), .CI(n_1_173), .CO(n_1_159), .S(n_424));
   FA_X1 i_1_160 (.A(n_251), .B(n_114), .CI(n_1_159), .CO(n_1_160), .S(n_425));
   FA_X1 i_1_161 (.A(n_252), .B(n_115), .CI(n_1_160), .CO(n_1_161), .S(n_426));
   FA_X1 i_1_162 (.A(n_253), .B(n_116), .CI(n_1_161), .CO(n_1_162), .S(n_427));
   FA_X1 i_1_163 (.A(n_254), .B(n_117), .CI(n_1_162), .CO(n_1_163), .S(n_428));
   FA_X1 i_1_164 (.A(n_255), .B(n_118), .CI(n_1_163), .CO(n_1_164), .S(n_429));
   FA_X1 i_1_165 (.A(n_256), .B(n_119), .CI(n_1_164), .CO(n_1_165), .S(n_430));
   HA_X1 i_1_166 (.A(B[0]), .B(n_189), .CO(n_1_166), .S(n_431));
   HA_X1 i_1_167 (.A(B[0]), .B(n_175), .CO(n_1_167), .S(n_432));
   HA_X1 i_1_168 (.A(B[0]), .B(n_162), .CO(n_1_168), .S(n_433));
   HA_X1 i_1_169 (.A(B[0]), .B(n_150), .CO(n_1_169), .S(n_434));
   HA_X1 i_1_170 (.A(B[0]), .B(n_139), .CO(n_1_170), .S(n_435));
   HA_X1 i_1_171 (.A(B[0]), .B(n_129), .CO(n_1_171), .S(n_436));
   HA_X1 i_1_172 (.A(B[0]), .B(n_120), .CO(n_1_172), .S(n_437));
   HA_X1 i_1_173 (.A(B[0]), .B(n_112), .CO(n_1_173), .S(n_438));
   XNOR2_X1 i_1_174 (.A(n_203), .B(n_1_174), .ZN(n_439));
   XNOR2_X1 i_1_175 (.A(n_263), .B(n_1_25), .ZN(n_1_174));
   XNOR2_X1 i_1_176 (.A(B[15]), .B(n_1_175), .ZN(n_440));
   XNOR2_X1 i_1_177 (.A(n_203), .B(n_1_14), .ZN(n_1_175));
endmodule

module multiplier_16bit(first_operand, second_operand, out, enable, overflow);
   input [15:0]first_operand;
   input [15:0]second_operand;
   output [15:0]out;
   input enable;
   output overflow;

   wire [31:0]temp_result_wire;
   wire n_0_0_4;
   wire n_0_0_6;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_5;
   wire n_0_0_7;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;

   booth_16bit_multiplier mult (.A({first_operand[12], uc_0, uc_1, uc_2, 
      first_operand[11], first_operand[10], first_operand[9], first_operand[8], 
      first_operand[7], first_operand[6], first_operand[5], first_operand[4], 
      first_operand[3], first_operand[2], first_operand[1], first_operand[0]}), 
      .B({second_operand[12], uc_3, uc_4, uc_5, second_operand[11], 
      second_operand[10], second_operand[9], second_operand[8], 
      second_operand[7], second_operand[6], second_operand[5], second_operand[4], 
      second_operand[3], second_operand[2], second_operand[1], second_operand[0]}), 
      .product({uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, 
      uc_16, uc_17, temp_result_wire[19], temp_result_wire[18], 
      temp_result_wire[17], temp_result_wire[16], temp_result_wire[15], 
      temp_result_wire[14], temp_result_wire[13], temp_result_wire[12], 
      temp_result_wire[11], temp_result_wire[10], temp_result_wire[9], 
      temp_result_wire[8], temp_result_wire[7], temp_result_wire[6], 
      temp_result_wire[5], temp_result_wire[4], temp_result_wire[3], 
      temp_result_wire[2], temp_result_wire[1], temp_result_wire[0]}));
   MUX2_X1 i_0_0_0 (.A(n_0_0_3), .B(n_0_0_4), .S(n_0_0_46), .Z(out[1]));
   MUX2_X1 i_0_0_1 (.A(n_0_0_4), .B(n_0_0_6), .S(n_0_0_46), .Z(out[2]));
   MUX2_X1 i_0_0_2 (.A(n_0_0_25), .B(n_0_0_9), .S(n_0_0_31), .Z(n_0_0_4));
   MUX2_X1 i_0_0_3 (.A(n_0_0_6), .B(n_0_0_8), .S(n_0_0_46), .Z(out[3]));
   MUX2_X1 i_0_0_4 (.A(n_0_0_7), .B(n_0_0_11), .S(n_0_0_31), .Z(n_0_0_6));
   MUX2_X1 i_0_0_5 (.A(n_0_0_8), .B(n_0_0_10), .S(n_0_0_46), .Z(out[4]));
   MUX2_X1 i_0_0_6 (.A(n_0_0_9), .B(n_0_0_13), .S(n_0_0_31), .Z(n_0_0_8));
   MUX2_X1 i_0_0_7 (.A(temp_result_wire[4]), .B(temp_result_wire[8]), .S(
      n_0_0_28), .Z(n_0_0_9));
   MUX2_X1 i_0_0_15 (.A(n_0_0_10), .B(n_0_0_12), .S(n_0_0_46), .Z(out[5]));
   MUX2_X1 i_0_0_8 (.A(n_0_0_11), .B(n_0_0_15), .S(n_0_0_31), .Z(n_0_0_10));
   MUX2_X1 i_0_0_9 (.A(temp_result_wire[5]), .B(temp_result_wire[9]), .S(
      n_0_0_28), .Z(n_0_0_11));
   MUX2_X1 i_0_0_18 (.A(n_0_0_12), .B(n_0_0_14), .S(n_0_0_46), .Z(out[6]));
   MUX2_X1 i_0_0_19 (.A(n_0_0_13), .B(n_0_0_17), .S(n_0_0_31), .Z(n_0_0_12));
   MUX2_X1 i_0_0_10 (.A(temp_result_wire[6]), .B(temp_result_wire[10]), .S(
      n_0_0_28), .Z(n_0_0_13));
   MUX2_X1 i_0_0_21 (.A(n_0_0_14), .B(n_0_0_16), .S(n_0_0_46), .Z(out[7]));
   MUX2_X1 i_0_0_22 (.A(n_0_0_15), .B(n_0_0_19), .S(n_0_0_31), .Z(n_0_0_14));
   MUX2_X1 i_0_0_11 (.A(temp_result_wire[7]), .B(temp_result_wire[11]), .S(
      n_0_0_28), .Z(n_0_0_15));
   MUX2_X1 i_0_0_24 (.A(n_0_0_16), .B(n_0_0_18), .S(n_0_0_46), .Z(out[8]));
   MUX2_X1 i_0_0_25 (.A(n_0_0_17), .B(n_0_0_21), .S(n_0_0_31), .Z(n_0_0_16));
   MUX2_X1 i_0_0_26 (.A(temp_result_wire[8]), .B(temp_result_wire[12]), .S(
      n_0_0_28), .Z(n_0_0_17));
   MUX2_X1 i_0_0_27 (.A(n_0_0_18), .B(n_0_0_20), .S(n_0_0_46), .Z(out[9]));
   MUX2_X1 i_0_0_28 (.A(n_0_0_19), .B(n_0_0_23), .S(n_0_0_31), .Z(n_0_0_18));
   MUX2_X1 i_0_0_29 (.A(temp_result_wire[9]), .B(temp_result_wire[13]), .S(
      n_0_0_28), .Z(n_0_0_19));
   MUX2_X1 i_0_0_30 (.A(n_0_0_20), .B(n_0_0_22), .S(n_0_0_46), .Z(out[10]));
   MUX2_X1 i_0_0_31 (.A(n_0_0_21), .B(n_0_0_63), .S(n_0_0_31), .Z(n_0_0_20));
   MUX2_X1 i_0_0_32 (.A(temp_result_wire[10]), .B(temp_result_wire[14]), 
      .S(n_0_0_28), .Z(n_0_0_21));
   MUX2_X1 i_0_0_12 (.A(n_0_0_22), .B(n_0_0_61), .S(n_0_0_46), .Z(out[11]));
   MUX2_X1 i_0_0_13 (.A(n_0_0_23), .B(n_0_0_58), .S(n_0_0_31), .Z(n_0_0_22));
   MUX2_X1 i_0_0_14 (.A(temp_result_wire[11]), .B(temp_result_wire[15]), 
      .S(n_0_0_28), .Z(n_0_0_23));
   AOI21_X1 i_0_0_16 (.A(n_0_0_40), .B1(n_0_0_37), .B2(n_0_0_52), .ZN(out[13]));
   NOR2_X1 i_0_0_17 (.A1(n_0_0_37), .A2(first_operand[13]), .ZN(n_0_0_40));
   AOI21_X1 i_0_0_55 (.A(n_0_0_41), .B1(n_0_0_37), .B2(n_0_0_53), .ZN(out[14]));
   NOR2_X1 i_0_0_56 (.A1(n_0_0_37), .A2(first_operand[14]), .ZN(n_0_0_41));
   OR2_X1 i_0_0_64 (.A1(second_operand[15]), .A2(first_operand[15]), .ZN(out[15]));
   INV_X1 i_0_0_20 (.A(n_0_0_0), .ZN(out[0]));
   AOI22_X1 i_0_0_23 (.A1(n_0_0_47), .A2(n_0_0_1), .B1(n_0_0_46), .B2(n_0_0_3), 
      .ZN(n_0_0_0));
   OAI22_X1 i_0_0_33 (.A1(n_0_0_31), .A2(n_0_0_2), .B1(n_0_0_30), .B2(n_0_0_26), 
      .ZN(n_0_0_1));
   AOI22_X1 i_0_0_34 (.A1(temp_result_wire[4]), .A2(n_0_0_28), .B1(
      temp_result_wire[0]), .B2(n_0_0_27), .ZN(n_0_0_2));
   AOI22_X1 i_0_0_35 (.A1(n_0_0_30), .A2(n_0_0_5), .B1(n_0_0_31), .B2(n_0_0_24), 
      .ZN(n_0_0_3));
   OAI22_X1 i_0_0_36 (.A1(temp_result_wire[5]), .A2(n_0_0_27), .B1(
      temp_result_wire[1]), .B2(n_0_0_28), .ZN(n_0_0_5));
   INV_X1 i_0_0_37 (.A(n_0_0_24), .ZN(n_0_0_7));
   OAI22_X1 i_0_0_38 (.A1(temp_result_wire[7]), .A2(n_0_0_27), .B1(
      temp_result_wire[3]), .B2(n_0_0_28), .ZN(n_0_0_24));
   INV_X1 i_0_0_39 (.A(n_0_0_26), .ZN(n_0_0_25));
   OAI22_X1 i_0_0_40 (.A1(temp_result_wire[6]), .A2(n_0_0_27), .B1(
      temp_result_wire[2]), .B2(n_0_0_28), .ZN(n_0_0_26));
   INV_X1 i_0_0_41 (.A(n_0_0_28), .ZN(n_0_0_27));
   OAI33_X1 i_0_0_42 (.A1(n_0_0_54), .A2(first_operand[15]), .A3(n_0_0_38), 
      .B1(n_0_0_45), .B2(n_0_0_39), .B3(n_0_0_29), .ZN(n_0_0_28));
   NOR2_X1 i_0_0_43 (.A1(n_0_0_48), .A2(n_0_0_42), .ZN(n_0_0_29));
   INV_X1 i_0_0_44 (.A(n_0_0_31), .ZN(n_0_0_30));
   OAI21_X1 i_0_0_45 (.A(n_0_0_32), .B1(n_0_0_36), .B2(n_0_0_33), .ZN(n_0_0_31));
   OAI221_X1 i_0_0_46 (.A(n_0_0_36), .B1(n_0_0_49), .B2(n_0_0_34), .C1(n_0_0_48), 
      .C2(n_0_0_35), .ZN(n_0_0_32));
   AOI22_X1 i_0_0_47 (.A1(n_0_0_51), .A2(n_0_0_34), .B1(n_0_0_50), .B2(n_0_0_35), 
      .ZN(n_0_0_33));
   INV_X1 i_0_0_48 (.A(n_0_0_35), .ZN(n_0_0_34));
   NOR2_X1 i_0_0_49 (.A1(n_0_0_42), .A2(n_0_0_39), .ZN(n_0_0_35));
   INV_X1 i_0_0_50 (.A(n_0_0_37), .ZN(n_0_0_36));
   OAI22_X1 i_0_0_51 (.A1(n_0_0_54), .A2(first_operand[15]), .B1(n_0_0_44), 
      .B2(n_0_0_38), .ZN(n_0_0_37));
   OAI21_X1 i_0_0_52 (.A(n_0_0_43), .B1(n_0_0_51), .B2(n_0_0_39), .ZN(n_0_0_38));
   NOR2_X1 i_0_0_53 (.A1(n_0_0_53), .A2(first_operand[14]), .ZN(n_0_0_39));
   INV_X1 i_0_0_54 (.A(n_0_0_43), .ZN(n_0_0_42));
   NAND2_X1 i_0_0_57 (.A1(n_0_0_53), .A2(first_operand[14]), .ZN(n_0_0_43));
   INV_X1 i_0_0_58 (.A(n_0_0_45), .ZN(n_0_0_44));
   NAND2_X1 i_0_0_59 (.A1(n_0_0_54), .A2(first_operand[15]), .ZN(n_0_0_45));
   INV_X1 i_0_0_60 (.A(n_0_0_47), .ZN(n_0_0_46));
   NOR2_X1 i_0_0_61 (.A1(n_0_0_50), .A2(n_0_0_49), .ZN(n_0_0_47));
   INV_X1 i_0_0_62 (.A(n_0_0_49), .ZN(n_0_0_48));
   NOR2_X1 i_0_0_63 (.A1(n_0_0_52), .A2(first_operand[13]), .ZN(n_0_0_49));
   INV_X1 i_0_0_65 (.A(n_0_0_51), .ZN(n_0_0_50));
   NAND2_X1 i_0_0_66 (.A1(n_0_0_52), .A2(first_operand[13]), .ZN(n_0_0_51));
   INV_X1 i_0_0_67 (.A(second_operand[13]), .ZN(n_0_0_52));
   INV_X1 i_0_0_68 (.A(second_operand[14]), .ZN(n_0_0_53));
   INV_X1 i_0_0_69 (.A(second_operand[15]), .ZN(n_0_0_54));
   OAI21_X1 i_0_0_70 (.A(n_0_0_55), .B1(n_0_0_46), .B2(n_0_0_60), .ZN(out[12]));
   NAND2_X1 i_0_0_71 (.A1(n_0_0_46), .A2(n_0_0_56), .ZN(n_0_0_55));
   OAI22_X1 i_0_0_72 (.A1(n_0_0_65), .A2(n_0_0_57), .B1(n_0_0_31), .B2(n_0_0_59), 
      .ZN(n_0_0_56));
   AOI22_X1 i_0_0_73 (.A1(n_0_0_66), .A2(temp_result_wire[15]), .B1(n_0_0_28), 
      .B2(temp_result_wire[19]), .ZN(n_0_0_57));
   INV_X1 i_0_0_74 (.A(n_0_0_59), .ZN(n_0_0_58));
   OAI22_X1 i_0_0_75 (.A1(n_0_0_28), .A2(temp_result_wire[13]), .B1(n_0_0_66), 
      .B2(temp_result_wire[17]), .ZN(n_0_0_59));
   INV_X1 i_0_0_76 (.A(n_0_0_61), .ZN(n_0_0_60));
   AOI22_X1 i_0_0_77 (.A1(n_0_0_31), .A2(n_0_0_62), .B1(n_0_0_65), .B2(n_0_0_64), 
      .ZN(n_0_0_61));
   OAI22_X1 i_0_0_78 (.A1(n_0_0_28), .A2(temp_result_wire[14]), .B1(n_0_0_66), 
      .B2(temp_result_wire[18]), .ZN(n_0_0_62));
   INV_X1 i_0_0_79 (.A(n_0_0_64), .ZN(n_0_0_63));
   OAI22_X1 i_0_0_80 (.A1(n_0_0_28), .A2(temp_result_wire[12]), .B1(n_0_0_66), 
      .B2(temp_result_wire[16]), .ZN(n_0_0_64));
   INV_X1 i_0_0_81 (.A(n_0_0_31), .ZN(n_0_0_65));
   INV_X1 i_0_0_82 (.A(n_0_0_28), .ZN(n_0_0_66));
endmodule

module Euler(INT, PROCESS, CLK, DONE, Interpolate_DONE, Interpolate_Enable, 
      RAM_DATA_RD1, RAM_DATA_RD2, RAM_ADD_RD1, RAM_ADD_RD2, RAM_ADD_WR, 
      RAM_DATA_WR, RAM_ENABLE_WR);
   input INT;
   input PROCESS;
   input CLK;
   output DONE;
   input Interpolate_DONE;
   output Interpolate_Enable;
   input [63:0]RAM_DATA_RD1;
   input [63:0]RAM_DATA_RD2;
   output [12:0]RAM_ADD_RD1;
   output [12:0]RAM_ADD_RD2;
   output [12:0]RAM_ADD_WR;
   output [63:0]RAM_DATA_WR;
   output RAM_ENABLE_WR;

   wire [15:0]NEW_MATRIX_ADD;
   wire [15:0]NEW_VECTOR2_ADD;
   wire [15:0]NEW_VECTOR_ADD;
   wire [15:0]NEW_RESULT_ADD;
   wire [15:0]h_VECTOR_RESULT;
   wire [15:0]Multiplication_Result;
   wire [19:0]MATRIX_CNT_adder_tempIn11;
   wire [19:0]FINAL_RESULT_adder_tempIn22;
   wire [19:0]FINAL_RESULT_adder_tempIn11;
   wire [15:0]FINAL_RESULT;
   wire FINAL_RESULT_adder_n_0;
   wire FINAL_RESULT_adder_n_1;
   wire FINAL_RESULT_adder_n_2;
   wire FINAL_RESULT_adder_n_3;
   wire FINAL_RESULT_adder_n_4;
   wire FINAL_RESULT_adder_n_0_0;
   wire FINAL_RESULT_adder_n_5;
   wire FINAL_RESULT_adder_n_0_1;
   wire FINAL_RESULT_adder_n_0_2;
   wire FINAL_RESULT_adder_n_0_3;
   wire FINAL_RESULT_adder_n_6;
   wire FINAL_RESULT_adder_n_0_4;
   wire FINAL_RESULT_adder_n_0_5;
   wire FINAL_RESULT_adder_n_0_6;
   wire FINAL_RESULT_adder_n_7;
   wire FINAL_RESULT_adder_n_0_7;
   wire FINAL_RESULT_adder_n_0_8;
   wire FINAL_RESULT_adder_n_0_9;
   wire FINAL_RESULT_adder_n_8;
   wire FINAL_RESULT_adder_n_0_10;
   wire FINAL_RESULT_adder_n_0_11;
   wire FINAL_RESULT_adder_n_0_12;
   wire FINAL_RESULT_adder_n_9;
   wire FINAL_RESULT_adder_n_0_13;
   wire FINAL_RESULT_adder_n_0_14;
   wire FINAL_RESULT_adder_n_0_15;
   wire FINAL_RESULT_adder_n_10;
   wire FINAL_RESULT_adder_n_0_16;
   wire FINAL_RESULT_adder_n_0_17;
   wire FINAL_RESULT_adder_n_0_18;
   wire FINAL_RESULT_adder_n_0_19;
   wire FINAL_RESULT_adder_n_11;
   wire FINAL_RESULT_adder_n_0_20;
   wire FINAL_RESULT_adder_n_0_21;
   wire FINAL_RESULT_adder_n_0_22;
   wire FINAL_RESULT_adder_n_0_23;
   wire FINAL_RESULT_adder_n_12;
   wire FINAL_RESULT_adder_n_0_24;
   wire FINAL_RESULT_adder_n_0_25;
   wire FINAL_RESULT_adder_n_0_26;
   wire FINAL_RESULT_adder_n_0_27;
   wire FINAL_RESULT_adder_n_0_28;
   wire FINAL_RESULT_adder_n_0_29;
   wire FINAL_RESULT_adder_n_0_30;
   wire FINAL_RESULT_adder_n_0_31;
   wire FINAL_RESULT_adder_n_0_32;
   wire FINAL_RESULT_adder_n_0_33;
   wire FINAL_RESULT_adder_n_14;
   wire FINAL_RESULT_adder_n_15;
   wire FINAL_RESULT_adder_n_16;
   wire FINAL_RESULT_adder_n_17;
   wire FINAL_RESULT_adder_n_18;
   wire FINAL_RESULT_adder_n_0_34;
   wire FINAL_RESULT_adder_n_19;
   wire FINAL_RESULT_adder_n_0_35;
   wire FINAL_RESULT_adder_n_0_36;
   wire FINAL_RESULT_adder_n_0_37;
   wire FINAL_RESULT_adder_n_20;
   wire FINAL_RESULT_adder_n_0_38;
   wire FINAL_RESULT_adder_n_0_39;
   wire FINAL_RESULT_adder_n_0_40;
   wire FINAL_RESULT_adder_n_21;
   wire FINAL_RESULT_adder_n_0_41;
   wire FINAL_RESULT_adder_n_0_42;
   wire FINAL_RESULT_adder_n_0_43;
   wire FINAL_RESULT_adder_n_22;
   wire FINAL_RESULT_adder_n_0_44;
   wire FINAL_RESULT_adder_n_0_45;
   wire FINAL_RESULT_adder_n_0_46;
   wire FINAL_RESULT_adder_n_23;
   wire FINAL_RESULT_adder_n_0_47;
   wire FINAL_RESULT_adder_n_0_48;
   wire FINAL_RESULT_adder_n_0_49;
   wire FINAL_RESULT_adder_n_24;
   wire FINAL_RESULT_adder_n_0_50;
   wire FINAL_RESULT_adder_n_0_51;
   wire FINAL_RESULT_adder_n_0_52;
   wire FINAL_RESULT_adder_n_0_53;
   wire FINAL_RESULT_adder_n_25;
   wire FINAL_RESULT_adder_n_0_54;
   wire FINAL_RESULT_adder_n_0_55;
   wire FINAL_RESULT_adder_n_0_56;
   wire FINAL_RESULT_adder_n_0_57;
   wire FINAL_RESULT_adder_n_26;
   wire FINAL_RESULT_adder_n_0_58;
   wire FINAL_RESULT_adder_n_0_59;
   wire FINAL_RESULT_adder_n_0_60;
   wire FINAL_RESULT_adder_n_0_61;
   wire FINAL_RESULT_adder_n_0_62;
   wire FINAL_RESULT_adder_n_0_63;
   wire FINAL_RESULT_adder_n_0_64;
   wire FINAL_RESULT_adder_n_0_65;
   wire FINAL_RESULT_adder_n_0_66;
   wire FINAL_RESULT_adder_n_0_67;
   wire FINAL_RESULT_adder_n_0_68;
   wire FINAL_RESULT_adder_n_0_69;
   wire FINAL_RESULT_adder_n_0_70;
   wire FINAL_RESULT_adder_n_27;
   wire FINAL_RESULT_adder_n_0_71;
   wire FINAL_RESULT_adder_n_0_72;
   wire FINAL_RESULT_adder_n_0_73;
   wire FINAL_RESULT_adder_n_0_74;
   wire FINAL_RESULT_adder_n_0_75;
   wire FINAL_RESULT_adder_n_0_76;
   wire FINAL_RESULT_adder_n_0_77;
   wire FINAL_RESULT_adder_n_0_78;
   wire FINAL_RESULT_adder_n_0_79;
   wire FINAL_RESULT_adder_n_0_80;
   wire FINAL_RESULT_adder_n_0_81;
   wire FINAL_RESULT_adder_n_13;
   wire FINAL_RESULT_adder_n_0_82;
   wire FINAL_RESULT_adder_n_0_83;
   wire FINAL_RESULT_adder_n_0_84;
   wire FINAL_RESULT_adder_n_0_85;
   wire FINAL_RESULT_adder_n_0_86;
   wire FINAL_RESULT_adder_n_0_87;
   wire FINAL_RESULT_adder_n_0_88;
   wire FINAL_RESULT_adder_n_0_89;
   wire FINAL_RESULT_adder_n_0_90;
   wire FINAL_RESULT_adder_n_0_91;
   wire FINAL_RESULT_adder_n_0_92;
   wire FINAL_RESULT_adder_n_0_93;
   wire FINAL_RESULT_adder_n_0_94;
   wire FINAL_RESULT_adder_n_1_0;
   wire FINAL_RESULT_adder_n_1_1;
   wire FINAL_RESULT_adder_n_1_3;
   wire FINAL_RESULT_adder_n_1_4;
   wire FINAL_RESULT_adder_n_1_5;
   wire FINAL_RESULT_adder_n_1_6;
   wire FINAL_RESULT_adder_n_1_7;
   wire FINAL_RESULT_adder_n_1_9;
   wire FINAL_RESULT_adder_n_1_10;
   wire FINAL_RESULT_adder_n_1_11;
   wire FINAL_RESULT_adder_n_1_12;
   wire FINAL_RESULT_adder_n_1_13;
   wire FINAL_RESULT_adder_n_1_14;
   wire FINAL_RESULT_adder_n_1_15;
   wire FINAL_RESULT_adder_n_1_16;
   wire FINAL_RESULT_adder_n_1_17;
   wire FINAL_RESULT_adder_n_1_18;
   wire FINAL_RESULT_adder_n_1_19;
   wire FINAL_RESULT_adder_n_1_34;
   wire FINAL_RESULT_adder_n_1_35;
   wire FINAL_RESULT_adder_n_1_36;
   wire FINAL_RESULT_adder_n_1_37;
   wire FINAL_RESULT_adder_n_1_45;
   wire FINAL_RESULT_adder_i_1_n_0;
   wire FINAL_RESULT_adder_n_1_38;
   wire FINAL_RESULT_adder_i_1_n_1;
   wire FINAL_RESULT_adder_n_1_40;
   wire FINAL_RESULT_adder_i_1_n_2;
   wire FINAL_RESULT_adder_n_1_43;
   wire FINAL_RESULT_adder_i_1_n_3;
   wire FINAL_RESULT_adder_i_1_n_4;
   wire FINAL_RESULT_adder_i_1_n_5;
   wire FINAL_RESULT_adder_n_1_20;
   wire FINAL_RESULT_adder_i_1_n_6;
   wire FINAL_RESULT_adder_n_1_23;
   wire FINAL_RESULT_adder_i_1_n_7;
   wire FINAL_RESULT_adder_i_1_n_8;
   wire FINAL_RESULT_adder_n_1_25;
   wire FINAL_RESULT_adder_i_1_n_9;
   wire FINAL_RESULT_adder_n_1_29;
   wire FINAL_RESULT_adder_i_1_n_10;
   wire FINAL_RESULT_adder_i_1_n_11;
   wire FINAL_RESULT_adder_n_1_32;
   wire FINAL_RESULT_adder_i_1_n_12;
   wire [19:0]VEC1_VEC2_adder_tempIn22;
   wire [19:0]VEC1_VEC2_adder_tempIn11;
   wire [15:0]Addition_Result;
   wire VEC1_VEC2_adder_n_0;
   wire VEC1_VEC2_adder_n_1;
   wire VEC1_VEC2_adder_n_2;
   wire VEC1_VEC2_adder_n_3;
   wire VEC1_VEC2_adder_n_4;
   wire VEC1_VEC2_adder_n_0_0;
   wire VEC1_VEC2_adder_n_5;
   wire VEC1_VEC2_adder_n_0_1;
   wire VEC1_VEC2_adder_n_0_2;
   wire VEC1_VEC2_adder_n_0_3;
   wire VEC1_VEC2_adder_n_6;
   wire VEC1_VEC2_adder_n_0_4;
   wire VEC1_VEC2_adder_n_0_5;
   wire VEC1_VEC2_adder_n_0_6;
   wire VEC1_VEC2_adder_n_7;
   wire VEC1_VEC2_adder_n_0_7;
   wire VEC1_VEC2_adder_n_0_8;
   wire VEC1_VEC2_adder_n_0_9;
   wire VEC1_VEC2_adder_n_8;
   wire VEC1_VEC2_adder_n_0_10;
   wire VEC1_VEC2_adder_n_0_11;
   wire VEC1_VEC2_adder_n_0_12;
   wire VEC1_VEC2_adder_n_9;
   wire VEC1_VEC2_adder_n_0_13;
   wire VEC1_VEC2_adder_n_0_14;
   wire VEC1_VEC2_adder_n_0_15;
   wire VEC1_VEC2_adder_n_10;
   wire VEC1_VEC2_adder_n_0_16;
   wire VEC1_VEC2_adder_n_0_17;
   wire VEC1_VEC2_adder_n_0_18;
   wire VEC1_VEC2_adder_n_0_19;
   wire VEC1_VEC2_adder_n_11;
   wire VEC1_VEC2_adder_n_0_20;
   wire VEC1_VEC2_adder_n_0_21;
   wire VEC1_VEC2_adder_n_0_22;
   wire VEC1_VEC2_adder_n_0_23;
   wire VEC1_VEC2_adder_n_12;
   wire VEC1_VEC2_adder_n_0_24;
   wire VEC1_VEC2_adder_n_0_25;
   wire VEC1_VEC2_adder_n_0_26;
   wire VEC1_VEC2_adder_n_0_27;
   wire VEC1_VEC2_adder_n_0_28;
   wire VEC1_VEC2_adder_n_0_29;
   wire VEC1_VEC2_adder_n_0_30;
   wire VEC1_VEC2_adder_n_0_31;
   wire VEC1_VEC2_adder_n_0_32;
   wire VEC1_VEC2_adder_n_0_33;
   wire VEC1_VEC2_adder_n_14;
   wire VEC1_VEC2_adder_n_15;
   wire VEC1_VEC2_adder_n_16;
   wire VEC1_VEC2_adder_n_17;
   wire VEC1_VEC2_adder_n_18;
   wire VEC1_VEC2_adder_n_0_34;
   wire VEC1_VEC2_adder_n_19;
   wire VEC1_VEC2_adder_n_0_35;
   wire VEC1_VEC2_adder_n_0_36;
   wire VEC1_VEC2_adder_n_0_37;
   wire VEC1_VEC2_adder_n_20;
   wire VEC1_VEC2_adder_n_0_38;
   wire VEC1_VEC2_adder_n_0_39;
   wire VEC1_VEC2_adder_n_0_40;
   wire VEC1_VEC2_adder_n_21;
   wire VEC1_VEC2_adder_n_0_41;
   wire VEC1_VEC2_adder_n_0_42;
   wire VEC1_VEC2_adder_n_0_43;
   wire VEC1_VEC2_adder_n_22;
   wire VEC1_VEC2_adder_n_0_44;
   wire VEC1_VEC2_adder_n_0_45;
   wire VEC1_VEC2_adder_n_0_46;
   wire VEC1_VEC2_adder_n_23;
   wire VEC1_VEC2_adder_n_0_47;
   wire VEC1_VEC2_adder_n_0_48;
   wire VEC1_VEC2_adder_n_0_49;
   wire VEC1_VEC2_adder_n_24;
   wire VEC1_VEC2_adder_n_0_50;
   wire VEC1_VEC2_adder_n_0_51;
   wire VEC1_VEC2_adder_n_0_52;
   wire VEC1_VEC2_adder_n_0_53;
   wire VEC1_VEC2_adder_n_25;
   wire VEC1_VEC2_adder_n_0_54;
   wire VEC1_VEC2_adder_n_0_55;
   wire VEC1_VEC2_adder_n_0_56;
   wire VEC1_VEC2_adder_n_0_57;
   wire VEC1_VEC2_adder_n_26;
   wire VEC1_VEC2_adder_n_0_58;
   wire VEC1_VEC2_adder_n_0_59;
   wire VEC1_VEC2_adder_n_0_60;
   wire VEC1_VEC2_adder_n_0_61;
   wire VEC1_VEC2_adder_n_0_62;
   wire VEC1_VEC2_adder_n_0_63;
   wire VEC1_VEC2_adder_n_0_64;
   wire VEC1_VEC2_adder_n_0_65;
   wire VEC1_VEC2_adder_n_0_66;
   wire VEC1_VEC2_adder_n_0_67;
   wire VEC1_VEC2_adder_n_0_68;
   wire VEC1_VEC2_adder_n_0_69;
   wire VEC1_VEC2_adder_n_0_70;
   wire VEC1_VEC2_adder_n_27;
   wire VEC1_VEC2_adder_n_0_71;
   wire VEC1_VEC2_adder_n_0_72;
   wire VEC1_VEC2_adder_n_0_73;
   wire VEC1_VEC2_adder_n_0_74;
   wire VEC1_VEC2_adder_n_0_75;
   wire VEC1_VEC2_adder_n_0_76;
   wire VEC1_VEC2_adder_n_0_77;
   wire VEC1_VEC2_adder_n_0_78;
   wire VEC1_VEC2_adder_n_0_79;
   wire VEC1_VEC2_adder_n_0_80;
   wire VEC1_VEC2_adder_n_0_81;
   wire VEC1_VEC2_adder_n_13;
   wire VEC1_VEC2_adder_n_0_82;
   wire VEC1_VEC2_adder_n_0_83;
   wire VEC1_VEC2_adder_n_0_84;
   wire VEC1_VEC2_adder_n_0_85;
   wire VEC1_VEC2_adder_n_0_86;
   wire VEC1_VEC2_adder_n_0_87;
   wire VEC1_VEC2_adder_n_0_88;
   wire VEC1_VEC2_adder_n_0_89;
   wire VEC1_VEC2_adder_n_0_90;
   wire VEC1_VEC2_adder_n_0_91;
   wire VEC1_VEC2_adder_n_0_92;
   wire VEC1_VEC2_adder_n_0_93;
   wire VEC1_VEC2_adder_n_0_94;
   wire VEC1_VEC2_adder_n_1_0;
   wire VEC1_VEC2_adder_n_1_1;
   wire VEC1_VEC2_adder_n_1_3;
   wire VEC1_VEC2_adder_n_1_4;
   wire VEC1_VEC2_adder_n_1_5;
   wire VEC1_VEC2_adder_n_1_6;
   wire VEC1_VEC2_adder_n_1_7;
   wire VEC1_VEC2_adder_n_1_9;
   wire VEC1_VEC2_adder_n_1_10;
   wire VEC1_VEC2_adder_n_1_11;
   wire VEC1_VEC2_adder_n_1_12;
   wire VEC1_VEC2_adder_n_1_13;
   wire VEC1_VEC2_adder_n_1_14;
   wire VEC1_VEC2_adder_n_1_15;
   wire VEC1_VEC2_adder_n_1_16;
   wire VEC1_VEC2_adder_n_1_17;
   wire VEC1_VEC2_adder_n_1_18;
   wire VEC1_VEC2_adder_n_1_19;
   wire VEC1_VEC2_adder_n_1_34;
   wire VEC1_VEC2_adder_n_1_35;
   wire VEC1_VEC2_adder_n_1_36;
   wire VEC1_VEC2_adder_n_1_37;
   wire VEC1_VEC2_adder_n_1_45;
   wire VEC1_VEC2_adder_i_1_n_0;
   wire VEC1_VEC2_adder_n_1_38;
   wire VEC1_VEC2_adder_i_1_n_1;
   wire VEC1_VEC2_adder_n_1_40;
   wire VEC1_VEC2_adder_i_1_n_2;
   wire VEC1_VEC2_adder_n_1_43;
   wire VEC1_VEC2_adder_i_1_n_3;
   wire VEC1_VEC2_adder_i_1_n_4;
   wire VEC1_VEC2_adder_i_1_n_5;
   wire VEC1_VEC2_adder_n_1_20;
   wire VEC1_VEC2_adder_i_1_n_6;
   wire VEC1_VEC2_adder_n_1_23;
   wire VEC1_VEC2_adder_i_1_n_7;
   wire VEC1_VEC2_adder_i_1_n_8;
   wire VEC1_VEC2_adder_n_1_25;
   wire VEC1_VEC2_adder_i_1_n_9;
   wire VEC1_VEC2_adder_n_1_29;
   wire VEC1_VEC2_adder_i_1_n_10;
   wire VEC1_VEC2_adder_i_1_n_11;
   wire VEC1_VEC2_adder_n_1_32;
   wire VEC1_VEC2_adder_i_1_n_12;
   wire [15:0]Element_Result;
   wire [15:0]RESULT_ADD;
   wire [15:0]VECTOR_ADD;
   wire [15:0]VECTOR2_ADD;
   wire [15:0]MATRIX_ADD;
   wire n_0_1;
   wire [15:0]MATRIX_CNT;
   wire [15:0]VECTOR_CNT;
   wire [2:0]state;
   wire [2:0]next;
   wire [1:0]counter;
   wire Matrix_Multiplication1_Enable;
   wire Matrix_Multiplication2_Enable;
   wire Final_Calc_Enable;
   wire Back;
   wire [63:0]n_val;
   wire [63:0]m_val;
   wire [19:0]ELEMENT_adder_tempIn22;
   wire [19:0]ELEMENT_adder_tempIn11;
   wire [15:0]NEW_Element_Result;
   wire ELEMENT_adder_n_0;
   wire ELEMENT_adder_n_1;
   wire ELEMENT_adder_n_2;
   wire ELEMENT_adder_n_3;
   wire ELEMENT_adder_n_4;
   wire ELEMENT_adder_n_0_0;
   wire ELEMENT_adder_n_5;
   wire ELEMENT_adder_n_0_1;
   wire ELEMENT_adder_n_0_2;
   wire ELEMENT_adder_n_0_3;
   wire ELEMENT_adder_n_6;
   wire ELEMENT_adder_n_0_4;
   wire ELEMENT_adder_n_0_5;
   wire ELEMENT_adder_n_0_6;
   wire ELEMENT_adder_n_7;
   wire ELEMENT_adder_n_0_7;
   wire ELEMENT_adder_n_0_8;
   wire ELEMENT_adder_n_0_9;
   wire ELEMENT_adder_n_8;
   wire ELEMENT_adder_n_0_10;
   wire ELEMENT_adder_n_0_11;
   wire ELEMENT_adder_n_0_12;
   wire ELEMENT_adder_n_9;
   wire ELEMENT_adder_n_0_13;
   wire ELEMENT_adder_n_0_14;
   wire ELEMENT_adder_n_0_15;
   wire ELEMENT_adder_n_10;
   wire ELEMENT_adder_n_0_16;
   wire ELEMENT_adder_n_0_17;
   wire ELEMENT_adder_n_0_18;
   wire ELEMENT_adder_n_0_19;
   wire ELEMENT_adder_n_11;
   wire ELEMENT_adder_n_0_20;
   wire ELEMENT_adder_n_0_21;
   wire ELEMENT_adder_n_0_22;
   wire ELEMENT_adder_n_0_23;
   wire ELEMENT_adder_n_12;
   wire ELEMENT_adder_n_0_24;
   wire ELEMENT_adder_n_0_25;
   wire ELEMENT_adder_n_0_26;
   wire ELEMENT_adder_n_0_27;
   wire ELEMENT_adder_n_0_28;
   wire ELEMENT_adder_n_0_29;
   wire ELEMENT_adder_n_0_30;
   wire ELEMENT_adder_n_0_31;
   wire ELEMENT_adder_n_0_32;
   wire ELEMENT_adder_n_0_33;
   wire ELEMENT_adder_n_14;
   wire ELEMENT_adder_n_15;
   wire ELEMENT_adder_n_16;
   wire ELEMENT_adder_n_17;
   wire ELEMENT_adder_n_18;
   wire ELEMENT_adder_n_0_34;
   wire ELEMENT_adder_n_19;
   wire ELEMENT_adder_n_0_35;
   wire ELEMENT_adder_n_0_36;
   wire ELEMENT_adder_n_0_37;
   wire ELEMENT_adder_n_20;
   wire ELEMENT_adder_n_0_38;
   wire ELEMENT_adder_n_0_39;
   wire ELEMENT_adder_n_0_40;
   wire ELEMENT_adder_n_21;
   wire ELEMENT_adder_n_0_41;
   wire ELEMENT_adder_n_0_42;
   wire ELEMENT_adder_n_0_43;
   wire ELEMENT_adder_n_22;
   wire ELEMENT_adder_n_0_44;
   wire ELEMENT_adder_n_0_45;
   wire ELEMENT_adder_n_0_46;
   wire ELEMENT_adder_n_23;
   wire ELEMENT_adder_n_0_47;
   wire ELEMENT_adder_n_0_48;
   wire ELEMENT_adder_n_0_49;
   wire ELEMENT_adder_n_24;
   wire ELEMENT_adder_n_0_50;
   wire ELEMENT_adder_n_0_51;
   wire ELEMENT_adder_n_0_52;
   wire ELEMENT_adder_n_0_53;
   wire ELEMENT_adder_n_25;
   wire ELEMENT_adder_n_0_54;
   wire ELEMENT_adder_n_0_55;
   wire ELEMENT_adder_n_0_56;
   wire ELEMENT_adder_n_0_57;
   wire ELEMENT_adder_n_26;
   wire ELEMENT_adder_n_0_58;
   wire ELEMENT_adder_n_0_59;
   wire ELEMENT_adder_n_0_60;
   wire ELEMENT_adder_n_0_61;
   wire ELEMENT_adder_n_0_62;
   wire ELEMENT_adder_n_0_63;
   wire ELEMENT_adder_n_0_64;
   wire ELEMENT_adder_n_0_65;
   wire ELEMENT_adder_n_0_66;
   wire ELEMENT_adder_n_0_67;
   wire ELEMENT_adder_n_0_68;
   wire ELEMENT_adder_n_0_69;
   wire ELEMENT_adder_n_0_70;
   wire ELEMENT_adder_n_27;
   wire ELEMENT_adder_n_0_71;
   wire ELEMENT_adder_n_0_72;
   wire ELEMENT_adder_n_0_73;
   wire ELEMENT_adder_n_0_74;
   wire ELEMENT_adder_n_0_75;
   wire ELEMENT_adder_n_0_76;
   wire ELEMENT_adder_n_0_77;
   wire ELEMENT_adder_n_0_78;
   wire ELEMENT_adder_n_0_79;
   wire ELEMENT_adder_n_0_80;
   wire ELEMENT_adder_n_0_81;
   wire ELEMENT_adder_n_13;
   wire ELEMENT_adder_n_0_82;
   wire ELEMENT_adder_n_0_83;
   wire ELEMENT_adder_n_0_84;
   wire ELEMENT_adder_n_0_85;
   wire ELEMENT_adder_n_0_86;
   wire ELEMENT_adder_n_0_87;
   wire ELEMENT_adder_n_0_88;
   wire ELEMENT_adder_n_0_89;
   wire ELEMENT_adder_n_0_90;
   wire ELEMENT_adder_n_0_91;
   wire ELEMENT_adder_n_0_92;
   wire ELEMENT_adder_n_0_93;
   wire ELEMENT_adder_n_0_94;
   wire ELEMENT_adder_n_1_0;
   wire ELEMENT_adder_n_1_1;
   wire ELEMENT_adder_n_1_3;
   wire ELEMENT_adder_n_1_4;
   wire ELEMENT_adder_n_1_5;
   wire ELEMENT_adder_n_1_6;
   wire ELEMENT_adder_n_1_7;
   wire ELEMENT_adder_n_1_9;
   wire ELEMENT_adder_n_1_10;
   wire ELEMENT_adder_n_1_11;
   wire ELEMENT_adder_n_1_12;
   wire ELEMENT_adder_n_1_13;
   wire ELEMENT_adder_n_1_14;
   wire ELEMENT_adder_n_1_15;
   wire ELEMENT_adder_n_1_16;
   wire ELEMENT_adder_n_1_17;
   wire ELEMENT_adder_n_1_18;
   wire ELEMENT_adder_n_1_19;
   wire ELEMENT_adder_n_1_34;
   wire ELEMENT_adder_n_1_35;
   wire ELEMENT_adder_n_1_36;
   wire ELEMENT_adder_n_1_37;
   wire ELEMENT_adder_n_1_45;
   wire ELEMENT_adder_i_1_n_0;
   wire ELEMENT_adder_n_1_38;
   wire ELEMENT_adder_i_1_n_1;
   wire ELEMENT_adder_n_1_40;
   wire ELEMENT_adder_i_1_n_2;
   wire ELEMENT_adder_n_1_43;
   wire ELEMENT_adder_i_1_n_3;
   wire ELEMENT_adder_i_1_n_4;
   wire ELEMENT_adder_i_1_n_5;
   wire ELEMENT_adder_n_1_20;
   wire ELEMENT_adder_i_1_n_6;
   wire ELEMENT_adder_n_1_23;
   wire ELEMENT_adder_i_1_n_7;
   wire ELEMENT_adder_i_1_n_8;
   wire ELEMENT_adder_n_1_25;
   wire ELEMENT_adder_i_1_n_9;
   wire ELEMENT_adder_n_1_29;
   wire ELEMENT_adder_i_1_n_10;
   wire ELEMENT_adder_i_1_n_11;
   wire ELEMENT_adder_n_1_32;
   wire ELEMENT_adder_i_1_n_12;
   wire [19:0]VECTOR_CNT_adder_tempIn11;
   wire n_0_0;
   wire VECTOR_CNT_adder_n_25;
   wire VECTOR_CNT_adder_n_26;
   wire n_0_0_0;
   wire VECTOR_CNT_adder_n_27;
   wire n_0_0_1;
   wire n_0_0_2;
   wire VECTOR_CNT_adder_n_29;
   wire n_0_0_6;
   wire n_0_0_8;
   wire VECTOR_CNT_adder_n_31;
   wire n_0_0_12;
   wire VECTOR_CNT_adder_n_19;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire VECTOR_CNT_adder_n_20;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire VECTOR_CNT_adder_n_21;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire VECTOR_CNT_adder_n_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire VECTOR_CNT_adder_n_23;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_2;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_3;
   wire n_0_0_46;
   wire n_0_5;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_6;
   wire n_0_7;
   wire n_0_0_70;
   wire n_0_8;
   wire n_0_0_71;
   wire n_0_9;
   wire n_0_0_72;
   wire n_0_10;
   wire n_0_0_73;
   wire n_0_11;
   wire n_0_0_74;
   wire n_0_12;
   wire n_0_0_75;
   wire n_0_13;
   wire n_0_0_76;
   wire n_0_14;
   wire n_0_0_77;
   wire n_0_15;
   wire n_0_0_78;
   wire n_0_16;
   wire n_0_0_79;
   wire n_0_17;
   wire n_0_0_80;
   wire n_0_18;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_23;
   wire n_0_22;
   wire n_0_4;
   wire n_0_25;
   wire n_0_24;
   wire n_0_26;
   wire n_0_0_92;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_0_93;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_0_94;
   wire n_0_39;
   wire n_0_0_95;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_45;
   wire n_0_44;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_0_120;
   wire n_0_56;
   wire n_0_0_121;
   wire n_0_57;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_58;
   wire n_0_0_125;
   wire n_0_59;
   wire n_0_0_126;
   wire n_0_60;
   wire n_0_0_127;
   wire n_0_61;
   wire n_0_0_128;
   wire n_0_62;
   wire n_0_0_129;
   wire n_0_63;
   wire n_0_0_130;
   wire n_0_64;
   wire n_0_0_131;
   wire n_0_65;
   wire n_0_0_132;
   wire n_0_66;
   wire n_0_0_133;
   wire n_0_67;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_68;
   wire n_0_69;
   wire n_0_0_136;
   wire n_0_70;
   wire n_0_0_137;
   wire n_0_71;
   wire n_0_0_138;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_0_139;
   wire n_0_75;
   wire n_0_0_140;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_0_141;
   wire n_0_103;
   wire n_0_104;
   wire n_0_0_142;
   wire n_0_105;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_0_145;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_0_146;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_118;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_119;
   wire n_0_0_156;
   wire n_0_120;
   wire n_0_0_157;
   wire n_0_121;
   wire n_0_0_158;
   wire n_0_122;
   wire n_0_0_159;
   wire n_0_123;
   wire n_0_0_160;
   wire n_0_124;
   wire n_0_0_161;
   wire n_0_125;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_126;
   wire n_0_0_164;
   wire n_0_127;
   wire n_0_0_165;
   wire n_0_128;
   wire n_0_0_166;
   wire n_0_129;
   wire n_0_0_167;
   wire n_0_130;
   wire n_0_0_168;
   wire n_0_131;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_132;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_0_187;
   wire n_0_136;
   wire n_0_0_188;
   wire n_0_137;
   wire n_0_138;
   wire n_0_0_189;
   wire n_0_139;
   wire n_0_0_190;
   wire n_0_140;
   wire n_0_141;
   wire n_0_0_191;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_0_192;
   wire n_0_149;
   wire n_0_0_193;
   wire n_0_150;
   wire n_0_151;
   wire n_0_0_194;
   wire n_0_152;
   wire n_0_0_195;
   wire n_0_153;
   wire n_0_154;
   wire n_0_0_196;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_46;
   wire n_0_0_197;
   wire n_0_0_199;
   wire n_0_164;
   wire n_0_0_205;
   wire n_0_165;
   wire n_0_0_206;
   wire n_0_166;
   wire n_0_0_207;
   wire n_0_167;
   wire n_0_0_208;
   wire n_0_168;
   wire n_0_0_209;
   wire n_0_169;
   wire n_0_0_210;
   wire n_0_170;
   wire n_0_0_211;
   wire n_0_171;
   wire n_0_0_212;
   wire n_0_172;
   wire n_0_0_213;
   wire n_0_173;
   wire n_0_0_214;
   wire n_0_174;
   wire n_0_0_215;
   wire n_0_175;
   wire n_0_0_216;
   wire n_0_176;
   wire n_0_0_217;
   wire n_0_177;
   wire n_0_0_218;
   wire n_0_178;
   wire n_0_0_219;
   wire n_0_179;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_180;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_47;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_242;
   wire n_0_0_246;
   wire n_0_181;
   wire n_0_0_247;
   wire n_0_182;
   wire n_0_0_248;
   wire n_0_183;
   wire n_0_0_249;
   wire n_0_184;
   wire n_0_0_250;
   wire n_0_185;
   wire n_0_0_251;
   wire n_0_186;
   wire n_0_0_252;
   wire n_0_187;
   wire n_0_0_253;
   wire n_0_188;
   wire n_0_0_254;
   wire n_0_189;
   wire n_0_0_255;
   wire n_0_190;
   wire n_0_0_256;
   wire n_0_191;
   wire n_0_0_257;
   wire n_0_192;
   wire n_0_0_258;
   wire n_0_193;
   wire n_0_0_259;
   wire n_0_194;
   wire n_0_0_260;
   wire n_0_195;
   wire n_0_0_261;
   wire n_0_196;
   wire n_0_0_262;
   wire n_0_197;
   wire n_0_0_263;
   wire n_0_198;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_343;
   wire n_0_0_370;
   wire n_0_0_373;
   wire n_0_0_377;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_0_385;
   wire n_0_0_388;
   wire n_0_0_393;
   wire n_0_199;
   wire n_0_0_394;
   wire n_0_0_396;
   wire n_0_0_397;
   wire n_0_52;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_0_401;
   wire MATRIX_CNT_adder_n_25;
   wire MATRIX_CNT_adder_n_26;
   wire n_0_0_402;
   wire MATRIX_CNT_adder_n_27;
   wire n_0_0_403;
   wire n_0_0_404;
   wire MATRIX_CNT_adder_n_29;
   wire n_0_0_408;
   wire n_0_0_409;
   wire MATRIX_CNT_adder_n_31;
   wire MATRIX_CNT_adder_n_19;
   wire n_0_0_416;
   wire n_0_0_417;
   wire n_0_0_418;
   wire MATRIX_CNT_adder_n_20;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_421;
   wire MATRIX_CNT_adder_n_21;
   wire n_0_0_422;
   wire n_0_0_423;
   wire n_0_0_424;
   wire MATRIX_CNT_adder_n_22;
   wire n_0_0_425;
   wire n_0_0_426;
   wire n_0_0_427;
   wire MATRIX_CNT_adder_n_23;
   wire n_0_0_428;
   wire n_0_0_429;
   wire n_0_0_430;
   wire MATRIX_CNT_adder_n_24;
   wire n_0_0_431;
   wire n_0_0_432;
   wire n_0_0_434;
   wire n_0_0_435;
   wire n_0_0_436;
   wire n_0_0_440;
   wire n_0_0_443;
   wire n_0_0_447;
   wire n_0_0_448;
   wire n_0_0_449;
   wire n_0_0_450;
   wire n_0_0_451;
   wire n_0_0_452;
   wire n_0_0_453;
   wire n_0_0_454;
   wire n_0_0_455;
   wire n_0_0_456;
   wire n_0_0_457;
   wire n_0_0_458;
   wire n_0_0_459;
   wire n_0_0_460;
   wire n_0_0_461;
   wire n_0_0_462;
   wire n_0_0_463;
   wire n_0_0_466;
   wire n_0_0_467;
   wire n_0_0_468;
   wire n_0_0_474;
   wire n_0_0_475;
   wire n_0_0_482;
   wire n_0_0_483;
   wire n_0_0_484;
   wire n_0_0_485;
   wire n_0_0_486;
   wire n_0_0_491;
   wire n_0_0_493;
   wire VECTOR_CNT_adder_n_28;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_7;
   wire n_0_0_9;
   wire VECTOR_CNT_adder_n_2;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_13;
   wire n_0_0_29;
   wire VECTOR_CNT_adder_n_30;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire VECTOR_CNT_adder_n_24;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_198;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_236;
   wire n_0_0_241;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_117;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_336;
   wire n_0_0_342;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_51;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_0_366;
   wire n_0_0_367;
   wire n_0_0_368;
   wire n_0_0_369;
   wire n_0_0_371;
   wire n_0_0_372;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_378;
   wire n_0_0_383;
   wire n_0_0_384;
   wire n_0_0_386;
   wire n_0_0_387;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_0_391;
   wire n_0_0_392;
   wire n_0_0_395;
   wire n_0_0_398;
   wire n_0_0_405;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_0_410;
   wire n_0_0_411;
   wire n_0_0_412;
   wire n_0_0_413;
   wire n_0_0_414;
   wire n_0_0_415;
   wire n_0_0_433;
   wire n_0_0_437;
   wire n_0_0_438;
   wire n_0_0_439;
   wire n_0_0_441;
   wire n_0_0_442;
   wire n_0_0_444;
   wire n_0_0_445;
   wire MATRIX_CNT_adder_n_28;
   wire n_0_0_446;
   wire n_0_0_464;
   wire n_0_0_465;
   wire n_0_0_469;
   wire n_0_0_470;
   wire n_0_0_471;
   wire MATRIX_CNT_adder_n_2;
   wire n_0_0_472;
   wire n_0_0_473;
   wire n_0_0_476;
   wire MATRIX_CNT_adder_n_30;
   wire n_0_0_477;
   wire n_0_0_478;
   wire n_0_0_479;
   wire n_0_0_480;
   wire n_0_0_481;
   wire n_0_0_487;
   wire n_0_0_488;
   wire n_0_0_489;
   wire n_0_0_490;
   wire n_0_0_492;

   assign DONE = 1'b0;
   assign RAM_DATA_WR[63] = 1'b0;
   assign RAM_DATA_WR[62] = 1'b0;
   assign RAM_DATA_WR[61] = 1'b0;
   assign RAM_DATA_WR[60] = 1'b0;
   assign RAM_DATA_WR[59] = 1'b0;
   assign RAM_DATA_WR[58] = 1'b0;
   assign RAM_DATA_WR[57] = 1'b0;
   assign RAM_DATA_WR[56] = 1'b0;
   assign RAM_DATA_WR[55] = 1'b0;
   assign RAM_DATA_WR[54] = 1'b0;
   assign RAM_DATA_WR[53] = 1'b0;
   assign RAM_DATA_WR[52] = 1'b0;
   assign RAM_DATA_WR[51] = 1'b0;
   assign RAM_DATA_WR[50] = 1'b0;
   assign RAM_DATA_WR[49] = 1'b0;
   assign RAM_DATA_WR[48] = 1'b0;
   assign RAM_DATA_WR[47] = 1'b0;
   assign RAM_DATA_WR[46] = 1'b0;
   assign RAM_DATA_WR[45] = 1'b0;
   assign RAM_DATA_WR[44] = 1'b0;
   assign RAM_DATA_WR[43] = 1'b0;
   assign RAM_DATA_WR[42] = 1'b0;
   assign RAM_DATA_WR[41] = 1'b0;
   assign RAM_DATA_WR[40] = 1'b0;
   assign RAM_DATA_WR[39] = 1'b0;
   assign RAM_DATA_WR[38] = 1'b0;
   assign RAM_DATA_WR[37] = 1'b0;
   assign RAM_DATA_WR[36] = 1'b0;
   assign RAM_DATA_WR[35] = 1'b0;
   assign RAM_DATA_WR[34] = 1'b0;
   assign RAM_DATA_WR[33] = 1'b0;
   assign RAM_DATA_WR[32] = 1'b0;
   assign RAM_DATA_WR[31] = 1'b0;
   assign RAM_DATA_WR[30] = 1'b0;
   assign RAM_DATA_WR[29] = 1'b0;
   assign RAM_DATA_WR[28] = 1'b0;
   assign RAM_DATA_WR[27] = 1'b0;
   assign RAM_DATA_WR[26] = 1'b0;
   assign RAM_DATA_WR[25] = 1'b0;
   assign RAM_DATA_WR[24] = 1'b0;
   assign RAM_DATA_WR[23] = 1'b0;
   assign RAM_DATA_WR[22] = 1'b0;
   assign RAM_DATA_WR[21] = 1'b0;
   assign RAM_DATA_WR[20] = 1'b0;
   assign RAM_DATA_WR[19] = 1'b0;
   assign RAM_DATA_WR[18] = 1'b0;
   assign RAM_DATA_WR[17] = 1'b0;
   assign RAM_DATA_WR[16] = 1'b0;

   add_sub_cla__0_283__GU MATRIX_ADD_adder (.enable(), .sub(), .in1(MATRIX_ADD), 
      .in2(), .cin(), .out({uc_0, uc_1, uc_2, NEW_MATRIX_ADD[12], 
      NEW_MATRIX_ADD[11], NEW_MATRIX_ADD[10], NEW_MATRIX_ADD[9], 
      NEW_MATRIX_ADD[8], NEW_MATRIX_ADD[7], NEW_MATRIX_ADD[6], NEW_MATRIX_ADD[5], 
      NEW_MATRIX_ADD[4], NEW_MATRIX_ADD[3], NEW_MATRIX_ADD[2], NEW_MATRIX_ADD[1], 
      NEW_MATRIX_ADD[0]}), .cout(), .invalid());
   add_sub_cla__0_254__GU VECTOR2_ADD_adder (.enable(), .sub(), .in1(VECTOR2_ADD), 
      .in2(), .cin(), .out({uc_3, uc_4, uc_5, NEW_VECTOR2_ADD[12], 
      NEW_VECTOR2_ADD[11], NEW_VECTOR2_ADD[10], NEW_VECTOR2_ADD[9], 
      NEW_VECTOR2_ADD[8], NEW_VECTOR2_ADD[7], NEW_VECTOR2_ADD[6], 
      NEW_VECTOR2_ADD[5], NEW_VECTOR2_ADD[4], NEW_VECTOR2_ADD[3], 
      NEW_VECTOR2_ADD[2], NEW_VECTOR2_ADD[1], NEW_VECTOR2_ADD[0]}), .cout(), 
      .invalid());
   add_sub_cla__GU VECTOR_ADD_adder (.enable(), .sub(), .in1(VECTOR_ADD), .in2(), 
      .cin(), .out({uc_6, uc_7, uc_8, NEW_VECTOR_ADD[12], NEW_VECTOR_ADD[11], 
      NEW_VECTOR_ADD[10], NEW_VECTOR_ADD[9], NEW_VECTOR_ADD[8], 
      NEW_VECTOR_ADD[7], NEW_VECTOR_ADD[6], NEW_VECTOR_ADD[5], NEW_VECTOR_ADD[4], 
      NEW_VECTOR_ADD[3], NEW_VECTOR_ADD[2], NEW_VECTOR_ADD[1], NEW_VECTOR_ADD[0]}), 
      .cout(), .invalid());
   add_sub_cla__0_312__GU RESULT_ADD_adder (.enable(), .sub(), .in1(RESULT_ADD), 
      .in2(), .cin(), .out({uc_9, uc_10, uc_11, NEW_RESULT_ADD[12], 
      NEW_RESULT_ADD[11], NEW_RESULT_ADD[10], NEW_RESULT_ADD[9], 
      NEW_RESULT_ADD[8], NEW_RESULT_ADD[7], NEW_RESULT_ADD[6], NEW_RESULT_ADD[5], 
      NEW_RESULT_ADD[4], NEW_RESULT_ADD[3], NEW_RESULT_ADD[2], NEW_RESULT_ADD[1], 
      NEW_RESULT_ADD[0]}), .cout(), .invalid());
   multiplier_16bit__0_313 h_MUL (.first_operand(Addition_Result), 
      .second_operand({n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, 
      n_11, n_12, n_13, n_14, n_15}), .out(h_VECTOR_RESULT), .enable(), 
      .overflow());
   multiplier_16bit MUL (.first_operand({RAM_DATA_RD1[15], RAM_DATA_RD1[14], 
      RAM_DATA_RD1[13], RAM_DATA_RD1[12], RAM_DATA_RD1[11], RAM_DATA_RD1[10], 
      RAM_DATA_RD1[9], RAM_DATA_RD1[8], RAM_DATA_RD1[7], RAM_DATA_RD1[6], 
      RAM_DATA_RD1[5], RAM_DATA_RD1[4], RAM_DATA_RD1[3], RAM_DATA_RD1[2], 
      RAM_DATA_RD1[1], RAM_DATA_RD1[0]}), .second_operand({RAM_DATA_RD2[15], 
      RAM_DATA_RD2[14], RAM_DATA_RD2[13], RAM_DATA_RD2[12], RAM_DATA_RD2[11], 
      RAM_DATA_RD2[10], RAM_DATA_RD2[9], RAM_DATA_RD2[8], RAM_DATA_RD2[7], 
      RAM_DATA_RD2[6], RAM_DATA_RD2[5], RAM_DATA_RD2[4], RAM_DATA_RD2[3], 
      RAM_DATA_RD2[2], RAM_DATA_RD2[1], RAM_DATA_RD2[0]}), .out(
      Multiplication_Result), .enable(), .overflow());
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[12]  (.D(MATRIX_CNT_adder_n_24), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[12]));
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[11]  (.D(MATRIX_CNT_adder_n_23), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[11]));
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[10]  (.D(MATRIX_CNT_adder_n_22), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[10]));
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[9]  (.D(MATRIX_CNT_adder_n_21), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[9]));
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[8]  (.D(MATRIX_CNT_adder_n_20), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[8]));
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[7]  (.D(MATRIX_CNT_adder_n_19), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[7]));
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[6]  (.D(MATRIX_CNT_adder_n_31), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[6]));
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[5]  (.D(MATRIX_CNT_adder_n_30), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[5]));
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[4]  (.D(MATRIX_CNT_adder_n_29), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[4]));
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[3]  (.D(MATRIX_CNT_adder_n_28), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[3]));
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[2]  (.D(MATRIX_CNT_adder_n_27), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[2]));
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[1]  (.D(MATRIX_CNT_adder_n_26), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[1]));
   DLH_X1 \MATRIX_CNT_adder_tempIn11_reg[0]  (.D(MATRIX_CNT_adder_n_25), 
      .G(MATRIX_CNT_adder_n_2), .Q(MATRIX_CNT_adder_tempIn11[0]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[12]  (.D(FINAL_RESULT_adder_n_26), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[12]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[11]  (.D(FINAL_RESULT_adder_n_25), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[11]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[10]  (.D(FINAL_RESULT_adder_n_24), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[10]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[9]  (.D(FINAL_RESULT_adder_n_23), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[9]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[8]  (.D(FINAL_RESULT_adder_n_22), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[8]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[7]  (.D(FINAL_RESULT_adder_n_21), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[7]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[6]  (.D(FINAL_RESULT_adder_n_20), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[6]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[5]  (.D(FINAL_RESULT_adder_n_19), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[5]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[4]  (.D(FINAL_RESULT_adder_n_18), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[4]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[3]  (.D(FINAL_RESULT_adder_n_17), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[3]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[2]  (.D(FINAL_RESULT_adder_n_16), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[2]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[1]  (.D(FINAL_RESULT_adder_n_15), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[1]));
   DLH_X1 \FINAL_RESULT_adder_tempIn22_reg[0]  (.D(FINAL_RESULT_adder_n_14), 
      .G(FINAL_RESULT_adder_n_27), .Q(FINAL_RESULT_adder_tempIn22[0]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[12]  (.D(FINAL_RESULT_adder_n_12), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[12]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[11]  (.D(FINAL_RESULT_adder_n_11), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[11]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[10]  (.D(FINAL_RESULT_adder_n_10), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[10]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[9]  (.D(FINAL_RESULT_adder_n_9), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[9]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[8]  (.D(FINAL_RESULT_adder_n_8), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[8]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[7]  (.D(FINAL_RESULT_adder_n_7), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[7]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[6]  (.D(FINAL_RESULT_adder_n_6), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[6]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[5]  (.D(FINAL_RESULT_adder_n_5), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[5]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[4]  (.D(FINAL_RESULT_adder_n_4), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[4]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[3]  (.D(FINAL_RESULT_adder_n_3), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[3]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[2]  (.D(FINAL_RESULT_adder_n_2), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[2]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[1]  (.D(FINAL_RESULT_adder_n_1), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[1]));
   DLH_X1 \FINAL_RESULT_adder_tempIn11_reg[0]  (.D(FINAL_RESULT_adder_n_0), 
      .G(FINAL_RESULT_adder_n_13), .Q(FINAL_RESULT_adder_tempIn11[0]));
   OAI22_X1 FINAL_RESULT_adder_i_0_0 (.A1(FINAL_RESULT_adder_n_0_89), .A2(
      FINAL_RESULT_adder_n_13), .B1(FINAL_RESULT_adder_n_0_93), .B2(
      FINAL_RESULT_adder_n_0_82), .ZN(FINAL_RESULT[13]));
   OAI22_X1 FINAL_RESULT_adder_i_0_1 (.A1(FINAL_RESULT_adder_n_0_90), .A2(
      FINAL_RESULT_adder_n_13), .B1(FINAL_RESULT_adder_n_0_94), .B2(
      FINAL_RESULT_adder_n_0_82), .ZN(FINAL_RESULT[14]));
   OR2_X1 FINAL_RESULT_adder_i_0_2 (.A1(Element_Result[15]), .A2(
      h_VECTOR_RESULT[15]), .ZN(FINAL_RESULT[15]));
   AND2_X1 FINAL_RESULT_adder_i_0_3 (.A1(h_VECTOR_RESULT[0]), .A2(
      FINAL_RESULT_adder_n_0_72), .ZN(FINAL_RESULT_adder_n_0));
   OAI22_X1 FINAL_RESULT_adder_i_0_4 (.A1(FINAL_RESULT_adder_n_0_3), .A2(
      FINAL_RESULT_adder_n_0_0), .B1(FINAL_RESULT_adder_n_0_75), .B2(
      FINAL_RESULT_adder_n_0_6), .ZN(FINAL_RESULT_adder_n_1));
   OAI22_X1 FINAL_RESULT_adder_i_0_5 (.A1(FINAL_RESULT_adder_n_0_75), .A2(
      FINAL_RESULT_adder_n_0_9), .B1(FINAL_RESULT_adder_n_0_6), .B2(
      FINAL_RESULT_adder_n_0_0), .ZN(FINAL_RESULT_adder_n_2));
   OAI22_X1 FINAL_RESULT_adder_i_0_6 (.A1(FINAL_RESULT_adder_n_0_75), .A2(
      FINAL_RESULT_adder_n_0_12), .B1(FINAL_RESULT_adder_n_0_9), .B2(
      FINAL_RESULT_adder_n_0_0), .ZN(FINAL_RESULT_adder_n_3));
   OAI22_X1 FINAL_RESULT_adder_i_0_7 (.A1(FINAL_RESULT_adder_n_0_78), .A2(
      FINAL_RESULT_adder_n_0_1), .B1(FINAL_RESULT_adder_n_0_12), .B2(
      FINAL_RESULT_adder_n_0_0), .ZN(FINAL_RESULT_adder_n_4));
   NAND2_X1 FINAL_RESULT_adder_i_0_8 (.A1(FINAL_RESULT_adder_n_0_78), .A2(
      FINAL_RESULT_adder_n_0_77), .ZN(FINAL_RESULT_adder_n_0_0));
   OAI22_X1 FINAL_RESULT_adder_i_0_9 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_1), .B1(FINAL_RESULT_adder_n_0_78), .B2(
      FINAL_RESULT_adder_n_0_4), .ZN(FINAL_RESULT_adder_n_5));
   INV_X1 FINAL_RESULT_adder_i_0_10 (.A(FINAL_RESULT_adder_n_0_2), .ZN(
      FINAL_RESULT_adder_n_0_1));
   OAI22_X1 FINAL_RESULT_adder_i_0_11 (.A1(FINAL_RESULT_adder_n_0_76), .A2(
      FINAL_RESULT_adder_n_0_15), .B1(FINAL_RESULT_adder_n_0_77), .B2(
      FINAL_RESULT_adder_n_0_3), .ZN(FINAL_RESULT_adder_n_0_2));
   NAND2_X1 FINAL_RESULT_adder_i_0_12 (.A1(h_VECTOR_RESULT[0]), .A2(
      FINAL_RESULT_adder_n_0_32), .ZN(FINAL_RESULT_adder_n_0_3));
   OAI22_X1 FINAL_RESULT_adder_i_0_13 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_4), .B1(FINAL_RESULT_adder_n_0_78), .B2(
      FINAL_RESULT_adder_n_0_7), .ZN(FINAL_RESULT_adder_n_6));
   INV_X1 FINAL_RESULT_adder_i_0_14 (.A(FINAL_RESULT_adder_n_0_5), .ZN(
      FINAL_RESULT_adder_n_0_4));
   OAI22_X1 FINAL_RESULT_adder_i_0_15 (.A1(FINAL_RESULT_adder_n_0_76), .A2(
      FINAL_RESULT_adder_n_0_18), .B1(FINAL_RESULT_adder_n_0_77), .B2(
      FINAL_RESULT_adder_n_0_6), .ZN(FINAL_RESULT_adder_n_0_5));
   NAND2_X1 FINAL_RESULT_adder_i_0_16 (.A1(h_VECTOR_RESULT[1]), .A2(
      FINAL_RESULT_adder_n_0_32), .ZN(FINAL_RESULT_adder_n_0_6));
   OAI22_X1 FINAL_RESULT_adder_i_0_17 (.A1(FINAL_RESULT_adder_n_0_78), .A2(
      FINAL_RESULT_adder_n_0_10), .B1(FINAL_RESULT_adder_n_0_79), .B2(
      FINAL_RESULT_adder_n_0_7), .ZN(FINAL_RESULT_adder_n_7));
   INV_X1 FINAL_RESULT_adder_i_0_18 (.A(FINAL_RESULT_adder_n_0_8), .ZN(
      FINAL_RESULT_adder_n_0_7));
   OAI22_X1 FINAL_RESULT_adder_i_0_19 (.A1(FINAL_RESULT_adder_n_0_77), .A2(
      FINAL_RESULT_adder_n_0_9), .B1(FINAL_RESULT_adder_n_0_76), .B2(
      FINAL_RESULT_adder_n_0_22), .ZN(FINAL_RESULT_adder_n_0_8));
   AOI22_X1 FINAL_RESULT_adder_i_0_20 (.A1(h_VECTOR_RESULT[2]), .A2(
      FINAL_RESULT_adder_n_0_32), .B1(h_VECTOR_RESULT[0]), .B2(
      FINAL_RESULT_adder_n_0_33), .ZN(FINAL_RESULT_adder_n_0_9));
   OAI22_X1 FINAL_RESULT_adder_i_0_21 (.A1(FINAL_RESULT_adder_n_0_78), .A2(
      FINAL_RESULT_adder_n_0_13), .B1(FINAL_RESULT_adder_n_0_79), .B2(
      FINAL_RESULT_adder_n_0_10), .ZN(FINAL_RESULT_adder_n_8));
   INV_X1 FINAL_RESULT_adder_i_0_22 (.A(FINAL_RESULT_adder_n_0_11), .ZN(
      FINAL_RESULT_adder_n_0_10));
   OAI22_X1 FINAL_RESULT_adder_i_0_23 (.A1(FINAL_RESULT_adder_n_0_77), .A2(
      FINAL_RESULT_adder_n_0_12), .B1(FINAL_RESULT_adder_n_0_76), .B2(
      FINAL_RESULT_adder_n_0_26), .ZN(FINAL_RESULT_adder_n_0_11));
   AOI22_X1 FINAL_RESULT_adder_i_0_24 (.A1(h_VECTOR_RESULT[3]), .A2(
      FINAL_RESULT_adder_n_0_32), .B1(h_VECTOR_RESULT[1]), .B2(
      FINAL_RESULT_adder_n_0_33), .ZN(FINAL_RESULT_adder_n_0_12));
   OAI22_X1 FINAL_RESULT_adder_i_0_25 (.A1(FINAL_RESULT_adder_n_0_78), .A2(
      FINAL_RESULT_adder_n_0_16), .B1(FINAL_RESULT_adder_n_0_79), .B2(
      FINAL_RESULT_adder_n_0_13), .ZN(FINAL_RESULT_adder_n_9));
   INV_X1 FINAL_RESULT_adder_i_0_26 (.A(FINAL_RESULT_adder_n_0_14), .ZN(
      FINAL_RESULT_adder_n_0_13));
   OAI22_X1 FINAL_RESULT_adder_i_0_27 (.A1(FINAL_RESULT_adder_n_0_77), .A2(
      FINAL_RESULT_adder_n_0_15), .B1(FINAL_RESULT_adder_n_0_76), .B2(
      FINAL_RESULT_adder_n_0_30), .ZN(FINAL_RESULT_adder_n_0_14));
   AOI22_X1 FINAL_RESULT_adder_i_0_28 (.A1(h_VECTOR_RESULT[4]), .A2(
      FINAL_RESULT_adder_n_0_32), .B1(h_VECTOR_RESULT[2]), .B2(
      FINAL_RESULT_adder_n_0_33), .ZN(FINAL_RESULT_adder_n_0_15));
   OAI22_X1 FINAL_RESULT_adder_i_0_29 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_16), .B1(FINAL_RESULT_adder_n_0_78), .B2(
      FINAL_RESULT_adder_n_0_20), .ZN(FINAL_RESULT_adder_n_10));
   INV_X1 FINAL_RESULT_adder_i_0_30 (.A(FINAL_RESULT_adder_n_0_17), .ZN(
      FINAL_RESULT_adder_n_0_16));
   OAI22_X1 FINAL_RESULT_adder_i_0_31 (.A1(FINAL_RESULT_adder_n_0_76), .A2(
      FINAL_RESULT_adder_n_0_19), .B1(FINAL_RESULT_adder_n_0_77), .B2(
      FINAL_RESULT_adder_n_0_18), .ZN(FINAL_RESULT_adder_n_0_17));
   AOI22_X1 FINAL_RESULT_adder_i_0_32 (.A1(h_VECTOR_RESULT[5]), .A2(
      FINAL_RESULT_adder_n_0_32), .B1(h_VECTOR_RESULT[3]), .B2(
      FINAL_RESULT_adder_n_0_33), .ZN(FINAL_RESULT_adder_n_0_18));
   AOI22_X1 FINAL_RESULT_adder_i_0_33 (.A1(h_VECTOR_RESULT[9]), .A2(
      FINAL_RESULT_adder_n_0_32), .B1(h_VECTOR_RESULT[7]), .B2(
      FINAL_RESULT_adder_n_0_33), .ZN(FINAL_RESULT_adder_n_0_19));
   OAI22_X1 FINAL_RESULT_adder_i_0_34 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_20), .B1(FINAL_RESULT_adder_n_0_78), .B2(
      FINAL_RESULT_adder_n_0_24), .ZN(FINAL_RESULT_adder_n_11));
   INV_X1 FINAL_RESULT_adder_i_0_35 (.A(FINAL_RESULT_adder_n_0_21), .ZN(
      FINAL_RESULT_adder_n_0_20));
   OAI22_X1 FINAL_RESULT_adder_i_0_36 (.A1(FINAL_RESULT_adder_n_0_76), .A2(
      FINAL_RESULT_adder_n_0_23), .B1(FINAL_RESULT_adder_n_0_77), .B2(
      FINAL_RESULT_adder_n_0_22), .ZN(FINAL_RESULT_adder_n_0_21));
   AOI22_X1 FINAL_RESULT_adder_i_0_37 (.A1(h_VECTOR_RESULT[6]), .A2(
      FINAL_RESULT_adder_n_0_32), .B1(h_VECTOR_RESULT[4]), .B2(
      FINAL_RESULT_adder_n_0_33), .ZN(FINAL_RESULT_adder_n_0_22));
   AOI22_X1 FINAL_RESULT_adder_i_0_38 (.A1(h_VECTOR_RESULT[10]), .A2(
      FINAL_RESULT_adder_n_0_32), .B1(h_VECTOR_RESULT[8]), .B2(
      FINAL_RESULT_adder_n_0_33), .ZN(FINAL_RESULT_adder_n_0_23));
   OAI22_X1 FINAL_RESULT_adder_i_0_39 (.A1(FINAL_RESULT_adder_n_0_78), .A2(
      FINAL_RESULT_adder_n_0_28), .B1(FINAL_RESULT_adder_n_0_79), .B2(
      FINAL_RESULT_adder_n_0_24), .ZN(FINAL_RESULT_adder_n_12));
   INV_X1 FINAL_RESULT_adder_i_0_40 (.A(FINAL_RESULT_adder_n_0_25), .ZN(
      FINAL_RESULT_adder_n_0_24));
   OAI22_X1 FINAL_RESULT_adder_i_0_41 (.A1(FINAL_RESULT_adder_n_0_76), .A2(
      FINAL_RESULT_adder_n_0_27), .B1(FINAL_RESULT_adder_n_0_77), .B2(
      FINAL_RESULT_adder_n_0_26), .ZN(FINAL_RESULT_adder_n_0_25));
   AOI22_X1 FINAL_RESULT_adder_i_0_42 (.A1(h_VECTOR_RESULT[7]), .A2(
      FINAL_RESULT_adder_n_0_32), .B1(h_VECTOR_RESULT[5]), .B2(
      FINAL_RESULT_adder_n_0_33), .ZN(FINAL_RESULT_adder_n_0_26));
   AOI22_X1 FINAL_RESULT_adder_i_0_43 (.A1(h_VECTOR_RESULT[9]), .A2(
      FINAL_RESULT_adder_n_0_33), .B1(h_VECTOR_RESULT[11]), .B2(
      FINAL_RESULT_adder_n_0_32), .ZN(FINAL_RESULT_adder_n_0_27));
   INV_X1 FINAL_RESULT_adder_i_0_44 (.A(FINAL_RESULT_adder_n_0_29), .ZN(
      FINAL_RESULT_adder_n_0_28));
   OAI22_X1 FINAL_RESULT_adder_i_0_45 (.A1(FINAL_RESULT_adder_n_0_76), .A2(
      FINAL_RESULT_adder_n_0_31), .B1(FINAL_RESULT_adder_n_0_77), .B2(
      FINAL_RESULT_adder_n_0_30), .ZN(FINAL_RESULT_adder_n_0_29));
   AOI22_X1 FINAL_RESULT_adder_i_0_46 (.A1(h_VECTOR_RESULT[8]), .A2(
      FINAL_RESULT_adder_n_0_32), .B1(h_VECTOR_RESULT[6]), .B2(
      FINAL_RESULT_adder_n_0_33), .ZN(FINAL_RESULT_adder_n_0_30));
   AOI22_X1 FINAL_RESULT_adder_i_0_47 (.A1(h_VECTOR_RESULT[10]), .A2(
      FINAL_RESULT_adder_n_0_33), .B1(h_VECTOR_RESULT[12]), .B2(
      FINAL_RESULT_adder_n_0_32), .ZN(FINAL_RESULT_adder_n_0_31));
   INV_X1 FINAL_RESULT_adder_i_0_48 (.A(FINAL_RESULT_adder_n_0_33), .ZN(
      FINAL_RESULT_adder_n_0_32));
   XOR2_X1 FINAL_RESULT_adder_i_0_49 (.A(FINAL_RESULT_adder_n_0_86), .B(
      FINAL_RESULT_adder_n_0_73), .Z(FINAL_RESULT_adder_n_0_33));
   AND2_X1 FINAL_RESULT_adder_i_0_50 (.A1(Element_Result[0]), .A2(
      FINAL_RESULT_adder_n_0_72), .ZN(FINAL_RESULT_adder_n_14));
   OAI22_X1 FINAL_RESULT_adder_i_0_51 (.A1(FINAL_RESULT_adder_n_0_37), .A2(
      FINAL_RESULT_adder_n_0_34), .B1(FINAL_RESULT_adder_n_0_92), .B2(
      FINAL_RESULT_adder_n_0_71), .ZN(FINAL_RESULT_adder_n_15));
   OAI33_X1 FINAL_RESULT_adder_i_0_52 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_69), .A3(FINAL_RESULT_adder_n_0_40), .B1(
      FINAL_RESULT_adder_n_0_78), .B2(FINAL_RESULT_adder_n_0_69), .B3(
      FINAL_RESULT_adder_n_0_43), .ZN(FINAL_RESULT_adder_n_16));
   OAI33_X1 FINAL_RESULT_adder_i_0_53 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_69), .A3(FINAL_RESULT_adder_n_0_43), .B1(
      FINAL_RESULT_adder_n_0_78), .B2(FINAL_RESULT_adder_n_0_69), .B3(
      FINAL_RESULT_adder_n_0_46), .ZN(FINAL_RESULT_adder_n_17));
   OAI22_X1 FINAL_RESULT_adder_i_0_54 (.A1(FINAL_RESULT_adder_n_0_46), .A2(
      FINAL_RESULT_adder_n_0_34), .B1(FINAL_RESULT_adder_n_0_78), .B2(
      FINAL_RESULT_adder_n_0_35), .ZN(FINAL_RESULT_adder_n_18));
   NAND2_X1 FINAL_RESULT_adder_i_0_55 (.A1(FINAL_RESULT_adder_n_0_78), .A2(
      FINAL_RESULT_adder_n_0_68), .ZN(FINAL_RESULT_adder_n_0_34));
   AOI22_X1 FINAL_RESULT_adder_i_0_56 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_38), .B1(FINAL_RESULT_adder_n_0_78), .B2(
      FINAL_RESULT_adder_n_0_35), .ZN(FINAL_RESULT_adder_n_19));
   INV_X1 FINAL_RESULT_adder_i_0_57 (.A(FINAL_RESULT_adder_n_0_36), .ZN(
      FINAL_RESULT_adder_n_0_35));
   OAI22_X1 FINAL_RESULT_adder_i_0_58 (.A1(FINAL_RESULT_adder_n_0_69), .A2(
      FINAL_RESULT_adder_n_0_49), .B1(FINAL_RESULT_adder_n_0_68), .B2(
      FINAL_RESULT_adder_n_0_37), .ZN(FINAL_RESULT_adder_n_0_36));
   NAND2_X1 FINAL_RESULT_adder_i_0_59 (.A1(Element_Result[0]), .A2(
      FINAL_RESULT_adder_n_0_67), .ZN(FINAL_RESULT_adder_n_0_37));
   OAI22_X1 FINAL_RESULT_adder_i_0_60 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_38), .B1(FINAL_RESULT_adder_n_0_78), .B2(
      FINAL_RESULT_adder_n_0_41), .ZN(FINAL_RESULT_adder_n_20));
   INV_X1 FINAL_RESULT_adder_i_0_61 (.A(FINAL_RESULT_adder_n_0_39), .ZN(
      FINAL_RESULT_adder_n_0_38));
   OAI22_X1 FINAL_RESULT_adder_i_0_62 (.A1(FINAL_RESULT_adder_n_0_69), .A2(
      FINAL_RESULT_adder_n_0_52), .B1(FINAL_RESULT_adder_n_0_68), .B2(
      FINAL_RESULT_adder_n_0_40), .ZN(FINAL_RESULT_adder_n_0_39));
   NAND2_X1 FINAL_RESULT_adder_i_0_63 (.A1(Element_Result[1]), .A2(
      FINAL_RESULT_adder_n_0_67), .ZN(FINAL_RESULT_adder_n_0_40));
   OAI22_X1 FINAL_RESULT_adder_i_0_64 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_41), .B1(FINAL_RESULT_adder_n_0_78), .B2(
      FINAL_RESULT_adder_n_0_44), .ZN(FINAL_RESULT_adder_n_21));
   INV_X1 FINAL_RESULT_adder_i_0_65 (.A(FINAL_RESULT_adder_n_0_42), .ZN(
      FINAL_RESULT_adder_n_0_41));
   OAI22_X1 FINAL_RESULT_adder_i_0_66 (.A1(FINAL_RESULT_adder_n_0_69), .A2(
      FINAL_RESULT_adder_n_0_56), .B1(FINAL_RESULT_adder_n_0_68), .B2(
      FINAL_RESULT_adder_n_0_43), .ZN(FINAL_RESULT_adder_n_0_42));
   AOI22_X1 FINAL_RESULT_adder_i_0_67 (.A1(Element_Result[2]), .A2(
      FINAL_RESULT_adder_n_0_67), .B1(Element_Result[0]), .B2(
      FINAL_RESULT_adder_n_0_66), .ZN(FINAL_RESULT_adder_n_0_43));
   OAI22_X1 FINAL_RESULT_adder_i_0_68 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_44), .B1(FINAL_RESULT_adder_n_0_78), .B2(
      FINAL_RESULT_adder_n_0_47), .ZN(FINAL_RESULT_adder_n_22));
   INV_X1 FINAL_RESULT_adder_i_0_69 (.A(FINAL_RESULT_adder_n_0_45), .ZN(
      FINAL_RESULT_adder_n_0_44));
   OAI22_X1 FINAL_RESULT_adder_i_0_70 (.A1(FINAL_RESULT_adder_n_0_69), .A2(
      FINAL_RESULT_adder_n_0_60), .B1(FINAL_RESULT_adder_n_0_68), .B2(
      FINAL_RESULT_adder_n_0_46), .ZN(FINAL_RESULT_adder_n_0_45));
   AOI22_X1 FINAL_RESULT_adder_i_0_71 (.A1(Element_Result[3]), .A2(
      FINAL_RESULT_adder_n_0_67), .B1(Element_Result[1]), .B2(
      FINAL_RESULT_adder_n_0_66), .ZN(FINAL_RESULT_adder_n_0_46));
   OAI22_X1 FINAL_RESULT_adder_i_0_72 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_47), .B1(FINAL_RESULT_adder_n_0_78), .B2(
      FINAL_RESULT_adder_n_0_50), .ZN(FINAL_RESULT_adder_n_23));
   INV_X1 FINAL_RESULT_adder_i_0_73 (.A(FINAL_RESULT_adder_n_0_48), .ZN(
      FINAL_RESULT_adder_n_0_47));
   OAI22_X1 FINAL_RESULT_adder_i_0_74 (.A1(FINAL_RESULT_adder_n_0_69), .A2(
      FINAL_RESULT_adder_n_0_64), .B1(FINAL_RESULT_adder_n_0_68), .B2(
      FINAL_RESULT_adder_n_0_49), .ZN(FINAL_RESULT_adder_n_0_48));
   AOI22_X1 FINAL_RESULT_adder_i_0_75 (.A1(Element_Result[4]), .A2(
      FINAL_RESULT_adder_n_0_67), .B1(Element_Result[2]), .B2(
      FINAL_RESULT_adder_n_0_66), .ZN(FINAL_RESULT_adder_n_0_49));
   OAI22_X1 FINAL_RESULT_adder_i_0_76 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_50), .B1(FINAL_RESULT_adder_n_0_78), .B2(
      FINAL_RESULT_adder_n_0_54), .ZN(FINAL_RESULT_adder_n_24));
   INV_X1 FINAL_RESULT_adder_i_0_77 (.A(FINAL_RESULT_adder_n_0_51), .ZN(
      FINAL_RESULT_adder_n_0_50));
   OAI22_X1 FINAL_RESULT_adder_i_0_78 (.A1(FINAL_RESULT_adder_n_0_69), .A2(
      FINAL_RESULT_adder_n_0_53), .B1(FINAL_RESULT_adder_n_0_68), .B2(
      FINAL_RESULT_adder_n_0_52), .ZN(FINAL_RESULT_adder_n_0_51));
   AOI22_X1 FINAL_RESULT_adder_i_0_79 (.A1(Element_Result[5]), .A2(
      FINAL_RESULT_adder_n_0_67), .B1(Element_Result[3]), .B2(
      FINAL_RESULT_adder_n_0_66), .ZN(FINAL_RESULT_adder_n_0_52));
   AOI22_X1 FINAL_RESULT_adder_i_0_80 (.A1(Element_Result[9]), .A2(
      FINAL_RESULT_adder_n_0_67), .B1(Element_Result[7]), .B2(
      FINAL_RESULT_adder_n_0_66), .ZN(FINAL_RESULT_adder_n_0_53));
   OAI22_X1 FINAL_RESULT_adder_i_0_81 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_54), .B1(FINAL_RESULT_adder_n_0_78), .B2(
      FINAL_RESULT_adder_n_0_58), .ZN(FINAL_RESULT_adder_n_25));
   INV_X1 FINAL_RESULT_adder_i_0_82 (.A(FINAL_RESULT_adder_n_0_55), .ZN(
      FINAL_RESULT_adder_n_0_54));
   OAI22_X1 FINAL_RESULT_adder_i_0_83 (.A1(FINAL_RESULT_adder_n_0_69), .A2(
      FINAL_RESULT_adder_n_0_57), .B1(FINAL_RESULT_adder_n_0_68), .B2(
      FINAL_RESULT_adder_n_0_56), .ZN(FINAL_RESULT_adder_n_0_55));
   AOI22_X1 FINAL_RESULT_adder_i_0_84 (.A1(Element_Result[6]), .A2(
      FINAL_RESULT_adder_n_0_67), .B1(Element_Result[4]), .B2(
      FINAL_RESULT_adder_n_0_66), .ZN(FINAL_RESULT_adder_n_0_56));
   AOI22_X1 FINAL_RESULT_adder_i_0_85 (.A1(Element_Result[10]), .A2(
      FINAL_RESULT_adder_n_0_67), .B1(Element_Result[8]), .B2(
      FINAL_RESULT_adder_n_0_66), .ZN(FINAL_RESULT_adder_n_0_57));
   OAI22_X1 FINAL_RESULT_adder_i_0_86 (.A1(FINAL_RESULT_adder_n_0_78), .A2(
      FINAL_RESULT_adder_n_0_62), .B1(FINAL_RESULT_adder_n_0_79), .B2(
      FINAL_RESULT_adder_n_0_58), .ZN(FINAL_RESULT_adder_n_26));
   INV_X1 FINAL_RESULT_adder_i_0_87 (.A(FINAL_RESULT_adder_n_0_59), .ZN(
      FINAL_RESULT_adder_n_0_58));
   OAI22_X1 FINAL_RESULT_adder_i_0_88 (.A1(FINAL_RESULT_adder_n_0_69), .A2(
      FINAL_RESULT_adder_n_0_61), .B1(FINAL_RESULT_adder_n_0_68), .B2(
      FINAL_RESULT_adder_n_0_60), .ZN(FINAL_RESULT_adder_n_0_59));
   AOI22_X1 FINAL_RESULT_adder_i_0_89 (.A1(Element_Result[7]), .A2(
      FINAL_RESULT_adder_n_0_67), .B1(Element_Result[5]), .B2(
      FINAL_RESULT_adder_n_0_66), .ZN(FINAL_RESULT_adder_n_0_60));
   AOI22_X1 FINAL_RESULT_adder_i_0_90 (.A1(Element_Result[9]), .A2(
      FINAL_RESULT_adder_n_0_66), .B1(Element_Result[11]), .B2(
      FINAL_RESULT_adder_n_0_67), .ZN(FINAL_RESULT_adder_n_0_61));
   INV_X1 FINAL_RESULT_adder_i_0_91 (.A(FINAL_RESULT_adder_n_0_63), .ZN(
      FINAL_RESULT_adder_n_0_62));
   OAI22_X1 FINAL_RESULT_adder_i_0_92 (.A1(FINAL_RESULT_adder_n_0_69), .A2(
      FINAL_RESULT_adder_n_0_65), .B1(FINAL_RESULT_adder_n_0_68), .B2(
      FINAL_RESULT_adder_n_0_64), .ZN(FINAL_RESULT_adder_n_0_63));
   AOI22_X1 FINAL_RESULT_adder_i_0_93 (.A1(Element_Result[8]), .A2(
      FINAL_RESULT_adder_n_0_67), .B1(Element_Result[6]), .B2(
      FINAL_RESULT_adder_n_0_66), .ZN(FINAL_RESULT_adder_n_0_64));
   AOI22_X1 FINAL_RESULT_adder_i_0_94 (.A1(Element_Result[10]), .A2(
      FINAL_RESULT_adder_n_0_66), .B1(Element_Result[12]), .B2(
      FINAL_RESULT_adder_n_0_67), .ZN(FINAL_RESULT_adder_n_0_65));
   INV_X1 FINAL_RESULT_adder_i_0_95 (.A(FINAL_RESULT_adder_n_0_67), .ZN(
      FINAL_RESULT_adder_n_0_66));
   OAI22_X1 FINAL_RESULT_adder_i_0_96 (.A1(FINAL_RESULT_adder_n_0_81), .A2(
      FINAL_RESULT_adder_n_0_73), .B1(FINAL_RESULT_adder_n_0_80), .B2(
      FINAL_RESULT_adder_n_0_74), .ZN(FINAL_RESULT_adder_n_0_67));
   INV_X1 FINAL_RESULT_adder_i_0_97 (.A(FINAL_RESULT_adder_n_0_69), .ZN(
      FINAL_RESULT_adder_n_0_68));
   XOR2_X1 FINAL_RESULT_adder_i_0_98 (.A(FINAL_RESULT_adder_n_0_83), .B(
      FINAL_RESULT_adder_n_0_70), .Z(FINAL_RESULT_adder_n_0_69));
   AOI21_X1 FINAL_RESULT_adder_i_0_99 (.A(FINAL_RESULT_adder_n_0_85), .B1(
      FINAL_RESULT_adder_n_0_87), .B2(FINAL_RESULT_adder_n_0_80), .ZN(
      FINAL_RESULT_adder_n_0_70));
   NAND2_X1 FINAL_RESULT_adder_i_0_100 (.A1(FINAL_RESULT_adder_n_13), .A2(
      FINAL_RESULT_adder_n_0_71), .ZN(FINAL_RESULT_adder_n_27));
   INV_X1 FINAL_RESULT_adder_i_0_101 (.A(FINAL_RESULT_adder_n_0_72), .ZN(
      FINAL_RESULT_adder_n_0_71));
   NOR2_X1 FINAL_RESULT_adder_i_0_102 (.A1(FINAL_RESULT_adder_n_0_75), .A2(
      FINAL_RESULT_adder_n_0_73), .ZN(FINAL_RESULT_adder_n_0_72));
   INV_X1 FINAL_RESULT_adder_i_0_103 (.A(FINAL_RESULT_adder_n_0_74), .ZN(
      FINAL_RESULT_adder_n_0_73));
   NOR2_X1 FINAL_RESULT_adder_i_0_104 (.A1(FINAL_RESULT_adder_n_0_88), .A2(
      FINAL_RESULT_adder_n_0_85), .ZN(FINAL_RESULT_adder_n_0_74));
   NAND2_X1 FINAL_RESULT_adder_i_0_105 (.A1(FINAL_RESULT_adder_n_0_79), .A2(
      FINAL_RESULT_adder_n_0_77), .ZN(FINAL_RESULT_adder_n_0_75));
   INV_X1 FINAL_RESULT_adder_i_0_106 (.A(FINAL_RESULT_adder_n_0_77), .ZN(
      FINAL_RESULT_adder_n_0_76));
   XOR2_X1 FINAL_RESULT_adder_i_0_107 (.A(FINAL_RESULT_adder_n_0_84), .B(
      FINAL_RESULT_adder_n_0_83), .Z(FINAL_RESULT_adder_n_0_77));
   INV_X1 FINAL_RESULT_adder_i_0_108 (.A(FINAL_RESULT_adder_n_0_79), .ZN(
      FINAL_RESULT_adder_n_0_78));
   NOR2_X1 FINAL_RESULT_adder_i_0_109 (.A1(FINAL_RESULT_adder_n_0_86), .A2(
      FINAL_RESULT_adder_n_0_81), .ZN(FINAL_RESULT_adder_n_0_79));
   INV_X1 FINAL_RESULT_adder_i_0_110 (.A(FINAL_RESULT_adder_n_0_81), .ZN(
      FINAL_RESULT_adder_n_0_80));
   NOR2_X1 FINAL_RESULT_adder_i_0_111 (.A1(FINAL_RESULT_adder_n_0_93), .A2(
      h_VECTOR_RESULT[13]), .ZN(FINAL_RESULT_adder_n_0_81));
   INV_X1 FINAL_RESULT_adder_i_0_112 (.A(FINAL_RESULT_adder_n_0_82), .ZN(
      FINAL_RESULT_adder_n_13));
   OAI22_X1 FINAL_RESULT_adder_i_0_113 (.A1(Element_Result[15]), .A2(
      FINAL_RESULT_adder_n_0_91), .B1(FINAL_RESULT_adder_n_0_84), .B2(
      FINAL_RESULT_adder_n_0_83), .ZN(FINAL_RESULT_adder_n_0_82));
   XNOR2_X1 FINAL_RESULT_adder_i_0_114 (.A(Element_Result[15]), .B(
      FINAL_RESULT_adder_n_0_91), .ZN(FINAL_RESULT_adder_n_0_83));
   OAI21_X1 FINAL_RESULT_adder_i_0_115 (.A(FINAL_RESULT_adder_n_0_87), .B1(
      FINAL_RESULT_adder_n_0_86), .B2(FINAL_RESULT_adder_n_0_85), .ZN(
      FINAL_RESULT_adder_n_0_84));
   NOR2_X1 FINAL_RESULT_adder_i_0_116 (.A1(Element_Result[14]), .A2(
      FINAL_RESULT_adder_n_0_90), .ZN(FINAL_RESULT_adder_n_0_85));
   NOR2_X1 FINAL_RESULT_adder_i_0_117 (.A1(Element_Result[13]), .A2(
      FINAL_RESULT_adder_n_0_89), .ZN(FINAL_RESULT_adder_n_0_86));
   INV_X1 FINAL_RESULT_adder_i_0_118 (.A(FINAL_RESULT_adder_n_0_88), .ZN(
      FINAL_RESULT_adder_n_0_87));
   NOR2_X1 FINAL_RESULT_adder_i_0_119 (.A1(FINAL_RESULT_adder_n_0_94), .A2(
      h_VECTOR_RESULT[14]), .ZN(FINAL_RESULT_adder_n_0_88));
   INV_X1 FINAL_RESULT_adder_i_0_120 (.A(h_VECTOR_RESULT[13]), .ZN(
      FINAL_RESULT_adder_n_0_89));
   INV_X1 FINAL_RESULT_adder_i_0_121 (.A(h_VECTOR_RESULT[14]), .ZN(
      FINAL_RESULT_adder_n_0_90));
   INV_X1 FINAL_RESULT_adder_i_0_122 (.A(h_VECTOR_RESULT[15]), .ZN(
      FINAL_RESULT_adder_n_0_91));
   INV_X1 FINAL_RESULT_adder_i_0_123 (.A(Element_Result[1]), .ZN(
      FINAL_RESULT_adder_n_0_92));
   INV_X1 FINAL_RESULT_adder_i_0_124 (.A(Element_Result[13]), .ZN(
      FINAL_RESULT_adder_n_0_93));
   INV_X1 FINAL_RESULT_adder_i_0_125 (.A(Element_Result[14]), .ZN(
      FINAL_RESULT_adder_n_0_94));
   XOR2_X1 FINAL_RESULT_adder_i_1_0 (.A(FINAL_RESULT_adder_tempIn22[0]), 
      .B(FINAL_RESULT_adder_tempIn11[0]), .Z(FINAL_RESULT[0]));
   XNOR2_X1 FINAL_RESULT_adder_i_1_1 (.A(FINAL_RESULT_adder_n_1_43), .B(
      FINAL_RESULT_adder_n_1_0), .ZN(FINAL_RESULT[1]));
   XOR2_X1 FINAL_RESULT_adder_i_1_2 (.A(FINAL_RESULT_adder_tempIn22[1]), 
      .B(FINAL_RESULT_adder_tempIn11[1]), .Z(FINAL_RESULT_adder_n_1_0));
   XNOR2_X1 FINAL_RESULT_adder_i_1_3 (.A(FINAL_RESULT_adder_n_1_40), .B(
      FINAL_RESULT_adder_n_1_1), .ZN(FINAL_RESULT[2]));
   XNOR2_X1 FINAL_RESULT_adder_i_1_4 (.A(FINAL_RESULT_adder_tempIn22[2]), 
      .B(FINAL_RESULT_adder_tempIn11[2]), .ZN(FINAL_RESULT_adder_n_1_1));
   XNOR2_X1 FINAL_RESULT_adder_i_1_7 (.A(FINAL_RESULT_adder_n_1_35), .B(
      FINAL_RESULT_adder_n_1_3), .ZN(FINAL_RESULT[4]));
   XNOR2_X1 FINAL_RESULT_adder_i_1_8 (.A(FINAL_RESULT_adder_tempIn22[4]), 
      .B(FINAL_RESULT_adder_tempIn11[4]), .ZN(FINAL_RESULT_adder_n_1_3));
   XNOR2_X1 FINAL_RESULT_adder_i_1_9 (.A(FINAL_RESULT_adder_n_1_32), .B(
      FINAL_RESULT_adder_n_1_4), .ZN(FINAL_RESULT[5]));
   XOR2_X1 FINAL_RESULT_adder_i_1_10 (.A(FINAL_RESULT_adder_tempIn22[5]), 
      .B(FINAL_RESULT_adder_tempIn11[5]), .Z(FINAL_RESULT_adder_n_1_4));
   XNOR2_X1 FINAL_RESULT_adder_i_1_11 (.A(FINAL_RESULT_adder_n_1_29), .B(
      FINAL_RESULT_adder_n_1_5), .ZN(FINAL_RESULT[6]));
   XNOR2_X1 FINAL_RESULT_adder_i_1_12 (.A(FINAL_RESULT_adder_tempIn22[6]), 
      .B(FINAL_RESULT_adder_tempIn11[6]), .ZN(FINAL_RESULT_adder_n_1_5));
   XNOR2_X1 FINAL_RESULT_adder_i_1_13 (.A(FINAL_RESULT_adder_n_1_25), .B(
      FINAL_RESULT_adder_n_1_6), .ZN(FINAL_RESULT[7]));
   XOR2_X1 FINAL_RESULT_adder_i_1_14 (.A(FINAL_RESULT_adder_tempIn22[7]), 
      .B(FINAL_RESULT_adder_tempIn11[7]), .Z(FINAL_RESULT_adder_n_1_6));
   XNOR2_X1 FINAL_RESULT_adder_i_1_15 (.A(FINAL_RESULT_adder_n_1_23), .B(
      FINAL_RESULT_adder_n_1_7), .ZN(FINAL_RESULT[8]));
   XNOR2_X1 FINAL_RESULT_adder_i_1_16 (.A(FINAL_RESULT_adder_tempIn22[8]), 
      .B(FINAL_RESULT_adder_tempIn11[8]), .ZN(FINAL_RESULT_adder_n_1_7));
   XNOR2_X1 FINAL_RESULT_adder_i_1_19 (.A(FINAL_RESULT_adder_n_1_17), .B(
      FINAL_RESULT_adder_n_1_9), .ZN(FINAL_RESULT[10]));
   XNOR2_X1 FINAL_RESULT_adder_i_1_20 (.A(FINAL_RESULT_adder_tempIn22[10]), 
      .B(FINAL_RESULT_adder_tempIn11[10]), .ZN(FINAL_RESULT_adder_n_1_9));
   XNOR2_X1 FINAL_RESULT_adder_i_1_21 (.A(FINAL_RESULT_adder_n_1_14), .B(
      FINAL_RESULT_adder_n_1_10), .ZN(FINAL_RESULT[11]));
   XOR2_X1 FINAL_RESULT_adder_i_1_22 (.A(FINAL_RESULT_adder_tempIn22[11]), 
      .B(FINAL_RESULT_adder_tempIn11[11]), .Z(FINAL_RESULT_adder_n_1_10));
   XNOR2_X1 FINAL_RESULT_adder_i_1_23 (.A(FINAL_RESULT_adder_n_1_45), .B(
      FINAL_RESULT_adder_n_1_11), .ZN(FINAL_RESULT[12]));
   OAI21_X1 FINAL_RESULT_adder_i_1_24 (.A(FINAL_RESULT_adder_n_1_12), .B1(
      FINAL_RESULT_adder_n_1_14), .B2(FINAL_RESULT_adder_n_1_13), .ZN(
      FINAL_RESULT_adder_n_1_11));
   NAND2_X1 FINAL_RESULT_adder_i_1_25 (.A1(FINAL_RESULT_adder_tempIn22[11]), 
      .A2(FINAL_RESULT_adder_tempIn11[11]), .ZN(FINAL_RESULT_adder_n_1_12));
   NOR2_X1 FINAL_RESULT_adder_i_1_26 (.A1(FINAL_RESULT_adder_tempIn22[11]), 
      .A2(FINAL_RESULT_adder_tempIn11[11]), .ZN(FINAL_RESULT_adder_n_1_13));
   OAI21_X1 FINAL_RESULT_adder_i_1_27 (.A(FINAL_RESULT_adder_n_1_15), .B1(
      FINAL_RESULT_adder_tempIn11[10]), .B2(FINAL_RESULT_adder_tempIn22[10]), 
      .ZN(FINAL_RESULT_adder_n_1_14));
   INV_X1 FINAL_RESULT_adder_i_1_28 (.A(FINAL_RESULT_adder_n_1_16), .ZN(
      FINAL_RESULT_adder_n_1_15));
   AOI21_X1 FINAL_RESULT_adder_i_1_29 (.A(FINAL_RESULT_adder_n_1_17), .B1(
      FINAL_RESULT_adder_tempIn11[10]), .B2(FINAL_RESULT_adder_tempIn22[10]), 
      .ZN(FINAL_RESULT_adder_n_1_16));
   AOI21_X1 FINAL_RESULT_adder_i_1_30 (.A(FINAL_RESULT_adder_n_1_18), .B1(
      FINAL_RESULT_adder_n_1_19), .B2(FINAL_RESULT_adder_n_1_20), .ZN(
      FINAL_RESULT_adder_n_1_17));
   NOR2_X1 FINAL_RESULT_adder_i_1_31 (.A1(FINAL_RESULT_adder_tempIn22[9]), 
      .A2(FINAL_RESULT_adder_tempIn11[9]), .ZN(FINAL_RESULT_adder_n_1_18));
   NAND2_X1 FINAL_RESULT_adder_i_1_32 (.A1(FINAL_RESULT_adder_tempIn22[9]), 
      .A2(FINAL_RESULT_adder_tempIn11[9]), .ZN(FINAL_RESULT_adder_n_1_19));
   AOI21_X1 FINAL_RESULT_adder_i_1_47 (.A(FINAL_RESULT_adder_n_1_35), .B1(
      FINAL_RESULT_adder_tempIn11[4]), .B2(FINAL_RESULT_adder_tempIn22[4]), 
      .ZN(FINAL_RESULT_adder_n_1_34));
   AOI21_X1 FINAL_RESULT_adder_i_1_48 (.A(FINAL_RESULT_adder_n_1_36), .B1(
      FINAL_RESULT_adder_n_1_37), .B2(FINAL_RESULT_adder_n_1_38), .ZN(
      FINAL_RESULT_adder_n_1_35));
   NOR2_X1 FINAL_RESULT_adder_i_1_49 (.A1(FINAL_RESULT_adder_tempIn22[3]), 
      .A2(FINAL_RESULT_adder_tempIn11[3]), .ZN(FINAL_RESULT_adder_n_1_36));
   NAND2_X1 FINAL_RESULT_adder_i_1_50 (.A1(FINAL_RESULT_adder_tempIn22[3]), 
      .A2(FINAL_RESULT_adder_tempIn11[3]), .ZN(FINAL_RESULT_adder_n_1_37));
   XNOR2_X1 FINAL_RESULT_adder_i_1_58 (.A(FINAL_RESULT_adder_tempIn22[12]), 
      .B(FINAL_RESULT_adder_tempIn11[12]), .ZN(FINAL_RESULT_adder_n_1_45));
   XOR2_X1 FINAL_RESULT_adder_i_1_5 (.A(FINAL_RESULT_adder_n_1_38), .B(
      FINAL_RESULT_adder_i_1_n_0), .Z(FINAL_RESULT[3]));
   XNOR2_X1 FINAL_RESULT_adder_i_1_6 (.A(FINAL_RESULT_adder_tempIn22[3]), 
      .B(FINAL_RESULT_adder_tempIn11[3]), .ZN(FINAL_RESULT_adder_i_1_n_0));
   OAI22_X1 FINAL_RESULT_adder_i_1_17 (.A1(FINAL_RESULT_adder_tempIn22[2]), 
      .A2(FINAL_RESULT_adder_tempIn11[2]), .B1(FINAL_RESULT_adder_n_1_40), 
      .B2(FINAL_RESULT_adder_i_1_n_1), .ZN(FINAL_RESULT_adder_n_1_38));
   AND2_X1 FINAL_RESULT_adder_i_1_18 (.A1(FINAL_RESULT_adder_tempIn22[2]), 
      .A2(FINAL_RESULT_adder_tempIn11[2]), .ZN(FINAL_RESULT_adder_i_1_n_1));
   OAI22_X1 FINAL_RESULT_adder_i_1_33 (.A1(FINAL_RESULT_adder_i_1_n_4), .A2(
      FINAL_RESULT_adder_i_1_n_3), .B1(FINAL_RESULT_adder_n_1_43), .B2(
      FINAL_RESULT_adder_i_1_n_2), .ZN(FINAL_RESULT_adder_n_1_40));
   NOR2_X1 FINAL_RESULT_adder_i_1_34 (.A1(FINAL_RESULT_adder_tempIn22[1]), 
      .A2(FINAL_RESULT_adder_tempIn11[1]), .ZN(FINAL_RESULT_adder_i_1_n_2));
   NAND2_X1 FINAL_RESULT_adder_i_1_35 (.A1(FINAL_RESULT_adder_tempIn22[0]), 
      .A2(FINAL_RESULT_adder_tempIn11[0]), .ZN(FINAL_RESULT_adder_n_1_43));
   INV_X1 FINAL_RESULT_adder_i_1_36 (.A(FINAL_RESULT_adder_tempIn11[1]), 
      .ZN(FINAL_RESULT_adder_i_1_n_3));
   INV_X1 FINAL_RESULT_adder_i_1_37 (.A(FINAL_RESULT_adder_tempIn22[1]), 
      .ZN(FINAL_RESULT_adder_i_1_n_4));
   XOR2_X1 FINAL_RESULT_adder_i_1_38 (.A(FINAL_RESULT_adder_n_1_20), .B(
      FINAL_RESULT_adder_i_1_n_5), .Z(FINAL_RESULT[9]));
   XNOR2_X1 FINAL_RESULT_adder_i_1_39 (.A(FINAL_RESULT_adder_tempIn22[9]), 
      .B(FINAL_RESULT_adder_tempIn11[9]), .ZN(FINAL_RESULT_adder_i_1_n_5));
   AOI22_X1 FINAL_RESULT_adder_i_1_40 (.A1(FINAL_RESULT_adder_tempIn22[8]), 
      .A2(FINAL_RESULT_adder_tempIn11[8]), .B1(FINAL_RESULT_adder_n_1_23), 
      .B2(FINAL_RESULT_adder_i_1_n_6), .ZN(FINAL_RESULT_adder_n_1_20));
   OR2_X1 FINAL_RESULT_adder_i_1_41 (.A1(FINAL_RESULT_adder_tempIn22[8]), 
      .A2(FINAL_RESULT_adder_tempIn11[8]), .ZN(FINAL_RESULT_adder_i_1_n_6));
   OAI21_X1 FINAL_RESULT_adder_i_1_42 (.A(FINAL_RESULT_adder_i_1_n_8), .B1(
      FINAL_RESULT_adder_n_1_25), .B2(FINAL_RESULT_adder_i_1_n_7), .ZN(
      FINAL_RESULT_adder_n_1_23));
   NOR2_X1 FINAL_RESULT_adder_i_1_43 (.A1(FINAL_RESULT_adder_tempIn22[7]), 
      .A2(FINAL_RESULT_adder_tempIn11[7]), .ZN(FINAL_RESULT_adder_i_1_n_7));
   NAND2_X1 FINAL_RESULT_adder_i_1_44 (.A1(FINAL_RESULT_adder_tempIn22[7]), 
      .A2(FINAL_RESULT_adder_tempIn11[7]), .ZN(FINAL_RESULT_adder_i_1_n_8));
   AOI22_X1 FINAL_RESULT_adder_i_1_45 (.A1(FINAL_RESULT_adder_tempIn22[6]), 
      .A2(FINAL_RESULT_adder_tempIn11[6]), .B1(FINAL_RESULT_adder_n_1_29), 
      .B2(FINAL_RESULT_adder_i_1_n_9), .ZN(FINAL_RESULT_adder_n_1_25));
   OR2_X1 FINAL_RESULT_adder_i_1_46 (.A1(FINAL_RESULT_adder_tempIn22[6]), 
      .A2(FINAL_RESULT_adder_tempIn11[6]), .ZN(FINAL_RESULT_adder_i_1_n_9));
   OAI21_X1 FINAL_RESULT_adder_i_1_51 (.A(FINAL_RESULT_adder_i_1_n_11), .B1(
      FINAL_RESULT_adder_n_1_32), .B2(FINAL_RESULT_adder_i_1_n_10), .ZN(
      FINAL_RESULT_adder_n_1_29));
   NOR2_X1 FINAL_RESULT_adder_i_1_52 (.A1(FINAL_RESULT_adder_tempIn22[5]), 
      .A2(FINAL_RESULT_adder_tempIn11[5]), .ZN(FINAL_RESULT_adder_i_1_n_10));
   NAND2_X1 FINAL_RESULT_adder_i_1_53 (.A1(FINAL_RESULT_adder_tempIn22[5]), 
      .A2(FINAL_RESULT_adder_tempIn11[5]), .ZN(FINAL_RESULT_adder_i_1_n_11));
   OAI21_X1 FINAL_RESULT_adder_i_1_54 (.A(FINAL_RESULT_adder_i_1_n_12), .B1(
      FINAL_RESULT_adder_tempIn22[4]), .B2(FINAL_RESULT_adder_tempIn11[4]), 
      .ZN(FINAL_RESULT_adder_n_1_32));
   INV_X1 FINAL_RESULT_adder_i_1_55 (.A(FINAL_RESULT_adder_n_1_34), .ZN(
      FINAL_RESULT_adder_i_1_n_12));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[12]  (.D(VEC1_VEC2_adder_n_26), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[12]));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[11]  (.D(VEC1_VEC2_adder_n_25), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[11]));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[10]  (.D(VEC1_VEC2_adder_n_24), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[10]));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[9]  (.D(VEC1_VEC2_adder_n_23), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[9]));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[8]  (.D(VEC1_VEC2_adder_n_22), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[8]));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[7]  (.D(VEC1_VEC2_adder_n_21), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[7]));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[6]  (.D(VEC1_VEC2_adder_n_20), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[6]));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[5]  (.D(VEC1_VEC2_adder_n_19), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[5]));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[4]  (.D(VEC1_VEC2_adder_n_18), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[4]));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[3]  (.D(VEC1_VEC2_adder_n_17), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[3]));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[2]  (.D(VEC1_VEC2_adder_n_16), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[2]));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[1]  (.D(VEC1_VEC2_adder_n_15), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[1]));
   DLH_X1 \VEC1_VEC2_adder_tempIn22_reg[0]  (.D(VEC1_VEC2_adder_n_14), .G(
      VEC1_VEC2_adder_n_27), .Q(VEC1_VEC2_adder_tempIn22[0]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[12]  (.D(VEC1_VEC2_adder_n_12), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[12]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[11]  (.D(VEC1_VEC2_adder_n_11), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[11]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[10]  (.D(VEC1_VEC2_adder_n_10), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[10]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[9]  (.D(VEC1_VEC2_adder_n_9), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[9]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[8]  (.D(VEC1_VEC2_adder_n_8), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[8]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[7]  (.D(VEC1_VEC2_adder_n_7), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[7]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[6]  (.D(VEC1_VEC2_adder_n_6), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[6]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[5]  (.D(VEC1_VEC2_adder_n_5), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[5]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[4]  (.D(VEC1_VEC2_adder_n_4), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[4]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[3]  (.D(VEC1_VEC2_adder_n_3), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[3]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[2]  (.D(VEC1_VEC2_adder_n_2), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[2]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[1]  (.D(VEC1_VEC2_adder_n_1), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[1]));
   DLH_X1 \VEC1_VEC2_adder_tempIn11_reg[0]  (.D(VEC1_VEC2_adder_n_0), .G(
      VEC1_VEC2_adder_n_13), .Q(VEC1_VEC2_adder_tempIn11[0]));
   OAI22_X1 VEC1_VEC2_adder_i_0_0 (.A1(VEC1_VEC2_adder_n_0_89), .A2(
      VEC1_VEC2_adder_n_13), .B1(VEC1_VEC2_adder_n_0_93), .B2(
      VEC1_VEC2_adder_n_0_82), .ZN(Addition_Result[13]));
   OAI22_X1 VEC1_VEC2_adder_i_0_1 (.A1(VEC1_VEC2_adder_n_0_90), .A2(
      VEC1_VEC2_adder_n_13), .B1(VEC1_VEC2_adder_n_0_94), .B2(
      VEC1_VEC2_adder_n_0_82), .ZN(Addition_Result[14]));
   OR2_X1 VEC1_VEC2_adder_i_0_2 (.A1(RAM_DATA_RD2[15]), .A2(RAM_DATA_RD1[15]), 
      .ZN(Addition_Result[15]));
   AND2_X1 VEC1_VEC2_adder_i_0_3 (.A1(RAM_DATA_RD1[0]), .A2(
      VEC1_VEC2_adder_n_0_72), .ZN(VEC1_VEC2_adder_n_0));
   OAI22_X1 VEC1_VEC2_adder_i_0_4 (.A1(VEC1_VEC2_adder_n_0_3), .A2(
      VEC1_VEC2_adder_n_0_0), .B1(VEC1_VEC2_adder_n_0_75), .B2(
      VEC1_VEC2_adder_n_0_6), .ZN(VEC1_VEC2_adder_n_1));
   OAI22_X1 VEC1_VEC2_adder_i_0_5 (.A1(VEC1_VEC2_adder_n_0_75), .A2(
      VEC1_VEC2_adder_n_0_9), .B1(VEC1_VEC2_adder_n_0_6), .B2(
      VEC1_VEC2_adder_n_0_0), .ZN(VEC1_VEC2_adder_n_2));
   OAI22_X1 VEC1_VEC2_adder_i_0_6 (.A1(VEC1_VEC2_adder_n_0_75), .A2(
      VEC1_VEC2_adder_n_0_12), .B1(VEC1_VEC2_adder_n_0_9), .B2(
      VEC1_VEC2_adder_n_0_0), .ZN(VEC1_VEC2_adder_n_3));
   OAI22_X1 VEC1_VEC2_adder_i_0_7 (.A1(VEC1_VEC2_adder_n_0_78), .A2(
      VEC1_VEC2_adder_n_0_1), .B1(VEC1_VEC2_adder_n_0_12), .B2(
      VEC1_VEC2_adder_n_0_0), .ZN(VEC1_VEC2_adder_n_4));
   NAND2_X1 VEC1_VEC2_adder_i_0_8 (.A1(VEC1_VEC2_adder_n_0_78), .A2(
      VEC1_VEC2_adder_n_0_77), .ZN(VEC1_VEC2_adder_n_0_0));
   OAI22_X1 VEC1_VEC2_adder_i_0_9 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_1), .B1(VEC1_VEC2_adder_n_0_78), .B2(
      VEC1_VEC2_adder_n_0_4), .ZN(VEC1_VEC2_adder_n_5));
   INV_X1 VEC1_VEC2_adder_i_0_10 (.A(VEC1_VEC2_adder_n_0_2), .ZN(
      VEC1_VEC2_adder_n_0_1));
   OAI22_X1 VEC1_VEC2_adder_i_0_11 (.A1(VEC1_VEC2_adder_n_0_76), .A2(
      VEC1_VEC2_adder_n_0_15), .B1(VEC1_VEC2_adder_n_0_77), .B2(
      VEC1_VEC2_adder_n_0_3), .ZN(VEC1_VEC2_adder_n_0_2));
   NAND2_X1 VEC1_VEC2_adder_i_0_12 (.A1(RAM_DATA_RD1[0]), .A2(
      VEC1_VEC2_adder_n_0_32), .ZN(VEC1_VEC2_adder_n_0_3));
   OAI22_X1 VEC1_VEC2_adder_i_0_13 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_4), .B1(VEC1_VEC2_adder_n_0_78), .B2(
      VEC1_VEC2_adder_n_0_7), .ZN(VEC1_VEC2_adder_n_6));
   INV_X1 VEC1_VEC2_adder_i_0_14 (.A(VEC1_VEC2_adder_n_0_5), .ZN(
      VEC1_VEC2_adder_n_0_4));
   OAI22_X1 VEC1_VEC2_adder_i_0_15 (.A1(VEC1_VEC2_adder_n_0_76), .A2(
      VEC1_VEC2_adder_n_0_18), .B1(VEC1_VEC2_adder_n_0_77), .B2(
      VEC1_VEC2_adder_n_0_6), .ZN(VEC1_VEC2_adder_n_0_5));
   NAND2_X1 VEC1_VEC2_adder_i_0_16 (.A1(RAM_DATA_RD1[1]), .A2(
      VEC1_VEC2_adder_n_0_32), .ZN(VEC1_VEC2_adder_n_0_6));
   OAI22_X1 VEC1_VEC2_adder_i_0_17 (.A1(VEC1_VEC2_adder_n_0_78), .A2(
      VEC1_VEC2_adder_n_0_10), .B1(VEC1_VEC2_adder_n_0_79), .B2(
      VEC1_VEC2_adder_n_0_7), .ZN(VEC1_VEC2_adder_n_7));
   INV_X1 VEC1_VEC2_adder_i_0_18 (.A(VEC1_VEC2_adder_n_0_8), .ZN(
      VEC1_VEC2_adder_n_0_7));
   OAI22_X1 VEC1_VEC2_adder_i_0_19 (.A1(VEC1_VEC2_adder_n_0_77), .A2(
      VEC1_VEC2_adder_n_0_9), .B1(VEC1_VEC2_adder_n_0_76), .B2(
      VEC1_VEC2_adder_n_0_22), .ZN(VEC1_VEC2_adder_n_0_8));
   AOI22_X1 VEC1_VEC2_adder_i_0_20 (.A1(RAM_DATA_RD1[2]), .A2(
      VEC1_VEC2_adder_n_0_32), .B1(RAM_DATA_RD1[0]), .B2(VEC1_VEC2_adder_n_0_33), 
      .ZN(VEC1_VEC2_adder_n_0_9));
   OAI22_X1 VEC1_VEC2_adder_i_0_21 (.A1(VEC1_VEC2_adder_n_0_78), .A2(
      VEC1_VEC2_adder_n_0_13), .B1(VEC1_VEC2_adder_n_0_79), .B2(
      VEC1_VEC2_adder_n_0_10), .ZN(VEC1_VEC2_adder_n_8));
   INV_X1 VEC1_VEC2_adder_i_0_22 (.A(VEC1_VEC2_adder_n_0_11), .ZN(
      VEC1_VEC2_adder_n_0_10));
   OAI22_X1 VEC1_VEC2_adder_i_0_23 (.A1(VEC1_VEC2_adder_n_0_77), .A2(
      VEC1_VEC2_adder_n_0_12), .B1(VEC1_VEC2_adder_n_0_76), .B2(
      VEC1_VEC2_adder_n_0_26), .ZN(VEC1_VEC2_adder_n_0_11));
   AOI22_X1 VEC1_VEC2_adder_i_0_24 (.A1(RAM_DATA_RD1[3]), .A2(
      VEC1_VEC2_adder_n_0_32), .B1(RAM_DATA_RD1[1]), .B2(VEC1_VEC2_adder_n_0_33), 
      .ZN(VEC1_VEC2_adder_n_0_12));
   OAI22_X1 VEC1_VEC2_adder_i_0_25 (.A1(VEC1_VEC2_adder_n_0_78), .A2(
      VEC1_VEC2_adder_n_0_16), .B1(VEC1_VEC2_adder_n_0_79), .B2(
      VEC1_VEC2_adder_n_0_13), .ZN(VEC1_VEC2_adder_n_9));
   INV_X1 VEC1_VEC2_adder_i_0_26 (.A(VEC1_VEC2_adder_n_0_14), .ZN(
      VEC1_VEC2_adder_n_0_13));
   OAI22_X1 VEC1_VEC2_adder_i_0_27 (.A1(VEC1_VEC2_adder_n_0_77), .A2(
      VEC1_VEC2_adder_n_0_15), .B1(VEC1_VEC2_adder_n_0_76), .B2(
      VEC1_VEC2_adder_n_0_30), .ZN(VEC1_VEC2_adder_n_0_14));
   AOI22_X1 VEC1_VEC2_adder_i_0_28 (.A1(RAM_DATA_RD1[4]), .A2(
      VEC1_VEC2_adder_n_0_32), .B1(RAM_DATA_RD1[2]), .B2(VEC1_VEC2_adder_n_0_33), 
      .ZN(VEC1_VEC2_adder_n_0_15));
   OAI22_X1 VEC1_VEC2_adder_i_0_29 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_16), .B1(VEC1_VEC2_adder_n_0_78), .B2(
      VEC1_VEC2_adder_n_0_20), .ZN(VEC1_VEC2_adder_n_10));
   INV_X1 VEC1_VEC2_adder_i_0_30 (.A(VEC1_VEC2_adder_n_0_17), .ZN(
      VEC1_VEC2_adder_n_0_16));
   OAI22_X1 VEC1_VEC2_adder_i_0_31 (.A1(VEC1_VEC2_adder_n_0_76), .A2(
      VEC1_VEC2_adder_n_0_19), .B1(VEC1_VEC2_adder_n_0_77), .B2(
      VEC1_VEC2_adder_n_0_18), .ZN(VEC1_VEC2_adder_n_0_17));
   AOI22_X1 VEC1_VEC2_adder_i_0_32 (.A1(RAM_DATA_RD1[5]), .A2(
      VEC1_VEC2_adder_n_0_32), .B1(RAM_DATA_RD1[3]), .B2(VEC1_VEC2_adder_n_0_33), 
      .ZN(VEC1_VEC2_adder_n_0_18));
   AOI22_X1 VEC1_VEC2_adder_i_0_33 (.A1(RAM_DATA_RD1[9]), .A2(
      VEC1_VEC2_adder_n_0_32), .B1(RAM_DATA_RD1[7]), .B2(VEC1_VEC2_adder_n_0_33), 
      .ZN(VEC1_VEC2_adder_n_0_19));
   OAI22_X1 VEC1_VEC2_adder_i_0_34 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_20), .B1(VEC1_VEC2_adder_n_0_78), .B2(
      VEC1_VEC2_adder_n_0_24), .ZN(VEC1_VEC2_adder_n_11));
   INV_X1 VEC1_VEC2_adder_i_0_35 (.A(VEC1_VEC2_adder_n_0_21), .ZN(
      VEC1_VEC2_adder_n_0_20));
   OAI22_X1 VEC1_VEC2_adder_i_0_36 (.A1(VEC1_VEC2_adder_n_0_76), .A2(
      VEC1_VEC2_adder_n_0_23), .B1(VEC1_VEC2_adder_n_0_77), .B2(
      VEC1_VEC2_adder_n_0_22), .ZN(VEC1_VEC2_adder_n_0_21));
   AOI22_X1 VEC1_VEC2_adder_i_0_37 (.A1(RAM_DATA_RD1[6]), .A2(
      VEC1_VEC2_adder_n_0_32), .B1(RAM_DATA_RD1[4]), .B2(VEC1_VEC2_adder_n_0_33), 
      .ZN(VEC1_VEC2_adder_n_0_22));
   AOI22_X1 VEC1_VEC2_adder_i_0_38 (.A1(RAM_DATA_RD1[10]), .A2(
      VEC1_VEC2_adder_n_0_32), .B1(RAM_DATA_RD1[8]), .B2(VEC1_VEC2_adder_n_0_33), 
      .ZN(VEC1_VEC2_adder_n_0_23));
   OAI22_X1 VEC1_VEC2_adder_i_0_39 (.A1(VEC1_VEC2_adder_n_0_78), .A2(
      VEC1_VEC2_adder_n_0_28), .B1(VEC1_VEC2_adder_n_0_79), .B2(
      VEC1_VEC2_adder_n_0_24), .ZN(VEC1_VEC2_adder_n_12));
   INV_X1 VEC1_VEC2_adder_i_0_40 (.A(VEC1_VEC2_adder_n_0_25), .ZN(
      VEC1_VEC2_adder_n_0_24));
   OAI22_X1 VEC1_VEC2_adder_i_0_41 (.A1(VEC1_VEC2_adder_n_0_76), .A2(
      VEC1_VEC2_adder_n_0_27), .B1(VEC1_VEC2_adder_n_0_77), .B2(
      VEC1_VEC2_adder_n_0_26), .ZN(VEC1_VEC2_adder_n_0_25));
   AOI22_X1 VEC1_VEC2_adder_i_0_42 (.A1(RAM_DATA_RD1[7]), .A2(
      VEC1_VEC2_adder_n_0_32), .B1(RAM_DATA_RD1[5]), .B2(VEC1_VEC2_adder_n_0_33), 
      .ZN(VEC1_VEC2_adder_n_0_26));
   AOI22_X1 VEC1_VEC2_adder_i_0_43 (.A1(RAM_DATA_RD1[9]), .A2(
      VEC1_VEC2_adder_n_0_33), .B1(RAM_DATA_RD1[11]), .B2(VEC1_VEC2_adder_n_0_32), 
      .ZN(VEC1_VEC2_adder_n_0_27));
   INV_X1 VEC1_VEC2_adder_i_0_44 (.A(VEC1_VEC2_adder_n_0_29), .ZN(
      VEC1_VEC2_adder_n_0_28));
   OAI22_X1 VEC1_VEC2_adder_i_0_45 (.A1(VEC1_VEC2_adder_n_0_76), .A2(
      VEC1_VEC2_adder_n_0_31), .B1(VEC1_VEC2_adder_n_0_77), .B2(
      VEC1_VEC2_adder_n_0_30), .ZN(VEC1_VEC2_adder_n_0_29));
   AOI22_X1 VEC1_VEC2_adder_i_0_46 (.A1(RAM_DATA_RD1[8]), .A2(
      VEC1_VEC2_adder_n_0_32), .B1(RAM_DATA_RD1[6]), .B2(VEC1_VEC2_adder_n_0_33), 
      .ZN(VEC1_VEC2_adder_n_0_30));
   AOI22_X1 VEC1_VEC2_adder_i_0_47 (.A1(RAM_DATA_RD1[10]), .A2(
      VEC1_VEC2_adder_n_0_33), .B1(RAM_DATA_RD1[12]), .B2(VEC1_VEC2_adder_n_0_32), 
      .ZN(VEC1_VEC2_adder_n_0_31));
   INV_X1 VEC1_VEC2_adder_i_0_48 (.A(VEC1_VEC2_adder_n_0_33), .ZN(
      VEC1_VEC2_adder_n_0_32));
   XOR2_X1 VEC1_VEC2_adder_i_0_49 (.A(VEC1_VEC2_adder_n_0_86), .B(
      VEC1_VEC2_adder_n_0_73), .Z(VEC1_VEC2_adder_n_0_33));
   AND2_X1 VEC1_VEC2_adder_i_0_50 (.A1(RAM_DATA_RD2[0]), .A2(
      VEC1_VEC2_adder_n_0_72), .ZN(VEC1_VEC2_adder_n_14));
   OAI22_X1 VEC1_VEC2_adder_i_0_51 (.A1(VEC1_VEC2_adder_n_0_37), .A2(
      VEC1_VEC2_adder_n_0_34), .B1(VEC1_VEC2_adder_n_0_92), .B2(
      VEC1_VEC2_adder_n_0_71), .ZN(VEC1_VEC2_adder_n_15));
   OAI33_X1 VEC1_VEC2_adder_i_0_52 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_69), .A3(VEC1_VEC2_adder_n_0_40), .B1(
      VEC1_VEC2_adder_n_0_78), .B2(VEC1_VEC2_adder_n_0_69), .B3(
      VEC1_VEC2_adder_n_0_43), .ZN(VEC1_VEC2_adder_n_16));
   OAI33_X1 VEC1_VEC2_adder_i_0_53 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_69), .A3(VEC1_VEC2_adder_n_0_43), .B1(
      VEC1_VEC2_adder_n_0_78), .B2(VEC1_VEC2_adder_n_0_69), .B3(
      VEC1_VEC2_adder_n_0_46), .ZN(VEC1_VEC2_adder_n_17));
   OAI22_X1 VEC1_VEC2_adder_i_0_54 (.A1(VEC1_VEC2_adder_n_0_46), .A2(
      VEC1_VEC2_adder_n_0_34), .B1(VEC1_VEC2_adder_n_0_78), .B2(
      VEC1_VEC2_adder_n_0_35), .ZN(VEC1_VEC2_adder_n_18));
   NAND2_X1 VEC1_VEC2_adder_i_0_55 (.A1(VEC1_VEC2_adder_n_0_78), .A2(
      VEC1_VEC2_adder_n_0_68), .ZN(VEC1_VEC2_adder_n_0_34));
   AOI22_X1 VEC1_VEC2_adder_i_0_56 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_38), .B1(VEC1_VEC2_adder_n_0_78), .B2(
      VEC1_VEC2_adder_n_0_35), .ZN(VEC1_VEC2_adder_n_19));
   INV_X1 VEC1_VEC2_adder_i_0_57 (.A(VEC1_VEC2_adder_n_0_36), .ZN(
      VEC1_VEC2_adder_n_0_35));
   OAI22_X1 VEC1_VEC2_adder_i_0_58 (.A1(VEC1_VEC2_adder_n_0_69), .A2(
      VEC1_VEC2_adder_n_0_49), .B1(VEC1_VEC2_adder_n_0_68), .B2(
      VEC1_VEC2_adder_n_0_37), .ZN(VEC1_VEC2_adder_n_0_36));
   NAND2_X1 VEC1_VEC2_adder_i_0_59 (.A1(RAM_DATA_RD2[0]), .A2(
      VEC1_VEC2_adder_n_0_67), .ZN(VEC1_VEC2_adder_n_0_37));
   OAI22_X1 VEC1_VEC2_adder_i_0_60 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_38), .B1(VEC1_VEC2_adder_n_0_78), .B2(
      VEC1_VEC2_adder_n_0_41), .ZN(VEC1_VEC2_adder_n_20));
   INV_X1 VEC1_VEC2_adder_i_0_61 (.A(VEC1_VEC2_adder_n_0_39), .ZN(
      VEC1_VEC2_adder_n_0_38));
   OAI22_X1 VEC1_VEC2_adder_i_0_62 (.A1(VEC1_VEC2_adder_n_0_69), .A2(
      VEC1_VEC2_adder_n_0_52), .B1(VEC1_VEC2_adder_n_0_68), .B2(
      VEC1_VEC2_adder_n_0_40), .ZN(VEC1_VEC2_adder_n_0_39));
   NAND2_X1 VEC1_VEC2_adder_i_0_63 (.A1(RAM_DATA_RD2[1]), .A2(
      VEC1_VEC2_adder_n_0_67), .ZN(VEC1_VEC2_adder_n_0_40));
   OAI22_X1 VEC1_VEC2_adder_i_0_64 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_41), .B1(VEC1_VEC2_adder_n_0_78), .B2(
      VEC1_VEC2_adder_n_0_44), .ZN(VEC1_VEC2_adder_n_21));
   INV_X1 VEC1_VEC2_adder_i_0_65 (.A(VEC1_VEC2_adder_n_0_42), .ZN(
      VEC1_VEC2_adder_n_0_41));
   OAI22_X1 VEC1_VEC2_adder_i_0_66 (.A1(VEC1_VEC2_adder_n_0_69), .A2(
      VEC1_VEC2_adder_n_0_56), .B1(VEC1_VEC2_adder_n_0_68), .B2(
      VEC1_VEC2_adder_n_0_43), .ZN(VEC1_VEC2_adder_n_0_42));
   AOI22_X1 VEC1_VEC2_adder_i_0_67 (.A1(RAM_DATA_RD2[2]), .A2(
      VEC1_VEC2_adder_n_0_67), .B1(RAM_DATA_RD2[0]), .B2(VEC1_VEC2_adder_n_0_66), 
      .ZN(VEC1_VEC2_adder_n_0_43));
   OAI22_X1 VEC1_VEC2_adder_i_0_68 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_44), .B1(VEC1_VEC2_adder_n_0_78), .B2(
      VEC1_VEC2_adder_n_0_47), .ZN(VEC1_VEC2_adder_n_22));
   INV_X1 VEC1_VEC2_adder_i_0_69 (.A(VEC1_VEC2_adder_n_0_45), .ZN(
      VEC1_VEC2_adder_n_0_44));
   OAI22_X1 VEC1_VEC2_adder_i_0_70 (.A1(VEC1_VEC2_adder_n_0_69), .A2(
      VEC1_VEC2_adder_n_0_60), .B1(VEC1_VEC2_adder_n_0_68), .B2(
      VEC1_VEC2_adder_n_0_46), .ZN(VEC1_VEC2_adder_n_0_45));
   AOI22_X1 VEC1_VEC2_adder_i_0_71 (.A1(RAM_DATA_RD2[3]), .A2(
      VEC1_VEC2_adder_n_0_67), .B1(RAM_DATA_RD2[1]), .B2(VEC1_VEC2_adder_n_0_66), 
      .ZN(VEC1_VEC2_adder_n_0_46));
   OAI22_X1 VEC1_VEC2_adder_i_0_72 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_47), .B1(VEC1_VEC2_adder_n_0_78), .B2(
      VEC1_VEC2_adder_n_0_50), .ZN(VEC1_VEC2_adder_n_23));
   INV_X1 VEC1_VEC2_adder_i_0_73 (.A(VEC1_VEC2_adder_n_0_48), .ZN(
      VEC1_VEC2_adder_n_0_47));
   OAI22_X1 VEC1_VEC2_adder_i_0_74 (.A1(VEC1_VEC2_adder_n_0_69), .A2(
      VEC1_VEC2_adder_n_0_64), .B1(VEC1_VEC2_adder_n_0_68), .B2(
      VEC1_VEC2_adder_n_0_49), .ZN(VEC1_VEC2_adder_n_0_48));
   AOI22_X1 VEC1_VEC2_adder_i_0_75 (.A1(RAM_DATA_RD2[4]), .A2(
      VEC1_VEC2_adder_n_0_67), .B1(RAM_DATA_RD2[2]), .B2(VEC1_VEC2_adder_n_0_66), 
      .ZN(VEC1_VEC2_adder_n_0_49));
   OAI22_X1 VEC1_VEC2_adder_i_0_76 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_50), .B1(VEC1_VEC2_adder_n_0_78), .B2(
      VEC1_VEC2_adder_n_0_54), .ZN(VEC1_VEC2_adder_n_24));
   INV_X1 VEC1_VEC2_adder_i_0_77 (.A(VEC1_VEC2_adder_n_0_51), .ZN(
      VEC1_VEC2_adder_n_0_50));
   OAI22_X1 VEC1_VEC2_adder_i_0_78 (.A1(VEC1_VEC2_adder_n_0_69), .A2(
      VEC1_VEC2_adder_n_0_53), .B1(VEC1_VEC2_adder_n_0_68), .B2(
      VEC1_VEC2_adder_n_0_52), .ZN(VEC1_VEC2_adder_n_0_51));
   AOI22_X1 VEC1_VEC2_adder_i_0_79 (.A1(RAM_DATA_RD2[5]), .A2(
      VEC1_VEC2_adder_n_0_67), .B1(RAM_DATA_RD2[3]), .B2(VEC1_VEC2_adder_n_0_66), 
      .ZN(VEC1_VEC2_adder_n_0_52));
   AOI22_X1 VEC1_VEC2_adder_i_0_80 (.A1(RAM_DATA_RD2[9]), .A2(
      VEC1_VEC2_adder_n_0_67), .B1(RAM_DATA_RD2[7]), .B2(VEC1_VEC2_adder_n_0_66), 
      .ZN(VEC1_VEC2_adder_n_0_53));
   OAI22_X1 VEC1_VEC2_adder_i_0_81 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_54), .B1(VEC1_VEC2_adder_n_0_78), .B2(
      VEC1_VEC2_adder_n_0_58), .ZN(VEC1_VEC2_adder_n_25));
   INV_X1 VEC1_VEC2_adder_i_0_82 (.A(VEC1_VEC2_adder_n_0_55), .ZN(
      VEC1_VEC2_adder_n_0_54));
   OAI22_X1 VEC1_VEC2_adder_i_0_83 (.A1(VEC1_VEC2_adder_n_0_69), .A2(
      VEC1_VEC2_adder_n_0_57), .B1(VEC1_VEC2_adder_n_0_68), .B2(
      VEC1_VEC2_adder_n_0_56), .ZN(VEC1_VEC2_adder_n_0_55));
   AOI22_X1 VEC1_VEC2_adder_i_0_84 (.A1(RAM_DATA_RD2[6]), .A2(
      VEC1_VEC2_adder_n_0_67), .B1(RAM_DATA_RD2[4]), .B2(VEC1_VEC2_adder_n_0_66), 
      .ZN(VEC1_VEC2_adder_n_0_56));
   AOI22_X1 VEC1_VEC2_adder_i_0_85 (.A1(RAM_DATA_RD2[10]), .A2(
      VEC1_VEC2_adder_n_0_67), .B1(RAM_DATA_RD2[8]), .B2(VEC1_VEC2_adder_n_0_66), 
      .ZN(VEC1_VEC2_adder_n_0_57));
   OAI22_X1 VEC1_VEC2_adder_i_0_86 (.A1(VEC1_VEC2_adder_n_0_78), .A2(
      VEC1_VEC2_adder_n_0_62), .B1(VEC1_VEC2_adder_n_0_79), .B2(
      VEC1_VEC2_adder_n_0_58), .ZN(VEC1_VEC2_adder_n_26));
   INV_X1 VEC1_VEC2_adder_i_0_87 (.A(VEC1_VEC2_adder_n_0_59), .ZN(
      VEC1_VEC2_adder_n_0_58));
   OAI22_X1 VEC1_VEC2_adder_i_0_88 (.A1(VEC1_VEC2_adder_n_0_69), .A2(
      VEC1_VEC2_adder_n_0_61), .B1(VEC1_VEC2_adder_n_0_68), .B2(
      VEC1_VEC2_adder_n_0_60), .ZN(VEC1_VEC2_adder_n_0_59));
   AOI22_X1 VEC1_VEC2_adder_i_0_89 (.A1(RAM_DATA_RD2[7]), .A2(
      VEC1_VEC2_adder_n_0_67), .B1(RAM_DATA_RD2[5]), .B2(VEC1_VEC2_adder_n_0_66), 
      .ZN(VEC1_VEC2_adder_n_0_60));
   AOI22_X1 VEC1_VEC2_adder_i_0_90 (.A1(RAM_DATA_RD2[9]), .A2(
      VEC1_VEC2_adder_n_0_66), .B1(RAM_DATA_RD2[11]), .B2(VEC1_VEC2_adder_n_0_67), 
      .ZN(VEC1_VEC2_adder_n_0_61));
   INV_X1 VEC1_VEC2_adder_i_0_91 (.A(VEC1_VEC2_adder_n_0_63), .ZN(
      VEC1_VEC2_adder_n_0_62));
   OAI22_X1 VEC1_VEC2_adder_i_0_92 (.A1(VEC1_VEC2_adder_n_0_69), .A2(
      VEC1_VEC2_adder_n_0_65), .B1(VEC1_VEC2_adder_n_0_68), .B2(
      VEC1_VEC2_adder_n_0_64), .ZN(VEC1_VEC2_adder_n_0_63));
   AOI22_X1 VEC1_VEC2_adder_i_0_93 (.A1(RAM_DATA_RD2[8]), .A2(
      VEC1_VEC2_adder_n_0_67), .B1(RAM_DATA_RD2[6]), .B2(VEC1_VEC2_adder_n_0_66), 
      .ZN(VEC1_VEC2_adder_n_0_64));
   AOI22_X1 VEC1_VEC2_adder_i_0_94 (.A1(RAM_DATA_RD2[10]), .A2(
      VEC1_VEC2_adder_n_0_66), .B1(RAM_DATA_RD2[12]), .B2(VEC1_VEC2_adder_n_0_67), 
      .ZN(VEC1_VEC2_adder_n_0_65));
   INV_X1 VEC1_VEC2_adder_i_0_95 (.A(VEC1_VEC2_adder_n_0_67), .ZN(
      VEC1_VEC2_adder_n_0_66));
   OAI22_X1 VEC1_VEC2_adder_i_0_96 (.A1(VEC1_VEC2_adder_n_0_81), .A2(
      VEC1_VEC2_adder_n_0_73), .B1(VEC1_VEC2_adder_n_0_80), .B2(
      VEC1_VEC2_adder_n_0_74), .ZN(VEC1_VEC2_adder_n_0_67));
   INV_X1 VEC1_VEC2_adder_i_0_97 (.A(VEC1_VEC2_adder_n_0_69), .ZN(
      VEC1_VEC2_adder_n_0_68));
   XOR2_X1 VEC1_VEC2_adder_i_0_98 (.A(VEC1_VEC2_adder_n_0_83), .B(
      VEC1_VEC2_adder_n_0_70), .Z(VEC1_VEC2_adder_n_0_69));
   AOI21_X1 VEC1_VEC2_adder_i_0_99 (.A(VEC1_VEC2_adder_n_0_85), .B1(
      VEC1_VEC2_adder_n_0_87), .B2(VEC1_VEC2_adder_n_0_80), .ZN(
      VEC1_VEC2_adder_n_0_70));
   NAND2_X1 VEC1_VEC2_adder_i_0_100 (.A1(VEC1_VEC2_adder_n_13), .A2(
      VEC1_VEC2_adder_n_0_71), .ZN(VEC1_VEC2_adder_n_27));
   INV_X1 VEC1_VEC2_adder_i_0_101 (.A(VEC1_VEC2_adder_n_0_72), .ZN(
      VEC1_VEC2_adder_n_0_71));
   NOR2_X1 VEC1_VEC2_adder_i_0_102 (.A1(VEC1_VEC2_adder_n_0_75), .A2(
      VEC1_VEC2_adder_n_0_73), .ZN(VEC1_VEC2_adder_n_0_72));
   INV_X1 VEC1_VEC2_adder_i_0_103 (.A(VEC1_VEC2_adder_n_0_74), .ZN(
      VEC1_VEC2_adder_n_0_73));
   NOR2_X1 VEC1_VEC2_adder_i_0_104 (.A1(VEC1_VEC2_adder_n_0_88), .A2(
      VEC1_VEC2_adder_n_0_85), .ZN(VEC1_VEC2_adder_n_0_74));
   NAND2_X1 VEC1_VEC2_adder_i_0_105 (.A1(VEC1_VEC2_adder_n_0_79), .A2(
      VEC1_VEC2_adder_n_0_77), .ZN(VEC1_VEC2_adder_n_0_75));
   INV_X1 VEC1_VEC2_adder_i_0_106 (.A(VEC1_VEC2_adder_n_0_77), .ZN(
      VEC1_VEC2_adder_n_0_76));
   XOR2_X1 VEC1_VEC2_adder_i_0_107 (.A(VEC1_VEC2_adder_n_0_84), .B(
      VEC1_VEC2_adder_n_0_83), .Z(VEC1_VEC2_adder_n_0_77));
   INV_X1 VEC1_VEC2_adder_i_0_108 (.A(VEC1_VEC2_adder_n_0_79), .ZN(
      VEC1_VEC2_adder_n_0_78));
   NOR2_X1 VEC1_VEC2_adder_i_0_109 (.A1(VEC1_VEC2_adder_n_0_86), .A2(
      VEC1_VEC2_adder_n_0_81), .ZN(VEC1_VEC2_adder_n_0_79));
   INV_X1 VEC1_VEC2_adder_i_0_110 (.A(VEC1_VEC2_adder_n_0_81), .ZN(
      VEC1_VEC2_adder_n_0_80));
   NOR2_X1 VEC1_VEC2_adder_i_0_111 (.A1(VEC1_VEC2_adder_n_0_93), .A2(
      RAM_DATA_RD1[13]), .ZN(VEC1_VEC2_adder_n_0_81));
   INV_X1 VEC1_VEC2_adder_i_0_112 (.A(VEC1_VEC2_adder_n_0_82), .ZN(
      VEC1_VEC2_adder_n_13));
   OAI22_X1 VEC1_VEC2_adder_i_0_113 (.A1(RAM_DATA_RD2[15]), .A2(
      VEC1_VEC2_adder_n_0_91), .B1(VEC1_VEC2_adder_n_0_84), .B2(
      VEC1_VEC2_adder_n_0_83), .ZN(VEC1_VEC2_adder_n_0_82));
   XNOR2_X1 VEC1_VEC2_adder_i_0_114 (.A(RAM_DATA_RD2[15]), .B(
      VEC1_VEC2_adder_n_0_91), .ZN(VEC1_VEC2_adder_n_0_83));
   OAI21_X1 VEC1_VEC2_adder_i_0_115 (.A(VEC1_VEC2_adder_n_0_87), .B1(
      VEC1_VEC2_adder_n_0_86), .B2(VEC1_VEC2_adder_n_0_85), .ZN(
      VEC1_VEC2_adder_n_0_84));
   NOR2_X1 VEC1_VEC2_adder_i_0_116 (.A1(RAM_DATA_RD2[14]), .A2(
      VEC1_VEC2_adder_n_0_90), .ZN(VEC1_VEC2_adder_n_0_85));
   NOR2_X1 VEC1_VEC2_adder_i_0_117 (.A1(RAM_DATA_RD2[13]), .A2(
      VEC1_VEC2_adder_n_0_89), .ZN(VEC1_VEC2_adder_n_0_86));
   INV_X1 VEC1_VEC2_adder_i_0_118 (.A(VEC1_VEC2_adder_n_0_88), .ZN(
      VEC1_VEC2_adder_n_0_87));
   NOR2_X1 VEC1_VEC2_adder_i_0_119 (.A1(VEC1_VEC2_adder_n_0_94), .A2(
      RAM_DATA_RD1[14]), .ZN(VEC1_VEC2_adder_n_0_88));
   INV_X1 VEC1_VEC2_adder_i_0_120 (.A(RAM_DATA_RD1[13]), .ZN(
      VEC1_VEC2_adder_n_0_89));
   INV_X1 VEC1_VEC2_adder_i_0_121 (.A(RAM_DATA_RD1[14]), .ZN(
      VEC1_VEC2_adder_n_0_90));
   INV_X1 VEC1_VEC2_adder_i_0_122 (.A(RAM_DATA_RD1[15]), .ZN(
      VEC1_VEC2_adder_n_0_91));
   INV_X1 VEC1_VEC2_adder_i_0_123 (.A(RAM_DATA_RD2[1]), .ZN(
      VEC1_VEC2_adder_n_0_92));
   INV_X1 VEC1_VEC2_adder_i_0_124 (.A(RAM_DATA_RD2[13]), .ZN(
      VEC1_VEC2_adder_n_0_93));
   INV_X1 VEC1_VEC2_adder_i_0_125 (.A(RAM_DATA_RD2[14]), .ZN(
      VEC1_VEC2_adder_n_0_94));
   XOR2_X1 VEC1_VEC2_adder_i_1_0 (.A(VEC1_VEC2_adder_tempIn22[0]), .B(
      VEC1_VEC2_adder_tempIn11[0]), .Z(Addition_Result[0]));
   XNOR2_X1 VEC1_VEC2_adder_i_1_1 (.A(VEC1_VEC2_adder_n_1_43), .B(
      VEC1_VEC2_adder_n_1_0), .ZN(Addition_Result[1]));
   XOR2_X1 VEC1_VEC2_adder_i_1_2 (.A(VEC1_VEC2_adder_tempIn22[1]), .B(
      VEC1_VEC2_adder_tempIn11[1]), .Z(VEC1_VEC2_adder_n_1_0));
   XNOR2_X1 VEC1_VEC2_adder_i_1_3 (.A(VEC1_VEC2_adder_n_1_40), .B(
      VEC1_VEC2_adder_n_1_1), .ZN(Addition_Result[2]));
   XNOR2_X1 VEC1_VEC2_adder_i_1_4 (.A(VEC1_VEC2_adder_tempIn22[2]), .B(
      VEC1_VEC2_adder_tempIn11[2]), .ZN(VEC1_VEC2_adder_n_1_1));
   XNOR2_X1 VEC1_VEC2_adder_i_1_7 (.A(VEC1_VEC2_adder_n_1_35), .B(
      VEC1_VEC2_adder_n_1_3), .ZN(Addition_Result[4]));
   XNOR2_X1 VEC1_VEC2_adder_i_1_8 (.A(VEC1_VEC2_adder_tempIn22[4]), .B(
      VEC1_VEC2_adder_tempIn11[4]), .ZN(VEC1_VEC2_adder_n_1_3));
   XNOR2_X1 VEC1_VEC2_adder_i_1_9 (.A(VEC1_VEC2_adder_n_1_32), .B(
      VEC1_VEC2_adder_n_1_4), .ZN(Addition_Result[5]));
   XOR2_X1 VEC1_VEC2_adder_i_1_10 (.A(VEC1_VEC2_adder_tempIn22[5]), .B(
      VEC1_VEC2_adder_tempIn11[5]), .Z(VEC1_VEC2_adder_n_1_4));
   XNOR2_X1 VEC1_VEC2_adder_i_1_11 (.A(VEC1_VEC2_adder_n_1_29), .B(
      VEC1_VEC2_adder_n_1_5), .ZN(Addition_Result[6]));
   XNOR2_X1 VEC1_VEC2_adder_i_1_12 (.A(VEC1_VEC2_adder_tempIn22[6]), .B(
      VEC1_VEC2_adder_tempIn11[6]), .ZN(VEC1_VEC2_adder_n_1_5));
   XNOR2_X1 VEC1_VEC2_adder_i_1_13 (.A(VEC1_VEC2_adder_n_1_25), .B(
      VEC1_VEC2_adder_n_1_6), .ZN(Addition_Result[7]));
   XOR2_X1 VEC1_VEC2_adder_i_1_14 (.A(VEC1_VEC2_adder_tempIn22[7]), .B(
      VEC1_VEC2_adder_tempIn11[7]), .Z(VEC1_VEC2_adder_n_1_6));
   XNOR2_X1 VEC1_VEC2_adder_i_1_15 (.A(VEC1_VEC2_adder_n_1_23), .B(
      VEC1_VEC2_adder_n_1_7), .ZN(Addition_Result[8]));
   XNOR2_X1 VEC1_VEC2_adder_i_1_16 (.A(VEC1_VEC2_adder_tempIn22[8]), .B(
      VEC1_VEC2_adder_tempIn11[8]), .ZN(VEC1_VEC2_adder_n_1_7));
   XNOR2_X1 VEC1_VEC2_adder_i_1_19 (.A(VEC1_VEC2_adder_n_1_17), .B(
      VEC1_VEC2_adder_n_1_9), .ZN(Addition_Result[10]));
   XNOR2_X1 VEC1_VEC2_adder_i_1_20 (.A(VEC1_VEC2_adder_tempIn22[10]), .B(
      VEC1_VEC2_adder_tempIn11[10]), .ZN(VEC1_VEC2_adder_n_1_9));
   XNOR2_X1 VEC1_VEC2_adder_i_1_21 (.A(VEC1_VEC2_adder_n_1_14), .B(
      VEC1_VEC2_adder_n_1_10), .ZN(Addition_Result[11]));
   XOR2_X1 VEC1_VEC2_adder_i_1_22 (.A(VEC1_VEC2_adder_tempIn22[11]), .B(
      VEC1_VEC2_adder_tempIn11[11]), .Z(VEC1_VEC2_adder_n_1_10));
   XNOR2_X1 VEC1_VEC2_adder_i_1_23 (.A(VEC1_VEC2_adder_n_1_45), .B(
      VEC1_VEC2_adder_n_1_11), .ZN(Addition_Result[12]));
   OAI21_X1 VEC1_VEC2_adder_i_1_24 (.A(VEC1_VEC2_adder_n_1_12), .B1(
      VEC1_VEC2_adder_n_1_14), .B2(VEC1_VEC2_adder_n_1_13), .ZN(
      VEC1_VEC2_adder_n_1_11));
   NAND2_X1 VEC1_VEC2_adder_i_1_25 (.A1(VEC1_VEC2_adder_tempIn22[11]), .A2(
      VEC1_VEC2_adder_tempIn11[11]), .ZN(VEC1_VEC2_adder_n_1_12));
   NOR2_X1 VEC1_VEC2_adder_i_1_26 (.A1(VEC1_VEC2_adder_tempIn22[11]), .A2(
      VEC1_VEC2_adder_tempIn11[11]), .ZN(VEC1_VEC2_adder_n_1_13));
   OAI21_X1 VEC1_VEC2_adder_i_1_27 (.A(VEC1_VEC2_adder_n_1_15), .B1(
      VEC1_VEC2_adder_tempIn11[10]), .B2(VEC1_VEC2_adder_tempIn22[10]), .ZN(
      VEC1_VEC2_adder_n_1_14));
   INV_X1 VEC1_VEC2_adder_i_1_28 (.A(VEC1_VEC2_adder_n_1_16), .ZN(
      VEC1_VEC2_adder_n_1_15));
   AOI21_X1 VEC1_VEC2_adder_i_1_29 (.A(VEC1_VEC2_adder_n_1_17), .B1(
      VEC1_VEC2_adder_tempIn11[10]), .B2(VEC1_VEC2_adder_tempIn22[10]), .ZN(
      VEC1_VEC2_adder_n_1_16));
   AOI21_X1 VEC1_VEC2_adder_i_1_30 (.A(VEC1_VEC2_adder_n_1_18), .B1(
      VEC1_VEC2_adder_n_1_19), .B2(VEC1_VEC2_adder_n_1_20), .ZN(
      VEC1_VEC2_adder_n_1_17));
   NOR2_X1 VEC1_VEC2_adder_i_1_31 (.A1(VEC1_VEC2_adder_tempIn22[9]), .A2(
      VEC1_VEC2_adder_tempIn11[9]), .ZN(VEC1_VEC2_adder_n_1_18));
   NAND2_X1 VEC1_VEC2_adder_i_1_32 (.A1(VEC1_VEC2_adder_tempIn22[9]), .A2(
      VEC1_VEC2_adder_tempIn11[9]), .ZN(VEC1_VEC2_adder_n_1_19));
   AOI21_X1 VEC1_VEC2_adder_i_1_47 (.A(VEC1_VEC2_adder_n_1_35), .B1(
      VEC1_VEC2_adder_tempIn11[4]), .B2(VEC1_VEC2_adder_tempIn22[4]), .ZN(
      VEC1_VEC2_adder_n_1_34));
   AOI21_X1 VEC1_VEC2_adder_i_1_48 (.A(VEC1_VEC2_adder_n_1_36), .B1(
      VEC1_VEC2_adder_n_1_37), .B2(VEC1_VEC2_adder_n_1_38), .ZN(
      VEC1_VEC2_adder_n_1_35));
   NOR2_X1 VEC1_VEC2_adder_i_1_49 (.A1(VEC1_VEC2_adder_tempIn22[3]), .A2(
      VEC1_VEC2_adder_tempIn11[3]), .ZN(VEC1_VEC2_adder_n_1_36));
   NAND2_X1 VEC1_VEC2_adder_i_1_50 (.A1(VEC1_VEC2_adder_tempIn22[3]), .A2(
      VEC1_VEC2_adder_tempIn11[3]), .ZN(VEC1_VEC2_adder_n_1_37));
   XNOR2_X1 VEC1_VEC2_adder_i_1_58 (.A(VEC1_VEC2_adder_tempIn22[12]), .B(
      VEC1_VEC2_adder_tempIn11[12]), .ZN(VEC1_VEC2_adder_n_1_45));
   XOR2_X1 VEC1_VEC2_adder_i_1_5 (.A(VEC1_VEC2_adder_n_1_38), .B(
      VEC1_VEC2_adder_i_1_n_0), .Z(Addition_Result[3]));
   XNOR2_X1 VEC1_VEC2_adder_i_1_6 (.A(VEC1_VEC2_adder_tempIn22[3]), .B(
      VEC1_VEC2_adder_tempIn11[3]), .ZN(VEC1_VEC2_adder_i_1_n_0));
   OAI22_X1 VEC1_VEC2_adder_i_1_17 (.A1(VEC1_VEC2_adder_tempIn22[2]), .A2(
      VEC1_VEC2_adder_tempIn11[2]), .B1(VEC1_VEC2_adder_n_1_40), .B2(
      VEC1_VEC2_adder_i_1_n_1), .ZN(VEC1_VEC2_adder_n_1_38));
   AND2_X1 VEC1_VEC2_adder_i_1_18 (.A1(VEC1_VEC2_adder_tempIn22[2]), .A2(
      VEC1_VEC2_adder_tempIn11[2]), .ZN(VEC1_VEC2_adder_i_1_n_1));
   OAI22_X1 VEC1_VEC2_adder_i_1_33 (.A1(VEC1_VEC2_adder_i_1_n_4), .A2(
      VEC1_VEC2_adder_i_1_n_3), .B1(VEC1_VEC2_adder_n_1_43), .B2(
      VEC1_VEC2_adder_i_1_n_2), .ZN(VEC1_VEC2_adder_n_1_40));
   NOR2_X1 VEC1_VEC2_adder_i_1_34 (.A1(VEC1_VEC2_adder_tempIn22[1]), .A2(
      VEC1_VEC2_adder_tempIn11[1]), .ZN(VEC1_VEC2_adder_i_1_n_2));
   NAND2_X1 VEC1_VEC2_adder_i_1_35 (.A1(VEC1_VEC2_adder_tempIn22[0]), .A2(
      VEC1_VEC2_adder_tempIn11[0]), .ZN(VEC1_VEC2_adder_n_1_43));
   INV_X1 VEC1_VEC2_adder_i_1_36 (.A(VEC1_VEC2_adder_tempIn11[1]), .ZN(
      VEC1_VEC2_adder_i_1_n_3));
   INV_X1 VEC1_VEC2_adder_i_1_37 (.A(VEC1_VEC2_adder_tempIn22[1]), .ZN(
      VEC1_VEC2_adder_i_1_n_4));
   XOR2_X1 VEC1_VEC2_adder_i_1_38 (.A(VEC1_VEC2_adder_n_1_20), .B(
      VEC1_VEC2_adder_i_1_n_5), .Z(Addition_Result[9]));
   XNOR2_X1 VEC1_VEC2_adder_i_1_39 (.A(VEC1_VEC2_adder_tempIn22[9]), .B(
      VEC1_VEC2_adder_tempIn11[9]), .ZN(VEC1_VEC2_adder_i_1_n_5));
   AOI22_X1 VEC1_VEC2_adder_i_1_40 (.A1(VEC1_VEC2_adder_tempIn22[8]), .A2(
      VEC1_VEC2_adder_tempIn11[8]), .B1(VEC1_VEC2_adder_n_1_23), .B2(
      VEC1_VEC2_adder_i_1_n_6), .ZN(VEC1_VEC2_adder_n_1_20));
   OR2_X1 VEC1_VEC2_adder_i_1_41 (.A1(VEC1_VEC2_adder_tempIn22[8]), .A2(
      VEC1_VEC2_adder_tempIn11[8]), .ZN(VEC1_VEC2_adder_i_1_n_6));
   OAI21_X1 VEC1_VEC2_adder_i_1_42 (.A(VEC1_VEC2_adder_i_1_n_8), .B1(
      VEC1_VEC2_adder_n_1_25), .B2(VEC1_VEC2_adder_i_1_n_7), .ZN(
      VEC1_VEC2_adder_n_1_23));
   NOR2_X1 VEC1_VEC2_adder_i_1_43 (.A1(VEC1_VEC2_adder_tempIn22[7]), .A2(
      VEC1_VEC2_adder_tempIn11[7]), .ZN(VEC1_VEC2_adder_i_1_n_7));
   NAND2_X1 VEC1_VEC2_adder_i_1_44 (.A1(VEC1_VEC2_adder_tempIn22[7]), .A2(
      VEC1_VEC2_adder_tempIn11[7]), .ZN(VEC1_VEC2_adder_i_1_n_8));
   AOI22_X1 VEC1_VEC2_adder_i_1_45 (.A1(VEC1_VEC2_adder_tempIn22[6]), .A2(
      VEC1_VEC2_adder_tempIn11[6]), .B1(VEC1_VEC2_adder_n_1_29), .B2(
      VEC1_VEC2_adder_i_1_n_9), .ZN(VEC1_VEC2_adder_n_1_25));
   OR2_X1 VEC1_VEC2_adder_i_1_46 (.A1(VEC1_VEC2_adder_tempIn22[6]), .A2(
      VEC1_VEC2_adder_tempIn11[6]), .ZN(VEC1_VEC2_adder_i_1_n_9));
   OAI21_X1 VEC1_VEC2_adder_i_1_51 (.A(VEC1_VEC2_adder_i_1_n_11), .B1(
      VEC1_VEC2_adder_n_1_32), .B2(VEC1_VEC2_adder_i_1_n_10), .ZN(
      VEC1_VEC2_adder_n_1_29));
   NOR2_X1 VEC1_VEC2_adder_i_1_52 (.A1(VEC1_VEC2_adder_tempIn22[5]), .A2(
      VEC1_VEC2_adder_tempIn11[5]), .ZN(VEC1_VEC2_adder_i_1_n_10));
   NAND2_X1 VEC1_VEC2_adder_i_1_53 (.A1(VEC1_VEC2_adder_tempIn22[5]), .A2(
      VEC1_VEC2_adder_tempIn11[5]), .ZN(VEC1_VEC2_adder_i_1_n_11));
   OAI21_X1 VEC1_VEC2_adder_i_1_54 (.A(VEC1_VEC2_adder_i_1_n_12), .B1(
      VEC1_VEC2_adder_tempIn22[4]), .B2(VEC1_VEC2_adder_tempIn11[4]), .ZN(
      VEC1_VEC2_adder_n_1_32));
   INV_X1 VEC1_VEC2_adder_i_1_55 (.A(VEC1_VEC2_adder_n_1_34), .ZN(
      VEC1_VEC2_adder_i_1_n_12));
   DLH_X1 RAM_ENABLE_WR_reg (.D(n_0_198), .G(n_0_199), .Q(RAM_ENABLE_WR));
   DLH_X1 \RAM_DATA_WR_reg[15]  (.D(n_0_197), .G(n_0_47), .Q(RAM_DATA_WR[15]));
   DLH_X1 \RAM_DATA_WR_reg[14]  (.D(n_0_196), .G(n_0_47), .Q(RAM_DATA_WR[14]));
   DLH_X1 \RAM_DATA_WR_reg[13]  (.D(n_0_195), .G(n_0_47), .Q(RAM_DATA_WR[13]));
   DLH_X1 \RAM_DATA_WR_reg[12]  (.D(n_0_194), .G(n_0_47), .Q(RAM_DATA_WR[12]));
   DLH_X1 \RAM_DATA_WR_reg[11]  (.D(n_0_193), .G(n_0_47), .Q(RAM_DATA_WR[11]));
   DLH_X1 \RAM_DATA_WR_reg[10]  (.D(n_0_192), .G(n_0_47), .Q(RAM_DATA_WR[10]));
   DLH_X1 \RAM_DATA_WR_reg[9]  (.D(n_0_191), .G(n_0_47), .Q(RAM_DATA_WR[9]));
   DLH_X1 \RAM_DATA_WR_reg[8]  (.D(n_0_190), .G(n_0_47), .Q(RAM_DATA_WR[8]));
   DLH_X1 \RAM_DATA_WR_reg[7]  (.D(n_0_189), .G(n_0_47), .Q(RAM_DATA_WR[7]));
   DLH_X1 \RAM_DATA_WR_reg[6]  (.D(n_0_188), .G(n_0_47), .Q(RAM_DATA_WR[6]));
   DLH_X1 \RAM_DATA_WR_reg[5]  (.D(n_0_187), .G(n_0_47), .Q(RAM_DATA_WR[5]));
   DLH_X1 \RAM_DATA_WR_reg[4]  (.D(n_0_186), .G(n_0_47), .Q(RAM_DATA_WR[4]));
   DLH_X1 \RAM_DATA_WR_reg[3]  (.D(n_0_185), .G(n_0_47), .Q(RAM_DATA_WR[3]));
   DLH_X1 \RAM_DATA_WR_reg[2]  (.D(n_0_184), .G(n_0_47), .Q(RAM_DATA_WR[2]));
   DLH_X1 \RAM_DATA_WR_reg[1]  (.D(n_0_183), .G(n_0_47), .Q(RAM_DATA_WR[1]));
   DLH_X1 \RAM_DATA_WR_reg[0]  (.D(n_0_182), .G(n_0_47), .Q(RAM_DATA_WR[0]));
   DLH_X1 \h_val_reg[15]  (.D(RAM_DATA_RD1[15]), .G(n_0_181), .Q(n_0));
   DLH_X1 \h_val_reg[14]  (.D(RAM_DATA_RD1[14]), .G(n_0_181), .Q(n_1));
   DLH_X1 \h_val_reg[13]  (.D(RAM_DATA_RD1[13]), .G(n_0_181), .Q(n_2));
   DLH_X1 \h_val_reg[12]  (.D(RAM_DATA_RD1[12]), .G(n_0_181), .Q(n_3));
   DLH_X1 \h_val_reg[11]  (.D(RAM_DATA_RD1[11]), .G(n_0_181), .Q(n_4));
   DLH_X1 \h_val_reg[10]  (.D(RAM_DATA_RD1[10]), .G(n_0_181), .Q(n_5));
   DLH_X1 \h_val_reg[9]  (.D(RAM_DATA_RD1[9]), .G(n_0_181), .Q(n_6));
   DLH_X1 \h_val_reg[8]  (.D(RAM_DATA_RD1[8]), .G(n_0_181), .Q(n_7));
   DLH_X1 \h_val_reg[7]  (.D(RAM_DATA_RD1[7]), .G(n_0_181), .Q(n_8));
   DLH_X1 \h_val_reg[6]  (.D(RAM_DATA_RD1[6]), .G(n_0_181), .Q(n_9));
   DLH_X1 \h_val_reg[5]  (.D(RAM_DATA_RD1[5]), .G(n_0_181), .Q(n_10));
   DLH_X1 \h_val_reg[4]  (.D(RAM_DATA_RD1[4]), .G(n_0_181), .Q(n_11));
   DLH_X1 \h_val_reg[3]  (.D(RAM_DATA_RD1[3]), .G(n_0_181), .Q(n_12));
   DLH_X1 \h_val_reg[2]  (.D(RAM_DATA_RD1[2]), .G(n_0_181), .Q(n_13));
   DLH_X1 \h_val_reg[1]  (.D(RAM_DATA_RD1[1]), .G(n_0_181), .Q(n_14));
   DLH_X1 \h_val_reg[0]  (.D(RAM_DATA_RD1[0]), .G(n_0_181), .Q(n_15));
   DLH_X1 \Element_Result_reg[15]  (.D(n_0_179), .G(n_0_180), .Q(
      Element_Result[15]));
   DLH_X1 \Element_Result_reg[14]  (.D(n_0_178), .G(n_0_180), .Q(
      Element_Result[14]));
   DLH_X1 \Element_Result_reg[13]  (.D(n_0_177), .G(n_0_180), .Q(
      Element_Result[13]));
   DLH_X1 \Element_Result_reg[12]  (.D(n_0_176), .G(n_0_180), .Q(
      Element_Result[12]));
   DLH_X1 \Element_Result_reg[11]  (.D(n_0_175), .G(n_0_180), .Q(
      Element_Result[11]));
   DLH_X1 \Element_Result_reg[10]  (.D(n_0_174), .G(n_0_180), .Q(
      Element_Result[10]));
   DLH_X1 \Element_Result_reg[9]  (.D(n_0_173), .G(n_0_180), .Q(
      Element_Result[9]));
   DLH_X1 \Element_Result_reg[8]  (.D(n_0_172), .G(n_0_180), .Q(
      Element_Result[8]));
   DLH_X1 \Element_Result_reg[7]  (.D(n_0_171), .G(n_0_180), .Q(
      Element_Result[7]));
   DLH_X1 \Element_Result_reg[6]  (.D(n_0_170), .G(n_0_180), .Q(
      Element_Result[6]));
   DLH_X1 \Element_Result_reg[5]  (.D(n_0_169), .G(n_0_180), .Q(
      Element_Result[5]));
   DLH_X1 \Element_Result_reg[4]  (.D(n_0_168), .G(n_0_180), .Q(
      Element_Result[4]));
   DLH_X1 \Element_Result_reg[3]  (.D(n_0_167), .G(n_0_180), .Q(
      Element_Result[3]));
   DLH_X1 \Element_Result_reg[2]  (.D(n_0_166), .G(n_0_180), .Q(
      Element_Result[2]));
   DLH_X1 \Element_Result_reg[1]  (.D(n_0_165), .G(n_0_180), .Q(
      Element_Result[1]));
   DLH_X1 \Element_Result_reg[0]  (.D(n_0_164), .G(n_0_180), .Q(
      Element_Result[0]));
   DLH_X1 \RAM_ADD_WR_reg[12]  (.D(n_0_146), .G(n_0_133), .Q(RAM_ADD_WR[12]));
   DLH_X1 \RAM_ADD_WR_reg[11]  (.D(n_0_145), .G(n_0_133), .Q(RAM_ADD_WR[11]));
   DLH_X1 \RAM_ADD_WR_reg[10]  (.D(n_0_144), .G(n_0_133), .Q(RAM_ADD_WR[10]));
   DLH_X1 \RAM_ADD_WR_reg[9]  (.D(n_0_143), .G(n_0_133), .Q(RAM_ADD_WR[9]));
   DLH_X1 \RAM_ADD_WR_reg[8]  (.D(n_0_142), .G(n_0_133), .Q(RAM_ADD_WR[8]));
   DLH_X1 \RAM_ADD_WR_reg[7]  (.D(n_0_141), .G(n_0_133), .Q(RAM_ADD_WR[7]));
   DLH_X1 \RAM_ADD_WR_reg[6]  (.D(n_0_140), .G(n_0_133), .Q(RAM_ADD_WR[6]));
   DLH_X1 \RAM_ADD_WR_reg[5]  (.D(n_0_139), .G(n_0_133), .Q(RAM_ADD_WR[5]));
   DLH_X1 \RAM_ADD_WR_reg[4]  (.D(n_0_138), .G(n_0_133), .Q(RAM_ADD_WR[4]));
   DLH_X1 \RAM_ADD_WR_reg[3]  (.D(n_0_137), .G(n_0_133), .Q(RAM_ADD_WR[3]));
   DLH_X1 \RAM_ADD_WR_reg[2]  (.D(n_0_136), .G(n_0_133), .Q(RAM_ADD_WR[2]));
   DLH_X1 \RAM_ADD_WR_reg[1]  (.D(n_0_135), .G(n_0_133), .Q(RAM_ADD_WR[1]));
   DLH_X1 \RAM_ADD_WR_reg[0]  (.D(n_0_134), .G(n_0_133), .Q(RAM_ADD_WR[0]));
   DLH_X1 \RESULT_ADD_reg[15]  (.D(n_0_162), .G(n_0_163), .Q(RESULT_ADD[15]));
   DLH_X1 \RESULT_ADD_reg[14]  (.D(n_0_161), .G(n_0_163), .Q(RESULT_ADD[14]));
   DLH_X1 \RESULT_ADD_reg[13]  (.D(n_0_160), .G(n_0_163), .Q(RESULT_ADD[13]));
   DLH_X1 \RESULT_ADD_reg[12]  (.D(n_0_159), .G(n_0_163), .Q(RESULT_ADD[12]));
   DLH_X1 \RESULT_ADD_reg[11]  (.D(n_0_158), .G(n_0_163), .Q(RESULT_ADD[11]));
   DLH_X1 \RESULT_ADD_reg[10]  (.D(n_0_157), .G(n_0_163), .Q(RESULT_ADD[10]));
   DLH_X1 \RESULT_ADD_reg[9]  (.D(n_0_156), .G(n_0_163), .Q(RESULT_ADD[9]));
   DLH_X1 \RESULT_ADD_reg[8]  (.D(n_0_155), .G(n_0_163), .Q(RESULT_ADD[8]));
   DLH_X1 \RESULT_ADD_reg[7]  (.D(n_0_154), .G(n_0_163), .Q(RESULT_ADD[7]));
   DLH_X1 \RESULT_ADD_reg[6]  (.D(n_0_153), .G(n_0_163), .Q(RESULT_ADD[6]));
   DLH_X1 \RESULT_ADD_reg[5]  (.D(n_0_152), .G(n_0_163), .Q(RESULT_ADD[5]));
   DLH_X1 \RESULT_ADD_reg[4]  (.D(n_0_151), .G(n_0_163), .Q(RESULT_ADD[4]));
   DLH_X1 \RESULT_ADD_reg[3]  (.D(n_0_150), .G(n_0_163), .Q(RESULT_ADD[3]));
   DLH_X1 \RESULT_ADD_reg[2]  (.D(n_0_149), .G(n_0_163), .Q(RESULT_ADD[2]));
   DLH_X1 \RESULT_ADD_reg[1]  (.D(n_0_148), .G(n_0_163), .Q(RESULT_ADD[1]));
   DLH_X1 \RESULT_ADD_reg[0]  (.D(n_0_147), .G(n_0_163), .Q(RESULT_ADD[0]));
   DLH_X1 \RAM_ADD_RD2_reg[12]  (.D(n_0_131), .G(n_0_132), .Q(RAM_ADD_RD2[12]));
   DLH_X1 \RAM_ADD_RD2_reg[11]  (.D(n_0_130), .G(n_0_132), .Q(RAM_ADD_RD2[11]));
   DLH_X1 \RAM_ADD_RD2_reg[10]  (.D(n_0_129), .G(n_0_132), .Q(RAM_ADD_RD2[10]));
   DLH_X1 \RAM_ADD_RD2_reg[9]  (.D(n_0_128), .G(n_0_132), .Q(RAM_ADD_RD2[9]));
   DLH_X1 \RAM_ADD_RD2_reg[8]  (.D(n_0_127), .G(n_0_132), .Q(RAM_ADD_RD2[8]));
   DLH_X1 \RAM_ADD_RD2_reg[7]  (.D(n_0_126), .G(n_0_132), .Q(RAM_ADD_RD2[7]));
   DLH_X1 \RAM_ADD_RD2_reg[6]  (.D(n_0_125), .G(n_0_132), .Q(RAM_ADD_RD2[6]));
   DLH_X1 \RAM_ADD_RD2_reg[5]  (.D(n_0_124), .G(n_0_132), .Q(RAM_ADD_RD2[5]));
   DLH_X1 \RAM_ADD_RD2_reg[4]  (.D(n_0_123), .G(n_0_132), .Q(RAM_ADD_RD2[4]));
   DLH_X1 \RAM_ADD_RD2_reg[3]  (.D(n_0_122), .G(n_0_132), .Q(RAM_ADD_RD2[3]));
   DLH_X1 \RAM_ADD_RD2_reg[2]  (.D(n_0_121), .G(n_0_132), .Q(RAM_ADD_RD2[2]));
   DLH_X1 \RAM_ADD_RD2_reg[1]  (.D(n_0_120), .G(n_0_132), .Q(RAM_ADD_RD2[1]));
   DLH_X1 \RAM_ADD_RD2_reg[0]  (.D(n_0_119), .G(n_0_132), .Q(RAM_ADD_RD2[0]));
   DLH_X1 \RAM_ADD_RD1_reg[12]  (.D(n_0_67), .G(n_0_118), .Q(RAM_ADD_RD1[12]));
   DLH_X1 \RAM_ADD_RD1_reg[11]  (.D(n_0_66), .G(n_0_118), .Q(RAM_ADD_RD1[11]));
   DLH_X1 \RAM_ADD_RD1_reg[10]  (.D(n_0_65), .G(n_0_118), .Q(RAM_ADD_RD1[10]));
   DLH_X1 \RAM_ADD_RD1_reg[9]  (.D(n_0_64), .G(n_0_118), .Q(RAM_ADD_RD1[9]));
   DLH_X1 \RAM_ADD_RD1_reg[8]  (.D(n_0_63), .G(n_0_118), .Q(RAM_ADD_RD1[8]));
   DLH_X1 \RAM_ADD_RD1_reg[7]  (.D(n_0_62), .G(n_0_118), .Q(RAM_ADD_RD1[7]));
   DLH_X1 \RAM_ADD_RD1_reg[6]  (.D(n_0_61), .G(n_0_118), .Q(RAM_ADD_RD1[6]));
   DLH_X1 \RAM_ADD_RD1_reg[5]  (.D(n_0_60), .G(n_0_118), .Q(RAM_ADD_RD1[5]));
   DLH_X1 \RAM_ADD_RD1_reg[4]  (.D(n_0_59), .G(n_0_118), .Q(RAM_ADD_RD1[4]));
   DLH_X1 \RAM_ADD_RD1_reg[3]  (.D(n_0_58), .G(n_0_118), .Q(RAM_ADD_RD1[3]));
   DLH_X1 \RAM_ADD_RD1_reg[2]  (.D(n_0_57), .G(n_0_118), .Q(RAM_ADD_RD1[2]));
   DLH_X1 \RAM_ADD_RD1_reg[1]  (.D(n_0_56), .G(n_0_118), .Q(RAM_ADD_RD1[1]));
   DLH_X1 \RAM_ADD_RD1_reg[0]  (.D(n_0_55), .G(n_0_118), .Q(RAM_ADD_RD1[0]));
   DLH_X1 \VECTOR_ADD_reg[15]  (.D(n_0_116), .G(n_0_117), .Q(VECTOR_ADD[15]));
   DLH_X1 \VECTOR_ADD_reg[14]  (.D(n_0_115), .G(n_0_117), .Q(VECTOR_ADD[14]));
   DLH_X1 \VECTOR_ADD_reg[13]  (.D(n_0_114), .G(n_0_117), .Q(VECTOR_ADD[13]));
   DLH_X1 \VECTOR_ADD_reg[12]  (.D(n_0_113), .G(n_0_117), .Q(VECTOR_ADD[12]));
   DLH_X1 \VECTOR_ADD_reg[11]  (.D(n_0_112), .G(n_0_117), .Q(VECTOR_ADD[11]));
   DLH_X1 \VECTOR_ADD_reg[10]  (.D(n_0_111), .G(n_0_117), .Q(VECTOR_ADD[10]));
   DLH_X1 \VECTOR_ADD_reg[9]  (.D(n_0_110), .G(n_0_117), .Q(VECTOR_ADD[9]));
   DLH_X1 \VECTOR_ADD_reg[8]  (.D(n_0_109), .G(n_0_117), .Q(VECTOR_ADD[8]));
   DLH_X1 \VECTOR_ADD_reg[7]  (.D(n_0_108), .G(n_0_117), .Q(VECTOR_ADD[7]));
   DLH_X1 \VECTOR_ADD_reg[6]  (.D(n_0_107), .G(n_0_117), .Q(VECTOR_ADD[6]));
   DLH_X1 \VECTOR_ADD_reg[5]  (.D(n_0_106), .G(n_0_117), .Q(VECTOR_ADD[5]));
   DLH_X1 \VECTOR_ADD_reg[4]  (.D(n_0_105), .G(n_0_117), .Q(VECTOR_ADD[4]));
   DLH_X1 \VECTOR_ADD_reg[3]  (.D(n_0_104), .G(n_0_117), .Q(VECTOR_ADD[3]));
   DLH_X1 \VECTOR_ADD_reg[2]  (.D(n_0_103), .G(n_0_117), .Q(VECTOR_ADD[2]));
   DLH_X1 \VECTOR_ADD_reg[1]  (.D(n_0_102), .G(n_0_117), .Q(VECTOR_ADD[1]));
   DLH_X1 \VECTOR_ADD_reg[0]  (.D(n_0_101), .G(n_0_117), .Q(VECTOR_ADD[0]));
   DLH_X1 \VECTOR2_ADD_reg[15]  (.D(n_0_99), .G(n_0_100), .Q(VECTOR2_ADD[15]));
   DLH_X1 \VECTOR2_ADD_reg[14]  (.D(n_0_98), .G(n_0_100), .Q(VECTOR2_ADD[14]));
   DLH_X1 \VECTOR2_ADD_reg[13]  (.D(n_0_97), .G(n_0_100), .Q(VECTOR2_ADD[13]));
   DLH_X1 \VECTOR2_ADD_reg[12]  (.D(n_0_96), .G(n_0_100), .Q(VECTOR2_ADD[12]));
   DLH_X1 \VECTOR2_ADD_reg[11]  (.D(n_0_95), .G(n_0_100), .Q(VECTOR2_ADD[11]));
   DLH_X1 \VECTOR2_ADD_reg[10]  (.D(n_0_94), .G(n_0_100), .Q(VECTOR2_ADD[10]));
   DLH_X1 \VECTOR2_ADD_reg[9]  (.D(n_0_93), .G(n_0_100), .Q(VECTOR2_ADD[9]));
   DLH_X1 \VECTOR2_ADD_reg[8]  (.D(n_0_92), .G(n_0_100), .Q(VECTOR2_ADD[8]));
   DLH_X1 \VECTOR2_ADD_reg[7]  (.D(n_0_91), .G(n_0_100), .Q(VECTOR2_ADD[7]));
   DLH_X1 \VECTOR2_ADD_reg[6]  (.D(n_0_90), .G(n_0_100), .Q(VECTOR2_ADD[6]));
   DLH_X1 \VECTOR2_ADD_reg[5]  (.D(n_0_89), .G(n_0_100), .Q(VECTOR2_ADD[5]));
   DLH_X1 \VECTOR2_ADD_reg[4]  (.D(n_0_88), .G(n_0_100), .Q(VECTOR2_ADD[4]));
   DLH_X1 \VECTOR2_ADD_reg[3]  (.D(n_0_87), .G(n_0_100), .Q(VECTOR2_ADD[3]));
   DLH_X1 \VECTOR2_ADD_reg[2]  (.D(n_0_86), .G(n_0_100), .Q(VECTOR2_ADD[2]));
   DLH_X1 \VECTOR2_ADD_reg[1]  (.D(n_0_85), .G(n_0_100), .Q(VECTOR2_ADD[1]));
   DLH_X1 \VECTOR2_ADD_reg[0]  (.D(n_0_84), .G(n_0_100), .Q(VECTOR2_ADD[0]));
   DLH_X1 \MATRIX_ADD_reg[15]  (.D(n_0_83), .G(n_0_46), .Q(MATRIX_ADD[15]));
   DLH_X1 \MATRIX_ADD_reg[14]  (.D(n_0_82), .G(n_0_46), .Q(MATRIX_ADD[14]));
   DLH_X1 \MATRIX_ADD_reg[13]  (.D(n_0_81), .G(n_0_46), .Q(MATRIX_ADD[13]));
   DLH_X1 \MATRIX_ADD_reg[12]  (.D(n_0_80), .G(n_0_46), .Q(MATRIX_ADD[12]));
   DLH_X1 \MATRIX_ADD_reg[11]  (.D(n_0_79), .G(n_0_46), .Q(MATRIX_ADD[11]));
   DLH_X1 \MATRIX_ADD_reg[10]  (.D(n_0_78), .G(n_0_46), .Q(MATRIX_ADD[10]));
   DLH_X1 \MATRIX_ADD_reg[9]  (.D(n_0_77), .G(n_0_46), .Q(MATRIX_ADD[9]));
   DLH_X1 \MATRIX_ADD_reg[8]  (.D(n_0_76), .G(n_0_46), .Q(MATRIX_ADD[8]));
   DLH_X1 \MATRIX_ADD_reg[7]  (.D(n_0_75), .G(n_0_46), .Q(MATRIX_ADD[7]));
   DLH_X1 \MATRIX_ADD_reg[6]  (.D(n_0_74), .G(n_0_46), .Q(MATRIX_ADD[6]));
   DLH_X1 \MATRIX_ADD_reg[5]  (.D(n_0_73), .G(n_0_46), .Q(MATRIX_ADD[5]));
   DLH_X1 \MATRIX_ADD_reg[4]  (.D(n_0_72), .G(n_0_46), .Q(MATRIX_ADD[4]));
   DLH_X1 \MATRIX_ADD_reg[3]  (.D(n_0_71), .G(n_0_46), .Q(MATRIX_ADD[3]));
   DLH_X1 \MATRIX_ADD_reg[2]  (.D(n_0_70), .G(n_0_46), .Q(MATRIX_ADD[2]));
   DLH_X1 \MATRIX_ADD_reg[1]  (.D(n_0_69), .G(n_0_46), .Q(MATRIX_ADD[1]));
   DLH_X1 \MATRIX_ADD_reg[0]  (.D(n_0_68), .G(n_0_46), .Q(MATRIX_ADD[0]));
   DLH_X1 Interpolate_Enable_reg (.D(n_0_0), .G(n_0_181), .Q(Interpolate_Enable));
   DLH_X1 DONE_reg (.D(Back), .G(n_0_54), .Q(n_0_1));
   DLH_X1 \MATRIX_CNT_reg[15]  (.D(n_0_21), .G(n_0_26), .Q(MATRIX_CNT[15]));
   DLH_X1 \MATRIX_CNT_reg[14]  (.D(n_0_20), .G(n_0_26), .Q(MATRIX_CNT[14]));
   DLH_X1 \MATRIX_CNT_reg[13]  (.D(n_0_19), .G(n_0_26), .Q(MATRIX_CNT[13]));
   DLH_X1 \MATRIX_CNT_reg[12]  (.D(n_0_18), .G(n_0_26), .Q(MATRIX_CNT[12]));
   DLH_X1 \MATRIX_CNT_reg[11]  (.D(n_0_17), .G(n_0_26), .Q(MATRIX_CNT[11]));
   DLH_X1 \MATRIX_CNT_reg[10]  (.D(n_0_16), .G(n_0_26), .Q(MATRIX_CNT[10]));
   DLH_X1 \MATRIX_CNT_reg[9]  (.D(n_0_15), .G(n_0_26), .Q(MATRIX_CNT[9]));
   DLH_X1 \MATRIX_CNT_reg[8]  (.D(n_0_14), .G(n_0_26), .Q(MATRIX_CNT[8]));
   DLH_X1 \MATRIX_CNT_reg[7]  (.D(n_0_13), .G(n_0_26), .Q(MATRIX_CNT[7]));
   DLH_X1 \MATRIX_CNT_reg[6]  (.D(n_0_12), .G(n_0_26), .Q(MATRIX_CNT[6]));
   DLH_X1 \MATRIX_CNT_reg[5]  (.D(n_0_11), .G(n_0_26), .Q(MATRIX_CNT[5]));
   DLH_X1 \MATRIX_CNT_reg[4]  (.D(n_0_10), .G(n_0_26), .Q(MATRIX_CNT[4]));
   DLH_X1 \MATRIX_CNT_reg[3]  (.D(n_0_9), .G(n_0_26), .Q(MATRIX_CNT[3]));
   DLH_X1 \MATRIX_CNT_reg[2]  (.D(n_0_8), .G(n_0_26), .Q(MATRIX_CNT[2]));
   DLH_X1 \MATRIX_CNT_reg[1]  (.D(n_0_7), .G(n_0_26), .Q(MATRIX_CNT[1]));
   DLH_X1 \MATRIX_CNT_reg[0]  (.D(n_0_6), .G(n_0_26), .Q(MATRIX_CNT[0]));
   DLH_X1 \VECTOR_CNT_reg[15]  (.D(n_0_42), .G(n_0_46), .Q(VECTOR_CNT[15]));
   DLH_X1 \VECTOR_CNT_reg[14]  (.D(n_0_41), .G(n_0_46), .Q(VECTOR_CNT[14]));
   DLH_X1 \VECTOR_CNT_reg[13]  (.D(n_0_40), .G(n_0_46), .Q(VECTOR_CNT[13]));
   DLH_X1 \VECTOR_CNT_reg[12]  (.D(n_0_39), .G(n_0_46), .Q(VECTOR_CNT[12]));
   DLH_X1 \VECTOR_CNT_reg[11]  (.D(n_0_38), .G(n_0_46), .Q(VECTOR_CNT[11]));
   DLH_X1 \VECTOR_CNT_reg[10]  (.D(n_0_37), .G(n_0_46), .Q(VECTOR_CNT[10]));
   DLH_X1 \VECTOR_CNT_reg[9]  (.D(n_0_36), .G(n_0_46), .Q(VECTOR_CNT[9]));
   DLH_X1 \VECTOR_CNT_reg[8]  (.D(n_0_35), .G(n_0_46), .Q(VECTOR_CNT[8]));
   DLH_X1 \VECTOR_CNT_reg[7]  (.D(n_0_34), .G(n_0_46), .Q(VECTOR_CNT[7]));
   DLH_X1 \VECTOR_CNT_reg[6]  (.D(n_0_33), .G(n_0_46), .Q(VECTOR_CNT[6]));
   DLH_X1 \VECTOR_CNT_reg[5]  (.D(n_0_32), .G(n_0_46), .Q(VECTOR_CNT[5]));
   DLH_X1 \VECTOR_CNT_reg[4]  (.D(n_0_31), .G(n_0_46), .Q(VECTOR_CNT[4]));
   DLH_X1 \VECTOR_CNT_reg[3]  (.D(n_0_30), .G(n_0_46), .Q(VECTOR_CNT[3]));
   DLH_X1 \VECTOR_CNT_reg[2]  (.D(n_0_29), .G(n_0_46), .Q(VECTOR_CNT[2]));
   DLH_X1 \VECTOR_CNT_reg[1]  (.D(n_0_28), .G(n_0_46), .Q(VECTOR_CNT[1]));
   DLH_X1 \VECTOR_CNT_reg[0]  (.D(n_0_27), .G(n_0_46), .Q(VECTOR_CNT[0]));
   DLH_X1 \state_reg[2]  (.D(next[2]), .G(n_0_51), .Q(state[2]));
   DLH_X1 \state_reg[1]  (.D(next[1]), .G(n_0_51), .Q(state[1]));
   DLH_X1 \state_reg[0]  (.D(next[0]), .G(n_0_51), .Q(state[0]));
   DLH_X1 \next_reg[2]  (.D(n_0_4), .G(n_0_5), .Q(next[2]));
   DLH_X1 \next_reg[1]  (.D(n_0_3), .G(n_0_5), .Q(next[1]));
   DLH_X1 \next_reg[0]  (.D(n_0_2), .G(n_0_5), .Q(next[0]));
   DLH_X1 \counter_reg[1]  (.D(n_0_49), .G(n_0_50), .Q(counter[1]));
   DLH_X1 \counter_reg[0]  (.D(n_0_48), .G(n_0_50), .Q(counter[0]));
   DLH_X1 Matrix_Multiplication1_Enable_reg (.D(n_0_22), .G(n_0_23), .Q(
      Matrix_Multiplication1_Enable));
   DLH_X1 Matrix_Multiplication2_Enable_reg (.D(n_0_24), .G(n_0_25), .Q(
      Matrix_Multiplication2_Enable));
   DLH_X1 Final_Calc_Enable_reg (.D(n_0_44), .G(n_0_45), .Q(Final_Calc_Enable));
   DLH_X1 Back_reg (.D(n_0_52), .G(n_0_53), .Q(Back));
   DLH_X1 \n_val_reg[63]  (.D(RAM_DATA_RD1[63]), .G(n_0_43), .Q(n_val[63]));
   DLH_X1 \n_val_reg[62]  (.D(RAM_DATA_RD1[62]), .G(n_0_43), .Q(n_val[62]));
   DLH_X1 \n_val_reg[61]  (.D(RAM_DATA_RD1[61]), .G(n_0_43), .Q(n_val[61]));
   DLH_X1 \n_val_reg[60]  (.D(RAM_DATA_RD1[60]), .G(n_0_43), .Q(n_val[60]));
   DLH_X1 \n_val_reg[59]  (.D(RAM_DATA_RD1[59]), .G(n_0_43), .Q(n_val[59]));
   DLH_X1 \n_val_reg[58]  (.D(RAM_DATA_RD1[58]), .G(n_0_43), .Q(n_val[58]));
   DLH_X1 \n_val_reg[57]  (.D(RAM_DATA_RD1[57]), .G(n_0_43), .Q(n_val[57]));
   DLH_X1 \n_val_reg[56]  (.D(RAM_DATA_RD1[56]), .G(n_0_43), .Q(n_val[56]));
   DLH_X1 \n_val_reg[55]  (.D(RAM_DATA_RD1[55]), .G(n_0_43), .Q(n_val[55]));
   DLH_X1 \n_val_reg[54]  (.D(RAM_DATA_RD1[54]), .G(n_0_43), .Q(n_val[54]));
   DLH_X1 \n_val_reg[53]  (.D(RAM_DATA_RD1[53]), .G(n_0_43), .Q(n_val[53]));
   DLH_X1 \n_val_reg[52]  (.D(RAM_DATA_RD1[52]), .G(n_0_43), .Q(n_val[52]));
   DLH_X1 \n_val_reg[51]  (.D(RAM_DATA_RD1[51]), .G(n_0_43), .Q(n_val[51]));
   DLH_X1 \n_val_reg[50]  (.D(RAM_DATA_RD1[50]), .G(n_0_43), .Q(n_val[50]));
   DLH_X1 \n_val_reg[49]  (.D(RAM_DATA_RD1[49]), .G(n_0_43), .Q(n_val[49]));
   DLH_X1 \n_val_reg[48]  (.D(RAM_DATA_RD1[48]), .G(n_0_43), .Q(n_val[48]));
   DLH_X1 \n_val_reg[47]  (.D(RAM_DATA_RD1[47]), .G(n_0_43), .Q(n_val[47]));
   DLH_X1 \n_val_reg[46]  (.D(RAM_DATA_RD1[46]), .G(n_0_43), .Q(n_val[46]));
   DLH_X1 \n_val_reg[45]  (.D(RAM_DATA_RD1[45]), .G(n_0_43), .Q(n_val[45]));
   DLH_X1 \n_val_reg[44]  (.D(RAM_DATA_RD1[44]), .G(n_0_43), .Q(n_val[44]));
   DLH_X1 \n_val_reg[43]  (.D(RAM_DATA_RD1[43]), .G(n_0_43), .Q(n_val[43]));
   DLH_X1 \n_val_reg[42]  (.D(RAM_DATA_RD1[42]), .G(n_0_43), .Q(n_val[42]));
   DLH_X1 \n_val_reg[41]  (.D(RAM_DATA_RD1[41]), .G(n_0_43), .Q(n_val[41]));
   DLH_X1 \n_val_reg[40]  (.D(RAM_DATA_RD1[40]), .G(n_0_43), .Q(n_val[40]));
   DLH_X1 \n_val_reg[39]  (.D(RAM_DATA_RD1[39]), .G(n_0_43), .Q(n_val[39]));
   DLH_X1 \n_val_reg[38]  (.D(RAM_DATA_RD1[38]), .G(n_0_43), .Q(n_val[38]));
   DLH_X1 \n_val_reg[37]  (.D(RAM_DATA_RD1[37]), .G(n_0_43), .Q(n_val[37]));
   DLH_X1 \n_val_reg[36]  (.D(RAM_DATA_RD1[36]), .G(n_0_43), .Q(n_val[36]));
   DLH_X1 \n_val_reg[35]  (.D(RAM_DATA_RD1[35]), .G(n_0_43), .Q(n_val[35]));
   DLH_X1 \n_val_reg[34]  (.D(RAM_DATA_RD1[34]), .G(n_0_43), .Q(n_val[34]));
   DLH_X1 \n_val_reg[33]  (.D(RAM_DATA_RD1[33]), .G(n_0_43), .Q(n_val[33]));
   DLH_X1 \n_val_reg[32]  (.D(RAM_DATA_RD1[32]), .G(n_0_43), .Q(n_val[32]));
   DLH_X1 \n_val_reg[31]  (.D(RAM_DATA_RD1[31]), .G(n_0_43), .Q(n_val[31]));
   DLH_X1 \n_val_reg[30]  (.D(RAM_DATA_RD1[30]), .G(n_0_43), .Q(n_val[30]));
   DLH_X1 \n_val_reg[29]  (.D(RAM_DATA_RD1[29]), .G(n_0_43), .Q(n_val[29]));
   DLH_X1 \n_val_reg[28]  (.D(RAM_DATA_RD1[28]), .G(n_0_43), .Q(n_val[28]));
   DLH_X1 \n_val_reg[27]  (.D(RAM_DATA_RD1[27]), .G(n_0_43), .Q(n_val[27]));
   DLH_X1 \n_val_reg[26]  (.D(RAM_DATA_RD1[26]), .G(n_0_43), .Q(n_val[26]));
   DLH_X1 \n_val_reg[25]  (.D(RAM_DATA_RD1[25]), .G(n_0_43), .Q(n_val[25]));
   DLH_X1 \n_val_reg[24]  (.D(RAM_DATA_RD1[24]), .G(n_0_43), .Q(n_val[24]));
   DLH_X1 \n_val_reg[23]  (.D(RAM_DATA_RD1[23]), .G(n_0_43), .Q(n_val[23]));
   DLH_X1 \n_val_reg[22]  (.D(RAM_DATA_RD1[22]), .G(n_0_43), .Q(n_val[22]));
   DLH_X1 \n_val_reg[21]  (.D(RAM_DATA_RD1[21]), .G(n_0_43), .Q(n_val[21]));
   DLH_X1 \n_val_reg[20]  (.D(RAM_DATA_RD1[20]), .G(n_0_43), .Q(n_val[20]));
   DLH_X1 \n_val_reg[19]  (.D(RAM_DATA_RD1[19]), .G(n_0_43), .Q(n_val[19]));
   DLH_X1 \n_val_reg[18]  (.D(RAM_DATA_RD1[18]), .G(n_0_43), .Q(n_val[18]));
   DLH_X1 \n_val_reg[17]  (.D(RAM_DATA_RD1[17]), .G(n_0_43), .Q(n_val[17]));
   DLH_X1 \n_val_reg[16]  (.D(RAM_DATA_RD1[16]), .G(n_0_43), .Q(n_val[16]));
   DLH_X1 \n_val_reg[15]  (.D(RAM_DATA_RD1[15]), .G(n_0_43), .Q(n_val[15]));
   DLH_X1 \n_val_reg[14]  (.D(RAM_DATA_RD1[14]), .G(n_0_43), .Q(n_val[14]));
   DLH_X1 \n_val_reg[13]  (.D(RAM_DATA_RD1[13]), .G(n_0_43), .Q(n_val[13]));
   DLH_X1 \n_val_reg[12]  (.D(RAM_DATA_RD1[12]), .G(n_0_43), .Q(n_val[12]));
   DLH_X1 \n_val_reg[11]  (.D(RAM_DATA_RD1[11]), .G(n_0_43), .Q(n_val[11]));
   DLH_X1 \n_val_reg[10]  (.D(RAM_DATA_RD1[10]), .G(n_0_43), .Q(n_val[10]));
   DLH_X1 \n_val_reg[9]  (.D(RAM_DATA_RD1[9]), .G(n_0_43), .Q(n_val[9]));
   DLH_X1 \n_val_reg[8]  (.D(RAM_DATA_RD1[8]), .G(n_0_43), .Q(n_val[8]));
   DLH_X1 \n_val_reg[7]  (.D(RAM_DATA_RD1[7]), .G(n_0_43), .Q(n_val[7]));
   DLH_X1 \n_val_reg[6]  (.D(RAM_DATA_RD1[6]), .G(n_0_43), .Q(n_val[6]));
   DLH_X1 \n_val_reg[5]  (.D(RAM_DATA_RD1[5]), .G(n_0_43), .Q(n_val[5]));
   DLH_X1 \n_val_reg[4]  (.D(RAM_DATA_RD1[4]), .G(n_0_43), .Q(n_val[4]));
   DLH_X1 \n_val_reg[3]  (.D(RAM_DATA_RD1[3]), .G(n_0_43), .Q(n_val[3]));
   DLH_X1 \n_val_reg[2]  (.D(RAM_DATA_RD1[2]), .G(n_0_43), .Q(n_val[2]));
   DLH_X1 \n_val_reg[1]  (.D(RAM_DATA_RD1[1]), .G(n_0_43), .Q(n_val[1]));
   DLH_X1 \n_val_reg[0]  (.D(RAM_DATA_RD1[0]), .G(n_0_43), .Q(n_val[0]));
   DLH_X1 \m_val_reg[63]  (.D(RAM_DATA_RD2[63]), .G(n_0_43), .Q(m_val[63]));
   DLH_X1 \m_val_reg[62]  (.D(RAM_DATA_RD2[62]), .G(n_0_43), .Q(m_val[62]));
   DLH_X1 \m_val_reg[61]  (.D(RAM_DATA_RD2[61]), .G(n_0_43), .Q(m_val[61]));
   DLH_X1 \m_val_reg[60]  (.D(RAM_DATA_RD2[60]), .G(n_0_43), .Q(m_val[60]));
   DLH_X1 \m_val_reg[59]  (.D(RAM_DATA_RD2[59]), .G(n_0_43), .Q(m_val[59]));
   DLH_X1 \m_val_reg[58]  (.D(RAM_DATA_RD2[58]), .G(n_0_43), .Q(m_val[58]));
   DLH_X1 \m_val_reg[57]  (.D(RAM_DATA_RD2[57]), .G(n_0_43), .Q(m_val[57]));
   DLH_X1 \m_val_reg[56]  (.D(RAM_DATA_RD2[56]), .G(n_0_43), .Q(m_val[56]));
   DLH_X1 \m_val_reg[55]  (.D(RAM_DATA_RD2[55]), .G(n_0_43), .Q(m_val[55]));
   DLH_X1 \m_val_reg[54]  (.D(RAM_DATA_RD2[54]), .G(n_0_43), .Q(m_val[54]));
   DLH_X1 \m_val_reg[53]  (.D(RAM_DATA_RD2[53]), .G(n_0_43), .Q(m_val[53]));
   DLH_X1 \m_val_reg[52]  (.D(RAM_DATA_RD2[52]), .G(n_0_43), .Q(m_val[52]));
   DLH_X1 \m_val_reg[51]  (.D(RAM_DATA_RD2[51]), .G(n_0_43), .Q(m_val[51]));
   DLH_X1 \m_val_reg[50]  (.D(RAM_DATA_RD2[50]), .G(n_0_43), .Q(m_val[50]));
   DLH_X1 \m_val_reg[49]  (.D(RAM_DATA_RD2[49]), .G(n_0_43), .Q(m_val[49]));
   DLH_X1 \m_val_reg[48]  (.D(RAM_DATA_RD2[48]), .G(n_0_43), .Q(m_val[48]));
   DLH_X1 \m_val_reg[47]  (.D(RAM_DATA_RD2[47]), .G(n_0_43), .Q(m_val[47]));
   DLH_X1 \m_val_reg[46]  (.D(RAM_DATA_RD2[46]), .G(n_0_43), .Q(m_val[46]));
   DLH_X1 \m_val_reg[45]  (.D(RAM_DATA_RD2[45]), .G(n_0_43), .Q(m_val[45]));
   DLH_X1 \m_val_reg[44]  (.D(RAM_DATA_RD2[44]), .G(n_0_43), .Q(m_val[44]));
   DLH_X1 \m_val_reg[43]  (.D(RAM_DATA_RD2[43]), .G(n_0_43), .Q(m_val[43]));
   DLH_X1 \m_val_reg[42]  (.D(RAM_DATA_RD2[42]), .G(n_0_43), .Q(m_val[42]));
   DLH_X1 \m_val_reg[41]  (.D(RAM_DATA_RD2[41]), .G(n_0_43), .Q(m_val[41]));
   DLH_X1 \m_val_reg[40]  (.D(RAM_DATA_RD2[40]), .G(n_0_43), .Q(m_val[40]));
   DLH_X1 \m_val_reg[39]  (.D(RAM_DATA_RD2[39]), .G(n_0_43), .Q(m_val[39]));
   DLH_X1 \m_val_reg[38]  (.D(RAM_DATA_RD2[38]), .G(n_0_43), .Q(m_val[38]));
   DLH_X1 \m_val_reg[37]  (.D(RAM_DATA_RD2[37]), .G(n_0_43), .Q(m_val[37]));
   DLH_X1 \m_val_reg[36]  (.D(RAM_DATA_RD2[36]), .G(n_0_43), .Q(m_val[36]));
   DLH_X1 \m_val_reg[35]  (.D(RAM_DATA_RD2[35]), .G(n_0_43), .Q(m_val[35]));
   DLH_X1 \m_val_reg[34]  (.D(RAM_DATA_RD2[34]), .G(n_0_43), .Q(m_val[34]));
   DLH_X1 \m_val_reg[33]  (.D(RAM_DATA_RD2[33]), .G(n_0_43), .Q(m_val[33]));
   DLH_X1 \m_val_reg[32]  (.D(RAM_DATA_RD2[32]), .G(n_0_43), .Q(m_val[32]));
   DLH_X1 \m_val_reg[31]  (.D(RAM_DATA_RD2[31]), .G(n_0_43), .Q(m_val[31]));
   DLH_X1 \m_val_reg[30]  (.D(RAM_DATA_RD2[30]), .G(n_0_43), .Q(m_val[30]));
   DLH_X1 \m_val_reg[29]  (.D(RAM_DATA_RD2[29]), .G(n_0_43), .Q(m_val[29]));
   DLH_X1 \m_val_reg[28]  (.D(RAM_DATA_RD2[28]), .G(n_0_43), .Q(m_val[28]));
   DLH_X1 \m_val_reg[27]  (.D(RAM_DATA_RD2[27]), .G(n_0_43), .Q(m_val[27]));
   DLH_X1 \m_val_reg[26]  (.D(RAM_DATA_RD2[26]), .G(n_0_43), .Q(m_val[26]));
   DLH_X1 \m_val_reg[25]  (.D(RAM_DATA_RD2[25]), .G(n_0_43), .Q(m_val[25]));
   DLH_X1 \m_val_reg[24]  (.D(RAM_DATA_RD2[24]), .G(n_0_43), .Q(m_val[24]));
   DLH_X1 \m_val_reg[23]  (.D(RAM_DATA_RD2[23]), .G(n_0_43), .Q(m_val[23]));
   DLH_X1 \m_val_reg[22]  (.D(RAM_DATA_RD2[22]), .G(n_0_43), .Q(m_val[22]));
   DLH_X1 \m_val_reg[21]  (.D(RAM_DATA_RD2[21]), .G(n_0_43), .Q(m_val[21]));
   DLH_X1 \m_val_reg[20]  (.D(RAM_DATA_RD2[20]), .G(n_0_43), .Q(m_val[20]));
   DLH_X1 \m_val_reg[19]  (.D(RAM_DATA_RD2[19]), .G(n_0_43), .Q(m_val[19]));
   DLH_X1 \m_val_reg[18]  (.D(RAM_DATA_RD2[18]), .G(n_0_43), .Q(m_val[18]));
   DLH_X1 \m_val_reg[17]  (.D(RAM_DATA_RD2[17]), .G(n_0_43), .Q(m_val[17]));
   DLH_X1 \m_val_reg[16]  (.D(RAM_DATA_RD2[16]), .G(n_0_43), .Q(m_val[16]));
   DLH_X1 \m_val_reg[15]  (.D(RAM_DATA_RD2[15]), .G(n_0_43), .Q(m_val[15]));
   DLH_X1 \m_val_reg[14]  (.D(RAM_DATA_RD2[14]), .G(n_0_43), .Q(m_val[14]));
   DLH_X1 \m_val_reg[13]  (.D(RAM_DATA_RD2[13]), .G(n_0_43), .Q(m_val[13]));
   DLH_X1 \m_val_reg[12]  (.D(RAM_DATA_RD2[12]), .G(n_0_43), .Q(m_val[12]));
   DLH_X1 \m_val_reg[11]  (.D(RAM_DATA_RD2[11]), .G(n_0_43), .Q(m_val[11]));
   DLH_X1 \m_val_reg[10]  (.D(RAM_DATA_RD2[10]), .G(n_0_43), .Q(m_val[10]));
   DLH_X1 \m_val_reg[9]  (.D(RAM_DATA_RD2[9]), .G(n_0_43), .Q(m_val[9]));
   DLH_X1 \m_val_reg[8]  (.D(RAM_DATA_RD2[8]), .G(n_0_43), .Q(m_val[8]));
   DLH_X1 \m_val_reg[7]  (.D(RAM_DATA_RD2[7]), .G(n_0_43), .Q(m_val[7]));
   DLH_X1 \m_val_reg[6]  (.D(RAM_DATA_RD2[6]), .G(n_0_43), .Q(m_val[6]));
   DLH_X1 \m_val_reg[5]  (.D(RAM_DATA_RD2[5]), .G(n_0_43), .Q(m_val[5]));
   DLH_X1 \m_val_reg[4]  (.D(RAM_DATA_RD2[4]), .G(n_0_43), .Q(m_val[4]));
   DLH_X1 \m_val_reg[3]  (.D(RAM_DATA_RD2[3]), .G(n_0_43), .Q(m_val[3]));
   DLH_X1 \m_val_reg[2]  (.D(RAM_DATA_RD2[2]), .G(n_0_43), .Q(m_val[2]));
   DLH_X1 \m_val_reg[1]  (.D(RAM_DATA_RD2[1]), .G(n_0_43), .Q(m_val[1]));
   DLH_X1 \m_val_reg[0]  (.D(RAM_DATA_RD2[0]), .G(n_0_43), .Q(m_val[0]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[12]  (.D(ELEMENT_adder_n_26), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[12]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[11]  (.D(ELEMENT_adder_n_25), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[11]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[10]  (.D(ELEMENT_adder_n_24), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[10]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[9]  (.D(ELEMENT_adder_n_23), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[9]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[8]  (.D(ELEMENT_adder_n_22), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[8]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[7]  (.D(ELEMENT_adder_n_21), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[7]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[6]  (.D(ELEMENT_adder_n_20), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[6]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[5]  (.D(ELEMENT_adder_n_19), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[5]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[4]  (.D(ELEMENT_adder_n_18), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[4]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[3]  (.D(ELEMENT_adder_n_17), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[3]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[2]  (.D(ELEMENT_adder_n_16), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[2]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[1]  (.D(ELEMENT_adder_n_15), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[1]));
   DLH_X1 \ELEMENT_adder_tempIn22_reg[0]  (.D(ELEMENT_adder_n_14), .G(
      ELEMENT_adder_n_27), .Q(ELEMENT_adder_tempIn22[0]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[12]  (.D(ELEMENT_adder_n_12), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[12]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[11]  (.D(ELEMENT_adder_n_11), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[11]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[10]  (.D(ELEMENT_adder_n_10), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[10]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[9]  (.D(ELEMENT_adder_n_9), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[9]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[8]  (.D(ELEMENT_adder_n_8), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[8]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[7]  (.D(ELEMENT_adder_n_7), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[7]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[6]  (.D(ELEMENT_adder_n_6), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[6]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[5]  (.D(ELEMENT_adder_n_5), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[5]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[4]  (.D(ELEMENT_adder_n_4), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[4]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[3]  (.D(ELEMENT_adder_n_3), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[3]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[2]  (.D(ELEMENT_adder_n_2), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[2]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[1]  (.D(ELEMENT_adder_n_1), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[1]));
   DLH_X1 \ELEMENT_adder_tempIn11_reg[0]  (.D(ELEMENT_adder_n_0), .G(
      ELEMENT_adder_n_13), .Q(ELEMENT_adder_tempIn11[0]));
   OAI22_X1 ELEMENT_adder_i_0_0 (.A1(ELEMENT_adder_n_0_89), .A2(
      ELEMENT_adder_n_13), .B1(ELEMENT_adder_n_0_93), .B2(ELEMENT_adder_n_0_82), 
      .ZN(NEW_Element_Result[13]));
   OAI22_X1 ELEMENT_adder_i_0_1 (.A1(ELEMENT_adder_n_0_90), .A2(
      ELEMENT_adder_n_13), .B1(ELEMENT_adder_n_0_94), .B2(ELEMENT_adder_n_0_82), 
      .ZN(NEW_Element_Result[14]));
   OR2_X1 ELEMENT_adder_i_0_2 (.A1(Multiplication_Result[15]), .A2(
      Element_Result[15]), .ZN(NEW_Element_Result[15]));
   AND2_X1 ELEMENT_adder_i_0_3 (.A1(Element_Result[0]), .A2(ELEMENT_adder_n_0_72), 
      .ZN(ELEMENT_adder_n_0));
   OAI22_X1 ELEMENT_adder_i_0_4 (.A1(ELEMENT_adder_n_0_3), .A2(
      ELEMENT_adder_n_0_0), .B1(ELEMENT_adder_n_0_75), .B2(ELEMENT_adder_n_0_6), 
      .ZN(ELEMENT_adder_n_1));
   OAI22_X1 ELEMENT_adder_i_0_5 (.A1(ELEMENT_adder_n_0_75), .A2(
      ELEMENT_adder_n_0_9), .B1(ELEMENT_adder_n_0_6), .B2(ELEMENT_adder_n_0_0), 
      .ZN(ELEMENT_adder_n_2));
   OAI22_X1 ELEMENT_adder_i_0_6 (.A1(ELEMENT_adder_n_0_75), .A2(
      ELEMENT_adder_n_0_12), .B1(ELEMENT_adder_n_0_9), .B2(ELEMENT_adder_n_0_0), 
      .ZN(ELEMENT_adder_n_3));
   OAI22_X1 ELEMENT_adder_i_0_7 (.A1(ELEMENT_adder_n_0_78), .A2(
      ELEMENT_adder_n_0_1), .B1(ELEMENT_adder_n_0_12), .B2(ELEMENT_adder_n_0_0), 
      .ZN(ELEMENT_adder_n_4));
   NAND2_X1 ELEMENT_adder_i_0_8 (.A1(ELEMENT_adder_n_0_78), .A2(
      ELEMENT_adder_n_0_77), .ZN(ELEMENT_adder_n_0_0));
   OAI22_X1 ELEMENT_adder_i_0_9 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_1), .B1(ELEMENT_adder_n_0_78), .B2(ELEMENT_adder_n_0_4), 
      .ZN(ELEMENT_adder_n_5));
   INV_X1 ELEMENT_adder_i_0_10 (.A(ELEMENT_adder_n_0_2), .ZN(ELEMENT_adder_n_0_1));
   OAI22_X1 ELEMENT_adder_i_0_11 (.A1(ELEMENT_adder_n_0_76), .A2(
      ELEMENT_adder_n_0_15), .B1(ELEMENT_adder_n_0_77), .B2(ELEMENT_adder_n_0_3), 
      .ZN(ELEMENT_adder_n_0_2));
   NAND2_X1 ELEMENT_adder_i_0_12 (.A1(Element_Result[0]), .A2(
      ELEMENT_adder_n_0_32), .ZN(ELEMENT_adder_n_0_3));
   OAI22_X1 ELEMENT_adder_i_0_13 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_4), .B1(ELEMENT_adder_n_0_78), .B2(ELEMENT_adder_n_0_7), 
      .ZN(ELEMENT_adder_n_6));
   INV_X1 ELEMENT_adder_i_0_14 (.A(ELEMENT_adder_n_0_5), .ZN(ELEMENT_adder_n_0_4));
   OAI22_X1 ELEMENT_adder_i_0_15 (.A1(ELEMENT_adder_n_0_76), .A2(
      ELEMENT_adder_n_0_18), .B1(ELEMENT_adder_n_0_77), .B2(ELEMENT_adder_n_0_6), 
      .ZN(ELEMENT_adder_n_0_5));
   NAND2_X1 ELEMENT_adder_i_0_16 (.A1(Element_Result[1]), .A2(
      ELEMENT_adder_n_0_32), .ZN(ELEMENT_adder_n_0_6));
   OAI22_X1 ELEMENT_adder_i_0_17 (.A1(ELEMENT_adder_n_0_78), .A2(
      ELEMENT_adder_n_0_10), .B1(ELEMENT_adder_n_0_79), .B2(ELEMENT_adder_n_0_7), 
      .ZN(ELEMENT_adder_n_7));
   INV_X1 ELEMENT_adder_i_0_18 (.A(ELEMENT_adder_n_0_8), .ZN(ELEMENT_adder_n_0_7));
   OAI22_X1 ELEMENT_adder_i_0_19 (.A1(ELEMENT_adder_n_0_77), .A2(
      ELEMENT_adder_n_0_9), .B1(ELEMENT_adder_n_0_76), .B2(ELEMENT_adder_n_0_22), 
      .ZN(ELEMENT_adder_n_0_8));
   AOI22_X1 ELEMENT_adder_i_0_20 (.A1(Element_Result[2]), .A2(
      ELEMENT_adder_n_0_32), .B1(Element_Result[0]), .B2(ELEMENT_adder_n_0_33), 
      .ZN(ELEMENT_adder_n_0_9));
   OAI22_X1 ELEMENT_adder_i_0_21 (.A1(ELEMENT_adder_n_0_78), .A2(
      ELEMENT_adder_n_0_13), .B1(ELEMENT_adder_n_0_79), .B2(ELEMENT_adder_n_0_10), 
      .ZN(ELEMENT_adder_n_8));
   INV_X1 ELEMENT_adder_i_0_22 (.A(ELEMENT_adder_n_0_11), .ZN(
      ELEMENT_adder_n_0_10));
   OAI22_X1 ELEMENT_adder_i_0_23 (.A1(ELEMENT_adder_n_0_77), .A2(
      ELEMENT_adder_n_0_12), .B1(ELEMENT_adder_n_0_76), .B2(ELEMENT_adder_n_0_26), 
      .ZN(ELEMENT_adder_n_0_11));
   AOI22_X1 ELEMENT_adder_i_0_24 (.A1(Element_Result[3]), .A2(
      ELEMENT_adder_n_0_32), .B1(Element_Result[1]), .B2(ELEMENT_adder_n_0_33), 
      .ZN(ELEMENT_adder_n_0_12));
   OAI22_X1 ELEMENT_adder_i_0_25 (.A1(ELEMENT_adder_n_0_78), .A2(
      ELEMENT_adder_n_0_16), .B1(ELEMENT_adder_n_0_79), .B2(ELEMENT_adder_n_0_13), 
      .ZN(ELEMENT_adder_n_9));
   INV_X1 ELEMENT_adder_i_0_26 (.A(ELEMENT_adder_n_0_14), .ZN(
      ELEMENT_adder_n_0_13));
   OAI22_X1 ELEMENT_adder_i_0_27 (.A1(ELEMENT_adder_n_0_77), .A2(
      ELEMENT_adder_n_0_15), .B1(ELEMENT_adder_n_0_76), .B2(ELEMENT_adder_n_0_30), 
      .ZN(ELEMENT_adder_n_0_14));
   AOI22_X1 ELEMENT_adder_i_0_28 (.A1(Element_Result[4]), .A2(
      ELEMENT_adder_n_0_32), .B1(Element_Result[2]), .B2(ELEMENT_adder_n_0_33), 
      .ZN(ELEMENT_adder_n_0_15));
   OAI22_X1 ELEMENT_adder_i_0_29 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_16), .B1(ELEMENT_adder_n_0_78), .B2(ELEMENT_adder_n_0_20), 
      .ZN(ELEMENT_adder_n_10));
   INV_X1 ELEMENT_adder_i_0_30 (.A(ELEMENT_adder_n_0_17), .ZN(
      ELEMENT_adder_n_0_16));
   OAI22_X1 ELEMENT_adder_i_0_31 (.A1(ELEMENT_adder_n_0_76), .A2(
      ELEMENT_adder_n_0_19), .B1(ELEMENT_adder_n_0_77), .B2(ELEMENT_adder_n_0_18), 
      .ZN(ELEMENT_adder_n_0_17));
   AOI22_X1 ELEMENT_adder_i_0_32 (.A1(Element_Result[5]), .A2(
      ELEMENT_adder_n_0_32), .B1(Element_Result[3]), .B2(ELEMENT_adder_n_0_33), 
      .ZN(ELEMENT_adder_n_0_18));
   AOI22_X1 ELEMENT_adder_i_0_33 (.A1(Element_Result[9]), .A2(
      ELEMENT_adder_n_0_32), .B1(Element_Result[7]), .B2(ELEMENT_adder_n_0_33), 
      .ZN(ELEMENT_adder_n_0_19));
   OAI22_X1 ELEMENT_adder_i_0_34 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_20), .B1(ELEMENT_adder_n_0_78), .B2(ELEMENT_adder_n_0_24), 
      .ZN(ELEMENT_adder_n_11));
   INV_X1 ELEMENT_adder_i_0_35 (.A(ELEMENT_adder_n_0_21), .ZN(
      ELEMENT_adder_n_0_20));
   OAI22_X1 ELEMENT_adder_i_0_36 (.A1(ELEMENT_adder_n_0_76), .A2(
      ELEMENT_adder_n_0_23), .B1(ELEMENT_adder_n_0_77), .B2(ELEMENT_adder_n_0_22), 
      .ZN(ELEMENT_adder_n_0_21));
   AOI22_X1 ELEMENT_adder_i_0_37 (.A1(Element_Result[6]), .A2(
      ELEMENT_adder_n_0_32), .B1(Element_Result[4]), .B2(ELEMENT_adder_n_0_33), 
      .ZN(ELEMENT_adder_n_0_22));
   AOI22_X1 ELEMENT_adder_i_0_38 (.A1(Element_Result[10]), .A2(
      ELEMENT_adder_n_0_32), .B1(Element_Result[8]), .B2(ELEMENT_adder_n_0_33), 
      .ZN(ELEMENT_adder_n_0_23));
   OAI22_X1 ELEMENT_adder_i_0_39 (.A1(ELEMENT_adder_n_0_78), .A2(
      ELEMENT_adder_n_0_28), .B1(ELEMENT_adder_n_0_79), .B2(ELEMENT_adder_n_0_24), 
      .ZN(ELEMENT_adder_n_12));
   INV_X1 ELEMENT_adder_i_0_40 (.A(ELEMENT_adder_n_0_25), .ZN(
      ELEMENT_adder_n_0_24));
   OAI22_X1 ELEMENT_adder_i_0_41 (.A1(ELEMENT_adder_n_0_76), .A2(
      ELEMENT_adder_n_0_27), .B1(ELEMENT_adder_n_0_77), .B2(ELEMENT_adder_n_0_26), 
      .ZN(ELEMENT_adder_n_0_25));
   AOI22_X1 ELEMENT_adder_i_0_42 (.A1(Element_Result[7]), .A2(
      ELEMENT_adder_n_0_32), .B1(Element_Result[5]), .B2(ELEMENT_adder_n_0_33), 
      .ZN(ELEMENT_adder_n_0_26));
   AOI22_X1 ELEMENT_adder_i_0_43 (.A1(Element_Result[9]), .A2(
      ELEMENT_adder_n_0_33), .B1(Element_Result[11]), .B2(ELEMENT_adder_n_0_32), 
      .ZN(ELEMENT_adder_n_0_27));
   INV_X1 ELEMENT_adder_i_0_44 (.A(ELEMENT_adder_n_0_29), .ZN(
      ELEMENT_adder_n_0_28));
   OAI22_X1 ELEMENT_adder_i_0_45 (.A1(ELEMENT_adder_n_0_76), .A2(
      ELEMENT_adder_n_0_31), .B1(ELEMENT_adder_n_0_77), .B2(ELEMENT_adder_n_0_30), 
      .ZN(ELEMENT_adder_n_0_29));
   AOI22_X1 ELEMENT_adder_i_0_46 (.A1(Element_Result[8]), .A2(
      ELEMENT_adder_n_0_32), .B1(Element_Result[6]), .B2(ELEMENT_adder_n_0_33), 
      .ZN(ELEMENT_adder_n_0_30));
   AOI22_X1 ELEMENT_adder_i_0_47 (.A1(Element_Result[10]), .A2(
      ELEMENT_adder_n_0_33), .B1(Element_Result[12]), .B2(ELEMENT_adder_n_0_32), 
      .ZN(ELEMENT_adder_n_0_31));
   INV_X1 ELEMENT_adder_i_0_48 (.A(ELEMENT_adder_n_0_33), .ZN(
      ELEMENT_adder_n_0_32));
   XOR2_X1 ELEMENT_adder_i_0_49 (.A(ELEMENT_adder_n_0_86), .B(
      ELEMENT_adder_n_0_73), .Z(ELEMENT_adder_n_0_33));
   AND2_X1 ELEMENT_adder_i_0_50 (.A1(Multiplication_Result[0]), .A2(
      ELEMENT_adder_n_0_72), .ZN(ELEMENT_adder_n_14));
   OAI22_X1 ELEMENT_adder_i_0_51 (.A1(ELEMENT_adder_n_0_37), .A2(
      ELEMENT_adder_n_0_34), .B1(ELEMENT_adder_n_0_92), .B2(ELEMENT_adder_n_0_71), 
      .ZN(ELEMENT_adder_n_15));
   OAI33_X1 ELEMENT_adder_i_0_52 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_69), .A3(ELEMENT_adder_n_0_40), .B1(ELEMENT_adder_n_0_78), 
      .B2(ELEMENT_adder_n_0_69), .B3(ELEMENT_adder_n_0_43), .ZN(
      ELEMENT_adder_n_16));
   OAI33_X1 ELEMENT_adder_i_0_53 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_69), .A3(ELEMENT_adder_n_0_43), .B1(ELEMENT_adder_n_0_78), 
      .B2(ELEMENT_adder_n_0_69), .B3(ELEMENT_adder_n_0_46), .ZN(
      ELEMENT_adder_n_17));
   OAI22_X1 ELEMENT_adder_i_0_54 (.A1(ELEMENT_adder_n_0_46), .A2(
      ELEMENT_adder_n_0_34), .B1(ELEMENT_adder_n_0_78), .B2(ELEMENT_adder_n_0_35), 
      .ZN(ELEMENT_adder_n_18));
   NAND2_X1 ELEMENT_adder_i_0_55 (.A1(ELEMENT_adder_n_0_78), .A2(
      ELEMENT_adder_n_0_68), .ZN(ELEMENT_adder_n_0_34));
   AOI22_X1 ELEMENT_adder_i_0_56 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_38), .B1(ELEMENT_adder_n_0_78), .B2(ELEMENT_adder_n_0_35), 
      .ZN(ELEMENT_adder_n_19));
   INV_X1 ELEMENT_adder_i_0_57 (.A(ELEMENT_adder_n_0_36), .ZN(
      ELEMENT_adder_n_0_35));
   OAI22_X1 ELEMENT_adder_i_0_58 (.A1(ELEMENT_adder_n_0_69), .A2(
      ELEMENT_adder_n_0_49), .B1(ELEMENT_adder_n_0_68), .B2(ELEMENT_adder_n_0_37), 
      .ZN(ELEMENT_adder_n_0_36));
   NAND2_X1 ELEMENT_adder_i_0_59 (.A1(Multiplication_Result[0]), .A2(
      ELEMENT_adder_n_0_67), .ZN(ELEMENT_adder_n_0_37));
   OAI22_X1 ELEMENT_adder_i_0_60 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_38), .B1(ELEMENT_adder_n_0_78), .B2(ELEMENT_adder_n_0_41), 
      .ZN(ELEMENT_adder_n_20));
   INV_X1 ELEMENT_adder_i_0_61 (.A(ELEMENT_adder_n_0_39), .ZN(
      ELEMENT_adder_n_0_38));
   OAI22_X1 ELEMENT_adder_i_0_62 (.A1(ELEMENT_adder_n_0_69), .A2(
      ELEMENT_adder_n_0_52), .B1(ELEMENT_adder_n_0_68), .B2(ELEMENT_adder_n_0_40), 
      .ZN(ELEMENT_adder_n_0_39));
   NAND2_X1 ELEMENT_adder_i_0_63 (.A1(Multiplication_Result[1]), .A2(
      ELEMENT_adder_n_0_67), .ZN(ELEMENT_adder_n_0_40));
   OAI22_X1 ELEMENT_adder_i_0_64 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_41), .B1(ELEMENT_adder_n_0_78), .B2(ELEMENT_adder_n_0_44), 
      .ZN(ELEMENT_adder_n_21));
   INV_X1 ELEMENT_adder_i_0_65 (.A(ELEMENT_adder_n_0_42), .ZN(
      ELEMENT_adder_n_0_41));
   OAI22_X1 ELEMENT_adder_i_0_66 (.A1(ELEMENT_adder_n_0_69), .A2(
      ELEMENT_adder_n_0_56), .B1(ELEMENT_adder_n_0_68), .B2(ELEMENT_adder_n_0_43), 
      .ZN(ELEMENT_adder_n_0_42));
   AOI22_X1 ELEMENT_adder_i_0_67 (.A1(Multiplication_Result[2]), .A2(
      ELEMENT_adder_n_0_67), .B1(Multiplication_Result[0]), .B2(
      ELEMENT_adder_n_0_66), .ZN(ELEMENT_adder_n_0_43));
   OAI22_X1 ELEMENT_adder_i_0_68 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_44), .B1(ELEMENT_adder_n_0_78), .B2(ELEMENT_adder_n_0_47), 
      .ZN(ELEMENT_adder_n_22));
   INV_X1 ELEMENT_adder_i_0_69 (.A(ELEMENT_adder_n_0_45), .ZN(
      ELEMENT_adder_n_0_44));
   OAI22_X1 ELEMENT_adder_i_0_70 (.A1(ELEMENT_adder_n_0_69), .A2(
      ELEMENT_adder_n_0_60), .B1(ELEMENT_adder_n_0_68), .B2(ELEMENT_adder_n_0_46), 
      .ZN(ELEMENT_adder_n_0_45));
   AOI22_X1 ELEMENT_adder_i_0_71 (.A1(Multiplication_Result[3]), .A2(
      ELEMENT_adder_n_0_67), .B1(Multiplication_Result[1]), .B2(
      ELEMENT_adder_n_0_66), .ZN(ELEMENT_adder_n_0_46));
   OAI22_X1 ELEMENT_adder_i_0_72 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_47), .B1(ELEMENT_adder_n_0_78), .B2(ELEMENT_adder_n_0_50), 
      .ZN(ELEMENT_adder_n_23));
   INV_X1 ELEMENT_adder_i_0_73 (.A(ELEMENT_adder_n_0_48), .ZN(
      ELEMENT_adder_n_0_47));
   OAI22_X1 ELEMENT_adder_i_0_74 (.A1(ELEMENT_adder_n_0_69), .A2(
      ELEMENT_adder_n_0_64), .B1(ELEMENT_adder_n_0_68), .B2(ELEMENT_adder_n_0_49), 
      .ZN(ELEMENT_adder_n_0_48));
   AOI22_X1 ELEMENT_adder_i_0_75 (.A1(Multiplication_Result[4]), .A2(
      ELEMENT_adder_n_0_67), .B1(Multiplication_Result[2]), .B2(
      ELEMENT_adder_n_0_66), .ZN(ELEMENT_adder_n_0_49));
   OAI22_X1 ELEMENT_adder_i_0_76 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_50), .B1(ELEMENT_adder_n_0_78), .B2(ELEMENT_adder_n_0_54), 
      .ZN(ELEMENT_adder_n_24));
   INV_X1 ELEMENT_adder_i_0_77 (.A(ELEMENT_adder_n_0_51), .ZN(
      ELEMENT_adder_n_0_50));
   OAI22_X1 ELEMENT_adder_i_0_78 (.A1(ELEMENT_adder_n_0_69), .A2(
      ELEMENT_adder_n_0_53), .B1(ELEMENT_adder_n_0_68), .B2(ELEMENT_adder_n_0_52), 
      .ZN(ELEMENT_adder_n_0_51));
   AOI22_X1 ELEMENT_adder_i_0_79 (.A1(Multiplication_Result[5]), .A2(
      ELEMENT_adder_n_0_67), .B1(Multiplication_Result[3]), .B2(
      ELEMENT_adder_n_0_66), .ZN(ELEMENT_adder_n_0_52));
   AOI22_X1 ELEMENT_adder_i_0_80 (.A1(Multiplication_Result[9]), .A2(
      ELEMENT_adder_n_0_67), .B1(Multiplication_Result[7]), .B2(
      ELEMENT_adder_n_0_66), .ZN(ELEMENT_adder_n_0_53));
   OAI22_X1 ELEMENT_adder_i_0_81 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_54), .B1(ELEMENT_adder_n_0_78), .B2(ELEMENT_adder_n_0_58), 
      .ZN(ELEMENT_adder_n_25));
   INV_X1 ELEMENT_adder_i_0_82 (.A(ELEMENT_adder_n_0_55), .ZN(
      ELEMENT_adder_n_0_54));
   OAI22_X1 ELEMENT_adder_i_0_83 (.A1(ELEMENT_adder_n_0_69), .A2(
      ELEMENT_adder_n_0_57), .B1(ELEMENT_adder_n_0_68), .B2(ELEMENT_adder_n_0_56), 
      .ZN(ELEMENT_adder_n_0_55));
   AOI22_X1 ELEMENT_adder_i_0_84 (.A1(Multiplication_Result[6]), .A2(
      ELEMENT_adder_n_0_67), .B1(Multiplication_Result[4]), .B2(
      ELEMENT_adder_n_0_66), .ZN(ELEMENT_adder_n_0_56));
   AOI22_X1 ELEMENT_adder_i_0_85 (.A1(Multiplication_Result[10]), .A2(
      ELEMENT_adder_n_0_67), .B1(Multiplication_Result[8]), .B2(
      ELEMENT_adder_n_0_66), .ZN(ELEMENT_adder_n_0_57));
   OAI22_X1 ELEMENT_adder_i_0_86 (.A1(ELEMENT_adder_n_0_78), .A2(
      ELEMENT_adder_n_0_62), .B1(ELEMENT_adder_n_0_79), .B2(ELEMENT_adder_n_0_58), 
      .ZN(ELEMENT_adder_n_26));
   INV_X1 ELEMENT_adder_i_0_87 (.A(ELEMENT_adder_n_0_59), .ZN(
      ELEMENT_adder_n_0_58));
   OAI22_X1 ELEMENT_adder_i_0_88 (.A1(ELEMENT_adder_n_0_69), .A2(
      ELEMENT_adder_n_0_61), .B1(ELEMENT_adder_n_0_68), .B2(ELEMENT_adder_n_0_60), 
      .ZN(ELEMENT_adder_n_0_59));
   AOI22_X1 ELEMENT_adder_i_0_89 (.A1(Multiplication_Result[7]), .A2(
      ELEMENT_adder_n_0_67), .B1(Multiplication_Result[5]), .B2(
      ELEMENT_adder_n_0_66), .ZN(ELEMENT_adder_n_0_60));
   AOI22_X1 ELEMENT_adder_i_0_90 (.A1(Multiplication_Result[9]), .A2(
      ELEMENT_adder_n_0_66), .B1(Multiplication_Result[11]), .B2(
      ELEMENT_adder_n_0_67), .ZN(ELEMENT_adder_n_0_61));
   INV_X1 ELEMENT_adder_i_0_91 (.A(ELEMENT_adder_n_0_63), .ZN(
      ELEMENT_adder_n_0_62));
   OAI22_X1 ELEMENT_adder_i_0_92 (.A1(ELEMENT_adder_n_0_69), .A2(
      ELEMENT_adder_n_0_65), .B1(ELEMENT_adder_n_0_68), .B2(ELEMENT_adder_n_0_64), 
      .ZN(ELEMENT_adder_n_0_63));
   AOI22_X1 ELEMENT_adder_i_0_93 (.A1(Multiplication_Result[8]), .A2(
      ELEMENT_adder_n_0_67), .B1(Multiplication_Result[6]), .B2(
      ELEMENT_adder_n_0_66), .ZN(ELEMENT_adder_n_0_64));
   AOI22_X1 ELEMENT_adder_i_0_94 (.A1(Multiplication_Result[10]), .A2(
      ELEMENT_adder_n_0_66), .B1(Multiplication_Result[12]), .B2(
      ELEMENT_adder_n_0_67), .ZN(ELEMENT_adder_n_0_65));
   INV_X1 ELEMENT_adder_i_0_95 (.A(ELEMENT_adder_n_0_67), .ZN(
      ELEMENT_adder_n_0_66));
   OAI22_X1 ELEMENT_adder_i_0_96 (.A1(ELEMENT_adder_n_0_81), .A2(
      ELEMENT_adder_n_0_73), .B1(ELEMENT_adder_n_0_80), .B2(ELEMENT_adder_n_0_74), 
      .ZN(ELEMENT_adder_n_0_67));
   INV_X1 ELEMENT_adder_i_0_97 (.A(ELEMENT_adder_n_0_69), .ZN(
      ELEMENT_adder_n_0_68));
   XOR2_X1 ELEMENT_adder_i_0_98 (.A(ELEMENT_adder_n_0_83), .B(
      ELEMENT_adder_n_0_70), .Z(ELEMENT_adder_n_0_69));
   AOI21_X1 ELEMENT_adder_i_0_99 (.A(ELEMENT_adder_n_0_85), .B1(
      ELEMENT_adder_n_0_87), .B2(ELEMENT_adder_n_0_80), .ZN(ELEMENT_adder_n_0_70));
   NAND2_X1 ELEMENT_adder_i_0_100 (.A1(ELEMENT_adder_n_13), .A2(
      ELEMENT_adder_n_0_71), .ZN(ELEMENT_adder_n_27));
   INV_X1 ELEMENT_adder_i_0_101 (.A(ELEMENT_adder_n_0_72), .ZN(
      ELEMENT_adder_n_0_71));
   NOR2_X1 ELEMENT_adder_i_0_102 (.A1(ELEMENT_adder_n_0_75), .A2(
      ELEMENT_adder_n_0_73), .ZN(ELEMENT_adder_n_0_72));
   INV_X1 ELEMENT_adder_i_0_103 (.A(ELEMENT_adder_n_0_74), .ZN(
      ELEMENT_adder_n_0_73));
   NOR2_X1 ELEMENT_adder_i_0_104 (.A1(ELEMENT_adder_n_0_88), .A2(
      ELEMENT_adder_n_0_85), .ZN(ELEMENT_adder_n_0_74));
   NAND2_X1 ELEMENT_adder_i_0_105 (.A1(ELEMENT_adder_n_0_79), .A2(
      ELEMENT_adder_n_0_77), .ZN(ELEMENT_adder_n_0_75));
   INV_X1 ELEMENT_adder_i_0_106 (.A(ELEMENT_adder_n_0_77), .ZN(
      ELEMENT_adder_n_0_76));
   XOR2_X1 ELEMENT_adder_i_0_107 (.A(ELEMENT_adder_n_0_84), .B(
      ELEMENT_adder_n_0_83), .Z(ELEMENT_adder_n_0_77));
   INV_X1 ELEMENT_adder_i_0_108 (.A(ELEMENT_adder_n_0_79), .ZN(
      ELEMENT_adder_n_0_78));
   NOR2_X1 ELEMENT_adder_i_0_109 (.A1(ELEMENT_adder_n_0_86), .A2(
      ELEMENT_adder_n_0_81), .ZN(ELEMENT_adder_n_0_79));
   INV_X1 ELEMENT_adder_i_0_110 (.A(ELEMENT_adder_n_0_81), .ZN(
      ELEMENT_adder_n_0_80));
   NOR2_X1 ELEMENT_adder_i_0_111 (.A1(ELEMENT_adder_n_0_93), .A2(
      Element_Result[13]), .ZN(ELEMENT_adder_n_0_81));
   INV_X1 ELEMENT_adder_i_0_112 (.A(ELEMENT_adder_n_0_82), .ZN(
      ELEMENT_adder_n_13));
   OAI22_X1 ELEMENT_adder_i_0_113 (.A1(Multiplication_Result[15]), .A2(
      ELEMENT_adder_n_0_91), .B1(ELEMENT_adder_n_0_84), .B2(ELEMENT_adder_n_0_83), 
      .ZN(ELEMENT_adder_n_0_82));
   XNOR2_X1 ELEMENT_adder_i_0_114 (.A(Multiplication_Result[15]), .B(
      ELEMENT_adder_n_0_91), .ZN(ELEMENT_adder_n_0_83));
   OAI21_X1 ELEMENT_adder_i_0_115 (.A(ELEMENT_adder_n_0_87), .B1(
      ELEMENT_adder_n_0_86), .B2(ELEMENT_adder_n_0_85), .ZN(ELEMENT_adder_n_0_84));
   NOR2_X1 ELEMENT_adder_i_0_116 (.A1(Multiplication_Result[14]), .A2(
      ELEMENT_adder_n_0_90), .ZN(ELEMENT_adder_n_0_85));
   NOR2_X1 ELEMENT_adder_i_0_117 (.A1(Multiplication_Result[13]), .A2(
      ELEMENT_adder_n_0_89), .ZN(ELEMENT_adder_n_0_86));
   INV_X1 ELEMENT_adder_i_0_118 (.A(ELEMENT_adder_n_0_88), .ZN(
      ELEMENT_adder_n_0_87));
   NOR2_X1 ELEMENT_adder_i_0_119 (.A1(ELEMENT_adder_n_0_94), .A2(
      Element_Result[14]), .ZN(ELEMENT_adder_n_0_88));
   INV_X1 ELEMENT_adder_i_0_120 (.A(Element_Result[13]), .ZN(
      ELEMENT_adder_n_0_89));
   INV_X1 ELEMENT_adder_i_0_121 (.A(Element_Result[14]), .ZN(
      ELEMENT_adder_n_0_90));
   INV_X1 ELEMENT_adder_i_0_122 (.A(Element_Result[15]), .ZN(
      ELEMENT_adder_n_0_91));
   INV_X1 ELEMENT_adder_i_0_123 (.A(Multiplication_Result[1]), .ZN(
      ELEMENT_adder_n_0_92));
   INV_X1 ELEMENT_adder_i_0_124 (.A(Multiplication_Result[13]), .ZN(
      ELEMENT_adder_n_0_93));
   INV_X1 ELEMENT_adder_i_0_125 (.A(Multiplication_Result[14]), .ZN(
      ELEMENT_adder_n_0_94));
   XOR2_X1 ELEMENT_adder_i_1_0 (.A(ELEMENT_adder_tempIn22[0]), .B(
      ELEMENT_adder_tempIn11[0]), .Z(NEW_Element_Result[0]));
   XNOR2_X1 ELEMENT_adder_i_1_1 (.A(ELEMENT_adder_n_1_43), .B(
      ELEMENT_adder_n_1_0), .ZN(NEW_Element_Result[1]));
   XOR2_X1 ELEMENT_adder_i_1_2 (.A(ELEMENT_adder_tempIn22[1]), .B(
      ELEMENT_adder_tempIn11[1]), .Z(ELEMENT_adder_n_1_0));
   XNOR2_X1 ELEMENT_adder_i_1_3 (.A(ELEMENT_adder_n_1_40), .B(
      ELEMENT_adder_n_1_1), .ZN(NEW_Element_Result[2]));
   XNOR2_X1 ELEMENT_adder_i_1_4 (.A(ELEMENT_adder_tempIn22[2]), .B(
      ELEMENT_adder_tempIn11[2]), .ZN(ELEMENT_adder_n_1_1));
   XNOR2_X1 ELEMENT_adder_i_1_5 (.A(ELEMENT_adder_n_1_35), .B(
      ELEMENT_adder_n_1_3), .ZN(NEW_Element_Result[4]));
   XNOR2_X1 ELEMENT_adder_i_1_6 (.A(ELEMENT_adder_tempIn22[4]), .B(
      ELEMENT_adder_tempIn11[4]), .ZN(ELEMENT_adder_n_1_3));
   XNOR2_X1 ELEMENT_adder_i_1_7 (.A(ELEMENT_adder_n_1_32), .B(
      ELEMENT_adder_n_1_4), .ZN(NEW_Element_Result[5]));
   XOR2_X1 ELEMENT_adder_i_1_8 (.A(ELEMENT_adder_tempIn22[5]), .B(
      ELEMENT_adder_tempIn11[5]), .Z(ELEMENT_adder_n_1_4));
   XNOR2_X1 ELEMENT_adder_i_1_9 (.A(ELEMENT_adder_n_1_29), .B(
      ELEMENT_adder_n_1_5), .ZN(NEW_Element_Result[6]));
   XNOR2_X1 ELEMENT_adder_i_1_10 (.A(ELEMENT_adder_tempIn22[6]), .B(
      ELEMENT_adder_tempIn11[6]), .ZN(ELEMENT_adder_n_1_5));
   XNOR2_X1 ELEMENT_adder_i_1_11 (.A(ELEMENT_adder_n_1_25), .B(
      ELEMENT_adder_n_1_6), .ZN(NEW_Element_Result[7]));
   XOR2_X1 ELEMENT_adder_i_1_12 (.A(ELEMENT_adder_tempIn22[7]), .B(
      ELEMENT_adder_tempIn11[7]), .Z(ELEMENT_adder_n_1_6));
   XNOR2_X1 ELEMENT_adder_i_1_13 (.A(ELEMENT_adder_n_1_23), .B(
      ELEMENT_adder_n_1_7), .ZN(NEW_Element_Result[8]));
   XNOR2_X1 ELEMENT_adder_i_1_14 (.A(ELEMENT_adder_tempIn22[8]), .B(
      ELEMENT_adder_tempIn11[8]), .ZN(ELEMENT_adder_n_1_7));
   XNOR2_X1 ELEMENT_adder_i_1_19 (.A(ELEMENT_adder_n_1_17), .B(
      ELEMENT_adder_n_1_9), .ZN(NEW_Element_Result[10]));
   XNOR2_X1 ELEMENT_adder_i_1_20 (.A(ELEMENT_adder_tempIn22[10]), .B(
      ELEMENT_adder_tempIn11[10]), .ZN(ELEMENT_adder_n_1_9));
   XNOR2_X1 ELEMENT_adder_i_1_21 (.A(ELEMENT_adder_n_1_14), .B(
      ELEMENT_adder_n_1_10), .ZN(NEW_Element_Result[11]));
   XOR2_X1 ELEMENT_adder_i_1_22 (.A(ELEMENT_adder_tempIn22[11]), .B(
      ELEMENT_adder_tempIn11[11]), .Z(ELEMENT_adder_n_1_10));
   XNOR2_X1 ELEMENT_adder_i_1_15 (.A(ELEMENT_adder_n_1_45), .B(
      ELEMENT_adder_n_1_11), .ZN(NEW_Element_Result[12]));
   OAI21_X1 ELEMENT_adder_i_1_16 (.A(ELEMENT_adder_n_1_12), .B1(
      ELEMENT_adder_n_1_14), .B2(ELEMENT_adder_n_1_13), .ZN(ELEMENT_adder_n_1_11));
   NAND2_X1 ELEMENT_adder_i_1_17 (.A1(ELEMENT_adder_tempIn22[11]), .A2(
      ELEMENT_adder_tempIn11[11]), .ZN(ELEMENT_adder_n_1_12));
   NOR2_X1 ELEMENT_adder_i_1_18 (.A1(ELEMENT_adder_tempIn22[11]), .A2(
      ELEMENT_adder_tempIn11[11]), .ZN(ELEMENT_adder_n_1_13));
   OAI21_X1 ELEMENT_adder_i_1_23 (.A(ELEMENT_adder_n_1_15), .B1(
      ELEMENT_adder_tempIn11[10]), .B2(ELEMENT_adder_tempIn22[10]), .ZN(
      ELEMENT_adder_n_1_14));
   INV_X1 ELEMENT_adder_i_1_24 (.A(ELEMENT_adder_n_1_16), .ZN(
      ELEMENT_adder_n_1_15));
   AOI21_X1 ELEMENT_adder_i_1_25 (.A(ELEMENT_adder_n_1_17), .B1(
      ELEMENT_adder_tempIn11[10]), .B2(ELEMENT_adder_tempIn22[10]), .ZN(
      ELEMENT_adder_n_1_16));
   AOI21_X1 ELEMENT_adder_i_1_26 (.A(ELEMENT_adder_n_1_18), .B1(
      ELEMENT_adder_n_1_19), .B2(ELEMENT_adder_n_1_20), .ZN(ELEMENT_adder_n_1_17));
   NOR2_X1 ELEMENT_adder_i_1_27 (.A1(ELEMENT_adder_tempIn22[9]), .A2(
      ELEMENT_adder_tempIn11[9]), .ZN(ELEMENT_adder_n_1_18));
   NAND2_X1 ELEMENT_adder_i_1_28 (.A1(ELEMENT_adder_tempIn22[9]), .A2(
      ELEMENT_adder_tempIn11[9]), .ZN(ELEMENT_adder_n_1_19));
   AOI21_X1 ELEMENT_adder_i_1_29 (.A(ELEMENT_adder_n_1_35), .B1(
      ELEMENT_adder_tempIn11[4]), .B2(ELEMENT_adder_tempIn22[4]), .ZN(
      ELEMENT_adder_n_1_34));
   AOI21_X1 ELEMENT_adder_i_1_30 (.A(ELEMENT_adder_n_1_36), .B1(
      ELEMENT_adder_n_1_37), .B2(ELEMENT_adder_n_1_38), .ZN(ELEMENT_adder_n_1_35));
   NOR2_X1 ELEMENT_adder_i_1_31 (.A1(ELEMENT_adder_tempIn22[3]), .A2(
      ELEMENT_adder_tempIn11[3]), .ZN(ELEMENT_adder_n_1_36));
   NAND2_X1 ELEMENT_adder_i_1_32 (.A1(ELEMENT_adder_tempIn22[3]), .A2(
      ELEMENT_adder_tempIn11[3]), .ZN(ELEMENT_adder_n_1_37));
   XNOR2_X1 ELEMENT_adder_i_1_33 (.A(ELEMENT_adder_tempIn22[12]), .B(
      ELEMENT_adder_tempIn11[12]), .ZN(ELEMENT_adder_n_1_45));
   XOR2_X1 ELEMENT_adder_i_1_34 (.A(ELEMENT_adder_n_1_38), .B(
      ELEMENT_adder_i_1_n_0), .Z(NEW_Element_Result[3]));
   XNOR2_X1 ELEMENT_adder_i_1_35 (.A(ELEMENT_adder_tempIn22[3]), .B(
      ELEMENT_adder_tempIn11[3]), .ZN(ELEMENT_adder_i_1_n_0));
   OAI22_X1 ELEMENT_adder_i_1_36 (.A1(ELEMENT_adder_tempIn22[2]), .A2(
      ELEMENT_adder_tempIn11[2]), .B1(ELEMENT_adder_n_1_40), .B2(
      ELEMENT_adder_i_1_n_1), .ZN(ELEMENT_adder_n_1_38));
   AND2_X1 ELEMENT_adder_i_1_37 (.A1(ELEMENT_adder_tempIn22[2]), .A2(
      ELEMENT_adder_tempIn11[2]), .ZN(ELEMENT_adder_i_1_n_1));
   OAI22_X1 ELEMENT_adder_i_1_38 (.A1(ELEMENT_adder_i_1_n_4), .A2(
      ELEMENT_adder_i_1_n_3), .B1(ELEMENT_adder_n_1_43), .B2(
      ELEMENT_adder_i_1_n_2), .ZN(ELEMENT_adder_n_1_40));
   NOR2_X1 ELEMENT_adder_i_1_39 (.A1(ELEMENT_adder_tempIn22[1]), .A2(
      ELEMENT_adder_tempIn11[1]), .ZN(ELEMENT_adder_i_1_n_2));
   NAND2_X1 ELEMENT_adder_i_1_40 (.A1(ELEMENT_adder_tempIn22[0]), .A2(
      ELEMENT_adder_tempIn11[0]), .ZN(ELEMENT_adder_n_1_43));
   INV_X1 ELEMENT_adder_i_1_41 (.A(ELEMENT_adder_tempIn11[1]), .ZN(
      ELEMENT_adder_i_1_n_3));
   INV_X1 ELEMENT_adder_i_1_42 (.A(ELEMENT_adder_tempIn22[1]), .ZN(
      ELEMENT_adder_i_1_n_4));
   XOR2_X1 ELEMENT_adder_i_1_43 (.A(ELEMENT_adder_n_1_20), .B(
      ELEMENT_adder_i_1_n_5), .Z(NEW_Element_Result[9]));
   XNOR2_X1 ELEMENT_adder_i_1_44 (.A(ELEMENT_adder_tempIn22[9]), .B(
      ELEMENT_adder_tempIn11[9]), .ZN(ELEMENT_adder_i_1_n_5));
   AOI22_X1 ELEMENT_adder_i_1_45 (.A1(ELEMENT_adder_tempIn22[8]), .A2(
      ELEMENT_adder_tempIn11[8]), .B1(ELEMENT_adder_n_1_23), .B2(
      ELEMENT_adder_i_1_n_6), .ZN(ELEMENT_adder_n_1_20));
   OR2_X1 ELEMENT_adder_i_1_46 (.A1(ELEMENT_adder_tempIn22[8]), .A2(
      ELEMENT_adder_tempIn11[8]), .ZN(ELEMENT_adder_i_1_n_6));
   OAI21_X1 ELEMENT_adder_i_1_47 (.A(ELEMENT_adder_i_1_n_8), .B1(
      ELEMENT_adder_n_1_25), .B2(ELEMENT_adder_i_1_n_7), .ZN(
      ELEMENT_adder_n_1_23));
   NOR2_X1 ELEMENT_adder_i_1_48 (.A1(ELEMENT_adder_tempIn22[7]), .A2(
      ELEMENT_adder_tempIn11[7]), .ZN(ELEMENT_adder_i_1_n_7));
   NAND2_X1 ELEMENT_adder_i_1_49 (.A1(ELEMENT_adder_tempIn22[7]), .A2(
      ELEMENT_adder_tempIn11[7]), .ZN(ELEMENT_adder_i_1_n_8));
   AOI22_X1 ELEMENT_adder_i_1_50 (.A1(ELEMENT_adder_tempIn22[6]), .A2(
      ELEMENT_adder_tempIn11[6]), .B1(ELEMENT_adder_n_1_29), .B2(
      ELEMENT_adder_i_1_n_9), .ZN(ELEMENT_adder_n_1_25));
   OR2_X1 ELEMENT_adder_i_1_51 (.A1(ELEMENT_adder_tempIn22[6]), .A2(
      ELEMENT_adder_tempIn11[6]), .ZN(ELEMENT_adder_i_1_n_9));
   OAI21_X1 ELEMENT_adder_i_1_52 (.A(ELEMENT_adder_i_1_n_11), .B1(
      ELEMENT_adder_n_1_32), .B2(ELEMENT_adder_i_1_n_10), .ZN(
      ELEMENT_adder_n_1_29));
   NOR2_X1 ELEMENT_adder_i_1_53 (.A1(ELEMENT_adder_tempIn22[5]), .A2(
      ELEMENT_adder_tempIn11[5]), .ZN(ELEMENT_adder_i_1_n_10));
   NAND2_X1 ELEMENT_adder_i_1_54 (.A1(ELEMENT_adder_tempIn22[5]), .A2(
      ELEMENT_adder_tempIn11[5]), .ZN(ELEMENT_adder_i_1_n_11));
   OAI21_X1 ELEMENT_adder_i_1_55 (.A(ELEMENT_adder_i_1_n_12), .B1(
      ELEMENT_adder_tempIn22[4]), .B2(ELEMENT_adder_tempIn11[4]), .ZN(
      ELEMENT_adder_n_1_32));
   INV_X1 ELEMENT_adder_i_1_56 (.A(ELEMENT_adder_n_1_34), .ZN(
      ELEMENT_adder_i_1_n_12));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[12]  (.D(VECTOR_CNT_adder_n_24), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[12]));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[11]  (.D(VECTOR_CNT_adder_n_23), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[11]));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[10]  (.D(VECTOR_CNT_adder_n_22), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[10]));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[9]  (.D(VECTOR_CNT_adder_n_21), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[9]));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[8]  (.D(VECTOR_CNT_adder_n_20), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[8]));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[7]  (.D(VECTOR_CNT_adder_n_19), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[7]));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[6]  (.D(VECTOR_CNT_adder_n_31), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[6]));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[5]  (.D(VECTOR_CNT_adder_n_30), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[5]));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[4]  (.D(VECTOR_CNT_adder_n_29), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[4]));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[3]  (.D(VECTOR_CNT_adder_n_28), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[3]));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[2]  (.D(VECTOR_CNT_adder_n_27), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[2]));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[1]  (.D(VECTOR_CNT_adder_n_26), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[1]));
   DLH_X1 \VECTOR_CNT_adder_tempIn11_reg[0]  (.D(VECTOR_CNT_adder_n_25), 
      .G(VECTOR_CNT_adder_n_2), .Q(VECTOR_CNT_adder_tempIn11[0]));
   INV_X1 i_0_70 (.A(n_0_22), .ZN(n_0_0));
   AND2_X1 i_0_0_0 (.A1(VECTOR_CNT[0]), .A2(VECTOR_CNT_adder_n_2), .ZN(
      VECTOR_CNT_adder_n_25));
   INV_X1 i_0_0_1 (.A(n_0_0_0), .ZN(VECTOR_CNT_adder_n_26));
   AOI22_X1 i_0_0_2 (.A1(VECTOR_CNT[1]), .A2(VECTOR_CNT_adder_n_2), .B1(n_0_0_9), 
      .B2(VECTOR_CNT[0]), .ZN(n_0_0_0));
   NAND2_X1 i_0_0_3 (.A1(n_0_0_1), .A2(n_0_0_2), .ZN(VECTOR_CNT_adder_n_27));
   AOI22_X1 i_0_0_4 (.A1(VECTOR_CNT[2]), .A2(VECTOR_CNT_adder_n_2), .B1(n_0_0_9), 
      .B2(VECTOR_CNT[1]), .ZN(n_0_0_1));
   NAND3_X1 i_0_0_5 (.A1(VECTOR_CNT[15]), .A2(VECTOR_CNT[0]), .A3(n_0_0_7), 
      .ZN(n_0_0_2));
   OAI211_X1 i_0_0_6 (.A(n_0_0_8), .B(n_0_0_6), .C1(VECTOR_CNT[13]), .C2(
      n_0_0_31), .ZN(VECTOR_CNT_adder_n_29));
   NAND3_X1 i_0_0_7 (.A1(VECTOR_CNT[15]), .A2(VECTOR_CNT[1]), .A3(n_0_0_5), 
      .ZN(n_0_0_6));
   NAND2_X1 i_0_0_8 (.A1(VECTOR_CNT[3]), .A2(n_0_0_9), .ZN(n_0_0_8));
   AOI21_X1 i_0_0_9 (.A(n_0_0_12), .B1(n_0_0_30), .B2(VECTOR_CNT[13]), .ZN(
      VECTOR_CNT_adder_n_31));
   NOR2_X1 i_0_0_10 (.A1(n_0_0_14), .A2(VECTOR_CNT[13]), .ZN(n_0_0_12));
   MUX2_X1 i_0_0_11 (.A(n_0_0_17), .B(n_0_0_14), .S(VECTOR_CNT[13]), .Z(
      VECTOR_CNT_adder_n_19));
   NAND2_X1 i_0_0_12 (.A1(n_0_0_16), .A2(n_0_0_15), .ZN(n_0_0_14));
   AOI22_X1 i_0_0_13 (.A1(n_0_0_33), .A2(VECTOR_CNT[6]), .B1(VECTOR_CNT[2]), 
      .B2(n_0_0_34), .ZN(n_0_0_15));
   AOI22_X1 i_0_0_14 (.A1(VECTOR_CNT[0]), .A2(n_0_0_47), .B1(n_0_0_32), .B2(
      VECTOR_CNT[4]), .ZN(n_0_0_16));
   MUX2_X1 i_0_0_15 (.A(n_0_0_20), .B(n_0_0_17), .S(VECTOR_CNT[13]), .Z(
      VECTOR_CNT_adder_n_20));
   NAND2_X1 i_0_0_16 (.A1(n_0_0_19), .A2(n_0_0_18), .ZN(n_0_0_17));
   AOI22_X1 i_0_0_17 (.A1(n_0_0_33), .A2(VECTOR_CNT[7]), .B1(VECTOR_CNT[3]), 
      .B2(n_0_0_34), .ZN(n_0_0_18));
   AOI22_X1 i_0_0_18 (.A1(VECTOR_CNT[1]), .A2(n_0_0_47), .B1(n_0_0_32), .B2(
      VECTOR_CNT[5]), .ZN(n_0_0_19));
   MUX2_X1 i_0_0_19 (.A(n_0_0_23), .B(n_0_0_20), .S(VECTOR_CNT[13]), .Z(
      VECTOR_CNT_adder_n_21));
   NAND2_X1 i_0_0_20 (.A1(n_0_0_22), .A2(n_0_0_21), .ZN(n_0_0_20));
   AOI22_X1 i_0_0_21 (.A1(VECTOR_CNT[2]), .A2(n_0_0_47), .B1(n_0_0_34), .B2(
      VECTOR_CNT[4]), .ZN(n_0_0_21));
   AOI22_X1 i_0_0_22 (.A1(VECTOR_CNT[8]), .A2(n_0_0_33), .B1(n_0_0_32), .B2(
      VECTOR_CNT[6]), .ZN(n_0_0_22));
   MUX2_X1 i_0_0_33 (.A(n_0_0_26), .B(n_0_0_23), .S(VECTOR_CNT[13]), .Z(
      VECTOR_CNT_adder_n_22));
   NAND2_X1 i_0_0_23 (.A1(n_0_0_25), .A2(n_0_0_24), .ZN(n_0_0_23));
   AOI22_X1 i_0_0_24 (.A1(n_0_0_33), .A2(VECTOR_CNT[9]), .B1(VECTOR_CNT[5]), 
      .B2(n_0_0_34), .ZN(n_0_0_24));
   AOI22_X1 i_0_0_25 (.A1(VECTOR_CNT[3]), .A2(n_0_0_47), .B1(n_0_0_32), .B2(
      VECTOR_CNT[7]), .ZN(n_0_0_25));
   MUX2_X1 i_0_0_37 (.A(n_0_0_41), .B(n_0_0_26), .S(VECTOR_CNT[13]), .Z(
      VECTOR_CNT_adder_n_23));
   NAND2_X1 i_0_0_38 (.A1(n_0_0_28), .A2(n_0_0_27), .ZN(n_0_0_26));
   AOI22_X1 i_0_0_39 (.A1(n_0_0_33), .A2(VECTOR_CNT[10]), .B1(VECTOR_CNT[6]), 
      .B2(n_0_0_34), .ZN(n_0_0_27));
   AOI22_X1 i_0_0_40 (.A1(VECTOR_CNT[4]), .A2(n_0_0_47), .B1(n_0_0_32), .B2(
      VECTOR_CNT[8]), .ZN(n_0_0_28));
   AND2_X1 i_0_0_26 (.A1(n_0_0_44), .A2(INT), .ZN(n_0_2));
   OAI33_X1 i_0_0_27 (.A1(n_0_1), .A2(PROCESS), .A3(n_0_0_119), .B1(n_0_0_322), 
      .B2(n_0_0_401), .B3(n_0_0_45), .ZN(n_0_0_44));
   NAND2_X1 i_0_0_28 (.A1(n_0_0_336), .A2(PROCESS), .ZN(n_0_0_45));
   NOR2_X1 i_0_0_29 (.A1(n_0_0_46), .A2(n_0_0_186), .ZN(n_0_3));
   AOI21_X1 i_0_0_30 (.A(n_0_0_400), .B1(n_0_0_324), .B2(state[0]), .ZN(n_0_0_46));
   OR2_X1 i_0_0_31 (.A1(n_0_0_66), .A2(n_0_0_48), .ZN(n_0_5));
   NAND2_X1 i_0_0_32 (.A1(n_0_0_96), .A2(n_0_0_67), .ZN(n_0_0_66));
   AOI211_X1 i_0_0_34 (.A(n_0_0_186), .B(n_0_0_68), .C1(state[0]), .C2(n_0_0_322), 
      .ZN(n_0_0_67));
   AOI21_X1 i_0_0_35 (.A(n_0_0_69), .B1(n_0_0_242), .B2(n_0_1), .ZN(n_0_0_68));
   OAI21_X1 i_0_0_36 (.A(n_0_0_342), .B1(n_0_0_247), .B2(Interpolate_DONE), 
      .ZN(n_0_0_69));
   NOR2_X1 i_0_0_41 (.A1(n_0_0_238), .A2(MATRIX_CNT_adder_tempIn11[0]), .ZN(
      n_0_6));
   AOI21_X1 i_0_0_42 (.A(n_0_0_70), .B1(MATRIX_CNT_adder_tempIn11[0]), .B2(
      MATRIX_CNT_adder_tempIn11[1]), .ZN(n_0_7));
   OAI21_X1 i_0_0_43 (.A(n_0_0_239), .B1(MATRIX_CNT_adder_tempIn11[0]), .B2(
      MATRIX_CNT_adder_tempIn11[1]), .ZN(n_0_0_70));
   NOR3_X1 i_0_0_44 (.A1(n_0_0_238), .A2(n_0_0_91), .A3(n_0_0_71), .ZN(n_0_8));
   AOI21_X1 i_0_0_45 (.A(MATRIX_CNT_adder_tempIn11[2]), .B1(
      MATRIX_CNT_adder_tempIn11[1]), .B2(MATRIX_CNT_adder_tempIn11[0]), .ZN(
      n_0_0_71));
   NOR3_X1 i_0_0_46 (.A1(n_0_0_238), .A2(n_0_0_90), .A3(n_0_0_72), .ZN(n_0_9));
   NOR2_X1 i_0_0_47 (.A1(MATRIX_CNT_adder_tempIn11[3]), .A2(n_0_0_91), .ZN(
      n_0_0_72));
   NOR2_X1 i_0_0_48 (.A1(n_0_0_89), .A2(n_0_0_73), .ZN(n_0_10));
   OAI21_X1 i_0_0_49 (.A(n_0_0_239), .B1(n_0_0_90), .B2(
      MATRIX_CNT_adder_tempIn11[4]), .ZN(n_0_0_73));
   NOR2_X1 i_0_0_50 (.A1(n_0_0_88), .A2(n_0_0_74), .ZN(n_0_11));
   OAI21_X1 i_0_0_51 (.A(n_0_0_239), .B1(n_0_0_89), .B2(
      MATRIX_CNT_adder_tempIn11[5]), .ZN(n_0_0_74));
   NOR2_X1 i_0_0_52 (.A1(n_0_0_87), .A2(n_0_0_75), .ZN(n_0_12));
   OAI21_X1 i_0_0_53 (.A(n_0_0_239), .B1(n_0_0_88), .B2(
      MATRIX_CNT_adder_tempIn11[6]), .ZN(n_0_0_75));
   NOR2_X1 i_0_0_54 (.A1(n_0_0_86), .A2(n_0_0_76), .ZN(n_0_13));
   OAI21_X1 i_0_0_55 (.A(n_0_0_239), .B1(n_0_0_87), .B2(
      MATRIX_CNT_adder_tempIn11[7]), .ZN(n_0_0_76));
   NOR2_X1 i_0_0_56 (.A1(n_0_0_85), .A2(n_0_0_77), .ZN(n_0_14));
   OAI21_X1 i_0_0_57 (.A(n_0_0_239), .B1(n_0_0_86), .B2(
      MATRIX_CNT_adder_tempIn11[8]), .ZN(n_0_0_77));
   NOR2_X1 i_0_0_58 (.A1(n_0_0_84), .A2(n_0_0_78), .ZN(n_0_15));
   OAI21_X1 i_0_0_59 (.A(n_0_0_239), .B1(n_0_0_85), .B2(
      MATRIX_CNT_adder_tempIn11[9]), .ZN(n_0_0_78));
   NOR2_X1 i_0_0_60 (.A1(n_0_0_83), .A2(n_0_0_79), .ZN(n_0_16));
   OAI21_X1 i_0_0_61 (.A(n_0_0_239), .B1(n_0_0_84), .B2(
      MATRIX_CNT_adder_tempIn11[10]), .ZN(n_0_0_79));
   AOI21_X1 i_0_0_62 (.A(n_0_0_80), .B1(n_0_0_83), .B2(
      MATRIX_CNT_adder_tempIn11[11]), .ZN(n_0_17));
   OAI21_X1 i_0_0_63 (.A(n_0_0_239), .B1(n_0_0_83), .B2(
      MATRIX_CNT_adder_tempIn11[11]), .ZN(n_0_0_80));
   NOR2_X1 i_0_0_64 (.A1(n_0_0_81), .A2(n_0_0_238), .ZN(n_0_18));
   XOR2_X1 i_0_0_65 (.A(MATRIX_CNT_adder_tempIn11[12]), .B(n_0_0_82), .Z(
      n_0_0_81));
   NAND2_X1 i_0_0_66 (.A1(MATRIX_CNT_adder_tempIn11[11]), .A2(n_0_0_83), 
      .ZN(n_0_0_82));
   AND2_X1 i_0_0_67 (.A1(MATRIX_CNT_adder_tempIn11[10]), .A2(n_0_0_84), .ZN(
      n_0_0_83));
   AND2_X1 i_0_0_68 (.A1(MATRIX_CNT_adder_tempIn11[9]), .A2(n_0_0_85), .ZN(
      n_0_0_84));
   AND2_X1 i_0_0_69 (.A1(MATRIX_CNT_adder_tempIn11[8]), .A2(n_0_0_86), .ZN(
      n_0_0_85));
   AND2_X1 i_0_0_70 (.A1(MATRIX_CNT_adder_tempIn11[7]), .A2(n_0_0_87), .ZN(
      n_0_0_86));
   AND2_X1 i_0_0_71 (.A1(MATRIX_CNT_adder_tempIn11[6]), .A2(n_0_0_88), .ZN(
      n_0_0_87));
   AND2_X1 i_0_0_72 (.A1(MATRIX_CNT_adder_tempIn11[5]), .A2(n_0_0_89), .ZN(
      n_0_0_88));
   AND2_X1 i_0_0_73 (.A1(MATRIX_CNT_adder_tempIn11[4]), .A2(n_0_0_90), .ZN(
      n_0_0_89));
   AND2_X1 i_0_0_74 (.A1(MATRIX_CNT_adder_tempIn11[3]), .A2(n_0_0_91), .ZN(
      n_0_0_90));
   AND3_X1 i_0_0_75 (.A1(MATRIX_CNT_adder_tempIn11[2]), .A2(
      MATRIX_CNT_adder_tempIn11[1]), .A3(MATRIX_CNT_adder_tempIn11[0]), .ZN(
      n_0_0_91));
   NOR2_X1 i_0_0_76 (.A1(n_0_0_472), .A2(n_0_0_238), .ZN(n_0_19));
   NOR2_X1 i_0_0_122 (.A1(n_0_0_473), .A2(n_0_0_238), .ZN(n_0_20));
   NOR2_X1 i_0_0_123 (.A1(n_0_0_476), .A2(n_0_0_238), .ZN(n_0_21));
   OR2_X1 i_0_0_77 (.A1(n_0_0_240), .A2(n_0_22), .ZN(n_0_23));
   AND3_X1 i_0_0_78 (.A1(state[1]), .A2(Interpolate_DONE), .A3(n_0_4), .ZN(
      n_0_22));
   NOR3_X1 i_0_0_79 (.A1(n_0_0_322), .A2(n_0_53), .A3(n_0_0_186), .ZN(n_0_4));
   OR2_X1 i_0_0_80 (.A1(n_0_0_316), .A2(n_0_24), .ZN(n_0_25));
   NOR3_X1 i_0_0_81 (.A1(n_0_0_96), .A2(state[0]), .A3(n_0_0_186), .ZN(n_0_24));
   INV_X1 i_0_0_82 (.A(n_0_0_92), .ZN(n_0_26));
   AOI21_X1 i_0_0_83 (.A(n_0_0_238), .B1(n_0_0_266), .B2(n_0_0_396), .ZN(
      n_0_0_92));
   NOR2_X1 i_0_0_84 (.A1(n_0_0_147), .A2(VECTOR_CNT_adder_tempIn11[0]), .ZN(
      n_0_27));
   NOR2_X1 i_0_0_132 (.A1(n_0_0_356), .A2(n_0_0_147), .ZN(n_0_28));
   NOR2_X1 i_0_0_133 (.A1(n_0_0_357), .A2(n_0_0_147), .ZN(n_0_29));
   AOI21_X1 i_0_0_134 (.A(n_0_0_93), .B1(n_0_0_358), .B2(
      VECTOR_CNT_adder_tempIn11[3]), .ZN(n_0_30));
   OAI21_X1 i_0_0_135 (.A(n_0_0_148), .B1(n_0_0_358), .B2(
      VECTOR_CNT_adder_tempIn11[3]), .ZN(n_0_0_93));
   NOR2_X1 i_0_0_136 (.A1(n_0_0_378), .A2(n_0_0_147), .ZN(n_0_31));
   NOR2_X1 i_0_0_137 (.A1(n_0_0_374), .A2(n_0_0_147), .ZN(n_0_32));
   NOR2_X1 i_0_0_138 (.A1(n_0_0_369), .A2(n_0_0_147), .ZN(n_0_33));
   NOR2_X1 i_0_0_139 (.A1(n_0_0_445), .A2(n_0_0_147), .ZN(n_0_34));
   NOR2_X1 i_0_0_140 (.A1(n_0_0_365), .A2(n_0_0_147), .ZN(n_0_35));
   NOR2_X1 i_0_0_141 (.A1(n_0_0_377), .A2(n_0_0_147), .ZN(n_0_36));
   NOR2_X1 i_0_0_142 (.A1(n_0_0_398), .A2(n_0_0_147), .ZN(n_0_37));
   NOR3_X1 i_0_0_143 (.A1(n_0_0_147), .A2(n_0_0_94), .A3(n_0_0_406), .ZN(n_0_38));
   NOR2_X1 i_0_0_144 (.A1(VECTOR_CNT_adder_tempIn11[11]), .A2(n_0_0_395), 
      .ZN(n_0_0_94));
   AOI21_X1 i_0_0_145 (.A(n_0_0_95), .B1(n_0_0_406), .B2(
      VECTOR_CNT_adder_tempIn11[12]), .ZN(n_0_39));
   OAI21_X1 i_0_0_146 (.A(n_0_0_148), .B1(n_0_0_406), .B2(
      VECTOR_CNT_adder_tempIn11[12]), .ZN(n_0_0_95));
   AND2_X1 i_0_0_147 (.A1(VECTOR_CNT[13]), .A2(n_0_0_148), .ZN(n_0_40));
   NOR2_X1 i_0_0_148 (.A1(n_0_0_13), .A2(n_0_0_147), .ZN(n_0_41));
   NOR2_X1 i_0_0_149 (.A1(n_0_0_29), .A2(n_0_0_147), .ZN(n_0_42));
   NOR3_X1 i_0_0_150 (.A1(n_0_0_298), .A2(state[0]), .A3(state[2]), .ZN(n_0_43));
   OR2_X1 i_0_0_151 (.A1(n_0_0_493), .A2(n_0_44), .ZN(n_0_45));
   NOR3_X1 i_0_0_152 (.A1(n_0_0_336), .A2(n_0_0_186), .A3(n_0_0_96), .ZN(n_0_44));
   OR4_X1 i_0_0_85 (.A1(n_0_0_181), .A2(n_0_0_116), .A3(n_0_0_111), .A4(n_0_0_97), 
      .ZN(n_0_0_96));
   NAND4_X1 i_0_0_86 (.A1(n_0_0_98), .A2(n_0_0_108), .A3(n_0_0_109), .A4(
      n_0_0_110), .ZN(n_0_0_97));
   NOR3_X1 i_0_0_87 (.A1(n_0_0_106), .A2(n_0_0_104), .A3(n_0_0_99), .ZN(n_0_0_98));
   NAND3_X1 i_0_0_88 (.A1(n_0_0_103), .A2(n_0_0_102), .A3(n_0_0_100), .ZN(
      n_0_0_99));
   AOI221_X1 i_0_0_89 (.A(n_0_0_101), .B1(n_val[5]), .B2(n_0_0_483), .C1(
      MATRIX_CNT[6]), .C2(n_0_0_474), .ZN(n_0_0_100));
   OAI22_X1 i_0_0_90 (.A1(MATRIX_CNT[6]), .A2(n_0_0_474), .B1(n_0_0_306), 
      .B2(MATRIX_CNT[1]), .ZN(n_0_0_101));
   XNOR2_X1 i_0_0_91 (.A(MATRIX_CNT[2]), .B(n_val[2]), .ZN(n_0_0_102));
   XNOR2_X1 i_0_0_92 (.A(MATRIX_CNT[9]), .B(n_val[9]), .ZN(n_0_0_103));
   OAI211_X1 i_0_0_93 (.A(n_0_0_324), .B(n_0_0_105), .C1(n_0_0_482), .C2(
      n_val[4]), .ZN(n_0_0_104));
   AOI22_X1 i_0_0_94 (.A1(n_0_0_482), .A2(n_val[4]), .B1(n_0_0_475), .B2(
      MATRIX_CNT[7]), .ZN(n_0_0_105));
   OAI221_X1 i_0_0_95 (.A(n_0_0_107), .B1(n_0_0_305), .B2(MATRIX_CNT[0]), 
      .C1(n_0_0_483), .C2(n_val[5]), .ZN(n_0_0_106));
   AOI22_X1 i_0_0_96 (.A1(n_0_0_484), .A2(n_val[7]), .B1(n_0_0_305), .B2(
      MATRIX_CNT[0]), .ZN(n_0_0_107));
   XNOR2_X1 i_0_0_97 (.A(MATRIX_CNT[8]), .B(n_val[8]), .ZN(n_0_0_108));
   XNOR2_X1 i_0_0_98 (.A(MATRIX_CNT[12]), .B(n_val[12]), .ZN(n_0_0_109));
   XNOR2_X1 i_0_0_99 (.A(MATRIX_CNT[14]), .B(n_val[14]), .ZN(n_0_0_110));
   NAND3_X1 i_0_0_100 (.A1(n_0_0_114), .A2(n_0_0_113), .A3(n_0_0_112), .ZN(
      n_0_0_111));
   AOI22_X1 i_0_0_101 (.A1(n_0_0_472), .A2(n_val[13]), .B1(n_0_0_307), .B2(
      MATRIX_CNT[3]), .ZN(n_0_0_112));
   AOI22_X1 i_0_0_102 (.A1(MATRIX_CNT[13]), .A2(n_0_0_313), .B1(n_0_0_306), 
      .B2(MATRIX_CNT[1]), .ZN(n_0_0_113));
   AOI221_X1 i_0_0_103 (.A(n_0_0_115), .B1(n_val[10]), .B2(n_0_0_486), .C1(
      n_0_0_476), .C2(n_val[15]), .ZN(n_0_0_114));
   OAI22_X1 i_0_0_104 (.A1(n_0_0_476), .A2(n_val[15]), .B1(n_0_0_307), .B2(
      MATRIX_CNT[3]), .ZN(n_0_0_115));
   OAI21_X1 i_0_0_105 (.A(n_0_0_117), .B1(n_0_0_311), .B2(MATRIX_CNT[11]), 
      .ZN(n_0_0_116));
   AOI22_X1 i_0_0_106 (.A1(MATRIX_CNT[11]), .A2(n_0_0_311), .B1(n_0_0_310), 
      .B2(MATRIX_CNT[10]), .ZN(n_0_0_117));
   AND2_X1 i_0_0_107 (.A1(n_0_0_118), .A2(n_0_0_326), .ZN(n_0_48));
   AND3_X1 i_0_0_108 (.A1(n_0_0_463), .A2(n_0_0_118), .A3(counter[0]), .ZN(
      n_0_49));
   OAI21_X1 i_0_0_109 (.A(n_0_0_118), .B1(n_0_0_327), .B2(CLK), .ZN(n_0_50));
   INV_X1 i_0_0_110 (.A(n_0_0_119), .ZN(n_0_0_118));
   NOR3_X1 i_0_0_111 (.A1(n_0_0_336), .A2(state[1]), .A3(state[2]), .ZN(
      n_0_0_119));
   AOI21_X1 i_0_0_112 (.A(state[2]), .B1(state[1]), .B2(state[0]), .ZN(n_0_53));
   AND2_X1 i_0_0_113 (.A1(Back), .A2(n_0_0_399), .ZN(n_0_54));
   OAI21_X1 i_0_0_182 (.A(n_0_0_315), .B1(n_0_0_185), .B2(n_0_0_120), .ZN(n_0_55));
   AOI222_X1 i_0_0_183 (.A1(NEW_MATRIX_ADD[0]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[0]), .C1(n_0_0_135), .C2(VECTOR_ADD[0]), .ZN(n_0_0_120));
   OAI21_X1 i_0_0_184 (.A(n_0_0_315), .B1(n_0_0_185), .B2(n_0_0_121), .ZN(n_0_56));
   AOI222_X1 i_0_0_185 (.A1(NEW_MATRIX_ADD[1]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[1]), .C1(n_0_0_135), .C2(VECTOR_ADD[1]), .ZN(n_0_0_121));
   OR2_X1 i_0_0_186 (.A1(n_0_0_122), .A2(n_0_0_199), .ZN(n_0_57));
   AOI21_X1 i_0_0_187 (.A(n_0_0_182), .B1(n_0_0_124), .B2(n_0_0_123), .ZN(
      n_0_0_122));
   AOI22_X1 i_0_0_188 (.A1(NEW_MATRIX_ADD[2]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[2]), .ZN(n_0_0_123));
   AOI21_X1 i_0_0_189 (.A(n_0_0_155), .B1(n_0_0_135), .B2(VECTOR_ADD[2]), 
      .ZN(n_0_0_124));
   OAI21_X1 i_0_0_190 (.A(n_0_0_323), .B1(n_0_0_125), .B2(n_0_0_182), .ZN(n_0_58));
   AOI222_X1 i_0_0_191 (.A1(NEW_MATRIX_ADD[3]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[3]), .C1(n_0_0_135), .C2(VECTOR_ADD[3]), .ZN(n_0_0_125));
   OAI21_X1 i_0_0_192 (.A(n_0_0_319), .B1(n_0_0_126), .B2(n_0_0_182), .ZN(n_0_59));
   AOI222_X1 i_0_0_193 (.A1(NEW_MATRIX_ADD[4]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[4]), .C1(n_0_0_135), .C2(VECTOR_ADD[4]), .ZN(n_0_0_126));
   NOR2_X1 i_0_0_194 (.A1(n_0_0_127), .A2(n_0_0_182), .ZN(n_0_60));
   AOI222_X1 i_0_0_195 (.A1(NEW_MATRIX_ADD[5]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[5]), .C1(n_0_0_135), .C2(VECTOR_ADD[5]), .ZN(n_0_0_127));
   OAI21_X1 i_0_0_196 (.A(n_0_0_347), .B1(n_0_0_128), .B2(n_0_0_182), .ZN(n_0_61));
   AOI222_X1 i_0_0_197 (.A1(NEW_MATRIX_ADD[6]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[6]), .C1(n_0_0_135), .C2(VECTOR_ADD[6]), .ZN(n_0_0_128));
   OAI21_X1 i_0_0_198 (.A(n_0_0_323), .B1(n_0_0_129), .B2(n_0_0_182), .ZN(n_0_62));
   AOI222_X1 i_0_0_199 (.A1(NEW_MATRIX_ADD[7]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[7]), .C1(n_0_0_135), .C2(VECTOR_ADD[7]), .ZN(n_0_0_129));
   OAI21_X1 i_0_0_200 (.A(n_0_0_323), .B1(n_0_0_130), .B2(n_0_0_182), .ZN(n_0_63));
   AOI222_X1 i_0_0_201 (.A1(NEW_MATRIX_ADD[8]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[8]), .C1(n_0_0_135), .C2(VECTOR_ADD[8]), .ZN(n_0_0_130));
   NOR2_X1 i_0_0_202 (.A1(n_0_0_131), .A2(n_0_0_182), .ZN(n_0_64));
   AOI222_X1 i_0_0_203 (.A1(NEW_MATRIX_ADD[9]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[9]), .C1(n_0_0_135), .C2(VECTOR_ADD[9]), .ZN(n_0_0_131));
   OAI21_X1 i_0_0_204 (.A(n_0_0_319), .B1(n_0_0_132), .B2(n_0_0_182), .ZN(n_0_65));
   AOI222_X1 i_0_0_205 (.A1(NEW_MATRIX_ADD[10]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[10]), .C1(n_0_0_135), .C2(VECTOR_ADD[10]), .ZN(n_0_0_132));
   OAI21_X1 i_0_0_206 (.A(n_0_0_323), .B1(n_0_0_133), .B2(n_0_0_182), .ZN(n_0_66));
   AOI222_X1 i_0_0_207 (.A1(NEW_MATRIX_ADD[11]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[11]), .C1(n_0_0_135), .C2(VECTOR_ADD[11]), .ZN(n_0_0_133));
   OAI21_X1 i_0_0_208 (.A(n_0_0_319), .B1(n_0_0_134), .B2(n_0_0_182), .ZN(n_0_67));
   AOI222_X1 i_0_0_209 (.A1(NEW_MATRIX_ADD[12]), .A2(n_0_0_329), .B1(n_0_0_325), 
      .B2(VECTOR2_ADD[12]), .C1(n_0_0_135), .C2(VECTOR_ADD[12]), .ZN(n_0_0_134));
   NOR2_X1 i_0_0_210 (.A1(n_0_0_327), .A2(n_0_0_326), .ZN(n_0_0_135));
   OR2_X1 i_0_0_211 (.A1(n_0_0_197), .A2(NEW_MATRIX_ADD[0]), .ZN(n_0_68));
   INV_X1 i_0_0_212 (.A(n_0_0_136), .ZN(n_0_69));
   AOI21_X1 i_0_0_213 (.A(n_0_0_238), .B1(n_0_0_319), .B2(NEW_MATRIX_ADD[1]), 
      .ZN(n_0_0_136));
   INV_X1 i_0_0_214 (.A(n_0_0_137), .ZN(n_0_70));
   AOI21_X1 i_0_0_215 (.A(n_0_0_199), .B1(n_0_0_323), .B2(NEW_MATRIX_ADD[2]), 
      .ZN(n_0_0_137));
   INV_X1 i_0_0_216 (.A(n_0_0_138), .ZN(n_0_71));
   AOI21_X1 i_0_0_217 (.A(n_0_0_318), .B1(n_0_0_317), .B2(NEW_MATRIX_ADD[3]), 
      .ZN(n_0_0_138));
   AND2_X1 i_0_0_218 (.A1(NEW_MATRIX_ADD[4]), .A2(n_0_0_315), .ZN(n_0_72));
   OAI21_X1 i_0_0_219 (.A(n_0_0_319), .B1(n_0_0_238), .B2(n_0_0_448), .ZN(n_0_73));
   INV_X1 i_0_0_220 (.A(n_0_0_139), .ZN(n_0_74));
   AOI21_X1 i_0_0_221 (.A(n_0_0_318), .B1(n_0_0_317), .B2(NEW_MATRIX_ADD[6]), 
      .ZN(n_0_0_139));
   INV_X1 i_0_0_222 (.A(n_0_0_140), .ZN(n_0_75));
   AOI21_X1 i_0_0_223 (.A(n_0_0_318), .B1(n_0_0_317), .B2(NEW_MATRIX_ADD[7]), 
      .ZN(n_0_0_140));
   OAI21_X1 i_0_0_224 (.A(n_0_0_323), .B1(n_0_0_199), .B2(n_0_0_449), .ZN(n_0_76));
   AND2_X1 i_0_0_114 (.A1(NEW_MATRIX_ADD[9]), .A2(n_0_0_315), .ZN(n_0_77));
   OAI21_X1 i_0_0_115 (.A(n_0_0_319), .B1(n_0_0_238), .B2(n_0_0_450), .ZN(n_0_78));
   OAI21_X1 i_0_0_116 (.A(n_0_0_323), .B1(n_0_0_199), .B2(n_0_0_451), .ZN(n_0_79));
   OAI21_X1 i_0_0_228 (.A(n_0_0_319), .B1(n_0_0_238), .B2(n_0_0_452), .ZN(n_0_80));
   AND2_X1 i_0_0_229 (.A1(MATRIX_ADD[13]), .A2(n_0_0_315), .ZN(n_0_81));
   AND2_X1 i_0_0_230 (.A1(MATRIX_ADD[14]), .A2(n_0_0_315), .ZN(n_0_82));
   AND2_X1 i_0_0_231 (.A1(MATRIX_ADD[15]), .A2(n_0_0_315), .ZN(n_0_83));
   OR2_X1 i_0_0_117 (.A1(NEW_VECTOR2_ADD[0]), .A2(n_0_0_493), .ZN(n_0_84));
   OR2_X1 i_0_0_233 (.A1(NEW_VECTOR2_ADD[1]), .A2(n_0_0_493), .ZN(n_0_85));
   OR2_X1 i_0_0_234 (.A1(NEW_VECTOR2_ADD[2]), .A2(n_0_0_493), .ZN(n_0_86));
   AND2_X1 i_0_0_235 (.A1(n_0_0_319), .A2(NEW_VECTOR2_ADD[3]), .ZN(n_0_87));
   OR2_X1 i_0_0_236 (.A1(NEW_VECTOR2_ADD[4]), .A2(n_0_0_493), .ZN(n_0_88));
   AND2_X1 i_0_0_237 (.A1(n_0_0_319), .A2(NEW_VECTOR2_ADD[5]), .ZN(n_0_89));
   OR2_X1 i_0_0_238 (.A1(NEW_VECTOR2_ADD[6]), .A2(n_0_0_493), .ZN(n_0_90));
   AND2_X1 i_0_0_239 (.A1(n_0_0_319), .A2(NEW_VECTOR2_ADD[7]), .ZN(n_0_91));
   AND2_X1 i_0_0_240 (.A1(n_0_0_319), .A2(NEW_VECTOR2_ADD[8]), .ZN(n_0_92));
   AND2_X1 i_0_0_241 (.A1(n_0_0_319), .A2(NEW_VECTOR2_ADD[9]), .ZN(n_0_93));
   OR2_X1 i_0_0_242 (.A1(NEW_VECTOR2_ADD[10]), .A2(n_0_0_493), .ZN(n_0_94));
   AND2_X1 i_0_0_243 (.A1(n_0_0_319), .A2(NEW_VECTOR2_ADD[11]), .ZN(n_0_95));
   OR2_X1 i_0_0_244 (.A1(NEW_VECTOR2_ADD[12]), .A2(n_0_0_493), .ZN(n_0_96));
   AND2_X1 i_0_0_245 (.A1(n_0_0_319), .A2(VECTOR2_ADD[13]), .ZN(n_0_97));
   AND2_X1 i_0_0_246 (.A1(n_0_0_319), .A2(VECTOR2_ADD[14]), .ZN(n_0_98));
   AND2_X1 i_0_0_247 (.A1(n_0_0_319), .A2(VECTOR2_ADD[15]), .ZN(n_0_99));
   NAND2_X1 i_0_0_248 (.A1(n_0_0_232), .A2(n_0_0_319), .ZN(n_0_100));
   OAI21_X1 i_0_0_249 (.A(n_0_0_146), .B1(n_0_0_147), .B2(n_0_0_453), .ZN(
      n_0_101));
   INV_X1 i_0_0_250 (.A(n_0_0_141), .ZN(n_0_102));
   AOI21_X1 i_0_0_251 (.A(n_0_0_144), .B1(n_0_0_148), .B2(NEW_VECTOR_ADD[1]), 
      .ZN(n_0_0_141));
   OAI21_X1 i_0_0_252 (.A(n_0_0_179), .B1(n_0_0_147), .B2(n_0_0_454), .ZN(
      n_0_103));
   INV_X1 i_0_0_253 (.A(n_0_0_142), .ZN(n_0_104));
   AOI21_X1 i_0_0_254 (.A(n_0_0_175), .B1(n_0_0_148), .B2(NEW_VECTOR_ADD[3]), 
      .ZN(n_0_0_142));
   INV_X1 i_0_0_255 (.A(n_0_0_143), .ZN(n_0_105));
   AOI21_X1 i_0_0_256 (.A(n_0_0_144), .B1(n_0_0_148), .B2(NEW_VECTOR_ADD[4]), 
      .ZN(n_0_0_143));
   NAND2_X1 i_0_0_257 (.A1(n_0_0_179), .A2(n_0_0_319), .ZN(n_0_0_144));
   OAI21_X1 i_0_0_258 (.A(n_0_0_319), .B1(n_0_0_147), .B2(n_0_0_455), .ZN(
      n_0_106));
   OAI21_X1 i_0_0_259 (.A(n_0_0_179), .B1(n_0_0_147), .B2(n_0_0_456), .ZN(
      n_0_107));
   INV_X1 i_0_0_260 (.A(n_0_0_145), .ZN(n_0_108));
   AOI21_X1 i_0_0_261 (.A(n_0_0_175), .B1(n_0_0_148), .B2(NEW_VECTOR_ADD[7]), 
      .ZN(n_0_0_145));
   AND2_X1 i_0_0_262 (.A1(NEW_VECTOR_ADD[8]), .A2(n_0_0_148), .ZN(n_0_109));
   AND2_X1 i_0_0_263 (.A1(NEW_VECTOR_ADD[9]), .A2(n_0_0_148), .ZN(n_0_110));
   OAI21_X1 i_0_0_264 (.A(n_0_0_146), .B1(n_0_0_147), .B2(n_0_0_457), .ZN(
      n_0_111));
   AND2_X1 i_0_0_265 (.A1(NEW_VECTOR_ADD[11]), .A2(n_0_0_148), .ZN(n_0_112));
   OAI21_X1 i_0_0_266 (.A(n_0_0_146), .B1(n_0_0_147), .B2(n_0_0_458), .ZN(
      n_0_113));
   NOR2_X1 i_0_0_267 (.A1(n_0_0_178), .A2(n_0_0_175), .ZN(n_0_0_146));
   AND2_X1 i_0_0_268 (.A1(VECTOR_ADD[13]), .A2(n_0_0_148), .ZN(n_0_114));
   AND2_X1 i_0_0_269 (.A1(VECTOR_ADD[14]), .A2(n_0_0_148), .ZN(n_0_115));
   AND2_X1 i_0_0_270 (.A1(VECTOR_ADD[15]), .A2(n_0_0_148), .ZN(n_0_116));
   OAI21_X1 i_0_0_118 (.A(n_0_0_315), .B1(n_0_0_172), .B2(n_0_0_328), .ZN(
      n_0_0_147));
   NOR2_X1 i_0_0_272 (.A1(n_0_0_149), .A2(n_0_0_197), .ZN(n_0_0_148));
   NOR2_X1 i_0_0_119 (.A1(n_0_0_328), .A2(n_0_0_172), .ZN(n_0_0_149));
   OAI21_X1 i_0_0_120 (.A(n_0_0_183), .B1(n_0_0_153), .B2(CLK), .ZN(n_0_118));
   AOI21_X1 i_0_0_121 (.A(n_0_0_155), .B1(n_0_0_154), .B2(next[2]), .ZN(
      n_0_0_153));
   OAI21_X1 i_0_0_124 (.A(next[1]), .B1(next[0]), .B2(counter[1]), .ZN(n_0_0_154));
   AND3_X1 i_0_0_125 (.A1(n_0_0_345), .A2(next[1]), .A3(next[0]), .ZN(n_0_0_155));
   NAND3_X1 i_0_0_126 (.A1(n_0_0_156), .A2(n_0_0_184), .A3(n_0_0_173), .ZN(
      n_0_119));
   AOI22_X1 i_0_0_127 (.A1(NEW_VECTOR_ADD[0]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[0]), .ZN(n_0_0_156));
   NAND2_X1 i_0_0_128 (.A1(n_0_0_157), .A2(n_0_0_177), .ZN(n_0_120));
   AOI22_X1 i_0_0_129 (.A1(NEW_VECTOR_ADD[1]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[1]), .ZN(n_0_0_157));
   NAND2_X1 i_0_0_130 (.A1(n_0_0_163), .A2(n_0_0_158), .ZN(n_0_121));
   AOI22_X1 i_0_0_131 (.A1(NEW_VECTOR_ADD[2]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[2]), .ZN(n_0_0_158));
   NAND2_X1 i_0_0_153 (.A1(n_0_0_174), .A2(n_0_0_159), .ZN(n_0_122));
   AOI22_X1 i_0_0_154 (.A1(NEW_VECTOR_ADD[3]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[3]), .ZN(n_0_0_159));
   NAND2_X1 i_0_0_290 (.A1(n_0_0_160), .A2(n_0_0_177), .ZN(n_0_123));
   AOI22_X1 i_0_0_291 (.A1(NEW_VECTOR_ADD[4]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[4]), .ZN(n_0_0_160));
   NAND2_X1 i_0_0_155 (.A1(n_0_0_161), .A2(n_0_0_319), .ZN(n_0_124));
   AOI22_X1 i_0_0_156 (.A1(NEW_VECTOR_ADD[5]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[5]), .ZN(n_0_0_161));
   NAND2_X1 i_0_0_294 (.A1(n_0_0_163), .A2(n_0_0_162), .ZN(n_0_125));
   AOI22_X1 i_0_0_295 (.A1(NEW_VECTOR_ADD[6]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[6]), .ZN(n_0_0_162));
   AOI21_X1 i_0_0_157 (.A(n_0_0_493), .B1(n_0_0_184), .B2(n_0_0_178), .ZN(
      n_0_0_163));
   NAND2_X1 i_0_0_297 (.A1(n_0_0_174), .A2(n_0_0_164), .ZN(n_0_126));
   AOI22_X1 i_0_0_298 (.A1(NEW_VECTOR_ADD[7]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[7]), .ZN(n_0_0_164));
   INV_X1 i_0_0_158 (.A(n_0_0_165), .ZN(n_0_127));
   AOI22_X1 i_0_0_159 (.A1(NEW_VECTOR_ADD[8]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[8]), .ZN(n_0_0_165));
   INV_X1 i_0_0_301 (.A(n_0_0_166), .ZN(n_0_128));
   AOI22_X1 i_0_0_302 (.A1(NEW_VECTOR_ADD[9]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[9]), .ZN(n_0_0_166));
   NAND2_X1 i_0_0_160 (.A1(n_0_0_173), .A2(n_0_0_167), .ZN(n_0_129));
   AOI22_X1 i_0_0_161 (.A1(NEW_VECTOR_ADD[10]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[10]), .ZN(n_0_0_167));
   INV_X1 i_0_0_305 (.A(n_0_0_168), .ZN(n_0_130));
   AOI22_X1 i_0_0_306 (.A1(NEW_VECTOR_ADD[11]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[11]), .ZN(n_0_0_168));
   NAND2_X1 i_0_0_307 (.A1(n_0_0_173), .A2(n_0_0_169), .ZN(n_0_131));
   AOI22_X1 i_0_0_308 (.A1(NEW_VECTOR_ADD[12]), .A2(n_0_0_171), .B1(n_0_0_170), 
      .B2(MATRIX_ADD[12]), .ZN(n_0_0_169));
   NOR2_X1 i_0_0_162 (.A1(n_0_0_327), .A2(n_0_0_182), .ZN(n_0_0_170));
   NOR3_X1 i_0_0_163 (.A1(n_0_0_397), .A2(n_0_0_266), .A3(n_0_0_182), .ZN(
      n_0_0_171));
   NOR2_X1 i_0_0_164 (.A1(n_0_0_397), .A2(n_0_0_266), .ZN(n_0_0_172));
   OAI21_X1 i_0_0_165 (.A(n_0_0_184), .B1(n_0_0_178), .B2(n_0_0_175), .ZN(
      n_0_0_173));
   NAND2_X1 i_0_0_166 (.A1(n_0_0_184), .A2(n_0_0_175), .ZN(n_0_0_174));
   NAND2_X1 i_0_0_167 (.A1(n_0_0_176), .A2(n_0_0_347), .ZN(n_0_0_175));
   NAND3_X1 i_0_0_168 (.A1(n_0_0_329), .A2(n_0_0_267), .A3(n_0_0_317), .ZN(
      n_0_0_176));
   NAND2_X1 i_0_0_169 (.A1(n_0_0_184), .A2(n_0_0_178), .ZN(n_0_0_177));
   INV_X1 i_0_0_170 (.A(n_0_0_179), .ZN(n_0_0_178));
   AOI21_X1 i_0_0_171 (.A(n_0_0_316), .B1(n_0_0_346), .B2(n_0_0_320), .ZN(
      n_0_0_179));
   NAND2_X1 i_0_0_172 (.A1(n_0_0_394), .A2(n_0_0_183), .ZN(n_0_132));
   NAND2_X1 i_0_0_173 (.A1(n_0_0_315), .A2(n_0_0_184), .ZN(n_0_0_182));
   NOR2_X1 i_0_0_174 (.A1(n_0_0_197), .A2(n_0_0_185), .ZN(n_0_0_183));
   INV_X1 i_0_0_175 (.A(n_0_0_185), .ZN(n_0_0_184));
   NOR3_X1 i_0_0_176 (.A1(n_0_52), .A2(n_0_0_186), .A3(n_0_1), .ZN(n_0_0_185));
   NAND2_X1 i_0_0_177 (.A1(INT), .A2(PROCESS), .ZN(n_0_0_186));
   NAND2_X1 i_0_0_178 (.A1(n_0_0_394), .A2(n_0_0_315), .ZN(n_0_133));
   OR2_X1 i_0_0_179 (.A1(n_0_0_197), .A2(RESULT_ADD[0]), .ZN(n_0_134));
   INV_X1 i_0_0_180 (.A(n_0_0_187), .ZN(n_0_135));
   AOI21_X1 i_0_0_181 (.A(n_0_0_318), .B1(n_0_0_317), .B2(RESULT_ADD[1]), 
      .ZN(n_0_0_187));
   INV_X1 i_0_0_225 (.A(n_0_0_188), .ZN(n_0_136));
   AOI21_X1 i_0_0_226 (.A(n_0_0_199), .B1(n_0_0_323), .B2(RESULT_ADD[2]), 
      .ZN(n_0_0_188));
   OR2_X1 i_0_0_333 (.A1(n_0_0_197), .A2(RESULT_ADD[3]), .ZN(n_0_137));
   INV_X1 i_0_0_334 (.A(n_0_0_189), .ZN(n_0_138));
   AOI21_X1 i_0_0_335 (.A(n_0_0_318), .B1(n_0_0_317), .B2(RESULT_ADD[4]), 
      .ZN(n_0_0_189));
   INV_X1 i_0_0_336 (.A(n_0_0_190), .ZN(n_0_139));
   AOI21_X1 i_0_0_337 (.A(n_0_0_238), .B1(n_0_0_319), .B2(RESULT_ADD[5]), 
      .ZN(n_0_0_190));
   OAI21_X1 i_0_0_227 (.A(n_0_0_317), .B1(n_0_0_318), .B2(n_0_0_459), .ZN(
      n_0_140));
   INV_X1 i_0_0_339 (.A(n_0_0_191), .ZN(n_0_141));
   AOI21_X1 i_0_0_340 (.A(n_0_0_238), .B1(n_0_0_319), .B2(RESULT_ADD[7]), 
      .ZN(n_0_0_191));
   OAI21_X1 i_0_0_232 (.A(n_0_0_319), .B1(n_0_0_238), .B2(n_0_0_460), .ZN(
      n_0_142));
   AND2_X1 i_0_0_342 (.A1(RESULT_ADD[9]), .A2(n_0_0_315), .ZN(n_0_143));
   OR2_X1 i_0_0_343 (.A1(n_0_0_197), .A2(RESULT_ADD[10]), .ZN(n_0_144));
   AND2_X1 i_0_0_344 (.A1(RESULT_ADD[11]), .A2(n_0_0_315), .ZN(n_0_145));
   OR2_X1 i_0_0_345 (.A1(n_0_0_197), .A2(RESULT_ADD[12]), .ZN(n_0_146));
   OR2_X1 i_0_0_346 (.A1(n_0_0_197), .A2(NEW_RESULT_ADD[0]), .ZN(n_0_147));
   INV_X1 i_0_0_347 (.A(n_0_0_192), .ZN(n_0_148));
   AOI21_X1 i_0_0_348 (.A(n_0_0_318), .B1(n_0_0_317), .B2(NEW_RESULT_ADD[1]), 
      .ZN(n_0_0_192));
   INV_X1 i_0_0_349 (.A(n_0_0_193), .ZN(n_0_149));
   AOI21_X1 i_0_0_350 (.A(n_0_0_199), .B1(n_0_0_323), .B2(NEW_RESULT_ADD[2]), 
      .ZN(n_0_0_193));
   OR2_X1 i_0_0_351 (.A1(n_0_0_197), .A2(NEW_RESULT_ADD[3]), .ZN(n_0_150));
   INV_X1 i_0_0_352 (.A(n_0_0_194), .ZN(n_0_151));
   AOI21_X1 i_0_0_353 (.A(n_0_0_318), .B1(n_0_0_317), .B2(NEW_RESULT_ADD[4]), 
      .ZN(n_0_0_194));
   INV_X1 i_0_0_354 (.A(n_0_0_195), .ZN(n_0_152));
   AOI21_X1 i_0_0_355 (.A(n_0_0_238), .B1(n_0_0_319), .B2(NEW_RESULT_ADD[5]), 
      .ZN(n_0_0_195));
   OAI21_X1 i_0_0_356 (.A(n_0_0_317), .B1(n_0_0_318), .B2(n_0_0_461), .ZN(
      n_0_153));
   INV_X1 i_0_0_357 (.A(n_0_0_196), .ZN(n_0_154));
   AOI21_X1 i_0_0_358 (.A(n_0_0_238), .B1(n_0_0_319), .B2(NEW_RESULT_ADD[7]), 
      .ZN(n_0_0_196));
   OAI21_X1 i_0_0_359 (.A(n_0_0_319), .B1(n_0_0_238), .B2(n_0_0_462), .ZN(
      n_0_155));
   AND2_X1 i_0_0_360 (.A1(NEW_RESULT_ADD[9]), .A2(n_0_0_315), .ZN(n_0_156));
   OR2_X1 i_0_0_361 (.A1(n_0_0_197), .A2(NEW_RESULT_ADD[10]), .ZN(n_0_157));
   AND2_X1 i_0_0_362 (.A1(NEW_RESULT_ADD[11]), .A2(n_0_0_315), .ZN(n_0_158));
   OR2_X1 i_0_0_363 (.A1(n_0_0_197), .A2(NEW_RESULT_ADD[12]), .ZN(n_0_159));
   AND2_X1 i_0_0_364 (.A1(RESULT_ADD[13]), .A2(n_0_0_315), .ZN(n_0_160));
   AND2_X1 i_0_0_365 (.A1(RESULT_ADD[14]), .A2(n_0_0_315), .ZN(n_0_161));
   AND2_X1 i_0_0_366 (.A1(RESULT_ADD[15]), .A2(n_0_0_315), .ZN(n_0_162));
   OAI21_X1 i_0_0_271 (.A(n_0_0_315), .B1(n_0_0_264), .B2(CLK), .ZN(n_0_163));
   OAI21_X1 i_0_0_273 (.A(n_0_0_315), .B1(n_0_0_265), .B2(CLK), .ZN(n_0_46));
   NAND2_X1 i_0_0_274 (.A1(n_0_0_347), .A2(n_0_0_317), .ZN(n_0_0_197));
   NAND2_X1 i_0_0_275 (.A1(n_0_0_317), .A2(n_0_0_319), .ZN(n_0_0_199));
   INV_X1 i_0_0_276 (.A(n_0_0_205), .ZN(n_0_164));
   AOI22_X1 i_0_0_277 (.A1(RAM_DATA_RD1[0]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[0]), .ZN(n_0_0_205));
   INV_X1 i_0_0_379 (.A(n_0_0_206), .ZN(n_0_165));
   AOI22_X1 i_0_0_380 (.A1(RAM_DATA_RD1[1]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[1]), .ZN(n_0_0_206));
   INV_X1 i_0_0_381 (.A(n_0_0_207), .ZN(n_0_166));
   AOI22_X1 i_0_0_382 (.A1(RAM_DATA_RD1[2]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[2]), .ZN(n_0_0_207));
   INV_X1 i_0_0_383 (.A(n_0_0_208), .ZN(n_0_167));
   AOI22_X1 i_0_0_384 (.A1(RAM_DATA_RD1[3]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[3]), .ZN(n_0_0_208));
   INV_X1 i_0_0_385 (.A(n_0_0_209), .ZN(n_0_168));
   AOI22_X1 i_0_0_386 (.A1(RAM_DATA_RD1[4]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[4]), .ZN(n_0_0_209));
   INV_X1 i_0_0_387 (.A(n_0_0_210), .ZN(n_0_169));
   AOI22_X1 i_0_0_388 (.A1(RAM_DATA_RD1[5]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[5]), .ZN(n_0_0_210));
   INV_X1 i_0_0_389 (.A(n_0_0_211), .ZN(n_0_170));
   AOI22_X1 i_0_0_390 (.A1(RAM_DATA_RD1[6]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[6]), .ZN(n_0_0_211));
   INV_X1 i_0_0_391 (.A(n_0_0_212), .ZN(n_0_171));
   AOI22_X1 i_0_0_392 (.A1(RAM_DATA_RD1[7]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[7]), .ZN(n_0_0_212));
   INV_X1 i_0_0_393 (.A(n_0_0_213), .ZN(n_0_172));
   AOI22_X1 i_0_0_394 (.A1(RAM_DATA_RD1[8]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[8]), .ZN(n_0_0_213));
   INV_X1 i_0_0_395 (.A(n_0_0_214), .ZN(n_0_173));
   AOI22_X1 i_0_0_396 (.A1(RAM_DATA_RD1[9]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[9]), .ZN(n_0_0_214));
   INV_X1 i_0_0_397 (.A(n_0_0_215), .ZN(n_0_174));
   AOI22_X1 i_0_0_398 (.A1(RAM_DATA_RD1[10]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[10]), .ZN(n_0_0_215));
   INV_X1 i_0_0_399 (.A(n_0_0_216), .ZN(n_0_175));
   AOI22_X1 i_0_0_400 (.A1(RAM_DATA_RD1[11]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[11]), .ZN(n_0_0_216));
   INV_X1 i_0_0_401 (.A(n_0_0_217), .ZN(n_0_176));
   AOI22_X1 i_0_0_402 (.A1(RAM_DATA_RD1[12]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[12]), .ZN(n_0_0_217));
   INV_X1 i_0_0_403 (.A(n_0_0_218), .ZN(n_0_177));
   AOI22_X1 i_0_0_404 (.A1(RAM_DATA_RD1[13]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[13]), .ZN(n_0_0_218));
   INV_X1 i_0_0_405 (.A(n_0_0_219), .ZN(n_0_178));
   AOI22_X1 i_0_0_406 (.A1(RAM_DATA_RD1[14]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[14]), .ZN(n_0_0_219));
   INV_X1 i_0_0_407 (.A(n_0_0_220), .ZN(n_0_179));
   AOI22_X1 i_0_0_408 (.A1(RAM_DATA_RD1[15]), .A2(n_0_0_222), .B1(n_0_0_221), 
      .B2(NEW_Element_Result[15]), .ZN(n_0_0_220));
   NOR3_X1 i_0_0_278 (.A1(n_0_0_328), .A2(n_0_0_224), .A3(n_0_0_238), .ZN(
      n_0_0_221));
   NOR3_X1 i_0_0_279 (.A1(n_0_0_224), .A2(n_0_0_238), .A3(n_0_0_327), .ZN(
      n_0_0_222));
   OAI21_X1 i_0_0_411 (.A(n_0_0_223), .B1(n_0_0_246), .B2(n_0_0_394), .ZN(
      n_0_180));
   NOR2_X1 i_0_0_412 (.A1(n_0_0_224), .A2(n_0_0_238), .ZN(n_0_0_223));
   AOI211_X1 i_0_0_280 (.A(n_0_0_225), .B(n_0_0_233), .C1(n_0_0_237), .C2(
      n_0_0_231), .ZN(n_0_0_224));
   OAI221_X1 i_0_0_281 (.A(n_0_0_324), .B1(n_0_47), .B2(n_0_0_226), .C1(
      VECTOR_CNT_adder_n_2), .C2(n_0_0_396), .ZN(n_0_0_225));
   NOR3_X1 i_0_0_282 (.A1(n_0_0_227), .A2(VECTOR_CNT[8]), .A3(VECTOR_CNT[9]), 
      .ZN(n_0_0_226));
   NAND3_X1 i_0_0_283 (.A1(n_0_0_230), .A2(n_0_0_229), .A3(n_0_0_228), .ZN(
      n_0_0_227));
   NOR3_X1 i_0_0_284 (.A1(VECTOR_CNT[5]), .A2(VECTOR_CNT[4]), .A3(VECTOR_CNT[1]), 
      .ZN(n_0_0_228));
   NOR4_X1 i_0_0_285 (.A1(VECTOR_CNT[12]), .A2(VECTOR_CNT[11]), .A3(
      VECTOR_CNT[10]), .A4(VECTOR_CNT[7]), .ZN(n_0_0_229));
   NOR4_X1 i_0_0_286 (.A1(VECTOR_CNT[6]), .A2(VECTOR_CNT[3]), .A3(VECTOR_CNT[2]), 
      .A4(VECTOR_CNT[0]), .ZN(n_0_0_230));
   INV_X1 i_0_0_287 (.A(n_0_0_232), .ZN(n_0_0_231));
   NAND2_X1 i_0_0_288 (.A1(next[1]), .A2(n_0_47), .ZN(n_0_0_232));
   NOR2_X1 i_0_0_289 (.A1(CLK), .A2(n_0_0_265), .ZN(n_0_47));
   NOR2_X1 i_0_0_292 (.A1(n_0_0_266), .A2(n_0_0_234), .ZN(n_0_0_233));
   OAI21_X1 i_0_0_293 (.A(n_0_0_396), .B1(n_0_0_237), .B2(n_0_0_235), .ZN(
      n_0_0_234));
   INV_X1 i_0_0_296 (.A(VECTOR_CNT_adder_n_2), .ZN(n_0_0_235));
   NAND2_X1 i_0_0_299 (.A1(VECTOR_CNT_adder_tempIn11[12]), .A2(n_0_0_406), 
      .ZN(n_0_0_237));
   NAND2_X1 i_0_0_300 (.A1(n_0_0_317), .A2(n_0_0_323), .ZN(n_0_0_238));
   NOR2_X1 i_0_0_303 (.A1(n_0_0_316), .A2(n_0_0_240), .ZN(n_0_0_239));
   INV_X1 i_0_0_304 (.A(n_0_0_323), .ZN(n_0_0_240));
   NOR2_X1 i_0_0_309 (.A1(state[1]), .A2(state[0]), .ZN(n_0_0_242));
   AOI21_X1 i_0_0_437 (.A(n_0_0_396), .B1(counter[0]), .B2(n_0_0_463), .ZN(
      n_0_0_246));
   NOR2_X1 i_0_0_310 (.A1(n_0_0_247), .A2(state[2]), .ZN(n_0_181));
   NAND2_X1 i_0_0_311 (.A1(state[1]), .A2(state[0]), .ZN(n_0_0_247));
   INV_X1 i_0_0_312 (.A(n_0_0_248), .ZN(n_0_182));
   AOI22_X1 i_0_0_313 (.A1(NEW_Element_Result[0]), .A2(n_0_0_329), .B1(n_0_0_328), 
      .B2(FINAL_RESULT[0]), .ZN(n_0_0_248));
   INV_X1 i_0_0_442 (.A(n_0_0_249), .ZN(n_0_183));
   AOI22_X1 i_0_0_443 (.A1(NEW_Element_Result[1]), .A2(n_0_0_329), .B1(n_0_0_328), 
      .B2(FINAL_RESULT[1]), .ZN(n_0_0_249));
   INV_X1 i_0_0_444 (.A(n_0_0_250), .ZN(n_0_184));
   AOI22_X1 i_0_0_445 (.A1(NEW_Element_Result[2]), .A2(n_0_0_329), .B1(n_0_0_328), 
      .B2(FINAL_RESULT[2]), .ZN(n_0_0_250));
   INV_X1 i_0_0_446 (.A(n_0_0_251), .ZN(n_0_185));
   AOI22_X1 i_0_0_447 (.A1(NEW_Element_Result[3]), .A2(n_0_0_329), .B1(n_0_0_328), 
      .B2(FINAL_RESULT[3]), .ZN(n_0_0_251));
   INV_X1 i_0_0_448 (.A(n_0_0_252), .ZN(n_0_186));
   AOI22_X1 i_0_0_449 (.A1(NEW_Element_Result[4]), .A2(n_0_0_329), .B1(n_0_0_328), 
      .B2(FINAL_RESULT[4]), .ZN(n_0_0_252));
   INV_X1 i_0_0_450 (.A(n_0_0_253), .ZN(n_0_187));
   AOI22_X1 i_0_0_451 (.A1(NEW_Element_Result[5]), .A2(n_0_0_329), .B1(n_0_0_328), 
      .B2(FINAL_RESULT[5]), .ZN(n_0_0_253));
   INV_X1 i_0_0_452 (.A(n_0_0_254), .ZN(n_0_188));
   AOI22_X1 i_0_0_453 (.A1(NEW_Element_Result[6]), .A2(n_0_0_329), .B1(n_0_0_328), 
      .B2(FINAL_RESULT[6]), .ZN(n_0_0_254));
   INV_X1 i_0_0_454 (.A(n_0_0_255), .ZN(n_0_189));
   AOI22_X1 i_0_0_455 (.A1(NEW_Element_Result[7]), .A2(n_0_0_329), .B1(n_0_0_328), 
      .B2(FINAL_RESULT[7]), .ZN(n_0_0_255));
   INV_X1 i_0_0_456 (.A(n_0_0_256), .ZN(n_0_190));
   AOI22_X1 i_0_0_457 (.A1(NEW_Element_Result[8]), .A2(n_0_0_329), .B1(n_0_0_328), 
      .B2(FINAL_RESULT[8]), .ZN(n_0_0_256));
   INV_X1 i_0_0_458 (.A(n_0_0_257), .ZN(n_0_191));
   AOI22_X1 i_0_0_459 (.A1(NEW_Element_Result[9]), .A2(n_0_0_329), .B1(n_0_0_328), 
      .B2(FINAL_RESULT[9]), .ZN(n_0_0_257));
   INV_X1 i_0_0_460 (.A(n_0_0_258), .ZN(n_0_192));
   AOI22_X1 i_0_0_461 (.A1(NEW_Element_Result[10]), .A2(n_0_0_329), .B1(
      n_0_0_328), .B2(FINAL_RESULT[10]), .ZN(n_0_0_258));
   INV_X1 i_0_0_462 (.A(n_0_0_259), .ZN(n_0_193));
   AOI22_X1 i_0_0_463 (.A1(NEW_Element_Result[11]), .A2(n_0_0_329), .B1(
      n_0_0_328), .B2(FINAL_RESULT[11]), .ZN(n_0_0_259));
   INV_X1 i_0_0_464 (.A(n_0_0_260), .ZN(n_0_194));
   AOI22_X1 i_0_0_465 (.A1(NEW_Element_Result[12]), .A2(n_0_0_329), .B1(
      n_0_0_328), .B2(FINAL_RESULT[12]), .ZN(n_0_0_260));
   INV_X1 i_0_0_466 (.A(n_0_0_261), .ZN(n_0_195));
   AOI22_X1 i_0_0_467 (.A1(NEW_Element_Result[13]), .A2(n_0_0_329), .B1(
      n_0_0_328), .B2(FINAL_RESULT[13]), .ZN(n_0_0_261));
   INV_X1 i_0_0_468 (.A(n_0_0_262), .ZN(n_0_196));
   AOI22_X1 i_0_0_469 (.A1(NEW_Element_Result[14]), .A2(n_0_0_329), .B1(
      n_0_0_328), .B2(FINAL_RESULT[14]), .ZN(n_0_0_262));
   INV_X1 i_0_0_470 (.A(n_0_0_263), .ZN(n_0_197));
   AOI22_X1 i_0_0_471 (.A1(NEW_Element_Result[15]), .A2(n_0_0_329), .B1(
      n_0_0_328), .B2(FINAL_RESULT[15]), .ZN(n_0_0_263));
   NOR2_X1 i_0_0_472 (.A1(n_0_0_264), .A2(n_0_0_399), .ZN(n_0_198));
   AOI21_X1 i_0_0_314 (.A(n_0_0_393), .B1(n_0_0_266), .B2(n_0_0_329), .ZN(
      n_0_0_264));
   NOR2_X1 i_0_0_315 (.A1(n_0_0_329), .A2(n_0_0_393), .ZN(n_0_0_265));
   OR2_X1 i_0_0_316 (.A1(n_0_0_320), .A2(n_0_0_267), .ZN(n_0_0_266));
   NOR3_X1 i_0_0_317 (.A1(n_0_0_433), .A2(n_0_0_361), .A3(n_0_0_268), .ZN(
      n_0_0_267));
   OAI21_X1 i_0_0_318 (.A(n_0_0_269), .B1(n_0_0_377), .B2(m_val[9]), .ZN(
      n_0_0_268));
   AOI21_X1 i_0_0_319 (.A(n_0_0_270), .B1(n_0_0_377), .B2(m_val[9]), .ZN(
      n_0_0_269));
   OAI21_X1 i_0_0_320 (.A(n_0_0_271), .B1(n_0_0_445), .B2(m_val[7]), .ZN(
      n_0_0_270));
   AOI21_X1 i_0_0_321 (.A(n_0_0_272), .B1(n_0_0_445), .B2(m_val[7]), .ZN(
      n_0_0_271));
   OAI211_X1 i_0_0_322 (.A(n_0_0_348), .B(n_0_0_273), .C1(m_val[6]), .C2(
      n_0_0_369), .ZN(n_0_0_272));
   NOR4_X1 i_0_0_323 (.A1(n_0_0_289), .A2(n_0_0_286), .A3(n_0_0_279), .A4(
      n_0_0_274), .ZN(n_0_0_273));
   NAND4_X1 i_0_0_324 (.A1(n_0_0_278), .A2(n_0_0_277), .A3(n_0_0_276), .A4(
      n_0_0_275), .ZN(n_0_0_274));
   NOR4_X1 i_0_0_325 (.A1(m_val[49]), .A2(m_val[48]), .A3(m_val[47]), .A4(
      m_val[46]), .ZN(n_0_0_275));
   NOR4_X1 i_0_0_326 (.A1(m_val[45]), .A2(m_val[44]), .A3(m_val[43]), .A4(
      m_val[42]), .ZN(n_0_0_276));
   NOR4_X1 i_0_0_327 (.A1(m_val[57]), .A2(m_val[56]), .A3(m_val[55]), .A4(
      m_val[54]), .ZN(n_0_0_277));
   NOR4_X1 i_0_0_328 (.A1(m_val[53]), .A2(m_val[52]), .A3(m_val[51]), .A4(
      m_val[50]), .ZN(n_0_0_278));
   NAND3_X1 i_0_0_329 (.A1(n_0_0_282), .A2(n_0_0_281), .A3(n_0_0_280), .ZN(
      n_0_0_279));
   NOR4_X1 i_0_0_330 (.A1(m_val[33]), .A2(m_val[32]), .A3(m_val[31]), .A4(
      m_val[30]), .ZN(n_0_0_280));
   NOR4_X1 i_0_0_331 (.A1(m_val[29]), .A2(m_val[28]), .A3(m_val[27]), .A4(
      m_val[26]), .ZN(n_0_0_281));
   AND3_X1 i_0_0_332 (.A1(n_0_0_285), .A2(n_0_0_284), .A3(n_0_0_283), .ZN(
      n_0_0_282));
   NOR4_X1 i_0_0_338 (.A1(m_val[41]), .A2(m_val[40]), .A3(m_val[39]), .A4(
      m_val[38]), .ZN(n_0_0_283));
   NOR2_X1 i_0_0_341 (.A1(m_val[35]), .A2(m_val[34]), .ZN(n_0_0_284));
   NOR2_X1 i_0_0_367 (.A1(m_val[37]), .A2(m_val[36]), .ZN(n_0_0_285));
   OAI211_X1 i_0_0_368 (.A(n_0_0_288), .B(n_0_0_287), .C1(VECTOR_CNT[13]), 
      .C2(n_0_0_466), .ZN(n_0_0_286));
   XNOR2_X1 i_0_0_369 (.A(m_val[0]), .B(n_0_0_447), .ZN(n_0_0_287));
   NAND2_X1 i_0_0_370 (.A1(n_0_0_359), .A2(n_0_0_491), .ZN(n_0_0_288));
   NAND4_X1 i_0_0_371 (.A1(n_0_0_293), .A2(n_0_0_292), .A3(n_0_0_291), .A4(
      n_0_0_290), .ZN(n_0_0_289));
   AOI211_X1 i_0_0_372 (.A(m_val[63]), .B(m_val[62]), .C1(n_0_0_466), .C2(
      VECTOR_CNT[13]), .ZN(n_0_0_290));
   NOR4_X1 i_0_0_373 (.A1(m_val[61]), .A2(m_val[60]), .A3(m_val[59]), .A4(
      m_val[58]), .ZN(n_0_0_291));
   AOI22_X1 i_0_0_374 (.A1(n_0_0_29), .A2(m_val[15]), .B1(n_0_0_13), .B2(
      m_val[14]), .ZN(n_0_0_292));
   AOI22_X1 i_0_0_375 (.A1(VECTOR_CNT[15]), .A2(n_0_0_468), .B1(n_0_0_467), 
      .B2(VECTOR_CNT[14]), .ZN(n_0_0_293));
   AND2_X1 i_0_0_376 (.A1(n_0_0_321), .A2(n_0_0_379), .ZN(n_0_0_320));
   AOI211_X1 i_0_0_377 (.A(n_0_0_330), .B(n_0_0_437), .C1(n_val[9]), .C2(
      n_0_0_377), .ZN(n_0_0_321));
   OAI21_X1 i_0_0_378 (.A(n_0_0_331), .B1(n_0_0_377), .B2(n_val[9]), .ZN(
      n_0_0_330));
   AOI211_X1 i_0_0_409 (.A(n_0_0_373), .B(n_0_0_332), .C1(n_val[4]), .C2(
      n_0_0_378), .ZN(n_0_0_331));
   NAND3_X1 i_0_0_410 (.A1(n_0_0_370), .A2(n_0_0_150), .A3(n_0_0_333), .ZN(
      n_0_0_332));
   AOI221_X1 i_0_0_413 (.A(n_0_0_334), .B1(n_0_0_357), .B2(n_val[2]), .C1(
      n_val[5]), .C2(n_0_0_374), .ZN(n_0_0_333));
   NAND4_X1 i_0_0_414 (.A1(n_0_0_337), .A2(next[0]), .A3(n_0_0_341), .A4(
      n_0_0_335), .ZN(n_0_0_334));
   NAND2_X1 i_0_0_415 (.A1(n_0_0_343), .A2(n_0_0_491), .ZN(n_0_0_335));
   OAI21_X1 i_0_0_416 (.A(n_0_0_338), .B1(n_0_0_339), .B2(n_0_0_340), .ZN(
      n_0_0_337));
   NAND3_X1 i_0_0_417 (.A1(n_val[0]), .A2(n_0_0_340), .A3(n_0_0_447), .ZN(
      n_0_0_338));
   NAND2_X1 i_0_0_418 (.A1(n_0_0_305), .A2(VECTOR_CNT_adder_tempIn11[0]), 
      .ZN(n_0_0_339));
   XNOR2_X1 i_0_0_419 (.A(n_val[1]), .B(VECTOR_CNT_adder_tempIn11[1]), .ZN(
      n_0_0_340));
   OR3_X1 i_0_0_420 (.A1(n_val[2]), .A2(n_0_0_343), .A3(n_0_0_360), .ZN(
      n_0_0_341));
   XNOR2_X1 i_0_0_421 (.A(n_0_0_307), .B(VECTOR_CNT_adder_tempIn11[3]), .ZN(
      n_0_0_343));
   XNOR2_X1 i_0_0_422 (.A(n_0_0_474), .B(n_0_0_369), .ZN(n_0_0_370));
   OAI22_X1 i_0_0_423 (.A1(n_0_0_374), .A2(n_val[5]), .B1(n_0_0_378), .B2(
      n_val[4]), .ZN(n_0_0_373));
   OAI21_X1 i_0_0_424 (.A(n_0_0_388), .B1(n_0_0_367), .B2(
      VECTOR_CNT_adder_tempIn11[9]), .ZN(n_0_0_377));
   OAI21_X1 i_0_0_425 (.A(n_0_0_385), .B1(n_0_0_380), .B2(n_0_0_444), .ZN(
      n_0_0_379));
   AOI211_X1 i_0_0_426 (.A(n_val[10]), .B(n_0_0_381), .C1(n_0_0_382), .C2(
      n_0_0_391), .ZN(n_0_0_380));
   NOR3_X1 i_0_0_427 (.A1(n_0_0_311), .A2(n_0_0_392), .A3(
      VECTOR_CNT_adder_tempIn11[11]), .ZN(n_0_0_381));
   INV_X1 i_0_0_428 (.A(n_0_0_442), .ZN(n_0_0_382));
   NAND4_X1 i_0_0_429 (.A1(VECTOR_CNT_adder_tempIn11[11]), .A2(n_0_0_395), 
      .A3(n_0_0_444), .A4(n_0_0_311), .ZN(n_0_0_385));
   INV_X1 i_0_0_430 (.A(n_0_0_390), .ZN(n_0_0_388));
   NOR3_X1 i_0_0_431 (.A1(n_0_0_463), .A2(n_0_0_327), .A3(counter[0]), .ZN(
      n_0_0_393));
   NAND2_X1 i_0_0_432 (.A1(n_0_0_394), .A2(n_0_52), .ZN(n_0_199));
   OAI21_X1 i_0_0_433 (.A(n_0_51), .B1(n_0_0_329), .B2(n_0_0_328), .ZN(n_0_0_394));
   NOR2_X1 i_0_0_434 (.A1(n_0_0_397), .A2(CLK), .ZN(n_0_0_396));
   NAND2_X1 i_0_0_435 (.A1(n_0_0_344), .A2(next[2]), .ZN(n_0_0_397));
   INV_X1 i_0_0_436 (.A(n_0_0_399), .ZN(n_0_52));
   NOR3_X1 i_0_0_438 (.A1(state[2]), .A2(state[1]), .A3(state[0]), .ZN(n_0_0_399));
   NOR2_X1 i_0_0_439 (.A1(state[2]), .A2(state[0]), .ZN(n_0_0_400));
   NOR2_X1 i_0_0_440 (.A1(state[2]), .A2(state[1]), .ZN(n_0_0_401));
   AND2_X1 i_0_0_613 (.A1(MATRIX_CNT[0]), .A2(MATRIX_CNT_adder_n_2), .ZN(
      MATRIX_CNT_adder_n_25));
   INV_X1 i_0_0_441 (.A(n_0_0_402), .ZN(MATRIX_CNT_adder_n_26));
   AOI22_X1 i_0_0_473 (.A1(MATRIX_CNT[1]), .A2(MATRIX_CNT_adder_n_2), .B1(
      n_0_0_470), .B2(MATRIX_CNT[0]), .ZN(n_0_0_402));
   NAND2_X1 i_0_0_474 (.A1(n_0_0_403), .A2(n_0_0_404), .ZN(MATRIX_CNT_adder_n_27));
   AOI22_X1 i_0_0_475 (.A1(MATRIX_CNT[2]), .A2(MATRIX_CNT_adder_n_2), .B1(
      n_0_0_470), .B2(MATRIX_CNT[1]), .ZN(n_0_0_403));
   NAND3_X1 i_0_0_476 (.A1(MATRIX_CNT[15]), .A2(MATRIX_CNT[0]), .A3(n_0_0_469), 
      .ZN(n_0_0_404));
   OAI211_X1 i_0_0_477 (.A(n_0_0_409), .B(n_0_0_408), .C1(MATRIX_CNT[13]), 
      .C2(n_0_0_477), .ZN(MATRIX_CNT_adder_n_29));
   NAND2_X1 i_0_0_478 (.A1(MATRIX_CNT[3]), .A2(n_0_0_470), .ZN(n_0_0_408));
   NAND3_X1 i_0_0_479 (.A1(MATRIX_CNT[15]), .A2(MATRIX_CNT[1]), .A3(n_0_0_465), 
      .ZN(n_0_0_409));
   MUX2_X1 i_0_0_480 (.A(n_0_0_416), .B(n_0_0_478), .S(MATRIX_CNT[13]), .Z(
      MATRIX_CNT_adder_n_31));
   MUX2_X1 i_0_0_481 (.A(n_0_0_416), .B(n_0_0_419), .S(n_0_0_472), .Z(
      MATRIX_CNT_adder_n_19));
   NAND2_X1 i_0_0_482 (.A1(n_0_0_418), .A2(n_0_0_417), .ZN(n_0_0_416));
   AOI22_X1 i_0_0_483 (.A1(MATRIX_CNT[2]), .A2(n_0_0_481), .B1(n_0_0_443), 
      .B2(MATRIX_CNT[0]), .ZN(n_0_0_417));
   AOI22_X1 i_0_0_484 (.A1(n_0_0_489), .A2(MATRIX_CNT[6]), .B1(MATRIX_CNT[4]), 
      .B2(n_0_0_480), .ZN(n_0_0_418));
   MUX2_X1 i_0_0_638 (.A(n_0_0_422), .B(n_0_0_419), .S(MATRIX_CNT[13]), .Z(
      MATRIX_CNT_adder_n_20));
   NAND2_X1 i_0_0_485 (.A1(n_0_0_421), .A2(n_0_0_420), .ZN(n_0_0_419));
   AOI22_X1 i_0_0_486 (.A1(MATRIX_CNT[1]), .A2(n_0_0_443), .B1(n_0_0_480), 
      .B2(MATRIX_CNT[5]), .ZN(n_0_0_420));
   AOI22_X1 i_0_0_487 (.A1(MATRIX_CNT[7]), .A2(n_0_0_489), .B1(n_0_0_481), 
      .B2(MATRIX_CNT[3]), .ZN(n_0_0_421));
   MUX2_X1 i_0_0_642 (.A(n_0_0_422), .B(n_0_0_425), .S(n_0_0_472), .Z(
      MATRIX_CNT_adder_n_21));
   NAND2_X1 i_0_0_643 (.A1(n_0_0_424), .A2(n_0_0_423), .ZN(n_0_0_422));
   AOI22_X1 i_0_0_644 (.A1(MATRIX_CNT[4]), .A2(n_0_0_481), .B1(n_0_0_443), 
      .B2(MATRIX_CNT[2]), .ZN(n_0_0_423));
   AOI22_X1 i_0_0_645 (.A1(n_0_0_489), .A2(MATRIX_CNT[8]), .B1(MATRIX_CNT[6]), 
      .B2(n_0_0_480), .ZN(n_0_0_424));
   MUX2_X1 i_0_0_488 (.A(n_0_0_428), .B(n_0_0_425), .S(MATRIX_CNT[13]), .Z(
      MATRIX_CNT_adder_n_22));
   NAND2_X1 i_0_0_489 (.A1(n_0_0_427), .A2(n_0_0_426), .ZN(n_0_0_425));
   AOI22_X1 i_0_0_490 (.A1(MATRIX_CNT[3]), .A2(n_0_0_443), .B1(n_0_0_480), 
      .B2(MATRIX_CNT[7]), .ZN(n_0_0_426));
   AOI22_X1 i_0_0_491 (.A1(MATRIX_CNT[9]), .A2(n_0_0_489), .B1(n_0_0_481), 
      .B2(MATRIX_CNT[5]), .ZN(n_0_0_427));
   MUX2_X1 i_0_0_492 (.A(n_0_0_435), .B(n_0_0_428), .S(MATRIX_CNT[13]), .Z(
      MATRIX_CNT_adder_n_23));
   NAND2_X1 i_0_0_493 (.A1(n_0_0_430), .A2(n_0_0_429), .ZN(n_0_0_428));
   AOI22_X1 i_0_0_494 (.A1(MATRIX_CNT[6]), .A2(n_0_0_481), .B1(n_0_0_480), 
      .B2(MATRIX_CNT[8]), .ZN(n_0_0_429));
   AOI22_X1 i_0_0_495 (.A1(n_0_0_489), .A2(MATRIX_CNT[10]), .B1(MATRIX_CNT[4]), 
      .B2(n_0_0_443), .ZN(n_0_0_430));
   OAI211_X1 i_0_0_496 (.A(n_0_0_431), .B(n_0_0_432), .C1(n_0_0_487), .C2(
      n_0_0_485), .ZN(MATRIX_CNT_adder_n_24));
   AOI22_X1 i_0_0_497 (.A1(n_0_0_435), .A2(MATRIX_CNT[13]), .B1(MATRIX_CNT[12]), 
      .B2(MATRIX_CNT_adder_n_2), .ZN(n_0_0_431));
   OAI211_X1 i_0_0_498 (.A(n_0_0_469), .B(n_0_0_434), .C1(MATRIX_CNT[6]), 
      .C2(MATRIX_CNT[15]), .ZN(n_0_0_432));
   NAND2_X1 i_0_0_499 (.A1(n_0_0_486), .A2(MATRIX_CNT[15]), .ZN(n_0_0_434));
   NAND2_X1 i_0_0_500 (.A1(n_0_0_440), .A2(n_0_0_436), .ZN(n_0_0_435));
   AOI22_X1 i_0_0_501 (.A1(MATRIX_CNT[7]), .A2(n_0_0_481), .B1(n_0_0_480), 
      .B2(MATRIX_CNT[9]), .ZN(n_0_0_436));
   AOI22_X1 i_0_0_502 (.A1(n_0_0_489), .A2(MATRIX_CNT[11]), .B1(MATRIX_CNT[5]), 
      .B2(n_0_0_443), .ZN(n_0_0_440));
   NOR3_X1 i_0_0_503 (.A1(MATRIX_CNT[15]), .A2(n_0_0_488), .A3(n_0_0_490), 
      .ZN(n_0_0_443));
   INV_X1 i_0_0_504 (.A(VECTOR_CNT_adder_tempIn11[0]), .ZN(n_0_0_447));
   INV_X1 i_0_0_673 (.A(NEW_MATRIX_ADD[5]), .ZN(n_0_0_448));
   INV_X1 i_0_0_674 (.A(NEW_MATRIX_ADD[8]), .ZN(n_0_0_449));
   INV_X1 i_0_0_505 (.A(NEW_MATRIX_ADD[10]), .ZN(n_0_0_450));
   INV_X1 i_0_0_506 (.A(NEW_MATRIX_ADD[11]), .ZN(n_0_0_451));
   INV_X1 i_0_0_677 (.A(NEW_MATRIX_ADD[12]), .ZN(n_0_0_452));
   INV_X1 i_0_0_678 (.A(NEW_VECTOR_ADD[0]), .ZN(n_0_0_453));
   INV_X1 i_0_0_679 (.A(NEW_VECTOR_ADD[2]), .ZN(n_0_0_454));
   INV_X1 i_0_0_680 (.A(NEW_VECTOR_ADD[5]), .ZN(n_0_0_455));
   INV_X1 i_0_0_681 (.A(NEW_VECTOR_ADD[6]), .ZN(n_0_0_456));
   INV_X1 i_0_0_682 (.A(NEW_VECTOR_ADD[10]), .ZN(n_0_0_457));
   INV_X1 i_0_0_683 (.A(NEW_VECTOR_ADD[12]), .ZN(n_0_0_458));
   INV_X1 i_0_0_507 (.A(RESULT_ADD[6]), .ZN(n_0_0_459));
   INV_X1 i_0_0_508 (.A(RESULT_ADD[8]), .ZN(n_0_0_460));
   INV_X1 i_0_0_686 (.A(NEW_RESULT_ADD[6]), .ZN(n_0_0_461));
   INV_X1 i_0_0_687 (.A(NEW_RESULT_ADD[8]), .ZN(n_0_0_462));
   INV_X1 i_0_0_509 (.A(counter[1]), .ZN(n_0_0_463));
   INV_X1 i_0_0_510 (.A(m_val[13]), .ZN(n_0_0_466));
   INV_X1 i_0_0_511 (.A(m_val[14]), .ZN(n_0_0_467));
   INV_X1 i_0_0_512 (.A(m_val[15]), .ZN(n_0_0_468));
   INV_X1 i_0_0_513 (.A(n_val[6]), .ZN(n_0_0_474));
   INV_X1 i_0_0_514 (.A(n_val[7]), .ZN(n_0_0_475));
   INV_X1 i_0_0_515 (.A(MATRIX_CNT[4]), .ZN(n_0_0_482));
   INV_X1 i_0_0_516 (.A(MATRIX_CNT[5]), .ZN(n_0_0_483));
   INV_X1 i_0_0_517 (.A(MATRIX_CNT[7]), .ZN(n_0_0_484));
   INV_X1 i_0_0_518 (.A(MATRIX_CNT[8]), .ZN(n_0_0_485));
   INV_X1 i_0_0_519 (.A(MATRIX_CNT[10]), .ZN(n_0_0_486));
   INV_X1 i_0_0_520 (.A(n_0_0_358), .ZN(n_0_0_491));
   INV_X1 i_0_0_521 (.A(n_0_0_319), .ZN(n_0_0_493));
   OAI21_X1 i_0_0_522 (.A(n_0_0_3), .B1(n_0_0_29), .B2(n_0_0_4), .ZN(
      VECTOR_CNT_adder_n_28));
   AOI22_X1 i_0_0_523 (.A1(VECTOR_CNT[3]), .A2(VECTOR_CNT_adder_n_2), .B1(
      VECTOR_CNT[2]), .B2(n_0_0_9), .ZN(n_0_0_3));
   AOI22_X1 i_0_0_524 (.A1(VECTOR_CNT[1]), .A2(n_0_0_7), .B1(VECTOR_CNT[0]), 
      .B2(n_0_0_5), .ZN(n_0_0_4));
   NOR2_X1 i_0_0_525 (.A1(VECTOR_CNT[14]), .A2(n_0_0_11), .ZN(n_0_0_5));
   NOR2_X1 i_0_0_526 (.A1(n_0_0_13), .A2(VECTOR_CNT[13]), .ZN(n_0_0_7));
   NOR3_X1 i_0_0_527 (.A1(n_0_0_29), .A2(n_0_0_11), .A3(n_0_0_13), .ZN(n_0_0_9));
   NOR2_X1 i_0_0_528 (.A1(VECTOR_CNT[15]), .A2(n_0_0_10), .ZN(
      VECTOR_CNT_adder_n_2));
   NAND2_X1 i_0_0_529 (.A1(n_0_0_13), .A2(n_0_0_11), .ZN(n_0_0_10));
   INV_X1 i_0_0_530 (.A(VECTOR_CNT[13]), .ZN(n_0_0_11));
   INV_X1 i_0_0_531 (.A(VECTOR_CNT[14]), .ZN(n_0_0_13));
   INV_X1 i_0_0_532 (.A(VECTOR_CNT[15]), .ZN(n_0_0_29));
   AOI22_X1 i_0_0_533 (.A1(n_0_0_37), .A2(n_0_0_30), .B1(VECTOR_CNT[13]), 
      .B2(n_0_0_31), .ZN(VECTOR_CNT_adder_n_30));
   AOI222_X1 i_0_0_534 (.A1(VECTOR_CNT[1]), .A2(n_0_0_34), .B1(VECTOR_CNT[5]), 
      .B2(n_0_0_33), .C1(VECTOR_CNT[3]), .C2(n_0_0_32), .ZN(n_0_0_30));
   AOI222_X1 i_0_0_535 (.A1(VECTOR_CNT[0]), .A2(n_0_0_34), .B1(VECTOR_CNT[4]), 
      .B2(n_0_0_33), .C1(VECTOR_CNT[2]), .C2(n_0_0_32), .ZN(n_0_0_31));
   AOI21_X1 i_0_0_536 (.A(n_0_0_35), .B1(VECTOR_CNT[14]), .B2(VECTOR_CNT[13]), 
      .ZN(n_0_0_32));
   OR2_X1 i_0_0_537 (.A1(VECTOR_CNT_adder_n_2), .A2(n_0_0_9), .ZN(n_0_0_33));
   AOI21_X1 i_0_0_538 (.A(n_0_0_36), .B1(VECTOR_CNT[15]), .B2(n_0_0_10), 
      .ZN(n_0_0_34));
   NAND2_X1 i_0_0_539 (.A1(VECTOR_CNT[15]), .A2(n_0_0_10), .ZN(n_0_0_35));
   AOI21_X1 i_0_0_540 (.A(VECTOR_CNT[15]), .B1(VECTOR_CNT[14]), .B2(
      VECTOR_CNT[13]), .ZN(n_0_0_36));
   INV_X1 i_0_0_541 (.A(VECTOR_CNT[13]), .ZN(n_0_0_37));
   OAI211_X1 i_0_0_542 (.A(n_0_0_40), .B(n_0_0_38), .C1(n_0_0_10), .C2(n_0_0_39), 
      .ZN(VECTOR_CNT_adder_n_24));
   AOI22_X1 i_0_0_543 (.A1(VECTOR_CNT[13]), .A2(n_0_0_41), .B1(VECTOR_CNT[12]), 
      .B2(VECTOR_CNT_adder_n_2), .ZN(n_0_0_38));
   NAND2_X1 i_0_0_544 (.A1(VECTOR_CNT[15]), .A2(VECTOR_CNT[8]), .ZN(n_0_0_39));
   OAI221_X1 i_0_0_545 (.A(n_0_0_7), .B1(VECTOR_CNT[10]), .B2(n_0_0_29), 
      .C1(VECTOR_CNT[15]), .C2(VECTOR_CNT[6]), .ZN(n_0_0_40));
   NAND2_X1 i_0_0_546 (.A1(n_0_0_43), .A2(n_0_0_42), .ZN(n_0_0_41));
   AOI22_X1 i_0_0_547 (.A1(VECTOR_CNT[5]), .A2(n_0_0_47), .B1(VECTOR_CNT[9]), 
      .B2(n_0_0_32), .ZN(n_0_0_42));
   AOI22_X1 i_0_0_548 (.A1(VECTOR_CNT[11]), .A2(n_0_0_33), .B1(VECTOR_CNT[7]), 
      .B2(n_0_0_34), .ZN(n_0_0_43));
   AND2_X1 i_0_0_549 (.A1(n_0_0_10), .A2(n_0_0_36), .ZN(n_0_0_47));
   AND4_X1 i_0_0_550 (.A1(n_0_0_64), .A2(n_0_0_59), .A3(n_0_0_49), .A4(n_0_0_150), 
      .ZN(n_0_0_48));
   NOR3_X1 i_0_0_551 (.A1(n_0_0_52), .A2(n_0_0_50), .A3(n_0_0_54), .ZN(n_0_0_49));
   OAI221_X1 i_0_0_552 (.A(n_0_0_51), .B1(n_val[4]), .B2(n_0_0_301), .C1(
      n_0_0_312), .C2(VECTOR_CNT[12]), .ZN(n_0_0_50));
   AOI22_X1 i_0_0_553 (.A1(n_0_0_312), .A2(VECTOR_CNT[12]), .B1(n_0_0_306), 
      .B2(VECTOR_CNT[1]), .ZN(n_0_0_51));
   OAI221_X1 i_0_0_554 (.A(n_0_0_53), .B1(n_0_0_311), .B2(VECTOR_CNT[11]), 
      .C1(n_val[11]), .C2(n_0_0_304), .ZN(n_0_0_52));
   AOI22_X1 i_0_0_555 (.A1(n_0_0_305), .A2(VECTOR_CNT[0]), .B1(n_0_0_309), 
      .B2(VECTOR_CNT[9]), .ZN(n_0_0_53));
   NAND4_X1 i_0_0_556 (.A1(n_0_0_58), .A2(n_0_0_57), .A3(n_0_0_56), .A4(n_0_0_55), 
      .ZN(n_0_0_54));
   XNOR2_X1 i_0_0_557 (.A(n_val[3]), .B(VECTOR_CNT[3]), .ZN(n_0_0_55));
   XNOR2_X1 i_0_0_558 (.A(n_val[10]), .B(VECTOR_CNT[10]), .ZN(n_0_0_56));
   AOI211_X1 i_0_0_559 (.A(n_0_0_298), .B(state[0]), .C1(n_val[4]), .C2(
      n_0_0_301), .ZN(n_0_0_57));
   XNOR2_X1 i_0_0_560 (.A(n_val[5]), .B(VECTOR_CNT[5]), .ZN(n_0_0_58));
   NOR2_X1 i_0_0_561 (.A1(n_0_0_62), .A2(n_0_0_60), .ZN(n_0_0_59));
   OAI221_X1 i_0_0_562 (.A(n_0_0_61), .B1(n_0_0_309), .B2(VECTOR_CNT[9]), 
      .C1(n_val[6]), .C2(n_0_0_302), .ZN(n_0_0_60));
   AOI22_X1 i_0_0_563 (.A1(n_val[6]), .A2(n_0_0_302), .B1(n_val[0]), .B2(
      n_0_0_299), .ZN(n_0_0_61));
   OAI221_X1 i_0_0_564 (.A(n_0_0_63), .B1(n_val[2]), .B2(n_0_0_300), .C1(
      n_0_0_308), .C2(VECTOR_CNT[7]), .ZN(n_0_0_62));
   AOI22_X1 i_0_0_565 (.A1(n_0_0_308), .A2(VECTOR_CNT[7]), .B1(n_val[8]), 
      .B2(n_0_0_303), .ZN(n_0_0_63));
   AOI21_X1 i_0_0_566 (.A(n_0_0_65), .B1(n_val[2]), .B2(n_0_0_300), .ZN(n_0_0_64));
   OAI22_X1 i_0_0_567 (.A1(n_val[8]), .A2(n_0_0_303), .B1(n_0_0_306), .B2(
      VECTOR_CNT[1]), .ZN(n_0_0_65));
   NOR4_X1 i_0_0_568 (.A1(n_0_0_152), .A2(n_0_0_151), .A3(n_0_0_180), .A4(
      n_0_0_181), .ZN(n_0_0_150));
   XOR2_X1 i_0_0_569 (.A(n_val[13]), .B(VECTOR_CNT[13]), .Z(n_0_0_151));
   XNOR2_X1 i_0_0_570 (.A(n_val[15]), .B(n_0_0_29), .ZN(n_0_0_152));
   XNOR2_X1 i_0_0_571 (.A(n_val[14]), .B(n_0_0_13), .ZN(n_0_0_180));
   OR3_X1 i_0_0_572 (.A1(n_0_0_245), .A2(n_0_0_204), .A3(n_0_0_198), .ZN(
      n_0_0_181));
   NAND4_X1 i_0_0_573 (.A1(n_0_0_203), .A2(n_0_0_202), .A3(n_0_0_201), .A4(
      n_0_0_200), .ZN(n_0_0_198));
   NOR4_X1 i_0_0_574 (.A1(n_val[55]), .A2(n_val[52]), .A3(n_val[50]), .A4(
      n_val[49]), .ZN(n_0_0_200));
   NOR4_X1 i_0_0_575 (.A1(n_val[62]), .A2(n_val[61]), .A3(n_val[59]), .A4(
      n_val[56]), .ZN(n_0_0_201));
   NOR4_X1 i_0_0_576 (.A1(n_val[35]), .A2(n_val[32]), .A3(n_val[38]), .A4(
      n_val[37]), .ZN(n_0_0_202));
   NOR4_X1 i_0_0_577 (.A1(n_val[42]), .A2(n_val[41]), .A3(n_val[47]), .A4(
      n_val[44]), .ZN(n_0_0_203));
   NAND4_X1 i_0_0_578 (.A1(n_0_0_244), .A2(n_0_0_243), .A3(n_0_0_236), .A4(
      n_0_0_241), .ZN(n_0_0_204));
   NOR4_X1 i_0_0_579 (.A1(n_val[63]), .A2(n_val[60]), .A3(n_val[58]), .A4(
      n_val[57]), .ZN(n_0_0_236));
   NOR4_X1 i_0_0_580 (.A1(n_val[54]), .A2(n_val[53]), .A3(n_val[51]), .A4(
      n_val[48]), .ZN(n_0_0_241));
   NOR4_X1 i_0_0_581 (.A1(n_val[39]), .A2(n_val[36]), .A3(n_val[34]), .A4(
      n_val[33]), .ZN(n_0_0_243));
   NOR4_X1 i_0_0_582 (.A1(n_val[46]), .A2(n_val[45]), .A3(n_val[43]), .A4(
      n_val[40]), .ZN(n_0_0_244));
   NAND4_X1 i_0_0_583 (.A1(n_0_0_297), .A2(n_0_0_296), .A3(n_0_0_295), .A4(
      n_0_0_294), .ZN(n_0_0_245));
   NOR4_X1 i_0_0_584 (.A1(n_val[18]), .A2(n_val[17]), .A3(n_val[23]), .A4(
      n_val[20]), .ZN(n_0_0_294));
   NOR4_X1 i_0_0_585 (.A1(n_val[27]), .A2(n_val[24]), .A3(n_val[30]), .A4(
      n_val[29]), .ZN(n_0_0_295));
   NOR4_X1 i_0_0_586 (.A1(n_val[19]), .A2(n_val[16]), .A3(n_val[22]), .A4(
      n_val[21]), .ZN(n_0_0_296));
   NOR4_X1 i_0_0_587 (.A1(n_val[26]), .A2(n_val[25]), .A3(n_val[31]), .A4(
      n_val[28]), .ZN(n_0_0_297));
   INV_X1 i_0_0_588 (.A(state[1]), .ZN(n_0_0_298));
   INV_X1 i_0_0_589 (.A(VECTOR_CNT[0]), .ZN(n_0_0_299));
   INV_X1 i_0_0_590 (.A(VECTOR_CNT[2]), .ZN(n_0_0_300));
   INV_X1 i_0_0_591 (.A(VECTOR_CNT[4]), .ZN(n_0_0_301));
   INV_X1 i_0_0_592 (.A(VECTOR_CNT[6]), .ZN(n_0_0_302));
   INV_X1 i_0_0_593 (.A(VECTOR_CNT[8]), .ZN(n_0_0_303));
   INV_X1 i_0_0_594 (.A(VECTOR_CNT[11]), .ZN(n_0_0_304));
   INV_X1 i_0_0_595 (.A(n_val[0]), .ZN(n_0_0_305));
   INV_X1 i_0_0_596 (.A(n_val[1]), .ZN(n_0_0_306));
   INV_X1 i_0_0_597 (.A(n_val[3]), .ZN(n_0_0_307));
   INV_X1 i_0_0_598 (.A(n_val[7]), .ZN(n_0_0_308));
   INV_X1 i_0_0_599 (.A(n_val[9]), .ZN(n_0_0_309));
   INV_X1 i_0_0_600 (.A(n_val[10]), .ZN(n_0_0_310));
   INV_X1 i_0_0_601 (.A(n_val[11]), .ZN(n_0_0_311));
   INV_X1 i_0_0_602 (.A(n_val[12]), .ZN(n_0_0_312));
   INV_X1 i_0_0_603 (.A(n_val[13]), .ZN(n_0_0_313));
   OAI21_X1 i_0_0_604 (.A(n_0_0_315), .B1(CLK), .B2(n_0_0_314), .ZN(n_0_117));
   NOR2_X1 i_0_0_605 (.A1(n_0_0_329), .A2(n_0_0_325), .ZN(n_0_0_314));
   NOR2_X1 i_0_0_606 (.A1(n_0_0_318), .A2(n_0_0_316), .ZN(n_0_0_315));
   INV_X1 i_0_0_607 (.A(n_0_0_317), .ZN(n_0_0_316));
   NAND3_X1 i_0_0_608 (.A1(state[0]), .A2(n_0_0_324), .A3(
      Matrix_Multiplication2_Enable), .ZN(n_0_0_317));
   NAND2_X1 i_0_0_609 (.A1(n_0_0_323), .A2(n_0_0_319), .ZN(n_0_0_318));
   NAND3_X1 i_0_0_610 (.A1(n_0_0_336), .A2(n_0_0_322), .A3(Final_Calc_Enable), 
      .ZN(n_0_0_319));
   NOR2_X1 i_0_0_611 (.A1(n_0_0_342), .A2(n_0_0_298), .ZN(n_0_0_322));
   NAND3_X1 i_0_0_612 (.A1(n_0_0_336), .A2(n_0_0_324), .A3(
      Matrix_Multiplication1_Enable), .ZN(n_0_0_323));
   NOR2_X1 i_0_0_614 (.A1(n_0_0_342), .A2(state[1]), .ZN(n_0_0_324));
   AND2_X1 i_0_0_615 (.A1(n_0_0_328), .A2(n_0_0_326), .ZN(n_0_0_325));
   NOR2_X1 i_0_0_616 (.A1(counter[1]), .A2(counter[0]), .ZN(n_0_0_326));
   INV_X1 i_0_0_617 (.A(n_0_0_328), .ZN(n_0_0_327));
   NOR3_X1 i_0_0_618 (.A1(n_0_0_345), .A2(next[0]), .A3(n_0_0_344), .ZN(
      n_0_0_328));
   NOR2_X1 i_0_0_619 (.A1(n_0_0_345), .A2(next[1]), .ZN(n_0_0_329));
   INV_X1 i_0_0_620 (.A(state[0]), .ZN(n_0_0_336));
   INV_X1 i_0_0_621 (.A(state[2]), .ZN(n_0_0_342));
   INV_X1 i_0_0_622 (.A(next[1]), .ZN(n_0_0_344));
   INV_X1 i_0_0_623 (.A(next[2]), .ZN(n_0_0_345));
   INV_X1 i_0_0_624 (.A(CLK), .ZN(n_0_51));
   AND2_X1 i_0_0_625 (.A1(n_0_0_347), .A2(n_0_0_329), .ZN(n_0_0_346));
   INV_X1 i_0_0_626 (.A(n_0_0_318), .ZN(n_0_0_347));
   NOR4_X1 i_0_0_627 (.A1(n_0_0_351), .A2(n_0_0_349), .A3(n_0_0_350), .A4(
      n_0_0_352), .ZN(n_0_0_348));
   NOR3_X1 i_0_0_628 (.A1(n_0_0_360), .A2(n_0_0_359), .A3(m_val[2]), .ZN(
      n_0_0_349));
   XNOR2_X1 i_0_0_629 (.A(m_val[1]), .B(n_0_0_356), .ZN(n_0_0_350));
   AND2_X1 i_0_0_630 (.A1(m_val[2]), .A2(n_0_0_357), .ZN(n_0_0_351));
   NAND3_X1 i_0_0_631 (.A1(n_0_0_355), .A2(n_0_0_353), .A3(n_0_0_354), .ZN(
      n_0_0_352));
   NOR4_X1 i_0_0_632 (.A1(m_val[21]), .A2(m_val[20]), .A3(m_val[19]), .A4(
      m_val[18]), .ZN(n_0_0_353));
   NOR4_X1 i_0_0_633 (.A1(m_val[25]), .A2(m_val[24]), .A3(m_val[23]), .A4(
      m_val[22]), .ZN(n_0_0_354));
   NOR3_X1 i_0_0_634 (.A1(m_val[17]), .A2(next[0]), .A3(m_val[16]), .ZN(
      n_0_0_355));
   XNOR2_X1 i_0_0_635 (.A(VECTOR_CNT_adder_tempIn11[1]), .B(
      VECTOR_CNT_adder_tempIn11[0]), .ZN(n_0_0_356));
   OR2_X1 i_0_0_636 (.A1(n_0_0_360), .A2(n_0_0_358), .ZN(n_0_0_357));
   AND3_X1 i_0_0_637 (.A1(VECTOR_CNT_adder_tempIn11[2]), .A2(
      VECTOR_CNT_adder_tempIn11[1]), .A3(VECTOR_CNT_adder_tempIn11[0]), .ZN(
      n_0_0_358));
   XOR2_X1 i_0_0_639 (.A(VECTOR_CNT_adder_tempIn11[3]), .B(m_val[3]), .Z(
      n_0_0_359));
   AOI21_X1 i_0_0_640 (.A(VECTOR_CNT_adder_tempIn11[2]), .B1(
      VECTOR_CNT_adder_tempIn11[1]), .B2(VECTOR_CNT_adder_tempIn11[0]), .ZN(
      n_0_0_360));
   OAI221_X1 i_0_0_641 (.A(n_0_0_362), .B1(n_0_0_387), .B2(n_0_0_366), .C1(
      m_val[8]), .C2(n_0_0_365), .ZN(n_0_0_361));
   AOI211_X1 i_0_0_646 (.A(n_0_0_363), .B(n_0_0_364), .C1(m_val[6]), .C2(
      n_0_0_369), .ZN(n_0_0_362));
   XNOR2_X1 i_0_0_647 (.A(m_val[5]), .B(n_0_0_374), .ZN(n_0_0_363));
   XNOR2_X1 i_0_0_648 (.A(m_val[4]), .B(n_0_0_378), .ZN(n_0_0_364));
   INV_X1 i_0_0_649 (.A(n_0_0_366), .ZN(n_0_0_365));
   AOI21_X1 i_0_0_650 (.A(n_0_0_367), .B1(n_0_0_389), .B2(n_0_0_368), .ZN(
      n_0_0_366));
   NOR2_X1 i_0_0_651 (.A1(n_0_0_389), .A2(n_0_0_368), .ZN(n_0_0_367));
   NAND2_X1 i_0_0_652 (.A1(VECTOR_CNT_adder_tempIn11[7]), .A2(n_0_0_371), 
      .ZN(n_0_0_368));
   OAI21_X1 i_0_0_653 (.A(n_0_0_372), .B1(VECTOR_CNT_adder_tempIn11[6]), 
      .B2(n_0_0_375), .ZN(n_0_0_369));
   INV_X1 i_0_0_654 (.A(n_0_0_372), .ZN(n_0_0_371));
   NAND2_X1 i_0_0_655 (.A1(VECTOR_CNT_adder_tempIn11[6]), .A2(n_0_0_375), 
      .ZN(n_0_0_372));
   OAI21_X1 i_0_0_656 (.A(n_0_0_376), .B1(VECTOR_CNT_adder_tempIn11[5]), 
      .B2(n_0_0_383), .ZN(n_0_0_374));
   INV_X1 i_0_0_657 (.A(n_0_0_376), .ZN(n_0_0_375));
   NAND2_X1 i_0_0_658 (.A1(VECTOR_CNT_adder_tempIn11[5]), .A2(n_0_0_383), 
      .ZN(n_0_0_376));
   OAI21_X1 i_0_0_659 (.A(n_0_0_384), .B1(VECTOR_CNT_adder_tempIn11[4]), 
      .B2(n_0_0_386), .ZN(n_0_0_378));
   INV_X1 i_0_0_660 (.A(n_0_0_384), .ZN(n_0_0_383));
   NAND2_X1 i_0_0_661 (.A1(VECTOR_CNT_adder_tempIn11[4]), .A2(n_0_0_386), 
      .ZN(n_0_0_384));
   AND2_X1 i_0_0_662 (.A1(VECTOR_CNT_adder_tempIn11[3]), .A2(n_0_0_358), 
      .ZN(n_0_0_386));
   INV_X1 i_0_0_663 (.A(m_val[8]), .ZN(n_0_0_387));
   INV_X1 i_0_0_664 (.A(VECTOR_CNT_adder_tempIn11[8]), .ZN(n_0_0_389));
   AND4_X1 i_0_0_665 (.A1(VECTOR_CNT_adder_tempIn11[9]), .A2(
      VECTOR_CNT_adder_tempIn11[8]), .A3(VECTOR_CNT_adder_tempIn11[7]), .A4(
      n_0_0_371), .ZN(n_0_0_390));
   NOR2_X1 i_0_0_666 (.A1(n_0_0_390), .A2(VECTOR_CNT_adder_tempIn11[10]), 
      .ZN(n_0_0_391));
   NAND2_X1 i_0_0_667 (.A1(n_0_0_390), .A2(VECTOR_CNT_adder_tempIn11[10]), 
      .ZN(n_0_0_392));
   INV_X1 i_0_0_668 (.A(n_0_0_392), .ZN(n_0_0_395));
   OR2_X1 i_0_0_669 (.A1(n_0_0_391), .A2(n_0_0_395), .ZN(n_0_0_398));
   INV_X1 i_0_0_670 (.A(VECTOR_CNT_adder_tempIn11[11]), .ZN(n_0_0_405));
   NOR2_X1 i_0_0_671 (.A1(n_0_0_392), .A2(n_0_0_405), .ZN(n_0_0_406));
   NAND2_X1 i_0_0_672 (.A1(n_0_0_405), .A2(m_val[11]), .ZN(n_0_0_407));
   OR3_X1 i_0_0_675 (.A1(n_0_0_392), .A2(m_val[10]), .A3(n_0_0_407), .ZN(
      n_0_0_410));
   OAI221_X1 i_0_0_676 (.A(n_0_0_407), .B1(n_0_0_405), .B2(m_val[11]), .C1(
      n_0_0_391), .C2(m_val[10]), .ZN(n_0_0_411));
   AND2_X1 i_0_0_684 (.A1(n_0_0_398), .A2(m_val[10]), .ZN(n_0_0_412));
   OAI21_X1 i_0_0_685 (.A(n_0_0_410), .B1(n_0_0_411), .B2(n_0_0_412), .ZN(
      n_0_0_413));
   XNOR2_X1 i_0_0_688 (.A(m_val[12]), .B(VECTOR_CNT_adder_tempIn11[12]), 
      .ZN(n_0_0_414));
   NOR3_X1 i_0_0_689 (.A1(n_0_0_414), .A2(m_val[10]), .A3(m_val[11]), .ZN(
      n_0_0_415));
   AOI22_X1 i_0_0_690 (.A1(n_0_0_413), .A2(n_0_0_414), .B1(n_0_0_406), .B2(
      n_0_0_415), .ZN(n_0_0_433));
   OAI221_X1 i_0_0_691 (.A(n_0_0_438), .B1(n_0_0_310), .B2(n_0_0_441), .C1(
      n_val[8]), .C2(n_0_0_365), .ZN(n_0_0_437));
   AOI221_X1 i_0_0_692 (.A(n_0_0_439), .B1(n_val[7]), .B2(n_0_0_445), .C1(
      n_val[8]), .C2(n_0_0_365), .ZN(n_0_0_438));
   NOR2_X1 i_0_0_693 (.A1(n_val[7]), .A2(n_0_0_445), .ZN(n_0_0_439));
   NOR3_X1 i_0_0_694 (.A1(n_0_0_444), .A2(n_0_0_442), .A3(n_0_0_398), .ZN(
      n_0_0_441));
   XNOR2_X1 i_0_0_695 (.A(VECTOR_CNT_adder_tempIn11[11]), .B(n_0_0_311), 
      .ZN(n_0_0_442));
   XOR2_X1 i_0_0_696 (.A(VECTOR_CNT_adder_tempIn11[12]), .B(n_val[12]), .Z(
      n_0_0_444));
   XNOR2_X1 i_0_0_697 (.A(VECTOR_CNT_adder_tempIn11[7]), .B(n_0_0_371), .ZN(
      n_0_0_445));
   OAI21_X1 i_0_0_698 (.A(n_0_0_446), .B1(n_0_0_476), .B2(n_0_0_464), .ZN(
      MATRIX_CNT_adder_n_28));
   AOI22_X1 i_0_0_699 (.A1(MATRIX_CNT[3]), .A2(MATRIX_CNT_adder_n_2), .B1(
      MATRIX_CNT[2]), .B2(n_0_0_470), .ZN(n_0_0_446));
   AOI22_X1 i_0_0_700 (.A1(MATRIX_CNT[1]), .A2(n_0_0_469), .B1(MATRIX_CNT[0]), 
      .B2(n_0_0_465), .ZN(n_0_0_464));
   NOR2_X1 i_0_0_701 (.A1(MATRIX_CNT[14]), .A2(n_0_0_472), .ZN(n_0_0_465));
   NOR2_X1 i_0_0_702 (.A1(n_0_0_473), .A2(MATRIX_CNT[13]), .ZN(n_0_0_469));
   NOR2_X1 i_0_0_703 (.A1(n_0_0_476), .A2(n_0_0_471), .ZN(n_0_0_470));
   NAND2_X1 i_0_0_704 (.A1(MATRIX_CNT[14]), .A2(MATRIX_CNT[13]), .ZN(n_0_0_471));
   NOR3_X1 i_0_0_705 (.A1(MATRIX_CNT[15]), .A2(MATRIX_CNT[13]), .A3(
      MATRIX_CNT[14]), .ZN(MATRIX_CNT_adder_n_2));
   INV_X1 i_0_0_706 (.A(MATRIX_CNT[13]), .ZN(n_0_0_472));
   INV_X1 i_0_0_707 (.A(MATRIX_CNT[14]), .ZN(n_0_0_473));
   INV_X1 i_0_0_708 (.A(MATRIX_CNT[15]), .ZN(n_0_0_476));
   OAI22_X1 i_0_0_709 (.A1(n_0_0_492), .A2(n_0_0_477), .B1(MATRIX_CNT[13]), 
      .B2(n_0_0_479), .ZN(MATRIX_CNT_adder_n_30));
   AOI222_X1 i_0_0_710 (.A1(MATRIX_CNT[0]), .A2(n_0_0_481), .B1(MATRIX_CNT[4]), 
      .B2(n_0_0_489), .C1(MATRIX_CNT[2]), .C2(n_0_0_480), .ZN(n_0_0_477));
   INV_X1 i_0_0_711 (.A(n_0_0_479), .ZN(n_0_0_478));
   AOI222_X1 i_0_0_712 (.A1(MATRIX_CNT[1]), .A2(n_0_0_481), .B1(MATRIX_CNT[5]), 
      .B2(n_0_0_489), .C1(MATRIX_CNT[3]), .C2(n_0_0_480), .ZN(n_0_0_479));
   NOR3_X1 i_0_0_713 (.A1(n_0_0_490), .A2(n_0_0_488), .A3(n_0_0_476), .ZN(
      n_0_0_480));
   OAI21_X1 i_0_0_714 (.A(n_0_0_487), .B1(MATRIX_CNT[15]), .B2(n_0_0_471), 
      .ZN(n_0_0_481));
   NAND2_X1 i_0_0_715 (.A1(MATRIX_CNT[15]), .A2(n_0_0_488), .ZN(n_0_0_487));
   NOR2_X1 i_0_0_716 (.A1(MATRIX_CNT[14]), .A2(MATRIX_CNT[13]), .ZN(n_0_0_488));
   OR2_X1 i_0_0_717 (.A1(MATRIX_CNT_adder_n_2), .A2(n_0_0_470), .ZN(n_0_0_489));
   INV_X1 i_0_0_718 (.A(n_0_0_471), .ZN(n_0_0_490));
   INV_X1 i_0_0_719 (.A(MATRIX_CNT[13]), .ZN(n_0_0_492));
endmodule
