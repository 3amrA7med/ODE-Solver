/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 22:22:10 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3240293018 */

module Division_CSA(reset, clk, dividend, divisor, Q, ready, overFlow, 
      divideByZero);
   input reset;
   input clk;
   input [15:0]dividend;
   input [15:0]divisor;
   output [15:0]Q;
   output ready;
   output overFlow;
   output divideByZero;

   wire csa0_n_0;
   wire csa0_n_1;
   wire csa1_n_0;
   wire n_0_0;
   wire n_0_1;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_2;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire [15:0]negated_second_operand_number;
   wire [15:0]second_operand_number;
   wire n_0_3;
   wire [4:0]number_of_bits_in_dividend;
   wire sign;
   wire n_0_6;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_0_0;
   wire n_0_57;
   wire n_0_0_1;
   wire n_0_58;
   wire n_0_0_2;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_76;
   wire n_0_0_7;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_77;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_78;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_79;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_80;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_81;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_82;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_83;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_84;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_85;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_86;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_87;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_71;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_89;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_90;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_101;
   wire n_0_0_103;
   wire n_0_0_112;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_124;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_154;
   wire n_0_93;
   wire n_0_0_155;
   wire n_0_94;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_95;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_96;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_97;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_98;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_99;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_100;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_101;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_102;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_103;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_104;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_105;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_106;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_107;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_247;
   wire n_0_0_72;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_281;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_53;
   wire n_0_0_283;
   wire n_0_74;
   wire n_0_75;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_287;
   wire n_0_60;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_4;
   wire n_0_5;
   wire n_0_0_291;
   wire n_0_7;
   wire n_0_8;
   wire n_0_0_292;
   wire n_0_9;
   wire n_0_10;
   wire n_0_0_293;
   wire n_0_11;
   wire n_0_12;
   wire n_0_0_294;
   wire n_0_13;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_126;
   wire n_0_124;
   wire n_0_0_331;
   wire n_0_0_342;
   wire n_0_118;
   wire n_0_0_360;
   wire n_0_0_366;
   wire n_0_0_372;
   wire n_0_0_376;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_385;
   wire n_0_0_387;
   wire n_0_0_394;
   wire n_0_0_395;
   wire n_0_0_396;
   wire n_0_0_399;
   wire n_0_0_411;
   wire n_0_0_412;
   wire n_0_0_426;
   wire n_0_0_427;
   wire n_0_0_428;
   wire n_0_0_429;
   wire n_0_0_435;
   wire n_0_0_436;
   wire n_0_0_437;
   wire n_0_0_438;
   wire n_0_0_439;
   wire n_0_0_440;
   wire n_0_0_441;
   wire n_0_0_442;
   wire n_0_0_443;
   wire n_0_0_444;
   wire n_0_0_448;
   wire n_0_0_451;
   wire n_0_0_452;
   wire n_0_0_453;
   wire n_0_0_460;
   wire n_0_0_461;
   wire n_0_0_462;
   wire n_0_0_463;
   wire n_0_0_464;
   wire n_0_0_465;
   wire n_0_0_472;
   wire n_0_0_474;
   wire n_0_0_480;
   wire n_0_0_321;
   wire n_0_0_367;
   wire n_0_0_373;
   wire n_0_0_3;
   wire n_0_117;
   wire n_0_123;
   wire n_0_0_4;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_102;
   wire n_0_0_450;
   wire n_0_0_392;
   wire n_0_116;
   wire n_0_0_368;
   wire n_0_0_322;
   wire n_0_0_377;
   wire n_0_115;
   wire n_0_114;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_361;
   wire n_0_0_353;
   wire n_0_0_352;
   wire n_0_119;
   wire n_0_0_343;
   wire n_0_0_334;
   wire n_0_0_333;
   wire n_0_121;
   wire n_0_0_328;
   wire n_0_0_317;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_123;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_136;
   wire n_0_0_311;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_304;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_122;
   wire n_0_0_286;
   wire n_0_0_459;
   wire n_0_0_135;
   wire n_0_0_309;
   wire n_0_0_113;
   wire n_0_0_139;
   wire n_0_0_310;
   wire n_0_0_140;
   wire n_0_0_282;
   wire n_0_0_449;
   wire n_0_88;
   wire n_0_0_312;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_323;
   wire n_0_0_85;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_88;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_335;
   wire n_0_0_125;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_64;
   wire n_0_0_152;
   wire n_0_91;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_344;
   wire n_0_0_100;
   wire n_0_0_345;
   wire n_0_0_104;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_350;
   wire n_0_92;
   wire n_0_0_351;
   wire n_0_0_280;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_0_362;
   wire n_0_0_114;
   wire n_0_0_363;
   wire n_0_0_116;
   wire n_0_0_364;
   wire n_0_0_115;
   wire n_0_0_365;
   wire n_0_0_369;
   wire n_0_0_370;
   wire n_0_0_371;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_0_142;
   wire n_0_0_141;
   wire n_0_0_383;
   wire n_0_0_143;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_391;
   wire n_0_0_401;
   wire n_0_0_405;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_0_417;
   wire n_0_0_418;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_423;
   wire n_0_0_446;
   wire n_0_0_445;
   wire n_0_0_447;
   wire n_0_0_475;
   wire n_0_0_476;
   wire n_0_0_477;
   wire n_0_0_481;
   wire n_0_0_145;
   wire n_0_0_144;
   wire n_0_0_482;
   wire n_0_0_483;
   wire n_0_0_484;
   wire n_0_0_149;
   wire n_0_0_148;
   wire n_0_0_153;
   wire n_0_0_485;
   wire n_0_0_486;
   wire n_0_127;
   wire n_0_0_487;
   wire n_0_0_488;
   wire n_0_0_489;
   wire n_0_0_490;
   wire n_0_0_491;
   wire n_0_0_393;
   wire n_0_0_492;
   wire n_0_128;
   wire n_0_129;
   wire n_0_0_493;
   wire n_0_0_494;
   wire n_0_0_495;
   wire n_0_0_496;
   wire n_0_0_497;
   wire n_0_0_498;
   wire n_0_0_499;
   wire n_0_0_500;
   wire n_0_0_501;
   wire n_0_0_424;
   wire n_0_0_502;
   wire n_0_0_503;
   wire n_0_0_504;
   wire n_0_122;
   wire n_0_120;
   wire n_0_0_505;
   wire n_0_0_506;
   wire n_0_0_507;
   wire n_0_0_508;
   wire n_0_0_509;
   wire n_0_0_510;
   wire n_0_0_511;
   wire n_0_0_512;
   wire n_0_0_513;
   wire n_0_0_514;
   wire n_0_0_515;
   wire n_0_0_516;
   wire n_0_0_329;
   wire n_0_0_517;
   wire n_0_0_518;
   wire n_0_0_519;
   wire n_0_0_520;
   wire n_0_0_521;
   wire n_0_0_522;
   wire n_0_0_523;
   wire n_0_0_524;
   wire n_0_0_525;
   wire n_0_0_526;
   wire n_0_0_527;
   wire n_0_0_528;
   wire n_0_0_529;
   wire n_0_0_336;
   wire n_0_0_530;
   wire n_0_0_330;
   wire n_0_0_332;
   wire n_0_0_397;
   wire n_0_0_305;
   wire n_0_59;
   wire n_0_0_531;
   wire n_0_113;
   wire n_0_0_532;
   wire n_0_0_533;
   wire n_0_20;
   wire n_0_14;
   wire n_0_0_534;
   wire n_0_0_316;
   wire n_0_0_535;
   wire n_0_15;
   wire n_0_0_536;
   wire n_0_0_537;
   wire n_0_125;
   wire n_0_16;
   wire n_0_0_538;
   wire n_0_0_539;
   wire n_0_0_540;
   wire n_0_17;
   wire n_0_0_541;
   wire n_0_0_542;
   wire n_0_0_543;
   wire n_0_0_303;
   wire n_0_0_544;
   wire n_0_18;
   wire n_0_0_545;
   wire n_0_0_546;
   wire n_0_0_547;
   wire n_0_19;
   wire n_0_0_548;
   wire n_0_0_549;
   wire n_0_0_550;
   wire n_0_0_551;
   wire n_0_0_552;
   wire n_0_0_553;
   wire n_0_0_554;
   wire n_0_0_555;
   wire n_0_0_556;
   wire n_0_0_557;
   wire n_0_0_558;
   wire n_0_0_559;
   wire n_0_0_560;
   wire n_0_0_561;
   wire n_0_0_562;
   wire n_0_0_563;
   wire n_0_0_564;
   wire n_0_0_565;
   wire n_0_0_384;
   wire n_0_0_566;
   wire n_0_0_567;
   wire n_0_0_568;
   wire n_0_0_569;
   wire n_0_0_570;
   wire n_0_0_386;
   wire n_0_0_571;
   wire n_0_0_572;
   wire n_0_0_573;
   wire n_0_0_574;
   wire n_0_0_575;
   wire n_0_0_576;
   wire n_0_0_577;
   wire n_0_0_578;
   wire n_0_0_579;
   wire n_0_0_580;
   wire n_0_0_581;
   wire n_0_0_403;
   wire n_0_0_404;
   wire n_0_0_582;
   wire n_0_0_583;
   wire n_0_0_584;
   wire n_0_0_585;
   wire n_0_0_586;
   wire n_0_0_587;
   wire n_0_0_588;
   wire n_0_0_589;
   wire n_0_0_590;
   wire n_0_0_382;
   wire n_0_0_591;
   wire n_0_0_592;
   wire n_0_0_593;
   wire n_0_0_594;
   wire n_0_0_595;
   wire n_0_0_596;
   wire n_0_0_597;
   wire n_0_0_598;
   wire n_0_0_599;
   wire n_0_0_600;
   wire n_0_0_601;
   wire n_0_0_602;
   wire n_0_0_603;
   wire n_0_0_604;
   wire n_0_0_605;
   wire n_0_0_606;
   wire n_0_0_607;
   wire n_0_0_608;
   wire n_0_0_609;
   wire n_0_0_610;
   wire n_0_0_611;
   wire n_0_0_612;
   wire n_0_0_613;
   wire n_0_0_614;
   wire n_0_0_615;
   wire n_0_0_616;
   wire n_0_0_617;
   wire n_0_0_618;
   wire n_0_0_619;
   wire n_0_0_620;
   wire n_0_0_621;
   wire n_0_0_622;
   wire n_0_0_623;
   wire n_0_0_349;
   wire n_0_0_624;
   wire n_0_0_625;
   wire n_0_0_626;
   wire n_0_0_627;
   wire n_0_0_628;
   wire n_0_0_629;
   wire n_0_0_630;
   wire n_0_0_631;
   wire n_0_0_632;
   wire n_0_0_633;
   wire n_0_0_634;
   wire n_0_0_635;
   wire n_0_0_636;
   wire n_0_0_637;
   wire n_0_0_638;
   wire n_0_0_639;
   wire n_0_0_640;
   wire n_0_0_641;
   wire n_0_0_642;
   wire n_0_0_643;
   wire n_0_0_644;
   wire n_0_0_645;
   wire n_0_0_646;
   wire n_0_0_647;
   wire n_0_0_648;
   wire n_0_0_649;
   wire n_0_0_650;
   wire n_0_0_651;
   wire n_0_0_652;
   wire n_0_0_653;
   wire n_0_0_654;
   wire n_0_0_655;
   wire n_0_0_656;
   wire n_0_0_657;
   wire n_0_0_658;
   wire n_0_0_659;
   wire n_0_0_660;
   wire n_0_0_661;
   wire n_0_0_662;
   wire n_0_0_663;
   wire n_0_0_664;
   wire n_0_0_398;
   wire n_0_0_665;
   wire n_0_0_666;
   wire n_0_0_667;
   wire n_0_0_668;
   wire n_0_0_669;
   wire n_0_0_670;
   wire n_0_0_671;
   wire n_0_0_672;
   wire n_0_0_673;
   wire n_0_0_674;
   wire n_0_0_675;
   wire n_0_0_676;
   wire n_0_0_409;
   wire n_0_0_677;
   wire n_0_0_678;
   wire n_0_0_679;
   wire n_0_0_680;
   wire n_0_0_402;
   wire n_0_0_681;
   wire n_0_0_682;
   wire n_0_0_408;
   wire n_0_0_683;
   wire n_0_0_684;
   wire n_0_0_685;
   wire n_0_0_686;
   wire n_0_0_687;
   wire n_0_0_688;
   wire n_0_0_689;
   wire n_0_0_690;
   wire n_0_0_691;
   wire n_0_0_414;
   wire n_0_0_413;
   wire n_0_0_692;
   wire n_0_0_693;
   wire n_0_0_694;
   wire n_0_0_695;
   wire n_0_0_696;
   wire n_0_0_697;
   wire n_0_0_479;
   wire n_0_0_698;
   wire n_0_0_699;
   wire n_0_0_416;
   wire n_0_0_700;
   wire n_0_0_400;
   wire n_0_0_701;
   wire n_0_0_702;
   wire n_0_0_703;
   wire n_0_0_704;
   wire n_0_0_705;
   wire n_0_0_706;
   wire n_0_0_707;
   wire n_0_0_708;
   wire n_0_0_709;
   wire n_0_0_710;
   wire n_0_0_410;
   wire n_0_0_711;
   wire n_0_0_473;
   wire n_0_0_712;
   wire n_0_0_713;
   wire n_0_0_714;
   wire n_0_0_715;
   wire n_0_0_716;
   wire n_0_0_717;
   wire n_0_0_718;
   wire n_0_0_478;
   wire n_0_0_390;
   wire n_0_0_719;
   wire n_0_0_720;
   wire n_0_0_721;
   wire n_0_0_722;
   wire n_0_0_723;
   wire n_0_0_724;
   wire n_0_0_415;
   wire n_0_0_725;
   wire n_0_0_726;
   wire n_0_0_727;
   wire n_0_0_728;
   wire n_0_0_729;
   wire n_0_0_730;
   wire n_0_0_731;
   wire n_0_0_732;
   wire n_0_0_733;
   wire n_0_0_734;
   wire n_0_0_735;
   wire n_0_0_421;
   wire n_0_0_422;
   wire n_0_0_736;
   wire n_0_0_8;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_246;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_318;
   wire n_0_0_425;
   wire n_0_0_430;
   wire n_0_0_431;
   wire n_0_0_432;
   wire n_0_0_433;
   wire n_0_0_434;
   wire n_0_0_454;
   wire n_0_0_455;
   wire n_0_0_456;
   wire n_0_0_457;
   wire n_0_0_458;
   wire n_0_0_466;
   wire n_0_0_467;
   wire n_0_0_468;
   wire n_0_0_469;
   wire n_0_0_470;
   wire n_0_0_471;
   wire n_0_111;
   wire n_0_112;

   assign Q[15] = 1'b0;
   assign Q[13] = Q[14];

   INV_X1 csa0_i_10 (.A(divisor[13]), .ZN(csa0_n_0));
   INV_X1 csa0_i_11 (.A(divisor[14]), .ZN(csa0_n_1));
   INV_X1 csa1_i_10 (.A(dividend[13]), .ZN(csa1_n_0));
   DFF_X1 divideByZero_reg (.D(n_0_113), .CK(n_0_6), .Q(divideByZero), .QN());
   DFF_X1 overFlow_reg (.D(n_0_111), .CK(clk), .Q(overFlow), .QN());
   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_0_110), .SE(1'b0), .GCK(n_0_0));
   DFF_X1 \Q_reg[14]  (.D(n_0_20), .CK(n_0_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_0_73), .CK(n_0_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_0_72), .CK(n_0_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_0_71), .CK(n_0_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_0_70), .CK(n_0_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_0_69), .CK(n_0_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_0_68), .CK(n_0_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_0_67), .CK(n_0_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_0_66), .CK(n_0_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_0_65), .CK(n_0_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_0_64), .CK(n_0_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_0_63), .CK(n_0_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_0_62), .CK(n_0_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0_61), .CK(n_0_0), .Q(Q[0]), .QN());
   CLKGATETST_X1 clk_gate_A_reg (.CK(clk), .E(n_0_109), .SE(1'b0), .GCK(n_0_1));
   DFF_X1 \A_reg[31]  (.D(n_0_107), .CK(n_0_1), .Q(n_0_21), .QN());
   DFF_X1 \A_reg[30]  (.D(n_0_106), .CK(n_0_1), .Q(n_0_22), .QN());
   DFF_X1 \A_reg[29]  (.D(n_0_105), .CK(n_0_1), .Q(n_0_23), .QN());
   DFF_X1 \A_reg[28]  (.D(n_0_104), .CK(n_0_1), .Q(n_0_24), .QN());
   DFF_X1 \A_reg[27]  (.D(n_0_103), .CK(n_0_1), .Q(n_0_25), .QN());
   DFF_X1 \A_reg[26]  (.D(n_0_102), .CK(n_0_1), .Q(n_0_26), .QN());
   DFF_X1 \A_reg[25]  (.D(n_0_101), .CK(n_0_1), .Q(n_0_27), .QN());
   DFF_X1 \A_reg[24]  (.D(n_0_100), .CK(n_0_1), .Q(n_0_28), .QN());
   DFF_X1 \A_reg[23]  (.D(n_0_99), .CK(n_0_1), .Q(n_0_29), .QN());
   DFF_X1 \A_reg[22]  (.D(n_0_98), .CK(n_0_1), .Q(n_0_30), .QN());
   DFF_X1 \A_reg[21]  (.D(n_0_97), .CK(n_0_1), .Q(n_0_31), .QN());
   DFF_X1 \A_reg[20]  (.D(n_0_96), .CK(n_0_1), .Q(n_0_32), .QN());
   DFF_X1 \A_reg[19]  (.D(n_0_95), .CK(n_0_1), .Q(n_0_33), .QN());
   DFF_X1 \A_reg[18]  (.D(n_0_94), .CK(n_0_1), .Q(n_0_34), .QN());
   DFF_X1 \A_reg[17]  (.D(n_0_93), .CK(n_0_1), .Q(n_0_35), .QN());
   DFF_X1 \A_reg[16]  (.D(n_0_92), .CK(n_0_1), .Q(n_0_36), .QN());
   CLKGATETST_X1 clk_gate_A_reg__15 (.CK(clk), .E(n_0_108), .SE(1'b0), .GCK(
      n_0_2));
   DFF_X1 \A_reg[15]  (.D(n_0_91), .CK(n_0_2), .Q(n_0_37), .QN());
   DFF_X1 \A_reg[14]  (.D(n_0_90), .CK(n_0_2), .Q(n_0_38), .QN());
   DFF_X1 \A_reg[13]  (.D(n_0_89), .CK(n_0_2), .Q(n_0_39), .QN());
   DFF_X1 \A_reg[12]  (.D(n_0_88), .CK(n_0_2), .Q(n_0_40), .QN());
   DFF_X1 \A_reg[11]  (.D(n_0_87), .CK(n_0_2), .Q(n_0_41), .QN());
   DFF_X1 \A_reg[10]  (.D(n_0_86), .CK(n_0_2), .Q(n_0_42), .QN());
   DFF_X1 \A_reg[9]  (.D(n_0_85), .CK(n_0_2), .Q(n_0_43), .QN());
   DFF_X1 \A_reg[8]  (.D(n_0_84), .CK(n_0_2), .Q(n_0_44), .QN());
   DFF_X1 \A_reg[7]  (.D(n_0_83), .CK(n_0_2), .Q(n_0_45), .QN());
   DFF_X1 \A_reg[6]  (.D(n_0_82), .CK(n_0_2), .Q(n_0_46), .QN());
   DFF_X1 \A_reg[5]  (.D(n_0_81), .CK(n_0_2), .Q(n_0_47), .QN());
   DFF_X1 \A_reg[4]  (.D(n_0_80), .CK(n_0_2), .Q(n_0_48), .QN());
   DFF_X1 \A_reg[3]  (.D(n_0_79), .CK(n_0_2), .Q(n_0_49), .QN());
   DFF_X1 \A_reg[2]  (.D(n_0_78), .CK(n_0_2), .Q(n_0_50), .QN());
   DFF_X1 \A_reg[1]  (.D(n_0_77), .CK(n_0_2), .Q(n_0_51), .QN());
   DFF_X1 \A_reg[0]  (.D(n_0_76), .CK(n_0_2), .Q(n_0_52), .QN());
   DFF_X1 \negated_second_operand_number_reg[15]  (.D(n_0_19), .CK(n_0_6), 
      .Q(negated_second_operand_number[15]), .QN());
   DFF_X1 \negated_second_operand_number_reg[14]  (.D(n_0_18), .CK(n_0_6), 
      .Q(negated_second_operand_number[14]), .QN());
   DFF_X1 \negated_second_operand_number_reg[13]  (.D(n_0_17), .CK(n_0_6), 
      .Q(negated_second_operand_number[13]), .QN());
   DFF_X1 \negated_second_operand_number_reg[12]  (.D(n_0_16), .CK(n_0_6), 
      .Q(negated_second_operand_number[12]), .QN());
   DFF_X1 \negated_second_operand_number_reg[11]  (.D(n_0_15), .CK(n_0_6), 
      .Q(negated_second_operand_number[11]), .QN());
   DFF_X1 \negated_second_operand_number_reg[10]  (.D(n_0_14), .CK(n_0_6), 
      .Q(negated_second_operand_number[10]), .QN());
   DFF_X1 \negated_second_operand_number_reg[9]  (.D(n_0_13), .CK(n_0_6), 
      .Q(negated_second_operand_number[9]), .QN());
   DFF_X1 \negated_second_operand_number_reg[8]  (.D(n_0_12), .CK(n_0_6), 
      .Q(negated_second_operand_number[8]), .QN());
   DFF_X1 \negated_second_operand_number_reg[7]  (.D(n_0_11), .CK(n_0_6), 
      .Q(negated_second_operand_number[7]), .QN());
   DFF_X1 \negated_second_operand_number_reg[6]  (.D(n_0_10), .CK(n_0_6), 
      .Q(negated_second_operand_number[6]), .QN());
   DFF_X1 \negated_second_operand_number_reg[5]  (.D(n_0_9), .CK(n_0_6), 
      .Q(negated_second_operand_number[5]), .QN());
   DFF_X1 \negated_second_operand_number_reg[4]  (.D(n_0_8), .CK(n_0_6), 
      .Q(negated_second_operand_number[4]), .QN());
   DFF_X1 \negated_second_operand_number_reg[3]  (.D(n_0_7), .CK(n_0_6), 
      .Q(negated_second_operand_number[3]), .QN());
   DFF_X1 \negated_second_operand_number_reg[2]  (.D(n_0_5), .CK(n_0_6), 
      .Q(negated_second_operand_number[2]), .QN());
   DFF_X1 \negated_second_operand_number_reg[1]  (.D(n_0_4), .CK(n_0_6), 
      .Q(negated_second_operand_number[1]), .QN());
   DFF_X1 \second_operand_number_reg[15]  (.D(n_0_129), .CK(n_0_6), .Q(
      second_operand_number[15]), .QN());
   DFF_X1 \second_operand_number_reg[14]  (.D(n_0_128), .CK(n_0_6), .Q(
      second_operand_number[14]), .QN());
   DFF_X1 \second_operand_number_reg[13]  (.D(n_0_127), .CK(n_0_6), .Q(
      second_operand_number[13]), .QN());
   DFF_X1 \second_operand_number_reg[12]  (.D(n_0_126), .CK(n_0_6), .Q(
      second_operand_number[12]), .QN());
   DFF_X1 \second_operand_number_reg[11]  (.D(n_0_125), .CK(n_0_6), .Q(
      second_operand_number[11]), .QN());
   DFF_X1 \second_operand_number_reg[10]  (.D(n_0_124), .CK(n_0_6), .Q(
      second_operand_number[10]), .QN());
   DFF_X1 \second_operand_number_reg[9]  (.D(n_0_123), .CK(n_0_6), .Q(
      second_operand_number[9]), .QN());
   DFF_X1 \second_operand_number_reg[8]  (.D(n_0_122), .CK(n_0_6), .Q(
      second_operand_number[8]), .QN());
   DFF_X1 \second_operand_number_reg[7]  (.D(n_0_121), .CK(n_0_6), .Q(
      second_operand_number[7]), .QN());
   DFF_X1 \second_operand_number_reg[6]  (.D(n_0_120), .CK(n_0_6), .Q(
      second_operand_number[6]), .QN());
   DFF_X1 \second_operand_number_reg[5]  (.D(n_0_119), .CK(n_0_6), .Q(
      second_operand_number[5]), .QN());
   DFF_X1 \second_operand_number_reg[4]  (.D(n_0_118), .CK(n_0_6), .Q(
      second_operand_number[4]), .QN());
   DFF_X1 \second_operand_number_reg[3]  (.D(n_0_117), .CK(n_0_6), .Q(
      second_operand_number[3]), .QN());
   DFF_X1 \second_operand_number_reg[2]  (.D(n_0_116), .CK(n_0_6), .Q(
      second_operand_number[2]), .QN());
   DFF_X1 \second_operand_number_reg[1]  (.D(n_0_115), .CK(n_0_6), .Q(
      second_operand_number[1]), .QN());
   DFF_X1 ready_reg (.D(n_0_112), .CK(clk), .Q(ready), .QN());
   CLKGATETST_X1 clk_gate_number_of_bits_in_dividend_reg (.CK(clk), .E(n_0_60), 
      .SE(1'b0), .GCK(n_0_3));
   DFF_X1 \number_of_bits_in_dividend_reg[4]  (.D(n_0_59), .CK(n_0_3), .Q(
      number_of_bits_in_dividend[4]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[3]  (.D(n_0_58), .CK(n_0_3), .Q(
      number_of_bits_in_dividend[3]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[2]  (.D(n_0_57), .CK(n_0_3), .Q(
      number_of_bits_in_dividend[2]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[1]  (.D(n_0_56), .CK(n_0_3), .Q(
      number_of_bits_in_dividend[1]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[0]  (.D(n_0_55), .CK(n_0_3), .Q(
      number_of_bits_in_dividend[0]), .QN());
   DFF_X1 sign_reg (.D(n_0_54), .CK(n_0_6), .Q(sign), .QN());
   CLKGATETST_X1 clk_gate_divideByZero_reg (.CK(clk), .E(reset), .SE(1'b0), 
      .GCK(n_0_6));
   DFF_X1 \negated_second_operand_number_reg[0]  (.D(n_0_114), .CK(n_0_6), 
      .Q(negated_second_operand_number[0]), .QN());
   OAI22_X1 i_0_0_0 (.A1(divisor[12]), .A2(n_0_0_449), .B1(n_0_0_479), .B2(
      dividend[12]), .ZN(n_0_54));
   NAND2_X1 i_0_0_1 (.A1(n_0_20), .A2(number_of_bits_in_dividend[0]), .ZN(n_0_55));
   OAI21_X1 i_0_0_2 (.A(n_0_0_0), .B1(number_of_bits_in_dividend[1]), .B2(
      number_of_bits_in_dividend[0]), .ZN(n_0_56));
   AOI21_X1 i_0_0_3 (.A(reset), .B1(number_of_bits_in_dividend[1]), .B2(
      number_of_bits_in_dividend[0]), .ZN(n_0_0_0));
   NAND3_X1 i_0_0_4 (.A1(n_0_20), .A2(n_0_0_6), .A3(n_0_0_1), .ZN(n_0_57));
   OAI21_X1 i_0_0_5 (.A(number_of_bits_in_dividend[2]), .B1(
      number_of_bits_in_dividend[1]), .B2(number_of_bits_in_dividend[0]), 
      .ZN(n_0_0_1));
   INV_X1 i_0_0_6 (.A(n_0_0_2), .ZN(n_0_58));
   AOI211_X1 i_0_0_7 (.A(reset), .B(n_0_0_5), .C1(number_of_bits_in_dividend[3]), 
      .C2(n_0_0_6), .ZN(n_0_0_2));
   NOR2_X1 i_0_0_11 (.A1(number_of_bits_in_dividend[3]), .A2(n_0_0_6), .ZN(
      n_0_0_5));
   OR3_X1 i_0_0_12 (.A1(number_of_bits_in_dividend[1]), .A2(
      number_of_bits_in_dividend[0]), .A3(number_of_bits_in_dividend[2]), 
      .ZN(n_0_0_6));
   AND2_X1 i_0_0_13 (.A1(n_0_52), .A2(n_0_20), .ZN(n_0_61));
   AND2_X1 i_0_0_14 (.A1(n_0_20), .A2(n_0_0_13), .ZN(n_0_62));
   AND2_X1 i_0_0_15 (.A1(n_0_20), .A2(n_0_0_15), .ZN(n_0_63));
   AND2_X1 i_0_0_16 (.A1(n_0_20), .A2(n_0_0_17), .ZN(n_0_64));
   AND2_X1 i_0_0_17 (.A1(n_0_20), .A2(n_0_0_19), .ZN(n_0_65));
   AND2_X1 i_0_0_18 (.A1(n_0_20), .A2(n_0_0_22), .ZN(n_0_66));
   AND2_X1 i_0_0_19 (.A1(n_0_20), .A2(n_0_0_29), .ZN(n_0_67));
   AND2_X1 i_0_0_20 (.A1(n_0_20), .A2(n_0_0_34), .ZN(n_0_68));
   AND2_X1 i_0_0_21 (.A1(n_0_20), .A2(n_0_0_40), .ZN(n_0_69));
   AND2_X1 i_0_0_22 (.A1(n_0_20), .A2(n_0_0_46), .ZN(n_0_70));
   AND2_X1 i_0_0_23 (.A1(n_0_20), .A2(n_0_0_52), .ZN(n_0_71));
   AND2_X1 i_0_0_24 (.A1(n_0_20), .A2(n_0_0_60), .ZN(n_0_72));
   AND2_X1 i_0_0_25 (.A1(n_0_20), .A2(n_0_0_74), .ZN(n_0_73));
   OAI21_X1 i_0_0_26 (.A(n_0_0_11), .B1(n_0_0_281), .B2(n_0_0_7), .ZN(n_0_76));
   AOI22_X1 i_0_0_27 (.A1(n_0_0_472), .A2(n_0_0_9), .B1(n_0_21), .B2(n_0_0_258), 
      .ZN(n_0_0_7));
   XNOR2_X1 i_0_0_28 (.A(negated_second_operand_number[15]), .B(n_0_0_10), 
      .ZN(n_0_0_9));
   OAI21_X1 i_0_0_29 (.A(n_0_0_213), .B1(n_0_0_444), .B2(n_0_0_212), .ZN(
      n_0_0_10));
   NAND2_X1 i_0_0_30 (.A1(n_0_52), .A2(n_0_0_282), .ZN(n_0_0_11));
   INV_X1 i_0_0_31 (.A(n_0_0_12), .ZN(n_0_77));
   AOI22_X1 i_0_0_32 (.A1(n_0_0_282), .A2(n_0_0_13), .B1(n_0_52), .B2(n_0_0_280), 
      .ZN(n_0_0_12));
   XNOR2_X1 i_0_0_33 (.A(n_0_51), .B(n_0_0_81), .ZN(n_0_0_13));
   OAI21_X1 i_0_0_34 (.A(n_0_0_14), .B1(n_0_0_452), .B2(n_0_0_281), .ZN(n_0_78));
   NAND2_X1 i_0_0_35 (.A1(n_0_0_282), .A2(n_0_0_15), .ZN(n_0_0_14));
   XOR2_X1 i_0_0_36 (.A(n_0_50), .B(n_0_0_80), .Z(n_0_0_15));
   INV_X1 i_0_0_37 (.A(n_0_0_16), .ZN(n_0_79));
   AOI22_X1 i_0_0_38 (.A1(n_0_50), .A2(n_0_0_280), .B1(n_0_0_282), .B2(n_0_0_17), 
      .ZN(n_0_0_16));
   XNOR2_X1 i_0_0_39 (.A(n_0_49), .B(n_0_0_79), .ZN(n_0_0_17));
   INV_X1 i_0_0_40 (.A(n_0_0_18), .ZN(n_0_80));
   AOI221_X1 i_0_0_41 (.A(n_0_0_20), .B1(n_0_49), .B2(n_0_0_280), .C1(n_0_0_282), 
      .C2(n_0_0_19), .ZN(n_0_0_18));
   XOR2_X1 i_0_0_42 (.A(n_0_48), .B(n_0_0_71), .Z(n_0_0_19));
   NOR3_X1 i_0_0_43 (.A1(n_0_0_445), .A2(n_0_20), .A3(n_0_0_142), .ZN(n_0_0_20));
   INV_X1 i_0_0_44 (.A(n_0_0_21), .ZN(n_0_81));
   AOI222_X1 i_0_0_45 (.A1(n_0_0_282), .A2(n_0_0_22), .B1(n_0_48), .B2(n_0_0_280), 
      .C1(reset), .C2(n_0_0_23), .ZN(n_0_0_21));
   XNOR2_X1 i_0_0_46 (.A(n_0_47), .B(n_0_0_251), .ZN(n_0_0_22));
   OAI22_X1 i_0_0_47 (.A1(n_0_0_142), .A2(n_0_0_68), .B1(n_0_0_445), .B2(
      n_0_0_24), .ZN(n_0_0_23));
   NAND2_X1 i_0_0_48 (.A1(n_0_0_393), .A2(n_0_0_28), .ZN(n_0_0_24));
   INV_X1 i_0_0_49 (.A(n_0_0_25), .ZN(n_0_82));
   AOI221_X1 i_0_0_50 (.A(n_0_0_26), .B1(n_0_47), .B2(n_0_0_280), .C1(n_0_0_282), 
      .C2(n_0_0_29), .ZN(n_0_0_25));
   AOI211_X1 i_0_0_51 (.A(n_0_20), .B(n_0_0_27), .C1(n_0_0_141), .C2(n_0_0_88), 
      .ZN(n_0_0_26));
   AOI221_X1 i_0_0_52 (.A(n_0_0_141), .B1(n_0_0_153), .B2(n_0_0_33), .C1(
      n_0_0_67), .C2(n_0_0_28), .ZN(n_0_0_27));
   AND2_X1 i_0_0_53 (.A1(n_0_0_152), .A2(n_0_0_143), .ZN(n_0_0_28));
   XOR2_X1 i_0_0_54 (.A(n_0_46), .B(n_0_0_250), .Z(n_0_0_29));
   INV_X1 i_0_0_55 (.A(n_0_0_30), .ZN(n_0_83));
   AOI221_X1 i_0_0_56 (.A(n_0_0_31), .B1(n_0_46), .B2(n_0_0_280), .C1(n_0_0_282), 
      .C2(n_0_0_34), .ZN(n_0_0_30));
   AOI211_X1 i_0_0_57 (.A(n_0_20), .B(n_0_0_32), .C1(n_0_0_141), .C2(n_0_0_97), 
      .ZN(n_0_0_31));
   AOI221_X1 i_0_0_58 (.A(n_0_0_141), .B1(n_0_0_152), .B2(n_0_0_33), .C1(
      n_0_0_153), .C2(n_0_0_38), .ZN(n_0_0_32));
   AND2_X1 i_0_0_59 (.A1(n_0_0_144), .A2(n_0_0_58), .ZN(n_0_0_33));
   XNOR2_X1 i_0_0_60 (.A(n_0_45), .B(n_0_0_248), .ZN(n_0_0_34));
   INV_X1 i_0_0_61 (.A(n_0_0_35), .ZN(n_0_84));
   AOI221_X1 i_0_0_62 (.A(n_0_0_36), .B1(n_0_45), .B2(n_0_0_280), .C1(n_0_0_282), 
      .C2(n_0_0_40), .ZN(n_0_0_35));
   AOI211_X1 i_0_0_63 (.A(n_0_20), .B(n_0_0_37), .C1(n_0_0_141), .C2(n_0_0_104), 
      .ZN(n_0_0_36));
   AOI221_X1 i_0_0_64 (.A(n_0_0_141), .B1(n_0_0_153), .B2(n_0_0_44), .C1(
      n_0_0_152), .C2(n_0_0_38), .ZN(n_0_0_37));
   OAI21_X1 i_0_0_65 (.A(n_0_0_39), .B1(n_0_0_68), .B2(n_0_0_59), .ZN(n_0_0_38));
   NAND2_X1 i_0_0_66 (.A1(n_0_0_143), .A2(n_0_0_96), .ZN(n_0_0_39));
   XOR2_X1 i_0_0_67 (.A(n_0_44), .B(n_0_0_246), .Z(n_0_0_40));
   INV_X1 i_0_0_68 (.A(n_0_0_41), .ZN(n_0_85));
   AOI221_X1 i_0_0_69 (.A(n_0_0_42), .B1(n_0_44), .B2(n_0_0_280), .C1(n_0_0_282), 
      .C2(n_0_0_46), .ZN(n_0_0_41));
   AOI211_X1 i_0_0_70 (.A(n_0_20), .B(n_0_0_43), .C1(n_0_0_141), .C2(n_0_0_115), 
      .ZN(n_0_0_42));
   AOI221_X1 i_0_0_71 (.A(n_0_0_141), .B1(n_0_0_153), .B2(n_0_0_50), .C1(
      n_0_0_152), .C2(n_0_0_44), .ZN(n_0_0_43));
   OAI21_X1 i_0_0_72 (.A(n_0_0_45), .B1(n_0_0_88), .B2(n_0_0_59), .ZN(n_0_0_44));
   AOI22_X1 i_0_0_73 (.A1(n_0_0_143), .A2(n_0_0_103), .B1(dividend[0]), .B2(
      n_0_0_140), .ZN(n_0_0_45));
   XNOR2_X1 i_0_0_74 (.A(n_0_43), .B(n_0_0_78), .ZN(n_0_0_46));
   INV_X1 i_0_0_75 (.A(n_0_0_47), .ZN(n_0_86));
   AOI221_X1 i_0_0_76 (.A(n_0_0_48), .B1(n_0_43), .B2(n_0_0_280), .C1(n_0_0_282), 
      .C2(n_0_0_52), .ZN(n_0_0_47));
   AOI211_X1 i_0_0_77 (.A(n_0_20), .B(n_0_0_49), .C1(n_0_0_141), .C2(n_0_0_125), 
      .ZN(n_0_0_48));
   AOI221_X1 i_0_0_78 (.A(n_0_0_141), .B1(n_0_0_152), .B2(n_0_0_50), .C1(
      n_0_0_153), .C2(n_0_0_56), .ZN(n_0_0_49));
   OAI21_X1 i_0_0_79 (.A(n_0_0_51), .B1(n_0_0_97), .B2(n_0_0_59), .ZN(n_0_0_50));
   NAND2_X1 i_0_0_80 (.A1(n_0_0_149), .A2(n_0_0_66), .ZN(n_0_0_51));
   XOR2_X1 i_0_0_81 (.A(n_0_42), .B(n_0_0_77), .Z(n_0_0_52));
   INV_X1 i_0_0_83 (.A(n_0_0_53), .ZN(n_0_87));
   AOI221_X1 i_0_0_84 (.A(n_0_0_54), .B1(n_0_42), .B2(n_0_0_280), .C1(n_0_0_282), 
      .C2(n_0_0_60), .ZN(n_0_0_53));
   AOI211_X1 i_0_0_85 (.A(n_0_20), .B(n_0_0_55), .C1(n_0_0_141), .C2(n_0_0_112), 
      .ZN(n_0_0_54));
   AOI221_X1 i_0_0_86 (.A(n_0_0_141), .B1(n_0_0_153), .B2(n_0_0_64), .C1(
      n_0_0_152), .C2(n_0_0_56), .ZN(n_0_0_55));
   OAI21_X1 i_0_0_82 (.A(n_0_0_57), .B1(n_0_0_104), .B2(n_0_0_59), .ZN(n_0_0_56));
   AOI22_X1 i_0_0_87 (.A1(n_0_0_143), .A2(n_0_0_124), .B1(n_0_0_145), .B2(
      n_0_0_58), .ZN(n_0_0_57));
   OAI22_X1 i_0_0_88 (.A1(n_0_0_445), .A2(n_0_0_149), .B1(n_0_0_148), .B2(
      n_0_0_88), .ZN(n_0_0_58));
   NAND2_X1 i_0_0_89 (.A1(n_0_0_148), .A2(n_0_0_144), .ZN(n_0_0_59));
   XNOR2_X1 i_0_0_90 (.A(n_0_41), .B(n_0_0_76), .ZN(n_0_0_60));
   NOR2_X1 i_0_0_97 (.A1(n_0_0_149), .A2(n_0_0_66), .ZN(n_0_0_65));
   OAI22_X1 i_0_0_91 (.A1(n_0_0_144), .A2(n_0_0_68), .B1(n_0_0_145), .B2(
      n_0_0_115), .ZN(n_0_0_66));
   INV_X1 i_0_0_92 (.A(n_0_0_68), .ZN(n_0_0_67));
   XNOR2_X1 i_0_0_95 (.A(dividend[1]), .B(n_0_0_139), .ZN(n_0_0_68));
   AOI21_X1 i_0_0_96 (.A(n_0_0_257), .B1(n_0_0_453), .B2(n_0_0_79), .ZN(n_0_0_71));
   OAI21_X1 i_0_0_98 (.A(sign), .B1(n_0_50), .B2(n_0_0_80), .ZN(n_0_0_79));
   AOI21_X1 i_0_0_99 (.A(n_0_0_257), .B1(n_0_0_452), .B2(n_0_0_81), .ZN(n_0_0_80));
   NAND2_X1 i_0_0_100 (.A1(n_0_52), .A2(sign), .ZN(n_0_0_81));
   OAI221_X1 i_0_0_101 (.A(n_0_0_283), .B1(n_0_0_256), .B2(n_0_0_281), .C1(
      n_0_0_84), .C2(n_0_0_82), .ZN(n_0_89));
   INV_X1 i_0_0_102 (.A(n_0_0_83), .ZN(n_0_0_82));
   AOI21_X1 i_0_0_103 (.A(n_0_20), .B1(n_0_0_141), .B2(n_0_0_116), .ZN(n_0_0_83));
   AOI221_X1 i_0_0_104 (.A(n_0_0_141), .B1(n_0_0_153), .B2(n_0_0_92), .C1(
      n_0_0_152), .C2(n_0_0_85), .ZN(n_0_0_84));
   OAI21_X1 i_0_0_122 (.A(n_0_0_89), .B1(n_0_20), .B2(n_0_0_90), .ZN(n_0_90));
   AOI21_X1 i_0_0_123 (.A(n_0_0_282), .B1(n_0_39), .B2(n_0_0_280), .ZN(n_0_0_89));
   AOI21_X1 i_0_0_124 (.A(n_0_0_91), .B1(n_0_0_141), .B2(n_0_0_121), .ZN(
      n_0_0_90));
   AOI221_X1 i_0_0_125 (.A(n_0_0_141), .B1(n_0_0_153), .B2(n_0_0_100), .C1(
      n_0_0_152), .C2(n_0_0_93), .ZN(n_0_0_91));
   INV_X1 i_0_0_105 (.A(n_0_0_93), .ZN(n_0_0_92));
   OAI21_X1 i_0_0_106 (.A(n_0_0_94), .B1(n_0_0_148), .B2(n_0_0_114), .ZN(
      n_0_0_93));
   NAND2_X1 i_0_0_107 (.A1(n_0_0_148), .A2(n_0_0_95), .ZN(n_0_0_94));
   OAI22_X1 i_0_0_108 (.A1(n_0_0_145), .A2(n_0_0_113), .B1(n_0_0_144), .B2(
      n_0_0_96), .ZN(n_0_0_95));
   INV_X1 i_0_0_109 (.A(n_0_0_97), .ZN(n_0_0_96));
   XNOR2_X1 i_0_0_110 (.A(dividend[3]), .B(n_0_0_135), .ZN(n_0_0_97));
   NOR2_X1 i_0_0_136 (.A1(n_0_0_148), .A2(n_0_0_120), .ZN(n_0_0_101));
   INV_X1 i_0_0_111 (.A(n_0_0_104), .ZN(n_0_0_103));
   INV_X1 i_0_0_148 (.A(n_0_0_113), .ZN(n_0_0_112));
   AOI22_X1 i_0_0_112 (.A1(n_0_0_144), .A2(n_0_0_121), .B1(n_0_0_145), .B2(
      n_0_0_124), .ZN(n_0_0_120));
   XOR2_X1 i_0_0_113 (.A(dividend[10]), .B(n_0_0_122), .Z(n_0_0_121));
   INV_X1 i_0_0_114 (.A(n_0_0_125), .ZN(n_0_0_124));
   OAI22_X1 i_0_0_115 (.A1(divisor[15]), .A2(n_0_0_451), .B1(n_0_0_480), 
      .B2(dividend[15]), .ZN(n_0_0_146));
   OAI21_X1 i_0_0_116 (.A(n_0_0_151), .B1(n_0_0_154), .B2(n_0_0_150), .ZN(
      n_0_0_147));
   OAI21_X1 i_0_0_117 (.A(n_0_0_151), .B1(divisor[14]), .B2(n_0_0_450), .ZN(
      n_0_0_150));
   NAND2_X1 i_0_0_118 (.A1(divisor[14]), .A2(n_0_0_450), .ZN(n_0_0_151));
   NOR2_X1 i_0_0_119 (.A1(divisor[13]), .A2(csa1_n_0), .ZN(n_0_0_154));
   OAI21_X1 i_0_0_120 (.A(n_0_0_155), .B1(n_0_0_460), .B2(n_0_0_286), .ZN(n_0_93));
   OAI211_X1 i_0_0_121 (.A(n_0_0_270), .B(n_0_0_280), .C1(n_0_36), .C2(
      negated_second_operand_number[0]), .ZN(n_0_0_155));
   OAI21_X1 i_0_0_126 (.A(n_0_0_156), .B1(n_0_0_461), .B2(n_0_0_286), .ZN(n_0_94));
   NAND2_X1 i_0_0_127 (.A1(n_0_0_280), .A2(n_0_0_157), .ZN(n_0_0_156));
   XNOR2_X1 i_0_0_128 (.A(n_0_0_159), .B(n_0_0_158), .ZN(n_0_0_157));
   AOI22_X1 i_0_0_129 (.A1(n_0_0_472), .A2(negated_second_operand_number[1]), 
      .B1(n_0_21), .B2(second_operand_number[1]), .ZN(n_0_0_158));
   AOI22_X1 i_0_0_130 (.A1(n_0_35), .A2(n_0_0_269), .B1(n_0_0_459), .B2(
      n_0_0_270), .ZN(n_0_0_159));
   OAI21_X1 i_0_0_131 (.A(n_0_0_160), .B1(n_0_0_462), .B2(n_0_0_286), .ZN(n_0_95));
   AOI22_X1 i_0_0_132 (.A1(n_0_0_278), .A2(n_0_0_162), .B1(n_0_0_209), .B2(
      n_0_0_161), .ZN(n_0_0_160));
   XOR2_X1 i_0_0_133 (.A(n_0_0_237), .B(n_0_0_235), .Z(n_0_0_161));
   XOR2_X1 i_0_0_134 (.A(n_0_0_267), .B(n_0_0_163), .Z(n_0_0_162));
   AOI22_X1 i_0_0_135 (.A1(n_0_0_460), .A2(n_0_0_426), .B1(n_0_34), .B2(
      second_operand_number[2]), .ZN(n_0_0_163));
   OAI21_X1 i_0_0_203 (.A(n_0_0_164), .B1(n_0_0_463), .B2(n_0_0_286), .ZN(n_0_96));
   AOI22_X1 i_0_0_204 (.A1(n_0_0_278), .A2(n_0_0_166), .B1(n_0_0_209), .B2(
      n_0_0_165), .ZN(n_0_0_164));
   XOR2_X1 i_0_0_205 (.A(n_0_0_234), .B(n_0_0_233), .Z(n_0_0_165));
   XOR2_X1 i_0_0_206 (.A(n_0_0_271), .B(n_0_0_265), .Z(n_0_0_166));
   OAI21_X1 i_0_0_207 (.A(n_0_0_167), .B1(n_0_0_464), .B2(n_0_0_286), .ZN(n_0_97));
   AOI22_X1 i_0_0_208 (.A1(n_0_0_278), .A2(n_0_0_170), .B1(n_0_0_209), .B2(
      n_0_0_168), .ZN(n_0_0_167));
   XNOR2_X1 i_0_0_209 (.A(n_0_0_232), .B(n_0_0_169), .ZN(n_0_0_168));
   OAI22_X1 i_0_0_210 (.A1(n_0_32), .A2(negated_second_operand_number[4]), 
      .B1(n_0_0_462), .B2(n_0_0_436), .ZN(n_0_0_169));
   XOR2_X1 i_0_0_211 (.A(n_0_0_264), .B(n_0_0_171), .Z(n_0_0_170));
   OAI22_X1 i_0_0_212 (.A1(n_0_32), .A2(second_operand_number[4]), .B1(n_0_0_462), 
      .B2(n_0_0_427), .ZN(n_0_0_171));
   OAI21_X1 i_0_0_213 (.A(n_0_0_172), .B1(n_0_0_465), .B2(n_0_0_286), .ZN(n_0_98));
   AOI22_X1 i_0_0_214 (.A1(n_0_0_278), .A2(n_0_0_174), .B1(n_0_0_209), .B2(
      n_0_0_173), .ZN(n_0_0_172));
   XOR2_X1 i_0_0_215 (.A(n_0_0_239), .B(n_0_0_230), .Z(n_0_0_173));
   XNOR2_X1 i_0_0_216 (.A(n_0_0_262), .B(n_0_0_175), .ZN(n_0_0_174));
   AOI22_X1 i_0_0_217 (.A1(n_0_0_463), .A2(n_0_0_428), .B1(n_0_31), .B2(
      second_operand_number[5]), .ZN(n_0_0_175));
   OAI21_X1 i_0_0_218 (.A(n_0_0_176), .B1(n_0_0_466), .B2(n_0_0_286), .ZN(n_0_99));
   AOI22_X1 i_0_0_219 (.A1(n_0_0_278), .A2(n_0_0_179), .B1(n_0_0_209), .B2(
      n_0_0_177), .ZN(n_0_0_176));
   XNOR2_X1 i_0_0_220 (.A(n_0_0_229), .B(n_0_0_178), .ZN(n_0_0_177));
   AOI22_X1 i_0_0_221 (.A1(n_0_0_464), .A2(n_0_0_437), .B1(n_0_30), .B2(
      negated_second_operand_number[6]), .ZN(n_0_0_178));
   XOR2_X1 i_0_0_222 (.A(n_0_0_273), .B(n_0_0_261), .Z(n_0_0_179));
   OAI21_X1 i_0_0_223 (.A(n_0_0_180), .B1(n_0_0_467), .B2(n_0_0_286), .ZN(
      n_0_100));
   AOI22_X1 i_0_0_224 (.A1(n_0_0_278), .A2(n_0_0_182), .B1(n_0_0_209), .B2(
      n_0_0_181), .ZN(n_0_0_180));
   XNOR2_X1 i_0_0_225 (.A(n_0_0_240), .B(n_0_0_227), .ZN(n_0_0_181));
   XNOR2_X1 i_0_0_226 (.A(n_0_0_260), .B(n_0_0_183), .ZN(n_0_0_182));
   AOI22_X1 i_0_0_227 (.A1(n_0_29), .A2(second_operand_number[7]), .B1(n_0_0_465), 
      .B2(n_0_0_429), .ZN(n_0_0_183));
   OAI21_X1 i_0_0_228 (.A(n_0_0_184), .B1(n_0_0_468), .B2(n_0_0_286), .ZN(
      n_0_101));
   AOI22_X1 i_0_0_229 (.A1(n_0_0_278), .A2(n_0_0_186), .B1(n_0_0_209), .B2(
      n_0_0_185), .ZN(n_0_0_184));
   XOR2_X1 i_0_0_230 (.A(n_0_0_241), .B(n_0_0_226), .Z(n_0_0_185));
   XNOR2_X1 i_0_0_231 (.A(n_0_0_433), .B(n_0_0_187), .ZN(n_0_0_186));
   AOI22_X1 i_0_0_232 (.A1(n_0_28), .A2(second_operand_number[8]), .B1(n_0_0_466), 
      .B2(n_0_0_455), .ZN(n_0_0_187));
   OAI21_X1 i_0_0_233 (.A(n_0_0_188), .B1(n_0_0_469), .B2(n_0_0_286), .ZN(
      n_0_102));
   AOI22_X1 i_0_0_234 (.A1(n_0_0_278), .A2(n_0_0_191), .B1(n_0_0_209), .B2(
      n_0_0_189), .ZN(n_0_0_188));
   XOR2_X1 i_0_0_235 (.A(n_0_0_224), .B(n_0_0_190), .Z(n_0_0_189));
   AOI22_X1 i_0_0_236 (.A1(n_0_27), .A2(negated_second_operand_number[9]), 
      .B1(n_0_0_467), .B2(n_0_0_440), .ZN(n_0_0_190));
   XOR2_X1 i_0_0_237 (.A(n_0_0_434), .B(n_0_0_431), .Z(n_0_0_191));
   OAI21_X1 i_0_0_238 (.A(n_0_0_192), .B1(n_0_0_470), .B2(n_0_0_286), .ZN(
      n_0_103));
   AOI22_X1 i_0_0_239 (.A1(n_0_0_278), .A2(n_0_0_195), .B1(n_0_0_209), .B2(
      n_0_0_193), .ZN(n_0_0_192));
   XNOR2_X1 i_0_0_240 (.A(n_0_0_223), .B(n_0_0_194), .ZN(n_0_0_193));
   AOI22_X1 i_0_0_241 (.A1(n_0_26), .A2(negated_second_operand_number[10]), 
      .B1(n_0_0_468), .B2(n_0_0_441), .ZN(n_0_0_194));
   XNOR2_X1 i_0_0_242 (.A(n_0_0_430), .B(n_0_0_196), .ZN(n_0_0_195));
   AOI22_X1 i_0_0_243 (.A1(n_0_0_468), .A2(n_0_0_456), .B1(n_0_26), .B2(
      second_operand_number[10]), .ZN(n_0_0_196));
   OAI21_X1 i_0_0_244 (.A(n_0_0_197), .B1(n_0_0_471), .B2(n_0_0_286), .ZN(
      n_0_104));
   AOI22_X1 i_0_0_138 (.A1(n_0_0_278), .A2(n_0_0_199), .B1(n_0_0_209), .B2(
      n_0_0_198), .ZN(n_0_0_197));
   XNOR2_X1 i_0_0_142 (.A(n_0_0_243), .B(n_0_0_221), .ZN(n_0_0_198));
   XNOR2_X1 i_0_0_143 (.A(n_0_0_318), .B(n_0_0_200), .ZN(n_0_0_199));
   AOI22_X1 i_0_0_152 (.A1(n_0_0_469), .A2(n_0_0_457), .B1(n_0_25), .B2(
      second_operand_number[11]), .ZN(n_0_0_200));
   INV_X1 i_0_0_153 (.A(n_0_0_201), .ZN(n_0_105));
   AOI221_X1 i_0_0_154 (.A(n_0_0_202), .B1(n_0_22), .B2(n_0_0_287), .C1(
      n_0_0_278), .C2(n_0_0_203), .ZN(n_0_0_201));
   AOI211_X1 i_0_0_156 (.A(n_0_0_217), .B(n_0_0_210), .C1(n_0_0_219), .C2(
      n_0_0_218), .ZN(n_0_0_202));
   XOR2_X1 i_0_0_157 (.A(n_0_0_454), .B(n_0_0_314), .Z(n_0_0_203));
   OAI21_X1 i_0_0_160 (.A(n_0_0_204), .B1(n_0_0_472), .B2(n_0_0_286), .ZN(
      n_0_106));
   AOI22_X1 i_0_0_162 (.A1(n_0_0_278), .A2(n_0_0_206), .B1(n_0_0_209), .B2(
      n_0_0_205), .ZN(n_0_0_204));
   XNOR2_X1 i_0_0_168 (.A(n_0_0_216), .B(n_0_0_215), .ZN(n_0_0_205));
   XNOR2_X1 i_0_0_170 (.A(n_0_0_313), .B(n_0_0_277), .ZN(n_0_0_206));
   NAND2_X1 i_0_0_257 (.A1(n_0_0_244), .A2(n_0_0_207), .ZN(n_0_107));
   OAI21_X1 i_0_0_258 (.A(n_0_0_208), .B1(n_0_0_444), .B2(n_0_0_211), .ZN(
      n_0_0_207));
   AOI21_X1 i_0_0_259 (.A(n_0_0_210), .B1(n_0_0_444), .B2(n_0_0_211), .ZN(
      n_0_0_208));
   INV_X1 i_0_0_171 (.A(n_0_0_210), .ZN(n_0_0_209));
   NAND2_X1 i_0_0_175 (.A1(n_0_0_472), .A2(n_0_0_280), .ZN(n_0_0_210));
   OAI21_X1 i_0_0_262 (.A(n_0_0_213), .B1(n_0_22), .B2(n_0_0_214), .ZN(n_0_0_211));
   NOR2_X1 i_0_0_176 (.A1(n_0_22), .A2(n_0_0_214), .ZN(n_0_0_212));
   NAND2_X1 i_0_0_177 (.A1(n_0_22), .A2(n_0_0_214), .ZN(n_0_0_213));
   AOI22_X1 i_0_0_182 (.A1(n_0_0_471), .A2(n_0_0_443), .B1(n_0_0_216), .B2(
      n_0_0_215), .ZN(n_0_0_214));
   AOI22_X1 i_0_0_183 (.A1(n_0_0_471), .A2(n_0_0_443), .B1(n_0_23), .B2(
      negated_second_operand_number[13]), .ZN(n_0_0_215));
   OAI22_X1 i_0_0_186 (.A1(n_0_24), .A2(n_0_0_220), .B1(
      negated_second_operand_number[12]), .B2(n_0_0_217), .ZN(n_0_0_216));
   NOR2_X1 i_0_0_187 (.A1(n_0_0_219), .A2(n_0_0_218), .ZN(n_0_0_217));
   XOR2_X1 i_0_0_188 (.A(n_0_0_470), .B(negated_second_operand_number[12]), 
      .Z(n_0_0_218));
   INV_X1 i_0_0_190 (.A(n_0_0_220), .ZN(n_0_0_219));
   AOI22_X1 i_0_0_191 (.A1(n_0_0_469), .A2(n_0_0_442), .B1(n_0_0_243), .B2(
      n_0_0_221), .ZN(n_0_0_220));
   OAI21_X1 i_0_0_192 (.A(n_0_0_222), .B1(n_0_26), .B2(
      negated_second_operand_number[10]), .ZN(n_0_0_221));
   OAI21_X1 i_0_0_193 (.A(n_0_0_223), .B1(n_0_0_468), .B2(n_0_0_441), .ZN(
      n_0_0_222));
   AOI22_X1 i_0_0_194 (.A1(n_0_27), .A2(negated_second_operand_number[9]), 
      .B1(n_0_0_242), .B2(n_0_0_224), .ZN(n_0_0_223));
   AOI22_X1 i_0_0_195 (.A1(n_0_0_466), .A2(n_0_0_439), .B1(n_0_0_241), .B2(
      n_0_0_225), .ZN(n_0_0_224));
   INV_X1 i_0_0_196 (.A(n_0_0_226), .ZN(n_0_0_225));
   AOI22_X1 i_0_0_197 (.A1(n_0_0_465), .A2(n_0_0_438), .B1(n_0_0_240), .B2(
      n_0_0_227), .ZN(n_0_0_226));
   AOI21_X1 i_0_0_198 (.A(n_0_0_228), .B1(n_0_30), .B2(
      negated_second_operand_number[6]), .ZN(n_0_0_227));
   AOI21_X1 i_0_0_199 (.A(n_0_0_229), .B1(n_0_0_464), .B2(n_0_0_437), .ZN(
      n_0_0_228));
   AOI22_X1 i_0_0_200 (.A1(n_0_31), .A2(negated_second_operand_number[5]), 
      .B1(n_0_0_239), .B2(n_0_0_230), .ZN(n_0_0_229));
   OAI21_X1 i_0_0_201 (.A(n_0_0_231), .B1(n_0_0_462), .B2(n_0_0_436), .ZN(
      n_0_0_230));
   OAI21_X1 i_0_0_282 (.A(n_0_0_232), .B1(n_0_32), .B2(
      negated_second_operand_number[4]), .ZN(n_0_0_231));
   OAI21_X1 i_0_0_283 (.A(n_0_0_238), .B1(n_0_0_234), .B2(n_0_0_233), .ZN(
      n_0_0_232));
   OAI21_X1 i_0_0_284 (.A(n_0_0_238), .B1(n_0_33), .B2(
      negated_second_operand_number[3]), .ZN(n_0_0_233));
   AOI22_X1 i_0_0_285 (.A1(n_0_34), .A2(negated_second_operand_number[2]), 
      .B1(n_0_0_237), .B2(n_0_0_235), .ZN(n_0_0_234));
   AOI21_X1 i_0_0_202 (.A(n_0_0_236), .B1(n_0_0_459), .B2(n_0_0_435), .ZN(
      n_0_0_235));
   AOI21_X1 i_0_0_245 (.A(n_0_0_269), .B1(n_0_35), .B2(
      negated_second_operand_number[1]), .ZN(n_0_0_236));
   XNOR2_X1 i_0_0_246 (.A(n_0_0_460), .B(negated_second_operand_number[2]), 
      .ZN(n_0_0_237));
   NAND2_X1 i_0_0_289 (.A1(n_0_33), .A2(negated_second_operand_number[3]), 
      .ZN(n_0_0_238));
   XNOR2_X1 i_0_0_247 (.A(n_0_0_463), .B(negated_second_operand_number[5]), 
      .ZN(n_0_0_239));
   AOI22_X1 i_0_0_248 (.A1(n_0_0_465), .A2(n_0_0_438), .B1(n_0_29), .B2(
      negated_second_operand_number[7]), .ZN(n_0_0_240));
   AOI22_X1 i_0_0_249 (.A1(n_0_0_466), .A2(n_0_0_439), .B1(n_0_28), .B2(
      negated_second_operand_number[8]), .ZN(n_0_0_241));
   NAND2_X1 i_0_0_250 (.A1(n_0_0_467), .A2(n_0_0_440), .ZN(n_0_0_242));
   AOI22_X1 i_0_0_251 (.A1(n_0_0_469), .A2(n_0_0_442), .B1(n_0_25), .B2(
      negated_second_operand_number[11]), .ZN(n_0_0_243));
   OAI21_X1 i_0_0_252 (.A(n_0_0_245), .B1(second_operand_number[14]), .B2(
      n_0_0_247), .ZN(n_0_0_244));
   AOI21_X1 i_0_0_253 (.A(n_0_0_279), .B1(second_operand_number[14]), .B2(
      n_0_0_247), .ZN(n_0_0_245));
   AOI21_X1 i_0_0_254 (.A(n_0_0_275), .B1(n_0_22), .B2(n_0_0_276), .ZN(n_0_0_247));
   OAI21_X1 i_0_0_255 (.A(n_0_0_260), .B1(n_0_0_465), .B2(n_0_0_429), .ZN(
      n_0_0_72));
   AOI22_X1 i_0_0_256 (.A1(n_0_30), .A2(second_operand_number[6]), .B1(n_0_0_273), 
      .B2(n_0_0_261), .ZN(n_0_0_260));
   AOI22_X1 i_0_0_260 (.A1(n_0_0_463), .A2(n_0_0_428), .B1(n_0_0_272), .B2(
      n_0_0_262), .ZN(n_0_0_261));
   AOI21_X1 i_0_0_261 (.A(n_0_0_263), .B1(n_0_32), .B2(second_operand_number[4]), 
      .ZN(n_0_0_262));
   AOI21_X1 i_0_0_263 (.A(n_0_0_264), .B1(n_0_0_462), .B2(n_0_0_427), .ZN(
      n_0_0_263));
   AOI22_X1 i_0_0_264 (.A1(n_0_33), .A2(second_operand_number[3]), .B1(n_0_0_271), 
      .B2(n_0_0_265), .ZN(n_0_0_264));
   OAI21_X1 i_0_0_265 (.A(n_0_0_266), .B1(n_0_0_460), .B2(n_0_0_426), .ZN(
      n_0_0_265));
   OAI21_X1 i_0_0_266 (.A(n_0_0_267), .B1(n_0_34), .B2(second_operand_number[2]), 
      .ZN(n_0_0_266));
   AOI21_X1 i_0_0_267 (.A(n_0_0_268), .B1(n_0_0_459), .B2(n_0_0_270), .ZN(
      n_0_0_267));
   AOI21_X1 i_0_0_268 (.A(second_operand_number[1]), .B1(n_0_35), .B2(n_0_0_269), 
      .ZN(n_0_0_268));
   INV_X1 i_0_0_269 (.A(n_0_0_270), .ZN(n_0_0_269));
   NAND2_X1 i_0_0_270 (.A1(n_0_36), .A2(negated_second_operand_number[0]), 
      .ZN(n_0_0_270));
   XNOR2_X1 i_0_0_271 (.A(n_0_0_461), .B(second_operand_number[3]), .ZN(
      n_0_0_271));
   NAND2_X1 i_0_0_272 (.A1(n_0_31), .A2(second_operand_number[5]), .ZN(n_0_0_272));
   XNOR2_X1 i_0_0_273 (.A(n_0_0_464), .B(second_operand_number[6]), .ZN(
      n_0_0_273));
   INV_X1 i_0_0_274 (.A(n_0_0_279), .ZN(n_0_0_278));
   NAND2_X1 i_0_0_275 (.A1(n_0_21), .A2(n_0_0_280), .ZN(n_0_0_279));
   NAND2_X1 i_0_0_276 (.A1(n_0_20), .A2(n_0_0_289), .ZN(n_0_0_281));
   AND2_X1 i_0_0_333 (.A1(n_0_0_284), .A2(n_0_109), .ZN(n_0_108));
   NAND2_X1 i_0_0_334 (.A1(ready), .A2(n_0_0_288), .ZN(n_0_109));
   NAND2_X1 i_0_0_335 (.A1(n_0_20), .A2(n_0_0_283), .ZN(n_0_110));
   NAND2_X1 i_0_0_277 (.A1(n_0_20), .A2(n_0_0_286), .ZN(n_0_53));
   NAND2_X1 i_0_0_278 (.A1(n_0_0_287), .A2(n_0_0_285), .ZN(n_0_0_283));
   NOR2_X1 i_0_0_339 (.A1(reset), .A2(n_0_0_285), .ZN(n_0_74));
   NAND2_X1 i_0_0_340 (.A1(n_0_20), .A2(n_0_0_284), .ZN(n_0_75));
   OR2_X1 i_0_0_341 (.A1(n_0_0_286), .A2(n_0_0_285), .ZN(n_0_0_284));
   NOR4_X1 i_0_0_279 (.A1(n_0_39), .A2(n_0_40), .A3(n_0_37), .A4(n_0_38), 
      .ZN(n_0_0_285));
   NOR2_X1 i_0_0_280 (.A1(ready), .A2(n_0_60), .ZN(n_0_0_287));
   INV_X1 i_0_0_281 (.A(n_0_0_288), .ZN(n_0_60));
   NOR2_X1 i_0_0_286 (.A1(reset), .A2(n_0_0_289), .ZN(n_0_0_288));
   NAND3_X1 i_0_0_287 (.A1(number_of_bits_in_dividend[4]), .A2(
      number_of_bits_in_dividend[2]), .A3(n_0_0_290), .ZN(n_0_0_289));
   AND3_X1 i_0_0_288 (.A1(number_of_bits_in_dividend[1]), .A2(
      number_of_bits_in_dividend[0]), .A3(number_of_bits_in_dividend[3]), 
      .ZN(n_0_0_290));
   AOI21_X1 i_0_0_350 (.A(n_0_0_373), .B1(divisor[0]), .B2(n_0_0_376), .ZN(n_0_4));
   INV_X1 i_0_0_351 (.A(n_0_0_291), .ZN(n_0_5));
   OAI21_X1 i_0_0_352 (.A(n_0_0_367), .B1(n_0_0_373), .B2(n_0_0_368), .ZN(
      n_0_0_291));
   AOI21_X1 i_0_0_353 (.A(n_0_0_361), .B1(n_0_0_367), .B2(n_0_117), .ZN(n_0_7));
   INV_X1 i_0_0_354 (.A(n_0_0_292), .ZN(n_0_8));
   OAI21_X1 i_0_0_355 (.A(n_0_0_352), .B1(n_0_0_361), .B2(n_0_0_353), .ZN(
      n_0_0_292));
   AOI21_X1 i_0_0_356 (.A(n_0_0_343), .B1(n_0_0_352), .B2(n_0_119), .ZN(n_0_9));
   INV_X1 i_0_0_290 (.A(n_0_0_293), .ZN(n_0_10));
   OAI21_X1 i_0_0_291 (.A(n_0_0_333), .B1(n_0_0_343), .B2(n_0_0_334), .ZN(
      n_0_0_293));
   AOI21_X1 i_0_0_359 (.A(n_0_0_328), .B1(n_0_0_333), .B2(n_0_121), .ZN(n_0_11));
   INV_X1 i_0_0_360 (.A(n_0_0_294), .ZN(n_0_12));
   OAI21_X1 i_0_0_361 (.A(n_0_0_321), .B1(n_0_0_328), .B2(n_0_0_322), .ZN(
      n_0_0_294));
   AOI21_X1 i_0_0_362 (.A(n_0_0_316), .B1(n_0_0_321), .B2(n_0_123), .ZN(n_0_13));
   NAND2_X1 i_0_0_292 (.A1(n_0_0_416), .A2(n_0_0_299), .ZN(n_0_0_298));
   AOI22_X1 i_0_0_293 (.A1(n_0_0_413), .A2(n_0_0_400), .B1(n_0_0_414), .B2(
      n_0_0_404), .ZN(n_0_0_299));
   INV_X1 i_0_0_379 (.A(n_0_0_303), .ZN(n_0_126));
   INV_X1 i_0_0_389 (.A(n_0_0_311), .ZN(n_0_124));
   OAI22_X1 i_0_0_294 (.A1(n_0_0_414), .A2(n_0_0_332), .B1(n_0_0_413), .B2(
      n_0_0_349), .ZN(n_0_0_331));
   OAI21_X1 i_0_0_295 (.A(divisor[12]), .B1(divisor[5]), .B2(n_0_0_409), 
      .ZN(n_0_0_342));
   INV_X1 i_0_0_437 (.A(n_0_0_353), .ZN(n_0_118));
   NOR2_X1 i_0_0_296 (.A1(n_0_0_479), .A2(n_0_0_410), .ZN(n_0_0_360));
   AOI21_X1 i_0_0_297 (.A(n_0_0_479), .B1(n_0_0_474), .B2(n_0_0_411), .ZN(
      n_0_0_366));
   NOR2_X1 i_0_0_298 (.A1(n_0_0_479), .A2(n_0_0_411), .ZN(n_0_0_372));
   INV_X1 i_0_0_464 (.A(n_0_0_377), .ZN(n_0_0_376));
   NOR2_X1 i_0_0_299 (.A1(n_0_0_479), .A2(n_0_0_473), .ZN(n_0_0_380));
   AOI22_X1 i_0_0_300 (.A1(n_0_0_414), .A2(n_0_0_384), .B1(n_0_0_412), .B2(
      n_0_0_382), .ZN(n_0_0_381));
   INV_X1 i_0_0_301 (.A(n_0_0_386), .ZN(n_0_0_385));
   NAND3_X1 i_0_0_302 (.A1(n_0_0_478), .A2(n_0_0_402), .A3(divisor[12]), 
      .ZN(n_0_0_387));
   AOI22_X1 i_0_0_303 (.A1(n_0_0_450), .A2(divisor[14]), .B1(n_0_0_451), 
      .B2(divisor[15]), .ZN(n_0_0_394));
   OAI21_X1 i_0_0_304 (.A(n_0_0_424), .B1(divisor[14]), .B2(n_0_0_450), .ZN(
      n_0_0_395));
   AOI22_X1 i_0_0_305 (.A1(n_0_0_412), .A2(n_0_0_403), .B1(n_0_0_414), .B2(
      n_0_0_397), .ZN(n_0_0_396));
   NOR2_X1 i_0_0_306 (.A1(n_0_0_479), .A2(n_0_0_408), .ZN(n_0_0_399));
   NOR2_X1 i_0_0_307 (.A1(divisor[1]), .A2(divisor[0]), .ZN(n_0_0_411));
   NOR2_X1 i_0_0_308 (.A1(n_0_0_415), .A2(n_0_0_414), .ZN(n_0_0_412));
   INV_X1 i_0_0_309 (.A(second_operand_number[2]), .ZN(n_0_0_426));
   INV_X1 i_0_0_310 (.A(second_operand_number[4]), .ZN(n_0_0_427));
   INV_X1 i_0_0_311 (.A(second_operand_number[5]), .ZN(n_0_0_428));
   INV_X1 i_0_0_312 (.A(second_operand_number[7]), .ZN(n_0_0_429));
   INV_X1 i_0_0_313 (.A(negated_second_operand_number[1]), .ZN(n_0_0_435));
   INV_X1 i_0_0_526 (.A(negated_second_operand_number[4]), .ZN(n_0_0_436));
   INV_X1 i_0_0_314 (.A(negated_second_operand_number[6]), .ZN(n_0_0_437));
   INV_X1 i_0_0_315 (.A(negated_second_operand_number[7]), .ZN(n_0_0_438));
   INV_X1 i_0_0_316 (.A(negated_second_operand_number[8]), .ZN(n_0_0_439));
   INV_X1 i_0_0_317 (.A(negated_second_operand_number[9]), .ZN(n_0_0_440));
   INV_X1 i_0_0_318 (.A(negated_second_operand_number[10]), .ZN(n_0_0_441));
   INV_X1 i_0_0_319 (.A(negated_second_operand_number[11]), .ZN(n_0_0_442));
   INV_X1 i_0_0_320 (.A(negated_second_operand_number[13]), .ZN(n_0_0_443));
   INV_X1 i_0_0_321 (.A(negated_second_operand_number[14]), .ZN(n_0_0_444));
   INV_X1 i_0_0_539 (.A(dividend[11]), .ZN(n_0_0_448));
   INV_X1 i_0_0_322 (.A(dividend[15]), .ZN(n_0_0_451));
   INV_X1 i_0_0_323 (.A(n_0_51), .ZN(n_0_0_452));
   INV_X1 i_0_0_324 (.A(n_0_49), .ZN(n_0_0_453));
   INV_X1 i_0_0_325 (.A(n_0_34), .ZN(n_0_0_460));
   INV_X1 i_0_0_326 (.A(n_0_33), .ZN(n_0_0_461));
   INV_X1 i_0_0_327 (.A(n_0_32), .ZN(n_0_0_462));
   INV_X1 i_0_0_328 (.A(n_0_31), .ZN(n_0_0_463));
   INV_X1 i_0_0_329 (.A(n_0_30), .ZN(n_0_0_464));
   INV_X1 i_0_0_330 (.A(n_0_29), .ZN(n_0_0_465));
   INV_X1 i_0_0_331 (.A(n_0_21), .ZN(n_0_0_472));
   INV_X1 i_0_0_332 (.A(divisor[2]), .ZN(n_0_0_474));
   INV_X1 i_0_0_336 (.A(divisor[15]), .ZN(n_0_0_480));
   NAND2_X1 i_0_0_8 (.A1(n_0_0_322), .A2(n_0_0_328), .ZN(n_0_0_321));
   INV_X1 i_0_0_9 (.A(n_0_0_106), .ZN(n_0_0_367));
   INV_X1 i_0_0_10 (.A(n_0_0_105), .ZN(n_0_0_373));
   NAND2_X1 i_0_0_337 (.A1(n_0_0_5), .A2(number_of_bits_in_dividend[4]), 
      .ZN(n_0_0_3));
   INV_X1 i_0_0_93 (.A(n_0_0_107), .ZN(n_0_117));
   INV_X1 i_0_0_94 (.A(n_0_0_317), .ZN(n_0_123));
   AOI21_X1 i_0_0_338 (.A(n_0_0_390), .B1(n_0_0_298), .B2(n_0_0_421), .ZN(
      n_0_0_4));
   NAND2_X1 i_0_0_342 (.A1(n_0_0_381), .A2(n_0_0_422), .ZN(n_0_0_61));
   NAND2_X1 i_0_0_343 (.A1(n_0_0_381), .A2(n_0_0_421), .ZN(n_0_0_62));
   INV_X1 i_0_0_344 (.A(n_0_0_396), .ZN(n_0_0_63));
   NAND2_X1 i_0_0_345 (.A1(n_0_0_396), .A2(n_0_0_421), .ZN(n_0_0_86));
   INV_X1 i_0_0_346 (.A(n_0_0_305), .ZN(n_0_0_87));
   INV_X1 i_0_0_347 (.A(divisor[3]), .ZN(n_0_0_98));
   INV_X1 i_0_0_348 (.A(divisor[2]), .ZN(n_0_0_99));
   BUF_X1 i_0_0_357 (.A(n_0_0_529), .Z(n_0_0_102));
   BUF_X1 i_0_0_358 (.A(n_0_0_123), .Z(n_0_0_450));
   BUF_X1 i_0_0_364 (.A(n_0_0_308), .Z(n_0_0_392));
   BUF_X1 i_0_0_137 (.A(n_0_0_296), .Z(n_0_116));
   BUF_X1 i_0_0_139 (.A(n_0_0_513), .Z(n_0_0_368));
   BUF_X1 i_0_0_140 (.A(n_0_0_118), .Z(n_0_0_322));
   BUF_X1 i_0_0_141 (.A(n_0_0_126), .Z(n_0_0_377));
   BUF_X1 i_0_0_365 (.A(n_0_0_127), .Z(n_0_115));
   BUF_X1 i_0_0_366 (.A(n_0_0_128), .Z(n_0_114));
   BUF_X1 i_0_0_144 (.A(n_0_0_129), .Z(n_0_0_105));
   BUF_X1 i_0_0_145 (.A(n_0_0_117), .Z(n_0_0_106));
   BUF_X1 i_0_0_146 (.A(n_0_0_295), .Z(n_0_0_107));
   BUF_X1 i_0_0_147 (.A(n_0_0_138), .Z(n_0_0_361));
   BUF_X1 i_0_0_149 (.A(n_0_0_131), .Z(n_0_0_353));
   BUF_X1 i_0_0_150 (.A(n_0_0_110), .Z(n_0_0_352));
   BUF_X1 i_0_0_151 (.A(n_0_0_130), .Z(n_0_119));
   BUF_X1 i_0_0_367 (.A(n_0_0_132), .Z(n_0_0_343));
   BUF_X1 i_0_0_368 (.A(n_0_0_133), .Z(n_0_0_334));
   BUF_X1 i_0_0_369 (.A(n_0_0_134), .Z(n_0_0_333));
   BUF_X1 i_0_0_155 (.A(n_0_0_119), .Z(n_0_121));
   BUF_X1 i_0_0_158 (.A(n_0_0_136), .Z(n_0_0_328));
   BUF_X1 i_0_0_159 (.A(n_0_0_137), .Z(n_0_0_317));
   INV_X1 i_0_0_161 (.A(n_0_0_510), .ZN(n_0_0_108));
   INV_X1 i_0_0_370 (.A(n_0_0_492), .ZN(n_0_0_109));
   NAND2_X1 i_0_0_163 (.A1(n_0_0_109), .A2(n_0_0_512), .ZN(n_0_0_110));
   INV_X1 i_0_0_164 (.A(n_0_0_513), .ZN(n_0_0_111));
   NOR2_X1 i_0_0_165 (.A1(n_0_0_111), .A2(n_0_0_108), .ZN(n_0_0_117));
   BUF_X1 i_0_0_166 (.A(n_0_0_307), .Z(n_0_0_118));
   BUF_X1 i_0_0_167 (.A(n_0_0_306), .Z(n_0_0_119));
   BUF_X1 i_0_0_371 (.A(n_0_0_502), .Z(n_0_0_123));
   BUF_X1 i_0_0_169 (.A(n_0_0_507), .Z(n_0_0_126));
   BUF_X1 i_0_0_372 (.A(n_0_0_509), .Z(n_0_0_127));
   BUF_X1 i_0_0_373 (.A(n_0_0_506), .Z(n_0_0_128));
   BUF_X1 i_0_0_172 (.A(n_0_0_108), .Z(n_0_0_129));
   BUF_X1 i_0_0_173 (.A(n_0_0_528), .Z(n_0_0_130));
   BUF_X1 i_0_0_174 (.A(n_0_0_512), .Z(n_0_0_131));
   BUF_X1 i_0_0_374 (.A(n_0_0_304), .Z(n_0_0_132));
   BUF_X1 i_0_0_375 (.A(n_0_0_302), .Z(n_0_0_133));
   BUF_X1 i_0_0_376 (.A(n_0_0_301), .Z(n_0_0_134));
   BUF_X1 i_0_0_178 (.A(n_0_0_300), .Z(n_0_0_136));
   BUF_X1 i_0_0_179 (.A(n_0_0_527), .Z(n_0_0_311));
   BUF_X1 i_0_0_180 (.A(n_0_0_576), .Z(n_0_0_137));
   BUF_X1 i_0_0_181 (.A(n_0_0_109), .Z(n_0_0_138));
   BUF_X1 i_0_0_184 (.A(n_0_0_505), .Z(n_0_0_295));
   BUF_X1 i_0_0_185 (.A(n_0_0_111), .Z(n_0_0_296));
   INV_X1 i_0_0_377 (.A(n_0_0_422), .ZN(n_0_0_297));
   INV_X1 i_0_0_189 (.A(n_0_0_517), .ZN(n_0_0_300));
   INV_X1 i_0_0_378 (.A(n_0_0_515), .ZN(n_0_0_301));
   INV_X1 i_0_0_381 (.A(n_0_120), .ZN(n_0_0_302));
   INV_X1 i_0_0_382 (.A(n_0_0_514), .ZN(n_0_0_304));
   NOR2_X1 i_0_0_349 (.A1(n_0_0_329), .A2(n_0_0_516), .ZN(n_0_0_306));
   INV_X1 i_0_0_363 (.A(n_0_122), .ZN(n_0_0_307));
   INV_X1 i_0_0_383 (.A(n_0_0_393), .ZN(n_0_0_308));
   NOR2_X1 i_0_0_384 (.A1(n_0_0_375), .A2(n_0_0_449), .ZN(n_0_0_122));
   INV_X1 i_0_0_385 (.A(n_0_0_287), .ZN(n_0_0_286));
   INV_X1 i_0_0_390 (.A(n_0_35), .ZN(n_0_0_459));
   INV_X1 i_0_0_391 (.A(n_0_0_309), .ZN(n_0_0_135));
   NAND2_X1 i_0_0_392 (.A1(n_0_0_446), .A2(dividend[12]), .ZN(n_0_0_309));
   INV_X1 i_0_0_393 (.A(n_0_0_369), .ZN(n_0_0_113));
   INV_X1 i_0_0_394 (.A(n_0_0_310), .ZN(n_0_0_139));
   NAND2_X1 i_0_0_395 (.A1(dividend[12]), .A2(dividend[0]), .ZN(n_0_0_310));
   INV_X1 i_0_0_396 (.A(n_0_0_481), .ZN(n_0_0_140));
   INV_X1 i_0_0_397 (.A(n_0_0_283), .ZN(n_0_0_282));
   INV_X1 i_0_0_398 (.A(dividend[12]), .ZN(n_0_0_449));
   OAI221_X1 i_0_0_380 (.A(n_0_0_312), .B1(n_0_0_283), .B2(n_0_0_73), .C1(
      n_0_0_320), .C2(n_0_0_319), .ZN(n_0_88));
   NAND2_X1 i_0_0_399 (.A1(n_0_0_280), .A2(n_0_41), .ZN(n_0_0_312));
   OAI21_X1 i_0_0_386 (.A(reset), .B1(n_0_0_142), .B2(n_0_0_405), .ZN(n_0_0_319));
   AOI211_X1 i_0_0_387 (.A(n_0_0_141), .B(n_0_0_323), .C1(n_0_0_64), .C2(
      n_0_0_152), .ZN(n_0_0_320));
   AND2_X1 i_0_0_388 (.A1(n_0_0_85), .A2(n_0_0_153), .ZN(n_0_0_323));
   MUX2_X1 i_0_0_401 (.A(n_0_0_324), .B(n_0_0_345), .S(n_0_0_149), .Z(n_0_0_85));
   NAND2_X1 i_0_0_408 (.A1(n_0_0_327), .A2(n_0_0_325), .ZN(n_0_0_324));
   OR2_X1 i_0_0_409 (.A1(n_0_0_144), .A2(n_0_0_88), .ZN(n_0_0_325));
   XNOR2_X1 i_0_0_410 (.A(n_0_0_326), .B(n_0_0_475), .ZN(n_0_0_88));
   OAI21_X1 i_0_0_411 (.A(dividend[12]), .B1(dividend[1]), .B2(dividend[0]), 
      .ZN(n_0_0_326));
   INV_X1 i_0_0_412 (.A(n_0_0_335), .ZN(n_0_0_327));
   NOR2_X1 i_0_0_413 (.A1(n_0_0_125), .A2(n_0_0_145), .ZN(n_0_0_335));
   INV_X1 i_0_0_417 (.A(n_0_0_337), .ZN(n_0_0_125));
   XNOR2_X1 i_0_0_425 (.A(n_0_0_338), .B(dividend[6]), .ZN(n_0_0_337));
   NAND2_X1 i_0_0_426 (.A1(n_0_0_418), .A2(dividend[12]), .ZN(n_0_0_338));
   AOI21_X1 i_0_0_400 (.A(n_0_0_65), .B1(n_0_0_95), .B2(n_0_0_149), .ZN(n_0_0_64));
   INV_X1 i_0_0_427 (.A(n_0_0_153), .ZN(n_0_0_152));
   OAI21_X1 i_0_0_402 (.A(n_0_0_350), .B1(n_0_0_341), .B2(n_0_0_339), .ZN(n_0_91));
   OAI21_X1 i_0_0_403 (.A(reset), .B1(n_0_0_340), .B2(n_0_0_142), .ZN(n_0_0_339));
   INV_X1 i_0_0_404 (.A(n_0_0_370), .ZN(n_0_0_340));
   AOI211_X1 i_0_0_405 (.A(n_0_0_141), .B(n_0_0_344), .C1(n_0_0_153), .C2(
      n_0_0_359), .ZN(n_0_0_341));
   NOR2_X1 i_0_0_406 (.A1(n_0_0_100), .A2(n_0_0_153), .ZN(n_0_0_344));
   AOI21_X1 i_0_0_407 (.A(n_0_0_101), .B1(n_0_0_148), .B2(n_0_0_345), .ZN(
      n_0_0_100));
   AOI21_X1 i_0_0_428 (.A(n_0_0_348), .B1(n_0_0_145), .B2(n_0_0_104), .ZN(
      n_0_0_345));
   INV_X1 i_0_0_429 (.A(n_0_0_346), .ZN(n_0_0_104));
   XNOR2_X1 i_0_0_430 (.A(n_0_0_347), .B(dividend[4]), .ZN(n_0_0_346));
   NAND2_X1 i_0_0_431 (.A1(n_0_0_423), .A2(dividend[12]), .ZN(n_0_0_347));
   NOR2_X1 i_0_0_432 (.A1(n_0_0_405), .A2(n_0_0_145), .ZN(n_0_0_348));
   NAND2_X1 i_0_0_414 (.A1(n_0_0_280), .A2(n_0_38), .ZN(n_0_0_350));
   NAND2_X1 i_0_0_415 (.A1(n_0_0_354), .A2(n_0_0_351), .ZN(n_0_92));
   AOI22_X1 i_0_0_416 (.A1(n_0_0_287), .A2(n_0_35), .B1(n_0_37), .B2(n_0_0_280), 
      .ZN(n_0_0_351));
   INV_X1 i_0_0_436 (.A(n_0_0_281), .ZN(n_0_0_280));
   OAI21_X1 i_0_0_418 (.A(n_0_0_355), .B1(n_0_0_391), .B2(n_0_0_357), .ZN(
      n_0_0_354));
   AOI21_X1 i_0_0_419 (.A(n_0_20), .B1(n_0_0_356), .B2(n_0_0_141), .ZN(n_0_0_355));
   NAND4_X1 i_0_0_420 (.A1(n_0_0_375), .A2(dividend[12]), .A3(n_0_0_379), 
      .A4(n_0_0_448), .ZN(n_0_0_356));
   OAI21_X1 i_0_0_421 (.A(n_0_0_142), .B1(n_0_0_358), .B2(n_0_0_153), .ZN(
      n_0_0_357));
   INV_X1 i_0_0_422 (.A(n_0_0_359), .ZN(n_0_0_358));
   OAI221_X1 i_0_0_423 (.A(n_0_0_362), .B1(n_0_0_481), .B2(n_0_0_369), .C1(
      n_0_0_370), .C2(n_0_0_388), .ZN(n_0_0_359));
   NAND2_X1 i_0_0_424 (.A1(n_0_0_114), .A2(n_0_0_148), .ZN(n_0_0_362));
   INV_X1 i_0_0_438 (.A(n_0_0_363), .ZN(n_0_0_114));
   MUX2_X1 i_0_0_440 (.A(n_0_0_116), .B(n_0_0_115), .S(n_0_0_145), .Z(n_0_0_363));
   XOR2_X1 i_0_0_441 (.A(dividend[9]), .B(n_0_0_364), .Z(n_0_0_116));
   NAND2_X1 i_0_0_442 (.A1(n_0_0_378), .A2(dividend[12]), .ZN(n_0_0_364));
   XNOR2_X1 i_0_0_443 (.A(n_0_0_365), .B(n_0_0_476), .ZN(n_0_0_115));
   NAND2_X1 i_0_0_444 (.A1(n_0_0_420), .A2(dividend[12]), .ZN(n_0_0_365));
   XNOR2_X1 i_0_0_445 (.A(n_0_0_417), .B(n_0_0_477), .ZN(n_0_0_369));
   XOR2_X1 i_0_0_433 (.A(dividend[11]), .B(n_0_0_371), .Z(n_0_0_370));
   NAND2_X1 i_0_0_434 (.A1(n_0_0_374), .A2(dividend[12]), .ZN(n_0_0_371));
   NAND2_X1 i_0_0_435 (.A1(n_0_0_375), .A2(n_0_0_379), .ZN(n_0_0_374));
   AOI21_X1 i_0_0_446 (.A(dividend[9]), .B1(n_0_0_378), .B2(dividend[12]), 
      .ZN(n_0_0_375));
   OR2_X1 i_0_0_447 (.A1(n_0_0_407), .A2(dividend[8]), .ZN(n_0_0_378));
   INV_X1 i_0_0_439 (.A(dividend[10]), .ZN(n_0_0_379));
   INV_X1 i_0_0_448 (.A(n_0_0_141), .ZN(n_0_0_142));
   NAND2_X1 i_0_0_449 (.A1(n_0_0_383), .A2(n_0_0_389), .ZN(n_0_0_141));
   NAND2_X1 i_0_0_450 (.A1(n_0_0_143), .A2(n_0_0_153), .ZN(n_0_0_383));
   INV_X1 i_0_0_451 (.A(n_0_0_388), .ZN(n_0_0_143));
   NAND2_X1 i_0_0_452 (.A1(n_0_0_144), .A2(n_0_0_149), .ZN(n_0_0_388));
   INV_X1 i_0_0_453 (.A(n_0_0_392), .ZN(n_0_0_389));
   AOI21_X1 i_0_0_454 (.A(n_0_0_401), .B1(n_0_0_120), .B2(n_0_0_150), .ZN(
      n_0_0_391));
   OAI21_X1 i_0_0_455 (.A(n_0_0_153), .B1(n_0_0_405), .B2(n_0_0_481), .ZN(
      n_0_0_401));
   XNOR2_X1 i_0_0_456 (.A(n_0_0_406), .B(dividend[8]), .ZN(n_0_0_405));
   NAND2_X1 i_0_0_457 (.A1(n_0_0_407), .A2(dividend[12]), .ZN(n_0_0_406));
   NAND2_X1 i_0_0_458 (.A1(n_0_0_417), .A2(n_0_0_477), .ZN(n_0_0_407));
   OAI21_X1 i_0_0_459 (.A(dividend[12]), .B1(n_0_0_418), .B2(dividend[6]), 
      .ZN(n_0_0_417));
   NAND2_X1 i_0_0_460 (.A1(n_0_0_419), .A2(n_0_0_476), .ZN(n_0_0_418));
   INV_X1 i_0_0_461 (.A(n_0_0_420), .ZN(n_0_0_419));
   OR2_X1 i_0_0_462 (.A1(n_0_0_423), .A2(dividend[4]), .ZN(n_0_0_420));
   OR2_X1 i_0_0_463 (.A1(n_0_0_446), .A2(dividend[3]), .ZN(n_0_0_423));
   NAND3_X1 i_0_0_465 (.A1(n_0_0_475), .A2(n_0_0_447), .A3(n_0_0_445), .ZN(
      n_0_0_446));
   INV_X1 i_0_0_466 (.A(dividend[0]), .ZN(n_0_0_445));
   INV_X1 i_0_0_467 (.A(dividend[1]), .ZN(n_0_0_447));
   INV_X1 i_0_0_468 (.A(dividend[2]), .ZN(n_0_0_475));
   INV_X1 i_0_0_469 (.A(dividend[5]), .ZN(n_0_0_476));
   INV_X1 i_0_0_470 (.A(dividend[7]), .ZN(n_0_0_477));
   NAND2_X1 i_0_0_471 (.A1(n_0_0_145), .A2(n_0_0_149), .ZN(n_0_0_481));
   INV_X1 i_0_0_472 (.A(n_0_0_144), .ZN(n_0_0_145));
   NAND2_X1 i_0_0_473 (.A1(n_0_0_483), .A2(n_0_0_482), .ZN(n_0_0_144));
   NAND2_X1 i_0_0_474 (.A1(n_0_0_484), .A2(n_0_0_146), .ZN(n_0_0_482));
   OR2_X1 i_0_0_475 (.A1(n_0_0_484), .A2(n_0_0_146), .ZN(n_0_0_483));
   INV_X1 i_0_0_476 (.A(n_0_0_147), .ZN(n_0_0_484));
   INV_X1 i_0_0_477 (.A(n_0_0_148), .ZN(n_0_0_149));
   XNOR2_X1 i_0_0_478 (.A(n_0_0_150), .B(n_0_0_486), .ZN(n_0_0_148));
   AND2_X1 i_0_0_479 (.A1(n_0_0_486), .A2(n_0_0_485), .ZN(n_0_0_153));
   NAND2_X1 i_0_0_480 (.A1(csa1_n_0), .A2(divisor[13]), .ZN(n_0_0_485));
   INV_X1 i_0_0_482 (.A(n_0_0_154), .ZN(n_0_0_486));
   INV_X1 i_0_0_481 (.A(n_0_0_562), .ZN(n_0_127));
   INV_X1 i_0_0_483 (.A(n_0_0_99), .ZN(n_0_0_487));
   INV_X1 i_0_0_484 (.A(n_0_0_98), .ZN(n_0_0_488));
   INV_X1 i_0_0_485 (.A(divisor[1]), .ZN(n_0_0_489));
   INV_X1 i_0_0_486 (.A(divisor[4]), .ZN(n_0_0_490));
   NAND2_X1 i_0_0_487 (.A1(n_0_0_398), .A2(n_0_0_390), .ZN(n_0_0_491));
   AOI22_X1 i_0_0_488 (.A1(n_0_0_395), .A2(n_0_0_394), .B1(dividend[15]), 
      .B2(n_0_0_480), .ZN(n_0_0_393));
   NAND2_X1 i_0_0_489 (.A1(n_0_0_511), .A2(n_0_0_513), .ZN(n_0_0_492));
   INV_X1 i_0_0_493 (.A(n_0_0_721), .ZN(n_0_128));
   INV_X1 i_0_0_494 (.A(n_0_0_559), .ZN(n_0_129));
   NAND3_X1 i_0_0_490 (.A1(n_0_0_495), .A2(n_0_0_722), .A3(n_0_0_494), .ZN(
      n_0_0_493));
   NAND2_X1 i_0_0_491 (.A1(n_0_0_336), .A2(n_0_0_422), .ZN(n_0_0_494));
   NAND2_X1 i_0_0_492 (.A1(n_0_0_330), .A2(n_0_0_421), .ZN(n_0_0_495));
   NAND2_X1 i_0_0_495 (.A1(n_0_0_390), .A2(n_0_0_497), .ZN(n_0_0_496));
   XNOR2_X1 i_0_0_496 (.A(n_0_0_372), .B(n_0_0_487), .ZN(n_0_0_497));
   OAI22_X1 i_0_0_497 (.A1(n_0_0_616), .A2(n_0_0_422), .B1(n_0_0_508), .B2(
      n_0_0_646), .ZN(n_0_0_498));
   NAND2_X1 i_0_0_498 (.A1(n_0_0_480), .A2(n_0_0_451), .ZN(n_0_0_499));
   NAND2_X1 i_0_0_499 (.A1(divisor[15]), .A2(dividend[15]), .ZN(n_0_0_500));
   INV_X1 i_0_0_500 (.A(n_0_0_424), .ZN(n_0_0_501));
   NAND2_X1 i_0_0_501 (.A1(csa0_n_0), .A2(dividend[13]), .ZN(n_0_0_424));
   BUF_X1 i_0_0_502 (.A(n_0_0_732), .Z(n_0_0_502));
   BUF_X1 i_0_0_503 (.A(n_0_0_719), .Z(n_0_0_503));
   BUF_X1 i_0_0_504 (.A(n_0_0_720), .Z(n_0_0_504));
   BUF_X1 i_0_0_510 (.A(n_0_0_649), .Z(n_0_122));
   BUF_X1 i_0_0_505 (.A(n_0_0_526), .Z(n_0_120));
   BUF_X1 i_0_0_512 (.A(n_0_0_613), .Z(n_0_0_505));
   BUF_X1 i_0_0_506 (.A(n_0_0_525), .Z(n_0_0_506));
   BUF_X1 i_0_0_514 (.A(n_0_0_611), .Z(n_0_0_507));
   BUF_X1 i_0_0_507 (.A(n_0_0_524), .Z(n_0_0_508));
   BUF_X1 i_0_0_508 (.A(n_0_0_523), .Z(n_0_0_509));
   BUF_X1 i_0_0_537 (.A(n_0_0_607), .Z(n_0_0_510));
   BUF_X1 i_0_0_509 (.A(n_0_0_521), .Z(n_0_0_511));
   BUF_X1 i_0_0_540 (.A(n_0_0_630), .Z(n_0_0_512));
   BUF_X1 i_0_0_511 (.A(n_0_0_606), .Z(n_0_0_513));
   BUF_X1 i_0_0_513 (.A(n_0_0_520), .Z(n_0_0_514));
   BUF_X1 i_0_0_515 (.A(n_0_0_552), .Z(n_0_0_515));
   BUF_X1 i_0_0_566 (.A(n_0_0_519), .Z(n_0_0_516));
   BUF_X1 i_0_0_567 (.A(n_0_0_518), .Z(n_0_0_329));
   BUF_X1 i_0_0_568 (.A(n_0_0_592), .Z(n_0_0_517));
   INV_X1 i_0_0_569 (.A(n_0_0_493), .ZN(n_0_0_518));
   INV_X1 i_0_0_570 (.A(n_0_0_491), .ZN(n_0_0_519));
   NAND2_X1 i_0_0_516 (.A1(n_0_0_602), .A2(n_0_0_630), .ZN(n_0_0_520));
   INV_X1 i_0_0_517 (.A(n_0_0_522), .ZN(n_0_0_521));
   NAND2_X1 i_0_0_518 (.A1(n_0_0_613), .A2(n_0_0_607), .ZN(n_0_0_522));
   NAND2_X1 i_0_0_519 (.A1(n_0_0_611), .A2(n_0_0_609), .ZN(n_0_0_523));
   NAND2_X1 i_0_0_520 (.A1(n_0_0_610), .A2(n_0_0_415), .ZN(n_0_0_524));
   INV_X1 i_0_0_521 (.A(n_0_0_612), .ZN(n_0_0_525));
   INV_X1 i_0_0_522 (.A(n_0_0_594), .ZN(n_0_0_526));
   AND2_X1 i_0_0_579 (.A1(n_0_0_582), .A2(n_0_0_590), .ZN(n_0_0_527));
   INV_X1 i_0_0_580 (.A(n_0_0_554), .ZN(n_0_0_528));
   INV_X1 i_0_0_523 (.A(n_0_0_497), .ZN(n_0_0_529));
   INV_X1 i_0_0_524 (.A(n_0_0_530), .ZN(n_0_0_336));
   NAND2_X1 i_0_0_525 (.A1(n_0_0_598), .A2(n_0_0_597), .ZN(n_0_0_530));
   INV_X1 i_0_0_527 (.A(n_0_0_331), .ZN(n_0_0_330));
   OAI21_X1 i_0_0_528 (.A(n_0_0_587), .B1(n_0_0_415), .B2(n_0_0_644), .ZN(
      n_0_0_332));
   AND2_X1 i_0_0_529 (.A1(n_0_0_663), .A2(n_0_0_664), .ZN(n_0_0_397));
   INV_X1 i_0_0_530 (.A(n_0_0_564), .ZN(n_0_0_305));
   NAND2_X1 i_0_0_531 (.A1(n_0_0_532), .A2(n_0_0_531), .ZN(n_0_59));
   OAI211_X1 i_0_0_532 (.A(n_0_20), .B(n_0_0_3), .C1(
      number_of_bits_in_dividend[4]), .C2(n_0_0_5), .ZN(n_0_0_531));
   INV_X1 i_0_0_533 (.A(n_0_0_532), .ZN(n_0_113));
   NAND3_X1 i_0_0_534 (.A1(n_0_0_572), .A2(n_0_0_560), .A3(n_0_0_533), .ZN(
      n_0_0_532));
   NOR3_X1 i_0_0_535 (.A1(n_0_0_547), .A2(n_0_20), .A3(n_0_0_558), .ZN(n_0_0_533));
   INV_X1 i_0_0_536 (.A(reset), .ZN(n_0_20));
   INV_X1 i_0_0_594 (.A(n_0_0_534), .ZN(n_0_14));
   OAI21_X1 i_0_0_595 (.A(n_0_0_551), .B1(n_0_0_316), .B2(n_0_0_311), .ZN(
      n_0_0_534));
   INV_X1 i_0_0_596 (.A(n_0_0_535), .ZN(n_0_0_316));
   NAND3_X1 i_0_0_597 (.A1(n_0_0_591), .A2(n_0_0_648), .A3(n_0_0_576), .ZN(
      n_0_0_535));
   INV_X1 i_0_0_598 (.A(n_0_0_536), .ZN(n_0_15));
   NAND2_X1 i_0_0_599 (.A1(n_0_0_537), .A2(n_0_0_573), .ZN(n_0_0_536));
   NAND2_X1 i_0_0_600 (.A1(n_0_0_551), .A2(n_0_125), .ZN(n_0_0_537));
   INV_X1 i_0_0_538 (.A(n_0_0_658), .ZN(n_0_125));
   INV_X1 i_0_0_541 (.A(n_0_0_538), .ZN(n_0_16));
   NAND2_X1 i_0_0_542 (.A1(n_0_0_540), .A2(n_0_0_539), .ZN(n_0_0_538));
   NAND2_X1 i_0_0_543 (.A1(n_0_0_573), .A2(n_0_0_544), .ZN(n_0_0_539));
   NAND2_X1 i_0_0_544 (.A1(n_0_0_572), .A2(n_0_0_303), .ZN(n_0_0_540));
   NAND2_X1 i_0_0_545 (.A1(n_0_0_541), .A2(n_0_0_542), .ZN(n_0_17));
   OAI21_X1 i_0_0_546 (.A(n_0_0_562), .B1(n_0_0_573), .B2(n_0_0_544), .ZN(
      n_0_0_541));
   NAND3_X1 i_0_0_547 (.A1(n_0_0_572), .A2(n_0_0_303), .A3(n_0_0_543), .ZN(
      n_0_0_542));
   INV_X1 i_0_0_548 (.A(n_0_0_562), .ZN(n_0_0_543));
   INV_X1 i_0_0_549 (.A(n_0_0_544), .ZN(n_0_0_303));
   NAND2_X1 i_0_0_550 (.A1(n_0_0_563), .A2(n_0_0_569), .ZN(n_0_0_544));
   INV_X1 i_0_0_612 (.A(n_0_0_545), .ZN(n_0_18));
   NAND2_X1 i_0_0_613 (.A1(n_0_0_546), .A2(n_0_0_549), .ZN(n_0_0_545));
   OAI21_X1 i_0_0_614 (.A(n_0_0_547), .B1(n_0_0_573), .B2(n_0_0_561), .ZN(
      n_0_0_546));
   INV_X1 i_0_0_551 (.A(n_0_0_721), .ZN(n_0_0_547));
   NAND2_X1 i_0_0_616 (.A1(n_0_0_548), .A2(n_0_0_557), .ZN(n_0_19));
   NAND2_X1 i_0_0_617 (.A1(n_0_0_549), .A2(n_0_0_559), .ZN(n_0_0_548));
   NAND4_X1 i_0_0_618 (.A1(n_0_0_550), .A2(n_0_0_721), .A3(n_0_0_658), .A4(
      n_0_0_560), .ZN(n_0_0_549));
   INV_X1 i_0_0_619 (.A(n_0_0_551), .ZN(n_0_0_550));
   NAND4_X1 i_0_0_620 (.A1(n_0_0_552), .A2(n_0_0_574), .A3(n_0_0_648), .A4(
      n_0_0_593), .ZN(n_0_0_551));
   INV_X1 i_0_0_552 (.A(n_0_0_553), .ZN(n_0_0_552));
   NAND4_X1 i_0_0_553 (.A1(n_0_0_554), .A2(n_0_0_594), .A3(n_0_0_630), .A4(
      n_0_0_604), .ZN(n_0_0_553));
   NAND2_X1 i_0_0_554 (.A1(n_0_0_555), .A2(n_0_0_628), .ZN(n_0_0_554));
   NAND2_X1 i_0_0_555 (.A1(n_0_0_556), .A2(n_0_0_722), .ZN(n_0_0_555));
   NAND2_X1 i_0_0_556 (.A1(n_0_0_620), .A2(n_0_0_626), .ZN(n_0_0_556));
   NAND4_X1 i_0_0_626 (.A1(n_0_0_572), .A2(n_0_0_721), .A3(n_0_0_560), .A4(
      n_0_0_558), .ZN(n_0_0_557));
   INV_X1 i_0_0_557 (.A(n_0_0_559), .ZN(n_0_0_558));
   NAND2_X1 i_0_0_558 (.A1(n_0_0_4), .A2(n_0_0_61), .ZN(n_0_0_559));
   INV_X1 i_0_0_559 (.A(n_0_0_561), .ZN(n_0_0_560));
   NAND3_X1 i_0_0_560 (.A1(n_0_0_563), .A2(n_0_0_569), .A3(n_0_0_562), .ZN(
      n_0_0_561));
   OAI211_X1 i_0_0_561 (.A(n_0_0_722), .B(n_0_0_86), .C1(n_0_0_87), .C2(
      n_0_0_297), .ZN(n_0_0_562));
   OAI211_X1 i_0_0_562 (.A(n_0_0_568), .B(n_0_0_722), .C1(n_0_0_422), .C2(
      n_0_0_564), .ZN(n_0_0_563));
   NAND2_X1 i_0_0_563 (.A1(n_0_0_565), .A2(n_0_0_567), .ZN(n_0_0_564));
   NAND2_X1 i_0_0_564 (.A1(n_0_0_384), .A2(n_0_0_413), .ZN(n_0_0_565));
   AOI21_X1 i_0_0_565 (.A(n_0_0_566), .B1(n_0_0_385), .B2(n_0_0_415), .ZN(
      n_0_0_384));
   AOI21_X1 i_0_0_571 (.A(n_0_0_415), .B1(n_0_0_697), .B2(n_0_0_696), .ZN(
      n_0_0_566));
   OAI21_X1 i_0_0_572 (.A(n_0_0_414), .B1(n_0_0_679), .B2(n_0_0_688), .ZN(
      n_0_0_567));
   NAND3_X1 i_0_0_573 (.A1(n_0_0_662), .A2(n_0_0_422), .A3(n_0_0_665), .ZN(
      n_0_0_568));
   NAND2_X1 i_0_0_574 (.A1(n_0_0_386), .A2(n_0_0_570), .ZN(n_0_0_569));
   NAND2_X1 i_0_0_575 (.A1(n_0_0_503), .A2(n_0_0_504), .ZN(n_0_0_570));
   INV_X1 i_0_0_576 (.A(n_0_0_571), .ZN(n_0_0_386));
   OR2_X1 i_0_0_577 (.A1(divisor[11]), .A2(n_0_0_387), .ZN(n_0_0_571));
   INV_X1 i_0_0_578 (.A(n_0_0_573), .ZN(n_0_0_572));
   NAND4_X1 i_0_0_581 (.A1(n_0_0_591), .A2(n_0_0_658), .A3(n_0_0_648), .A4(
      n_0_0_574), .ZN(n_0_0_573));
   INV_X1 i_0_0_582 (.A(n_0_0_575), .ZN(n_0_0_574));
   NAND3_X1 i_0_0_583 (.A1(n_0_0_576), .A2(n_0_0_582), .A3(n_0_0_590), .ZN(
      n_0_0_575));
   AOI21_X1 i_0_0_584 (.A(n_0_0_580), .B1(n_0_0_579), .B2(n_0_0_577), .ZN(
      n_0_0_576));
   AOI21_X1 i_0_0_585 (.A(n_0_0_390), .B1(n_0_0_578), .B2(n_0_0_422), .ZN(
      n_0_0_577));
   NAND2_X1 i_0_0_586 (.A1(n_0_0_653), .A2(n_0_0_654), .ZN(n_0_0_578));
   NAND2_X1 i_0_0_587 (.A1(n_0_0_584), .A2(n_0_0_421), .ZN(n_0_0_579));
   INV_X1 i_0_0_588 (.A(n_0_0_581), .ZN(n_0_0_580));
   NAND2_X1 i_0_0_589 (.A1(n_0_0_403), .A2(n_0_0_390), .ZN(n_0_0_581));
   INV_X1 i_0_0_590 (.A(n_0_0_404), .ZN(n_0_0_403));
   NAND2_X1 i_0_0_591 (.A1(n_0_0_673), .A2(n_0_0_672), .ZN(n_0_0_404));
   NAND3_X1 i_0_0_592 (.A1(n_0_0_589), .A2(n_0_0_722), .A3(n_0_0_583), .ZN(
      n_0_0_582));
   NAND2_X1 i_0_0_593 (.A1(n_0_0_584), .A2(n_0_0_422), .ZN(n_0_0_583));
   NAND2_X1 i_0_0_601 (.A1(n_0_0_585), .A2(n_0_0_586), .ZN(n_0_0_584));
   NAND3_X1 i_0_0_602 (.A1(n_0_0_671), .A2(n_0_0_413), .A3(n_0_0_667), .ZN(
      n_0_0_585));
   OAI211_X1 i_0_0_603 (.A(n_0_0_587), .B(n_0_0_414), .C1(n_0_0_415), .C2(
      n_0_0_644), .ZN(n_0_0_586));
   NAND2_X1 i_0_0_604 (.A1(n_0_0_415), .A2(n_0_0_588), .ZN(n_0_0_587));
   INV_X1 i_0_0_605 (.A(n_0_0_398), .ZN(n_0_0_588));
   NAND3_X1 i_0_0_606 (.A1(n_0_0_678), .A2(n_0_0_421), .A3(n_0_0_691), .ZN(
      n_0_0_589));
   NAND2_X1 i_0_0_607 (.A1(n_0_0_382), .A2(n_0_0_390), .ZN(n_0_0_590));
   NAND2_X1 i_0_0_608 (.A1(n_0_0_680), .A2(n_0_0_681), .ZN(n_0_0_382));
   INV_X1 i_0_0_609 (.A(n_0_0_592), .ZN(n_0_0_591));
   NAND4_X1 i_0_0_610 (.A1(n_0_0_602), .A2(n_0_0_630), .A3(n_0_0_594), .A4(
      n_0_0_593), .ZN(n_0_0_592));
   NAND2_X1 i_0_0_611 (.A1(n_0_0_491), .A2(n_0_0_493), .ZN(n_0_0_593));
   NAND2_X1 i_0_0_615 (.A1(n_0_0_595), .A2(n_0_0_601), .ZN(n_0_0_594));
   OAI211_X1 i_0_0_621 (.A(n_0_0_596), .B(n_0_0_722), .C1(n_0_0_599), .C2(
      n_0_0_421), .ZN(n_0_0_595));
   NAND3_X1 i_0_0_622 (.A1(n_0_0_598), .A2(n_0_0_597), .A3(n_0_0_421), .ZN(
      n_0_0_596));
   NAND3_X1 i_0_0_623 (.A1(n_0_0_637), .A2(n_0_0_414), .A3(n_0_0_640), .ZN(
      n_0_0_597));
   OAI211_X1 i_0_0_624 (.A(n_0_0_655), .B(n_0_0_413), .C1(n_0_0_656), .C2(
      n_0_0_415), .ZN(n_0_0_598));
   AOI21_X1 i_0_0_625 (.A(n_0_0_600), .B1(n_0_0_349), .B2(n_0_0_413), .ZN(
      n_0_0_599));
   INV_X1 i_0_0_627 (.A(n_0_0_621), .ZN(n_0_0_600));
   OR2_X1 i_0_0_628 (.A1(n_0_0_722), .A2(n_0_0_690), .ZN(n_0_0_601));
   INV_X1 i_0_0_629 (.A(n_0_0_603), .ZN(n_0_0_602));
   OAI21_X1 i_0_0_630 (.A(n_0_0_604), .B1(n_0_0_619), .B2(n_0_0_627), .ZN(
      n_0_0_603));
   INV_X1 i_0_0_631 (.A(n_0_0_605), .ZN(n_0_0_604));
   NAND3_X1 i_0_0_632 (.A1(n_0_0_613), .A2(n_0_0_607), .A3(n_0_0_606), .ZN(
      n_0_0_605));
   OAI21_X1 i_0_0_633 (.A(n_0_0_496), .B1(n_0_0_390), .B2(n_0_0_498), .ZN(
      n_0_0_606));
   INV_X1 i_0_0_634 (.A(n_0_0_608), .ZN(n_0_0_607));
   NAND3_X1 i_0_0_635 (.A1(n_0_0_612), .A2(n_0_0_611), .A3(n_0_0_609), .ZN(
      n_0_0_608));
   NAND4_X1 i_0_0_636 (.A1(n_0_0_610), .A2(divisor[0]), .A3(n_0_0_720), .A4(
      n_0_0_415), .ZN(n_0_0_609));
   NOR2_X1 i_0_0_637 (.A1(n_0_0_414), .A2(n_0_0_421), .ZN(n_0_0_610));
   NAND2_X1 i_0_0_638 (.A1(n_0_0_390), .A2(n_0_0_647), .ZN(n_0_0_611));
   NAND2_X1 i_0_0_639 (.A1(n_0_0_390), .A2(divisor[0]), .ZN(n_0_0_612));
   NAND2_X1 i_0_0_640 (.A1(n_0_0_614), .A2(n_0_0_618), .ZN(n_0_0_613));
   OAI211_X1 i_0_0_641 (.A(n_0_0_722), .B(n_0_0_615), .C1(n_0_0_616), .C2(
      n_0_0_421), .ZN(n_0_0_614));
   NAND4_X1 i_0_0_642 (.A1(n_0_0_645), .A2(n_0_0_415), .A3(n_0_0_421), .A4(
      n_0_0_643), .ZN(n_0_0_615));
   OAI211_X1 i_0_0_643 (.A(n_0_0_415), .B(n_0_0_617), .C1(divisor[0]), .C2(
      n_0_0_413), .ZN(n_0_0_616));
   NAND2_X1 i_0_0_644 (.A1(n_0_0_413), .A2(n_0_0_497), .ZN(n_0_0_617));
   NAND2_X1 i_0_0_645 (.A1(n_0_0_390), .A2(n_0_0_644), .ZN(n_0_0_618));
   AOI21_X1 i_0_0_646 (.A(n_0_0_390), .B1(n_0_0_620), .B2(n_0_0_626), .ZN(
      n_0_0_619));
   NAND3_X1 i_0_0_647 (.A1(n_0_0_623), .A2(n_0_0_421), .A3(n_0_0_621), .ZN(
      n_0_0_620));
   NAND3_X1 i_0_0_648 (.A1(n_0_0_415), .A2(n_0_0_414), .A3(n_0_0_622), .ZN(
      n_0_0_621));
   INV_X1 i_0_0_649 (.A(n_0_0_644), .ZN(n_0_0_622));
   NAND2_X1 i_0_0_650 (.A1(n_0_0_349), .A2(n_0_0_413), .ZN(n_0_0_623));
   NAND2_X1 i_0_0_651 (.A1(n_0_0_624), .A2(n_0_0_625), .ZN(n_0_0_349));
   OAI21_X1 i_0_0_652 (.A(n_0_0_415), .B1(n_0_0_668), .B2(n_0_0_670), .ZN(
      n_0_0_624));
   NAND2_X1 i_0_0_653 (.A1(n_0_0_416), .A2(n_0_0_647), .ZN(n_0_0_625));
   NAND2_X1 i_0_0_654 (.A1(n_0_0_633), .A2(n_0_0_422), .ZN(n_0_0_626));
   INV_X1 i_0_0_655 (.A(n_0_0_628), .ZN(n_0_0_627));
   NAND2_X1 i_0_0_656 (.A1(n_0_0_390), .A2(n_0_0_629), .ZN(n_0_0_628));
   NOR2_X1 i_0_0_657 (.A1(n_0_0_668), .A2(n_0_0_670), .ZN(n_0_0_629));
   OAI21_X1 i_0_0_658 (.A(n_0_0_631), .B1(n_0_0_632), .B2(n_0_0_390), .ZN(
      n_0_0_630));
   OR2_X1 i_0_0_659 (.A1(n_0_0_722), .A2(n_0_0_699), .ZN(n_0_0_631));
   AOI21_X1 i_0_0_660 (.A(n_0_0_641), .B1(n_0_0_633), .B2(n_0_0_421), .ZN(
      n_0_0_632));
   NOR2_X1 i_0_0_661 (.A1(n_0_0_636), .A2(n_0_0_634), .ZN(n_0_0_633));
   INV_X1 i_0_0_662 (.A(n_0_0_635), .ZN(n_0_0_634));
   NAND3_X1 i_0_0_663 (.A1(n_0_0_415), .A2(n_0_0_102), .A3(n_0_0_414), .ZN(
      n_0_0_635));
   AOI21_X1 i_0_0_664 (.A(n_0_0_414), .B1(n_0_0_637), .B2(n_0_0_640), .ZN(
      n_0_0_636));
   OAI21_X1 i_0_0_665 (.A(n_0_0_699), .B1(n_0_0_639), .B2(n_0_0_638), .ZN(
      n_0_0_637));
   AOI21_X1 i_0_0_666 (.A(n_0_0_728), .B1(n_0_0_730), .B2(n_0_0_734), .ZN(
      n_0_0_638));
   INV_X1 i_0_0_667 (.A(n_0_0_727), .ZN(n_0_0_639));
   NAND3_X1 i_0_0_668 (.A1(n_0_0_725), .A2(divisor[0]), .A3(n_0_0_727), .ZN(
      n_0_0_640));
   AOI21_X1 i_0_0_669 (.A(n_0_0_421), .B1(n_0_0_642), .B2(n_0_0_415), .ZN(
      n_0_0_641));
   AND2_X1 i_0_0_670 (.A1(n_0_0_645), .A2(n_0_0_643), .ZN(n_0_0_642));
   NAND2_X1 i_0_0_671 (.A1(n_0_0_413), .A2(n_0_0_644), .ZN(n_0_0_643));
   XNOR2_X1 i_0_0_672 (.A(n_0_0_366), .B(n_0_0_488), .ZN(n_0_0_644));
   NAND2_X1 i_0_0_673 (.A1(n_0_0_414), .A2(n_0_0_646), .ZN(n_0_0_645));
   INV_X1 i_0_0_674 (.A(n_0_0_647), .ZN(n_0_0_646));
   XNOR2_X1 i_0_0_675 (.A(n_0_0_380), .B(n_0_0_489), .ZN(n_0_0_647));
   INV_X1 i_0_0_676 (.A(n_0_0_649), .ZN(n_0_0_648));
   AOI22_X1 i_0_0_677 (.A1(n_0_0_652), .A2(n_0_0_650), .B1(n_0_0_390), .B2(
      n_0_0_657), .ZN(n_0_0_649));
   INV_X1 i_0_0_678 (.A(n_0_0_651), .ZN(n_0_0_650));
   OAI21_X1 i_0_0_679 (.A(n_0_0_722), .B1(n_0_0_331), .B2(n_0_0_421), .ZN(
      n_0_0_651));
   NAND3_X1 i_0_0_680 (.A1(n_0_0_653), .A2(n_0_0_421), .A3(n_0_0_654), .ZN(
      n_0_0_652));
   NAND3_X1 i_0_0_681 (.A1(n_0_0_695), .A2(n_0_0_698), .A3(n_0_0_413), .ZN(
      n_0_0_653));
   OAI211_X1 i_0_0_682 (.A(n_0_0_655), .B(n_0_0_414), .C1(n_0_0_656), .C2(
      n_0_0_415), .ZN(n_0_0_654));
   NAND2_X1 i_0_0_683 (.A1(n_0_0_415), .A2(n_0_0_690), .ZN(n_0_0_655));
   INV_X1 i_0_0_684 (.A(n_0_0_102), .ZN(n_0_0_656));
   NAND2_X1 i_0_0_685 (.A1(n_0_0_697), .A2(n_0_0_696), .ZN(n_0_0_657));
   OAI21_X1 i_0_0_686 (.A(n_0_0_700), .B1(n_0_0_659), .B2(n_0_0_390), .ZN(
      n_0_0_658));
   INV_X1 i_0_0_687 (.A(n_0_0_660), .ZN(n_0_0_659));
   NAND2_X1 i_0_0_688 (.A1(n_0_0_661), .A2(n_0_0_677), .ZN(n_0_0_660));
   NAND3_X1 i_0_0_689 (.A1(n_0_0_662), .A2(n_0_0_421), .A3(n_0_0_665), .ZN(
      n_0_0_661));
   NAND3_X1 i_0_0_690 (.A1(n_0_0_663), .A2(n_0_0_413), .A3(n_0_0_664), .ZN(
      n_0_0_662));
   OAI21_X1 i_0_0_691 (.A(n_0_0_415), .B1(n_0_0_701), .B2(n_0_0_703), .ZN(
      n_0_0_663));
   NAND2_X1 i_0_0_692 (.A1(n_0_0_416), .A2(n_0_0_398), .ZN(n_0_0_664));
   XNOR2_X1 i_0_0_693 (.A(divisor[7]), .B(n_0_0_399), .ZN(n_0_0_398));
   NAND2_X1 i_0_0_694 (.A1(n_0_0_666), .A2(n_0_0_414), .ZN(n_0_0_665));
   NAND2_X1 i_0_0_695 (.A1(n_0_0_671), .A2(n_0_0_667), .ZN(n_0_0_666));
   OAI21_X1 i_0_0_696 (.A(n_0_0_416), .B1(n_0_0_670), .B2(n_0_0_668), .ZN(
      n_0_0_667));
   INV_X1 i_0_0_697 (.A(n_0_0_669), .ZN(n_0_0_668));
   NAND3_X1 i_0_0_698 (.A1(n_0_0_409), .A2(divisor[12]), .A3(n_0_0_709), 
      .ZN(n_0_0_669));
   AOI21_X1 i_0_0_699 (.A(n_0_0_709), .B1(n_0_0_409), .B2(divisor[12]), .ZN(
      n_0_0_670));
   NAND3_X1 i_0_0_700 (.A1(n_0_0_673), .A2(n_0_0_415), .A3(n_0_0_672), .ZN(
      n_0_0_671));
   NAND3_X1 i_0_0_701 (.A1(n_0_0_675), .A2(divisor[12]), .A3(divisor[9]), 
      .ZN(n_0_0_672));
   OAI21_X1 i_0_0_702 (.A(n_0_0_718), .B1(n_0_0_674), .B2(n_0_0_479), .ZN(
      n_0_0_673));
   INV_X1 i_0_0_703 (.A(n_0_0_675), .ZN(n_0_0_674));
   NAND4_X1 i_0_0_704 (.A1(n_0_0_676), .A2(n_0_0_717), .A3(n_0_0_716), .A4(
      n_0_0_707), .ZN(n_0_0_675));
   INV_X1 i_0_0_705 (.A(n_0_0_409), .ZN(n_0_0_676));
   NAND3_X1 i_0_0_706 (.A1(n_0_0_686), .A2(n_0_0_684), .A3(n_0_0_715), .ZN(
      n_0_0_409));
   NAND3_X1 i_0_0_707 (.A1(n_0_0_678), .A2(n_0_0_422), .A3(n_0_0_691), .ZN(
      n_0_0_677));
   OAI21_X1 i_0_0_708 (.A(n_0_0_413), .B1(n_0_0_679), .B2(n_0_0_688), .ZN(
      n_0_0_678));
   AOI21_X1 i_0_0_709 (.A(n_0_0_416), .B1(n_0_0_680), .B2(n_0_0_681), .ZN(
      n_0_0_679));
   OAI21_X1 i_0_0_710 (.A(divisor[10]), .B1(n_0_0_402), .B2(n_0_0_479), .ZN(
      n_0_0_680));
   INV_X1 i_0_0_711 (.A(n_0_0_682), .ZN(n_0_0_402));
   NAND3_X1 i_0_0_712 (.A1(n_0_0_682), .A2(divisor[12]), .A3(n_0_0_478), 
      .ZN(n_0_0_681));
   NAND4_X1 i_0_0_713 (.A1(n_0_0_408), .A2(n_0_0_718), .A3(n_0_0_717), .A4(
      n_0_0_716), .ZN(n_0_0_682));
   INV_X1 i_0_0_714 (.A(n_0_0_683), .ZN(n_0_0_408));
   NAND4_X1 i_0_0_715 (.A1(n_0_0_686), .A2(n_0_0_684), .A3(n_0_0_707), .A4(
      n_0_0_715), .ZN(n_0_0_683));
   INV_X1 i_0_0_716 (.A(n_0_0_685), .ZN(n_0_0_684));
   NAND2_X1 i_0_0_717 (.A1(n_0_0_712), .A2(n_0_0_473), .ZN(n_0_0_685));
   INV_X1 i_0_0_718 (.A(n_0_0_687), .ZN(n_0_0_686));
   NAND2_X1 i_0_0_719 (.A1(n_0_0_714), .A2(n_0_0_713), .ZN(n_0_0_687));
   INV_X1 i_0_0_720 (.A(n_0_0_689), .ZN(n_0_0_688));
   NAND2_X1 i_0_0_721 (.A1(n_0_0_416), .A2(n_0_0_690), .ZN(n_0_0_689));
   XNOR2_X1 i_0_0_722 (.A(divisor[6]), .B(n_0_0_342), .ZN(n_0_0_690));
   NAND2_X1 i_0_0_723 (.A1(n_0_0_694), .A2(n_0_0_414), .ZN(n_0_0_691));
   INV_X1 i_0_0_724 (.A(n_0_0_413), .ZN(n_0_0_414));
   NAND2_X1 i_0_0_725 (.A1(n_0_0_692), .A2(n_0_0_730), .ZN(n_0_0_413));
   NAND3_X1 i_0_0_726 (.A1(n_0_0_693), .A2(n_0_0_69), .A3(n_0_0_8), .ZN(
      n_0_0_692));
   NAND2_X1 i_0_0_727 (.A1(n_0_0_731), .A2(n_0_0_733), .ZN(n_0_0_693));
   NAND2_X1 i_0_0_728 (.A1(n_0_0_695), .A2(n_0_0_698), .ZN(n_0_0_694));
   NAND3_X1 i_0_0_729 (.A1(n_0_0_697), .A2(n_0_0_415), .A3(n_0_0_696), .ZN(
      n_0_0_695));
   NAND3_X1 i_0_0_730 (.A1(n_0_0_706), .A2(divisor[12]), .A3(divisor[8]), 
      .ZN(n_0_0_696));
   OAI21_X1 i_0_0_731 (.A(n_0_0_717), .B1(n_0_0_705), .B2(n_0_0_479), .ZN(
      n_0_0_697));
   INV_X1 i_0_0_732 (.A(divisor[12]), .ZN(n_0_0_479));
   NAND2_X1 i_0_0_733 (.A1(n_0_0_416), .A2(n_0_0_699), .ZN(n_0_0_698));
   XNOR2_X1 i_0_0_734 (.A(n_0_0_360), .B(n_0_0_490), .ZN(n_0_0_699));
   INV_X1 i_0_0_735 (.A(n_0_0_415), .ZN(n_0_0_416));
   NAND2_X1 i_0_0_736 (.A1(n_0_0_400), .A2(n_0_0_390), .ZN(n_0_0_700));
   OR2_X1 i_0_0_737 (.A1(n_0_0_701), .A2(n_0_0_703), .ZN(n_0_0_400));
   INV_X1 i_0_0_738 (.A(n_0_0_702), .ZN(n_0_0_701));
   NAND3_X1 i_0_0_739 (.A1(n_0_0_704), .A2(divisor[12]), .A3(divisor[11]), 
      .ZN(n_0_0_702));
   AOI21_X1 i_0_0_740 (.A(divisor[11]), .B1(n_0_0_704), .B2(divisor[12]), 
      .ZN(n_0_0_703));
   NAND4_X1 i_0_0_741 (.A1(n_0_0_705), .A2(n_0_0_478), .A3(n_0_0_718), .A4(
      n_0_0_717), .ZN(n_0_0_704));
   INV_X1 i_0_0_742 (.A(n_0_0_706), .ZN(n_0_0_705));
   NAND4_X1 i_0_0_743 (.A1(n_0_0_410), .A2(n_0_0_716), .A3(n_0_0_715), .A4(
      n_0_0_707), .ZN(n_0_0_706));
   INV_X1 i_0_0_744 (.A(n_0_0_708), .ZN(n_0_0_707));
   NAND2_X1 i_0_0_745 (.A1(n_0_0_710), .A2(n_0_0_709), .ZN(n_0_0_708));
   INV_X1 i_0_0_746 (.A(divisor[5]), .ZN(n_0_0_709));
   INV_X1 i_0_0_747 (.A(divisor[6]), .ZN(n_0_0_710));
   INV_X1 i_0_0_748 (.A(n_0_0_711), .ZN(n_0_0_410));
   NAND4_X1 i_0_0_749 (.A1(n_0_0_714), .A2(n_0_0_713), .A3(n_0_0_712), .A4(
      n_0_0_473), .ZN(n_0_0_711));
   INV_X1 i_0_0_750 (.A(divisor[0]), .ZN(n_0_0_473));
   INV_X1 i_0_0_751 (.A(divisor[1]), .ZN(n_0_0_712));
   INV_X1 i_0_0_752 (.A(divisor[2]), .ZN(n_0_0_713));
   INV_X1 i_0_0_753 (.A(divisor[3]), .ZN(n_0_0_714));
   INV_X1 i_0_0_754 (.A(divisor[4]), .ZN(n_0_0_715));
   INV_X1 i_0_0_755 (.A(divisor[7]), .ZN(n_0_0_716));
   INV_X1 i_0_0_756 (.A(divisor[8]), .ZN(n_0_0_717));
   INV_X1 i_0_0_757 (.A(divisor[9]), .ZN(n_0_0_718));
   INV_X1 i_0_0_758 (.A(divisor[10]), .ZN(n_0_0_478));
   NAND2_X1 i_0_0_759 (.A1(n_0_0_719), .A2(n_0_0_720), .ZN(n_0_0_390));
   NAND2_X1 i_0_0_760 (.A1(n_0_0_415), .A2(n_0_0_723), .ZN(n_0_0_719));
   INV_X1 i_0_0_761 (.A(n_0_0_393), .ZN(n_0_0_720));
   OAI211_X1 i_0_0_762 (.A(n_0_0_722), .B(n_0_0_62), .C1(n_0_0_63), .C2(
      n_0_0_421), .ZN(n_0_0_721));
   AOI21_X1 i_0_0_763 (.A(n_0_0_393), .B1(n_0_0_415), .B2(n_0_0_723), .ZN(
      n_0_0_722));
   INV_X1 i_0_0_764 (.A(n_0_0_724), .ZN(n_0_0_723));
   NAND3_X1 i_0_0_765 (.A1(n_0_0_421), .A2(n_0_0_733), .A3(n_0_0_731), .ZN(
      n_0_0_724));
   NAND2_X1 i_0_0_766 (.A1(n_0_0_725), .A2(n_0_0_727), .ZN(n_0_0_415));
   NAND2_X1 i_0_0_767 (.A1(n_0_0_726), .A2(n_0_0_729), .ZN(n_0_0_725));
   NAND2_X1 i_0_0_768 (.A1(n_0_0_730), .A2(n_0_0_734), .ZN(n_0_0_726));
   NAND3_X1 i_0_0_769 (.A1(n_0_0_730), .A2(n_0_0_734), .A3(n_0_0_728), .ZN(
      n_0_0_727));
   INV_X1 i_0_0_770 (.A(n_0_0_729), .ZN(n_0_0_728));
   NAND2_X1 i_0_0_771 (.A1(n_0_0_499), .A2(n_0_0_500), .ZN(n_0_0_729));
   NAND3_X1 i_0_0_772 (.A1(n_0_0_736), .A2(n_0_0_731), .A3(n_0_0_733), .ZN(
      n_0_0_730));
   NAND2_X1 i_0_0_773 (.A1(n_0_0_732), .A2(divisor[14]), .ZN(n_0_0_731));
   INV_X1 i_0_0_774 (.A(dividend[14]), .ZN(n_0_0_732));
   NAND2_X1 i_0_0_775 (.A1(dividend[14]), .A2(csa0_n_1), .ZN(n_0_0_733));
   NAND2_X1 i_0_0_776 (.A1(n_0_0_735), .A2(dividend[14]), .ZN(n_0_0_734));
   INV_X1 i_0_0_777 (.A(divisor[14]), .ZN(n_0_0_735));
   INV_X1 i_0_0_778 (.A(n_0_0_422), .ZN(n_0_0_421));
   NAND2_X1 i_0_0_779 (.A1(n_0_0_736), .A2(n_0_0_70), .ZN(n_0_0_422));
   NAND2_X1 i_0_0_780 (.A1(n_0_0_69), .A2(n_0_0_8), .ZN(n_0_0_736));
   INV_X1 i_0_0_781 (.A(csa0_n_0), .ZN(n_0_0_8));
   INV_X1 i_0_0_782 (.A(dividend[13]), .ZN(n_0_0_69));
   INV_X1 i_0_0_783 (.A(n_0_0_501), .ZN(n_0_0_70));
   INV_X1 i_0_0_784 (.A(n_0_0_74), .ZN(n_0_0_73));
   XOR2_X1 i_0_0_785 (.A(n_0_40), .B(n_0_0_75), .Z(n_0_0_74));
   OAI21_X1 i_0_0_786 (.A(n_0_0_76), .B1(n_0_0_257), .B2(n_0_0_255), .ZN(
      n_0_0_75));
   OAI21_X1 i_0_0_787 (.A(sign), .B1(n_0_42), .B2(n_0_0_77), .ZN(n_0_0_76));
   AOI21_X1 i_0_0_788 (.A(n_0_0_257), .B1(n_0_0_254), .B2(n_0_0_78), .ZN(
      n_0_0_77));
   OAI21_X1 i_0_0_789 (.A(sign), .B1(n_0_44), .B2(n_0_0_246), .ZN(n_0_0_78));
   AOI21_X1 i_0_0_790 (.A(n_0_0_257), .B1(n_0_0_253), .B2(n_0_0_248), .ZN(
      n_0_0_246));
   NAND2_X1 i_0_0_791 (.A1(sign), .A2(n_0_0_249), .ZN(n_0_0_248));
   OR4_X1 i_0_0_792 (.A1(n_0_48), .A2(n_0_0_71), .A3(n_0_47), .A4(n_0_46), 
      .ZN(n_0_0_249));
   AOI21_X1 i_0_0_793 (.A(n_0_0_257), .B1(n_0_0_252), .B2(n_0_0_251), .ZN(
      n_0_0_250));
   OAI21_X1 i_0_0_794 (.A(sign), .B1(n_0_48), .B2(n_0_0_71), .ZN(n_0_0_251));
   INV_X1 i_0_0_795 (.A(n_0_47), .ZN(n_0_0_252));
   INV_X1 i_0_0_796 (.A(n_0_45), .ZN(n_0_0_253));
   INV_X1 i_0_0_797 (.A(n_0_43), .ZN(n_0_0_254));
   INV_X1 i_0_0_798 (.A(n_0_41), .ZN(n_0_0_255));
   INV_X1 i_0_0_799 (.A(n_0_40), .ZN(n_0_0_256));
   INV_X1 i_0_0_800 (.A(sign), .ZN(n_0_0_257));
   XNOR2_X1 i_0_0_801 (.A(second_operand_number[15]), .B(n_0_0_259), .ZN(
      n_0_0_258));
   AOI22_X1 i_0_0_802 (.A1(n_0_22), .A2(n_0_0_276), .B1(
      second_operand_number[14]), .B2(n_0_0_274), .ZN(n_0_0_259));
   INV_X1 i_0_0_803 (.A(n_0_0_275), .ZN(n_0_0_274));
   NOR2_X1 i_0_0_804 (.A1(n_0_22), .A2(n_0_0_276), .ZN(n_0_0_275));
   AOI22_X1 i_0_0_805 (.A1(n_0_0_471), .A2(n_0_0_458), .B1(n_0_0_313), .B2(
      n_0_0_277), .ZN(n_0_0_276));
   AOI22_X1 i_0_0_806 (.A1(n_0_0_471), .A2(n_0_0_458), .B1(n_0_23), .B2(
      second_operand_number[13]), .ZN(n_0_0_277));
   AOI22_X1 i_0_0_807 (.A1(n_0_24), .A2(second_operand_number[12]), .B1(
      n_0_0_454), .B2(n_0_0_314), .ZN(n_0_0_313));
   OAI22_X1 i_0_0_808 (.A1(n_0_0_469), .A2(n_0_0_457), .B1(n_0_0_318), .B2(
      n_0_0_315), .ZN(n_0_0_314));
   NOR2_X1 i_0_0_809 (.A1(n_0_25), .A2(second_operand_number[11]), .ZN(n_0_0_315));
   AOI21_X1 i_0_0_810 (.A(n_0_0_425), .B1(n_0_26), .B2(second_operand_number[10]), 
      .ZN(n_0_0_318));
   AOI21_X1 i_0_0_811 (.A(n_0_0_430), .B1(n_0_0_468), .B2(n_0_0_456), .ZN(
      n_0_0_425));
   AOI22_X1 i_0_0_812 (.A1(n_0_27), .A2(second_operand_number[9]), .B1(n_0_0_434), 
      .B2(n_0_0_431), .ZN(n_0_0_430));
   OAI22_X1 i_0_0_813 (.A1(n_0_0_466), .A2(n_0_0_455), .B1(n_0_0_433), .B2(
      n_0_0_432), .ZN(n_0_0_431));
   NOR2_X1 i_0_0_814 (.A1(n_0_28), .A2(second_operand_number[8]), .ZN(n_0_0_432));
   OAI21_X1 i_0_0_815 (.A(n_0_0_72), .B1(n_0_29), .B2(second_operand_number[7]), 
      .ZN(n_0_0_433));
   XOR2_X1 i_0_0_816 (.A(n_0_27), .B(second_operand_number[9]), .Z(n_0_0_434));
   XOR2_X1 i_0_0_817 (.A(n_0_24), .B(second_operand_number[12]), .Z(n_0_0_454));
   INV_X1 i_0_0_818 (.A(second_operand_number[8]), .ZN(n_0_0_455));
   INV_X1 i_0_0_819 (.A(second_operand_number[10]), .ZN(n_0_0_456));
   INV_X1 i_0_0_820 (.A(second_operand_number[11]), .ZN(n_0_0_457));
   INV_X1 i_0_0_821 (.A(second_operand_number[13]), .ZN(n_0_0_458));
   INV_X1 i_0_0_822 (.A(n_0_28), .ZN(n_0_0_466));
   INV_X1 i_0_0_823 (.A(n_0_27), .ZN(n_0_0_467));
   INV_X1 i_0_0_824 (.A(n_0_26), .ZN(n_0_0_468));
   INV_X1 i_0_0_825 (.A(n_0_25), .ZN(n_0_0_469));
   INV_X1 i_0_0_826 (.A(n_0_24), .ZN(n_0_0_470));
   INV_X1 i_0_0_827 (.A(n_0_23), .ZN(n_0_0_471));
   MUX2_X1 overFlow_reg_enable_mux_0 (.A(overFlow), .B(n_0_74), .S(n_0_75), 
      .Z(n_0_111));
   MUX2_X1 ready_reg_enable_mux_0 (.A(ready), .B(n_0_20), .S(n_0_53), .Z(n_0_112));
endmodule
