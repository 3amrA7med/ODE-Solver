/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 22:11:50 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 797789819 */

module Division_CLHA(reset, clk, dividend, divisor, Q, ready, overFlow, 
      divideByZero);
   input reset;
   input clk;
   input [15:0]dividend;
   input [15:0]divisor;
   output [15:0]Q;
   output ready;
   output overFlow;
   output divideByZero;

   wire cla0_n_0;
   wire cla0_n_1;
   wire cla0_n_2;
   wire cla1_n_0;
   wire n_0_0;
   wire n_0_1;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_2;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire [15:0]negated_second_operand_number;
   wire [15:0]second_operand_number;
   wire n_0_3;
   wire [4:0]number_of_bits_in_dividend;
   wire sign;
   wire n_0_6;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_0_0;
   wire n_0_57;
   wire n_0_0_1;
   wire n_0_58;
   wire n_0_0_2;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_53;
   wire n_0_76;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_77;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_78;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_79;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_80;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_81;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_82;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_83;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_84;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_85;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_86;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_87;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_88;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_89;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_90;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_91;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_92;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_93;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_94;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_95;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_96;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_97;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_98;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_99;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_100;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_101;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_102;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_103;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_104;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_105;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_106;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_107;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_108;
   wire n_0_109;
   wire n_0_60;
   wire n_0_0_312;
   wire n_0_110;
   wire n_0_74;
   wire n_0_75;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_4;
   wire n_0_5;
   wire n_0_7;
   wire n_0_0_318;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_334;
   wire n_0_0_337;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_120;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_358;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_366;
   wire n_0_0_367;
   wire n_0_0_370;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_128;
   wire n_0_0_384;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_0_391;
   wire n_0_0_392;
   wire n_0_0_393;
   wire n_0_0_397;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_0_402;
   wire n_0_0_403;
   wire n_0_0_404;
   wire n_0_0_405;
   wire n_0_0_412;
   wire n_0_0_413;
   wire n_0_0_426;
   wire n_0_0_428;
   wire n_0_0_429;
   wire n_0_0_430;
   wire n_0_0_431;
   wire n_0_0_433;
   wire n_0_0_435;
   wire n_0_0_436;
   wire n_0_0_438;
   wire n_0_0_440;
   wire n_0_0_441;
   wire n_0_0_442;
   wire n_0_0_411;
   wire n_0_0_351;
   wire n_0_0_344;
   wire n_0_0_365;
   wire n_0_0_329;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_117;
   wire n_0_121;
   wire n_0_122;
   wire n_0_124;
   wire n_0_127;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_317;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_348;
   wire n_0_0_371;
   wire n_0_0_386;
   wire n_0_0_387;
   wire n_0_0_395;
   wire n_0_0_396;
   wire n_0_0_406;
   wire n_0_0_417;
   wire n_0_0_408;
   wire n_0_0_437;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_421;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_0_360;
   wire n_0_16;
   wire n_0_126;
   wire n_0_0_377;
   wire n_0_0_425;
   wire n_0_0_427;
   wire n_0_0_359;
   wire n_0_0_434;
   wire n_0_0_368;
   wire n_0_0_443;
   wire n_0_0_394;
   wire n_0_0_444;
   wire n_0_0_445;
   wire n_0_0_414;
   wire n_0_0_415;
   wire n_0_0_446;
   wire n_0_0_416;
   wire n_0_0_447;
   wire n_0_0_448;
   wire n_0_0_449;
   wire n_0_0_450;
   wire n_0_0_369;
   wire n_0_0_361;
   wire n_0_0_451;
   wire n_0_0_452;
   wire n_0_0_418;
   wire n_0_0_453;
   wire n_0_0_454;
   wire n_0_0_455;
   wire n_0_0_456;
   wire n_0_0_457;
   wire n_0_0_458;
   wire n_0_0_459;
   wire n_0_0_460;
   wire n_0_0_461;
   wire n_0_0_385;
   wire n_0_0_372;
   wire n_0_59;
   wire n_0_0_462;
   wire n_0_20;
   wire n_0_113;
   wire n_0_0_463;
   wire n_0_114;
   wire n_0_115;
   wire n_0_118;
   wire n_0_17;
   wire n_0_0_464;
   wire n_0_0_465;
   wire n_0_0_466;
   wire n_0_18;
   wire n_0_0_467;
   wire n_0_0_468;
   wire n_0_0_469;
   wire n_0_0_330;
   wire n_0_0_470;
   wire n_0_0_335;
   wire n_0_19;
   wire n_0_0_471;
   wire n_0_0_472;
   wire n_0_0_473;
   wire n_0_0_474;
   wire n_0_0_475;
   wire n_0_0_383;
   wire n_0_0_476;
   wire n_0_0_477;
   wire n_0_0_478;
   wire n_0_0_479;
   wire n_0_0_480;
   wire n_0_129;
   wire n_0_0_481;
   wire n_0_0_482;
   wire n_0_0_483;
   wire n_0_125;
   wire n_0_0_484;
   wire n_0_0_485;
   wire n_0_0_486;
   wire n_0_0_328;
   wire n_0_0_487;
   wire n_0_0_488;
   wire n_0_0_489;
   wire n_0_0_490;
   wire n_0_0_491;
   wire n_0_0_492;
   wire n_0_0_493;
   wire n_0_0_494;
   wire n_0_123;
   wire n_0_0_495;
   wire n_0_0_496;
   wire n_0_0_497;
   wire n_0_0_498;
   wire n_0_0_499;
   wire n_0_0_500;
   wire n_0_0_501;
   wire n_0_0_502;
   wire n_0_0_503;
   wire n_0_0_333;
   wire n_0_0_504;
   wire n_0_0_505;
   wire n_0_0_506;
   wire n_0_0_507;
   wire n_0_0_508;
   wire n_0_0_509;
   wire n_0_0_510;
   wire n_0_0_511;
   wire n_0_119;
   wire n_0_0_512;
   wire n_0_0_336;
   wire n_0_0_513;
   wire n_0_0_514;
   wire n_0_0_357;
   wire n_0_0_515;
   wire n_0_0_516;
   wire n_0_0_517;
   wire n_0_0_518;
   wire n_0_0_519;
   wire n_0_0_520;
   wire n_0_0_521;
   wire n_0_0_522;
   wire n_0_0_523;
   wire n_0_0_524;
   wire n_0_0_525;
   wire n_0_116;
   wire n_0_0_526;
   wire n_0_0_527;
   wire n_0_0_528;
   wire n_0_0_422;
   wire n_0_0_529;
   wire n_0_0_388;
   wire n_0_0_530;
   wire n_0_0_531;
   wire n_0_0_532;
   wire n_0_0_533;
   wire n_0_0_534;
   wire n_0_0_535;
   wire n_0_0_439;
   wire n_0_0_536;
   wire n_0_0_537;
   wire n_0_0_538;
   wire n_0_0_539;
   wire n_0_0_407;
   wire n_0_0_540;
   wire n_0_0_541;
   wire n_0_0_542;
   wire n_0_0_543;
   wire n_0_0_544;
   wire n_0_0_545;
   wire n_0_0_546;
   wire n_0_0_547;
   wire n_0_0_548;
   wire n_0_0_549;
   wire n_0_0_550;
   wire n_0_0_551;
   wire n_0_0_552;
   wire n_0_0_553;
   wire n_0_0_554;
   wire n_0_0_555;
   wire n_0_0_556;
   wire n_0_0_557;
   wire n_0_0_558;
   wire n_0_0_432;
   wire n_0_0_559;
   wire n_0_0_560;
   wire n_0_111;
   wire n_0_112;

   assign Q[15] = 1'b0;
   assign Q[13] = Q[14];

   INV_X1 cla0_i_5 (.A(divisor[13]), .ZN(cla0_n_0));
   INV_X1 cla0_i_6 (.A(divisor[14]), .ZN(cla0_n_1));
   INV_X1 cla0_i_7 (.A(divisor[15]), .ZN(cla0_n_2));
   INV_X1 cla1_i_5 (.A(dividend[13]), .ZN(cla1_n_0));
   DFF_X1 divideByZero_reg (.D(n_0_113), .CK(n_0_6), .Q(divideByZero), .QN());
   DFF_X1 overFlow_reg (.D(n_0_111), .CK(clk), .Q(overFlow), .QN());
   CLKGATETST_X1 clk_gate_Q_reg (.CK(clk), .E(n_0_110), .SE(1'b0), .GCK(n_0_0));
   DFF_X1 \Q_reg[14]  (.D(n_0_20), .CK(n_0_0), .Q(Q[14]), .QN());
   DFF_X1 \Q_reg[12]  (.D(n_0_73), .CK(n_0_0), .Q(Q[12]), .QN());
   DFF_X1 \Q_reg[11]  (.D(n_0_72), .CK(n_0_0), .Q(Q[11]), .QN());
   DFF_X1 \Q_reg[10]  (.D(n_0_71), .CK(n_0_0), .Q(Q[10]), .QN());
   DFF_X1 \Q_reg[9]  (.D(n_0_70), .CK(n_0_0), .Q(Q[9]), .QN());
   DFF_X1 \Q_reg[8]  (.D(n_0_69), .CK(n_0_0), .Q(Q[8]), .QN());
   DFF_X1 \Q_reg[7]  (.D(n_0_68), .CK(n_0_0), .Q(Q[7]), .QN());
   DFF_X1 \Q_reg[6]  (.D(n_0_67), .CK(n_0_0), .Q(Q[6]), .QN());
   DFF_X1 \Q_reg[5]  (.D(n_0_66), .CK(n_0_0), .Q(Q[5]), .QN());
   DFF_X1 \Q_reg[4]  (.D(n_0_65), .CK(n_0_0), .Q(Q[4]), .QN());
   DFF_X1 \Q_reg[3]  (.D(n_0_64), .CK(n_0_0), .Q(Q[3]), .QN());
   DFF_X1 \Q_reg[2]  (.D(n_0_63), .CK(n_0_0), .Q(Q[2]), .QN());
   DFF_X1 \Q_reg[1]  (.D(n_0_62), .CK(n_0_0), .Q(Q[1]), .QN());
   DFF_X1 \Q_reg[0]  (.D(n_0_61), .CK(n_0_0), .Q(Q[0]), .QN());
   CLKGATETST_X1 clk_gate_A_reg (.CK(clk), .E(n_0_109), .SE(1'b0), .GCK(n_0_1));
   DFF_X1 \A_reg[31]  (.D(n_0_107), .CK(n_0_1), .Q(n_0_21), .QN());
   DFF_X1 \A_reg[30]  (.D(n_0_106), .CK(n_0_1), .Q(n_0_22), .QN());
   DFF_X1 \A_reg[29]  (.D(n_0_105), .CK(n_0_1), .Q(n_0_23), .QN());
   DFF_X1 \A_reg[28]  (.D(n_0_104), .CK(n_0_1), .Q(n_0_24), .QN());
   DFF_X1 \A_reg[27]  (.D(n_0_103), .CK(n_0_1), .Q(n_0_25), .QN());
   DFF_X1 \A_reg[26]  (.D(n_0_102), .CK(n_0_1), .Q(n_0_26), .QN());
   DFF_X1 \A_reg[25]  (.D(n_0_101), .CK(n_0_1), .Q(n_0_27), .QN());
   DFF_X1 \A_reg[24]  (.D(n_0_100), .CK(n_0_1), .Q(n_0_28), .QN());
   DFF_X1 \A_reg[23]  (.D(n_0_99), .CK(n_0_1), .Q(n_0_29), .QN());
   DFF_X1 \A_reg[22]  (.D(n_0_98), .CK(n_0_1), .Q(n_0_30), .QN());
   DFF_X1 \A_reg[21]  (.D(n_0_97), .CK(n_0_1), .Q(n_0_31), .QN());
   DFF_X1 \A_reg[20]  (.D(n_0_96), .CK(n_0_1), .Q(n_0_32), .QN());
   DFF_X1 \A_reg[19]  (.D(n_0_95), .CK(n_0_1), .Q(n_0_33), .QN());
   DFF_X1 \A_reg[18]  (.D(n_0_94), .CK(n_0_1), .Q(n_0_34), .QN());
   DFF_X1 \A_reg[17]  (.D(n_0_93), .CK(n_0_1), .Q(n_0_35), .QN());
   DFF_X1 \A_reg[16]  (.D(n_0_92), .CK(n_0_1), .Q(n_0_36), .QN());
   CLKGATETST_X1 clk_gate_A_reg__15 (.CK(clk), .E(n_0_108), .SE(1'b0), .GCK(
      n_0_2));
   DFF_X1 \A_reg[15]  (.D(n_0_91), .CK(n_0_2), .Q(n_0_37), .QN());
   DFF_X1 \A_reg[14]  (.D(n_0_90), .CK(n_0_2), .Q(n_0_38), .QN());
   DFF_X1 \A_reg[13]  (.D(n_0_89), .CK(n_0_2), .Q(n_0_39), .QN());
   DFF_X1 \A_reg[12]  (.D(n_0_88), .CK(n_0_2), .Q(n_0_40), .QN());
   DFF_X1 \A_reg[11]  (.D(n_0_87), .CK(n_0_2), .Q(n_0_41), .QN());
   DFF_X1 \A_reg[10]  (.D(n_0_86), .CK(n_0_2), .Q(n_0_42), .QN());
   DFF_X1 \A_reg[9]  (.D(n_0_85), .CK(n_0_2), .Q(n_0_43), .QN());
   DFF_X1 \A_reg[8]  (.D(n_0_84), .CK(n_0_2), .Q(n_0_44), .QN());
   DFF_X1 \A_reg[7]  (.D(n_0_83), .CK(n_0_2), .Q(n_0_45), .QN());
   DFF_X1 \A_reg[6]  (.D(n_0_82), .CK(n_0_2), .Q(n_0_46), .QN());
   DFF_X1 \A_reg[5]  (.D(n_0_81), .CK(n_0_2), .Q(n_0_47), .QN());
   DFF_X1 \A_reg[4]  (.D(n_0_80), .CK(n_0_2), .Q(n_0_48), .QN());
   DFF_X1 \A_reg[3]  (.D(n_0_79), .CK(n_0_2), .Q(n_0_49), .QN());
   DFF_X1 \A_reg[2]  (.D(n_0_78), .CK(n_0_2), .Q(n_0_50), .QN());
   DFF_X1 \A_reg[1]  (.D(n_0_77), .CK(n_0_2), .Q(n_0_51), .QN());
   DFF_X1 \A_reg[0]  (.D(n_0_76), .CK(n_0_2), .Q(n_0_52), .QN());
   DFF_X1 \negated_second_operand_number_reg[15]  (.D(n_0_19), .CK(n_0_6), 
      .Q(negated_second_operand_number[15]), .QN());
   DFF_X1 \negated_second_operand_number_reg[14]  (.D(n_0_18), .CK(n_0_6), 
      .Q(negated_second_operand_number[14]), .QN());
   DFF_X1 \negated_second_operand_number_reg[13]  (.D(n_0_17), .CK(n_0_6), 
      .Q(negated_second_operand_number[13]), .QN());
   DFF_X1 \negated_second_operand_number_reg[12]  (.D(n_0_16), .CK(n_0_6), 
      .Q(negated_second_operand_number[12]), .QN());
   DFF_X1 \negated_second_operand_number_reg[11]  (.D(n_0_15), .CK(n_0_6), 
      .Q(negated_second_operand_number[11]), .QN());
   DFF_X1 \negated_second_operand_number_reg[10]  (.D(n_0_14), .CK(n_0_6), 
      .Q(negated_second_operand_number[10]), .QN());
   DFF_X1 \negated_second_operand_number_reg[9]  (.D(n_0_13), .CK(n_0_6), 
      .Q(negated_second_operand_number[9]), .QN());
   DFF_X1 \negated_second_operand_number_reg[8]  (.D(n_0_12), .CK(n_0_6), 
      .Q(negated_second_operand_number[8]), .QN());
   DFF_X1 \negated_second_operand_number_reg[7]  (.D(n_0_11), .CK(n_0_6), 
      .Q(negated_second_operand_number[7]), .QN());
   DFF_X1 \negated_second_operand_number_reg[6]  (.D(n_0_10), .CK(n_0_6), 
      .Q(negated_second_operand_number[6]), .QN());
   DFF_X1 \negated_second_operand_number_reg[5]  (.D(n_0_9), .CK(n_0_6), 
      .Q(negated_second_operand_number[5]), .QN());
   DFF_X1 \negated_second_operand_number_reg[4]  (.D(n_0_8), .CK(n_0_6), 
      .Q(negated_second_operand_number[4]), .QN());
   DFF_X1 \negated_second_operand_number_reg[3]  (.D(n_0_7), .CK(n_0_6), 
      .Q(negated_second_operand_number[3]), .QN());
   DFF_X1 \negated_second_operand_number_reg[2]  (.D(n_0_5), .CK(n_0_6), 
      .Q(negated_second_operand_number[2]), .QN());
   DFF_X1 \negated_second_operand_number_reg[1]  (.D(n_0_4), .CK(n_0_6), 
      .Q(negated_second_operand_number[1]), .QN());
   DFF_X1 \second_operand_number_reg[15]  (.D(n_0_129), .CK(n_0_6), .Q(
      second_operand_number[15]), .QN());
   DFF_X1 \second_operand_number_reg[14]  (.D(n_0_128), .CK(n_0_6), .Q(
      second_operand_number[14]), .QN());
   DFF_X1 \second_operand_number_reg[13]  (.D(n_0_127), .CK(n_0_6), .Q(
      second_operand_number[13]), .QN());
   DFF_X1 \second_operand_number_reg[12]  (.D(n_0_126), .CK(n_0_6), .Q(
      second_operand_number[12]), .QN());
   DFF_X1 \second_operand_number_reg[11]  (.D(n_0_125), .CK(n_0_6), .Q(
      second_operand_number[11]), .QN());
   DFF_X1 \second_operand_number_reg[10]  (.D(n_0_124), .CK(n_0_6), .Q(
      second_operand_number[10]), .QN());
   DFF_X1 \second_operand_number_reg[9]  (.D(n_0_123), .CK(n_0_6), .Q(
      second_operand_number[9]), .QN());
   DFF_X1 \second_operand_number_reg[8]  (.D(n_0_122), .CK(n_0_6), .Q(
      second_operand_number[8]), .QN());
   DFF_X1 \second_operand_number_reg[7]  (.D(n_0_121), .CK(n_0_6), .Q(
      second_operand_number[7]), .QN());
   DFF_X1 \second_operand_number_reg[6]  (.D(n_0_120), .CK(n_0_6), .Q(
      second_operand_number[6]), .QN());
   DFF_X1 \second_operand_number_reg[5]  (.D(n_0_119), .CK(n_0_6), .Q(
      second_operand_number[5]), .QN());
   DFF_X1 \second_operand_number_reg[4]  (.D(n_0_118), .CK(n_0_6), .Q(
      second_operand_number[4]), .QN());
   DFF_X1 \second_operand_number_reg[3]  (.D(n_0_117), .CK(n_0_6), .Q(
      second_operand_number[3]), .QN());
   DFF_X1 \second_operand_number_reg[2]  (.D(n_0_116), .CK(n_0_6), .Q(
      second_operand_number[2]), .QN());
   DFF_X1 \second_operand_number_reg[1]  (.D(n_0_115), .CK(n_0_6), .Q(
      second_operand_number[1]), .QN());
   DFF_X1 ready_reg (.D(n_0_112), .CK(clk), .Q(ready), .QN());
   CLKGATETST_X1 clk_gate_number_of_bits_in_dividend_reg (.CK(clk), .E(n_0_60), 
      .SE(1'b0), .GCK(n_0_3));
   DFF_X1 \number_of_bits_in_dividend_reg[4]  (.D(n_0_59), .CK(n_0_3), .Q(
      number_of_bits_in_dividend[4]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[3]  (.D(n_0_58), .CK(n_0_3), .Q(
      number_of_bits_in_dividend[3]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[2]  (.D(n_0_57), .CK(n_0_3), .Q(
      number_of_bits_in_dividend[2]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[1]  (.D(n_0_56), .CK(n_0_3), .Q(
      number_of_bits_in_dividend[1]), .QN());
   DFF_X1 \number_of_bits_in_dividend_reg[0]  (.D(n_0_55), .CK(n_0_3), .Q(
      number_of_bits_in_dividend[0]), .QN());
   DFF_X1 sign_reg (.D(n_0_54), .CK(n_0_6), .Q(sign), .QN());
   CLKGATETST_X1 clk_gate_divideByZero_reg (.CK(clk), .E(reset), .SE(1'b0), 
      .GCK(n_0_6));
   DFF_X1 \negated_second_operand_number_reg[0]  (.D(n_0_114), .CK(n_0_6), 
      .Q(negated_second_operand_number[0]), .QN());
   XNOR2_X1 i_0_0_0 (.A(n_0_0_437), .B(dividend[12]), .ZN(n_0_54));
   NAND2_X1 i_0_0_1 (.A1(n_0_20), .A2(number_of_bits_in_dividend[0]), .ZN(n_0_55));
   NAND2_X1 i_0_0_2 (.A1(n_0_20), .A2(n_0_0_0), .ZN(n_0_56));
   XOR2_X1 i_0_0_3 (.A(number_of_bits_in_dividend[1]), .B(
      number_of_bits_in_dividend[0]), .Z(n_0_0_0));
   NAND3_X1 i_0_0_4 (.A1(n_0_20), .A2(n_0_0_6), .A3(n_0_0_1), .ZN(n_0_57));
   OAI21_X1 i_0_0_5 (.A(number_of_bits_in_dividend[2]), .B1(
      number_of_bits_in_dividend[1]), .B2(number_of_bits_in_dividend[0]), 
      .ZN(n_0_0_1));
   NAND3_X1 i_0_0_6 (.A1(n_0_20), .A2(n_0_0_5), .A3(n_0_0_2), .ZN(n_0_58));
   NAND2_X1 i_0_0_7 (.A1(n_0_0_6), .A2(number_of_bits_in_dividend[3]), .ZN(
      n_0_0_2));
   OR2_X1 i_0_0_8 (.A1(n_0_0_6), .A2(number_of_bits_in_dividend[3]), .ZN(n_0_0_5));
   OR3_X1 i_0_0_9 (.A1(number_of_bits_in_dividend[2]), .A2(
      number_of_bits_in_dividend[1]), .A3(number_of_bits_in_dividend[0]), 
      .ZN(n_0_0_6));
   AND2_X1 i_0_0_10 (.A1(n_0_20), .A2(n_0_52), .ZN(n_0_61));
   NOR2_X1 i_0_0_11 (.A1(reset), .A2(n_0_0_17), .ZN(n_0_62));
   NOR2_X1 i_0_0_12 (.A1(reset), .A2(n_0_0_19), .ZN(n_0_63));
   NOR2_X1 i_0_0_13 (.A1(reset), .A2(n_0_0_23), .ZN(n_0_64));
   NOR2_X1 i_0_0_14 (.A1(reset), .A2(n_0_0_27), .ZN(n_0_65));
   NOR2_X1 i_0_0_15 (.A1(reset), .A2(n_0_0_32), .ZN(n_0_66));
   AND2_X1 i_0_0_16 (.A1(n_0_20), .A2(n_0_0_36), .ZN(n_0_67));
   NOR2_X1 i_0_0_17 (.A1(reset), .A2(n_0_0_38), .ZN(n_0_68));
   NOR2_X1 i_0_0_18 (.A1(reset), .A2(n_0_0_43), .ZN(n_0_69));
   NOR2_X1 i_0_0_19 (.A1(reset), .A2(n_0_0_48), .ZN(n_0_70));
   NOR2_X1 i_0_0_20 (.A1(reset), .A2(n_0_0_58), .ZN(n_0_71));
   NOR2_X1 i_0_0_21 (.A1(reset), .A2(n_0_0_65), .ZN(n_0_72));
   NOR2_X1 i_0_0_22 (.A1(reset), .A2(n_0_0_71), .ZN(n_0_73));
   NAND2_X1 i_0_0_23 (.A1(n_0_20), .A2(n_0_0_314), .ZN(n_0_53));
   OAI21_X1 i_0_0_24 (.A(n_0_0_7), .B1(n_0_0_12), .B2(n_0_0_264), .ZN(n_0_76));
   AOI22_X1 i_0_0_25 (.A1(n_0_0_8), .A2(n_0_0_309), .B1(n_0_52), .B2(n_0_0_96), 
      .ZN(n_0_0_7));
   XNOR2_X1 i_0_0_26 (.A(negated_second_operand_number[15]), .B(n_0_0_9), 
      .ZN(n_0_0_8));
   OAI21_X1 i_0_0_27 (.A(n_0_0_11), .B1(n_0_0_267), .B2(n_0_0_10), .ZN(n_0_0_9));
   NOR2_X1 i_0_0_28 (.A1(n_0_22), .A2(negated_second_operand_number[14]), 
      .ZN(n_0_0_10));
   NAND2_X1 i_0_0_29 (.A1(n_0_22), .A2(negated_second_operand_number[14]), 
      .ZN(n_0_0_11));
   XNOR2_X1 i_0_0_30 (.A(second_operand_number[15]), .B(n_0_0_13), .ZN(n_0_0_12));
   OAI21_X1 i_0_0_31 (.A(n_0_0_14), .B1(n_0_0_227), .B2(n_0_0_15), .ZN(n_0_0_13));
   NAND2_X1 i_0_0_32 (.A1(n_0_22), .A2(second_operand_number[14]), .ZN(n_0_0_14));
   NOR2_X1 i_0_0_33 (.A1(n_0_22), .A2(second_operand_number[14]), .ZN(n_0_0_15));
   OAI21_X1 i_0_0_34 (.A(n_0_0_16), .B1(n_0_0_95), .B2(n_0_0_17), .ZN(n_0_77));
   NAND2_X1 i_0_0_35 (.A1(n_0_52), .A2(n_0_0_311), .ZN(n_0_0_16));
   XOR2_X1 i_0_0_36 (.A(n_0_51), .B(n_0_0_21), .Z(n_0_0_17));
   OAI21_X1 i_0_0_37 (.A(n_0_0_18), .B1(n_0_0_95), .B2(n_0_0_19), .ZN(n_0_78));
   NAND2_X1 i_0_0_38 (.A1(n_0_51), .A2(n_0_0_311), .ZN(n_0_0_18));
   XOR2_X1 i_0_0_39 (.A(n_0_50), .B(n_0_0_20), .Z(n_0_0_19));
   NAND2_X1 i_0_0_40 (.A1(n_0_0_82), .A2(sign), .ZN(n_0_0_20));
   NAND2_X1 i_0_0_41 (.A1(n_0_52), .A2(sign), .ZN(n_0_0_21));
   OAI21_X1 i_0_0_42 (.A(n_0_0_22), .B1(n_0_0_95), .B2(n_0_0_23), .ZN(n_0_79));
   NAND2_X1 i_0_0_43 (.A1(n_0_50), .A2(n_0_0_311), .ZN(n_0_0_22));
   OAI211_X1 i_0_0_44 (.A(n_0_0_81), .B(n_0_0_24), .C1(n_0_49), .C2(sign), 
      .ZN(n_0_0_23));
   OAI211_X1 i_0_0_45 (.A(n_0_49), .B(sign), .C1(n_0_0_82), .C2(n_0_50), 
      .ZN(n_0_0_24));
   INV_X1 i_0_0_46 (.A(n_0_0_25), .ZN(n_0_80));
   AOI221_X1 i_0_0_47 (.A(n_0_0_26), .B1(n_0_0_107), .B2(dividend[0]), .C1(
      n_0_49), .C2(n_0_0_311), .ZN(n_0_0_25));
   NOR2_X1 i_0_0_48 (.A1(n_0_0_27), .A2(n_0_0_95), .ZN(n_0_0_26));
   XOR2_X1 i_0_0_49 (.A(n_0_48), .B(n_0_0_28), .Z(n_0_0_27));
   NAND2_X1 i_0_0_50 (.A1(n_0_0_81), .A2(sign), .ZN(n_0_0_28));
   OAI211_X1 i_0_0_51 (.A(n_0_0_29), .B(n_0_0_31), .C1(n_0_0_32), .C2(n_0_0_95), 
      .ZN(n_0_81));
   AOI22_X1 i_0_0_52 (.A1(n_0_48), .A2(n_0_0_311), .B1(n_0_0_119), .B2(n_0_0_30), 
      .ZN(n_0_0_29));
   AND2_X1 i_0_0_53 (.A1(dividend[0]), .A2(n_0_0_127), .ZN(n_0_0_30));
   NAND2_X1 i_0_0_54 (.A1(n_0_0_107), .A2(n_0_0_69), .ZN(n_0_0_31));
   OAI211_X1 i_0_0_55 (.A(n_0_0_80), .B(n_0_0_33), .C1(n_0_47), .C2(sign), 
      .ZN(n_0_0_32));
   OAI211_X1 i_0_0_56 (.A(n_0_47), .B(sign), .C1(n_0_0_81), .C2(n_0_48), 
      .ZN(n_0_0_33));
   OAI211_X1 i_0_0_60 (.A(n_0_0_34), .B(n_0_0_35), .C1(n_0_0_40), .C2(n_0_0_116), 
      .ZN(n_0_82));
   AOI222_X1 i_0_0_61 (.A1(n_0_0_36), .A2(n_0_0_96), .B1(n_0_0_107), .B2(
      n_0_0_86), .C1(n_0_47), .C2(n_0_0_311), .ZN(n_0_0_34));
   NAND3_X1 i_0_0_62 (.A1(n_0_0_127), .A2(n_0_0_119), .A3(n_0_0_69), .ZN(
      n_0_0_35));
   XNOR2_X1 i_0_0_57 (.A(n_0_46), .B(n_0_0_79), .ZN(n_0_0_36));
   OAI221_X1 i_0_0_64 (.A(n_0_0_37), .B1(n_0_0_38), .B2(n_0_0_95), .C1(n_0_0_118), 
      .C2(n_0_0_40), .ZN(n_0_83));
   AOI221_X1 i_0_0_65 (.A(n_0_0_41), .B1(n_0_0_92), .B2(n_0_0_107), .C1(n_0_46), 
      .C2(n_0_0_311), .ZN(n_0_0_37));
   XOR2_X1 i_0_0_58 (.A(n_0_45), .B(n_0_0_39), .Z(n_0_0_38));
   OAI21_X1 i_0_0_59 (.A(sign), .B1(n_0_0_80), .B2(n_0_46), .ZN(n_0_0_39));
   AOI22_X1 i_0_0_68 (.A1(n_0_0_127), .A2(n_0_0_86), .B1(n_0_0_57), .B2(
      dividend[0]), .ZN(n_0_0_40));
   NOR2_X1 i_0_0_69 (.A1(n_0_0_116), .A2(n_0_0_47), .ZN(n_0_0_41));
   OAI211_X1 i_0_0_70 (.A(n_0_0_45), .B(n_0_0_42), .C1(n_0_0_43), .C2(n_0_0_95), 
      .ZN(n_0_84));
   NAND2_X1 i_0_0_71 (.A1(n_0_0_107), .A2(n_0_0_103), .ZN(n_0_0_42));
   OAI211_X1 i_0_0_63 (.A(n_0_0_76), .B(n_0_0_44), .C1(n_0_44), .C2(sign), 
      .ZN(n_0_0_43));
   NAND3_X1 i_0_0_66 (.A1(n_0_0_77), .A2(sign), .A3(n_0_44), .ZN(n_0_0_44));
   AOI21_X1 i_0_0_74 (.A(n_0_0_46), .B1(n_0_0_311), .B2(n_0_45), .ZN(n_0_0_45));
   OAI22_X1 i_0_0_75 (.A1(n_0_0_52), .A2(n_0_0_116), .B1(n_0_0_118), .B2(
      n_0_0_47), .ZN(n_0_0_46));
   AOI22_X1 i_0_0_76 (.A1(n_0_0_127), .A2(n_0_0_92), .B1(n_0_0_57), .B2(n_0_0_69), 
      .ZN(n_0_0_47));
   OAI221_X1 i_0_0_77 (.A(n_0_0_50), .B1(n_0_0_48), .B2(n_0_0_95), .C1(n_0_0_56), 
      .C2(n_0_0_116), .ZN(n_0_85));
   OAI211_X1 i_0_0_67 (.A(n_0_0_75), .B(n_0_0_49), .C1(n_0_43), .C2(sign), 
      .ZN(n_0_0_48));
   NAND3_X1 i_0_0_72 (.A1(n_0_0_76), .A2(sign), .A3(n_0_43), .ZN(n_0_0_49));
   AOI221_X1 i_0_0_80 (.A(n_0_0_51), .B1(n_0_0_107), .B2(n_0_0_138), .C1(n_0_44), 
      .C2(n_0_0_311), .ZN(n_0_0_50));
   NOR2_X1 i_0_0_81 (.A1(n_0_0_52), .A2(n_0_0_118), .ZN(n_0_0_51));
   AOI22_X1 i_0_0_82 (.A1(n_0_0_151), .A2(n_0_0_63), .B1(n_0_0_57), .B2(n_0_0_86), 
      .ZN(n_0_0_52));
   OAI21_X1 i_0_0_83 (.A(n_0_0_53), .B1(n_0_0_58), .B2(n_0_0_95), .ZN(n_0_86));
   AOI21_X1 i_0_0_84 (.A(n_0_0_54), .B1(n_0_0_62), .B2(n_0_0_117), .ZN(n_0_0_53));
   OAI21_X1 i_0_0_85 (.A(n_0_0_55), .B1(n_0_0_56), .B2(n_0_0_118), .ZN(n_0_0_54));
   AOI22_X1 i_0_0_86 (.A1(n_0_0_112), .A2(n_0_0_107), .B1(n_0_43), .B2(n_0_0_311), 
      .ZN(n_0_0_55));
   AOI22_X1 i_0_0_87 (.A1(n_0_0_151), .A2(n_0_0_68), .B1(n_0_0_57), .B2(n_0_0_92), 
      .ZN(n_0_0_56));
   NOR2_X1 i_0_0_88 (.A1(n_0_0_151), .A2(n_0_0_148), .ZN(n_0_0_57));
   XOR2_X1 i_0_0_73 (.A(n_0_42), .B(n_0_0_59), .Z(n_0_0_58));
   NAND2_X1 i_0_0_78 (.A1(n_0_0_75), .A2(sign), .ZN(n_0_0_59));
   OAI211_X1 i_0_0_91 (.A(n_0_0_61), .B(n_0_0_60), .C1(n_0_0_95), .C2(n_0_0_65), 
      .ZN(n_0_87));
   NAND2_X1 i_0_0_92 (.A1(n_0_0_67), .A2(n_0_0_117), .ZN(n_0_0_60));
   AOI222_X1 i_0_0_93 (.A1(n_0_0_119), .A2(n_0_0_62), .B1(n_0_0_107), .B2(
      n_0_0_130), .C1(n_0_42), .C2(n_0_0_311), .ZN(n_0_0_61));
   MUX2_X1 i_0_0_94 (.A(n_0_0_63), .B(n_0_0_85), .S(n_0_0_151), .Z(n_0_0_62));
   OAI21_X1 i_0_0_95 (.A(n_0_0_64), .B1(n_0_0_102), .B2(n_0_0_148), .ZN(n_0_0_63));
   NAND2_X1 i_0_0_96 (.A1(dividend[0]), .A2(n_0_0_148), .ZN(n_0_0_64));
   XOR2_X1 i_0_0_79 (.A(n_0_41), .B(n_0_0_74), .Z(n_0_0_65));
   OAI221_X1 i_0_0_98 (.A(n_0_0_66), .B1(n_0_0_71), .B2(n_0_0_95), .C1(n_0_0_116), 
      .C2(n_0_0_83), .ZN(n_0_88));
   AOI222_X1 i_0_0_89 (.A1(n_0_0_119), .A2(n_0_0_67), .B1(n_0_0_107), .B2(
      n_0_0_109), .C1(n_0_0_311), .C2(n_0_41), .ZN(n_0_0_66));
   MUX2_X1 i_0_0_90 (.A(n_0_0_68), .B(n_0_0_91), .S(n_0_0_151), .Z(n_0_0_67));
   MUX2_X1 i_0_0_97 (.A(n_0_0_138), .B(n_0_0_69), .S(n_0_0_148), .Z(n_0_0_68));
   XNOR2_X1 i_0_0_99 (.A(dividend[1]), .B(n_0_0_70), .ZN(n_0_0_69));
   NAND2_X1 i_0_0_100 (.A1(dividend[12]), .A2(dividend[0]), .ZN(n_0_0_70));
   XNOR2_X1 i_0_0_101 (.A(n_0_40), .B(n_0_0_72), .ZN(n_0_0_71));
   NAND2_X1 i_0_0_102 (.A1(n_0_0_74), .A2(n_0_0_73), .ZN(n_0_0_72));
   NAND2_X1 i_0_0_103 (.A1(n_0_41), .A2(sign), .ZN(n_0_0_73));
   OAI21_X1 i_0_0_104 (.A(sign), .B1(n_0_0_75), .B2(n_0_42), .ZN(n_0_0_74));
   OR2_X1 i_0_0_105 (.A1(n_0_0_76), .A2(n_0_43), .ZN(n_0_0_75));
   OR2_X1 i_0_0_106 (.A1(n_0_0_77), .A2(n_0_44), .ZN(n_0_0_76));
   NAND2_X1 i_0_0_107 (.A1(n_0_0_79), .A2(n_0_0_78), .ZN(n_0_0_77));
   NOR2_X1 i_0_0_108 (.A1(n_0_45), .A2(n_0_46), .ZN(n_0_0_78));
   NAND2_X1 i_0_0_109 (.A1(n_0_0_80), .A2(sign), .ZN(n_0_0_79));
   OR3_X1 i_0_0_110 (.A1(n_0_0_81), .A2(n_0_48), .A3(n_0_47), .ZN(n_0_0_80));
   OR3_X1 i_0_0_111 (.A1(n_0_0_82), .A2(n_0_50), .A3(n_0_49), .ZN(n_0_0_81));
   OR2_X1 i_0_0_112 (.A1(n_0_51), .A2(n_0_52), .ZN(n_0_0_82));
   OAI221_X1 i_0_0_116 (.A(n_0_0_88), .B1(n_0_0_83), .B2(n_0_0_118), .C1(
      n_0_0_89), .C2(n_0_0_116), .ZN(n_0_89));
   AOI21_X1 i_0_0_117 (.A(n_0_0_84), .B1(n_0_0_85), .B2(n_0_0_150), .ZN(n_0_0_83));
   NOR2_X1 i_0_0_118 (.A1(n_0_0_150), .A2(n_0_0_100), .ZN(n_0_0_84));
   MUX2_X1 i_0_0_119 (.A(n_0_0_112), .B(n_0_0_86), .S(n_0_0_148), .Z(n_0_0_85));
   XNOR2_X1 i_0_0_120 (.A(dividend[2]), .B(n_0_0_87), .ZN(n_0_0_86));
   NAND2_X1 i_0_0_121 (.A1(n_0_0_147), .A2(dividend[12]), .ZN(n_0_0_87));
   AOI221_X1 i_0_0_122 (.A(n_0_0_96), .B1(n_0_0_311), .B2(n_0_40), .C1(n_0_0_140), 
      .C2(n_0_0_107), .ZN(n_0_0_88));
   OAI221_X1 i_0_0_123 (.A(n_0_0_94), .B1(n_0_0_89), .B2(n_0_0_118), .C1(
      n_0_0_98), .C2(n_0_0_116), .ZN(n_0_90));
   AOI21_X1 i_0_0_124 (.A(n_0_0_90), .B1(n_0_0_91), .B2(n_0_0_150), .ZN(n_0_0_89));
   NOR2_X1 i_0_0_125 (.A1(n_0_0_150), .A2(n_0_0_135), .ZN(n_0_0_90));
   MUX2_X1 i_0_0_113 (.A(n_0_0_130), .B(n_0_0_92), .S(n_0_0_148), .Z(n_0_0_91));
   XNOR2_X1 i_0_0_114 (.A(dividend[3]), .B(n_0_0_93), .ZN(n_0_0_92));
   OAI21_X1 i_0_0_115 (.A(dividend[12]), .B1(n_0_0_147), .B2(dividend[2]), 
      .ZN(n_0_0_93));
   AOI221_X1 i_0_0_129 (.A(n_0_0_96), .B1(n_0_0_311), .B2(n_0_39), .C1(n_0_0_114), 
      .C2(n_0_0_107), .ZN(n_0_0_94));
   NAND2_X1 i_0_0_126 (.A1(n_0_0_313), .A2(n_0_0_222), .ZN(n_0_0_95));
   NOR3_X1 i_0_0_127 (.A1(n_0_60), .A2(ready), .A3(n_0_0_442), .ZN(n_0_0_96));
   OAI221_X1 i_0_0_132 (.A(n_0_0_97), .B1(n_0_0_98), .B2(n_0_0_118), .C1(
      n_0_0_124), .C2(n_0_0_116), .ZN(n_0_91));
   AOI22_X1 i_0_0_133 (.A1(n_0_0_132), .A2(n_0_0_107), .B1(n_0_38), .B2(
      n_0_0_311), .ZN(n_0_0_97));
   AOI21_X1 i_0_0_134 (.A(n_0_0_99), .B1(n_0_0_111), .B2(n_0_0_151), .ZN(
      n_0_0_98));
   NOR2_X1 i_0_0_135 (.A1(n_0_0_100), .A2(n_0_0_151), .ZN(n_0_0_99));
   OAI21_X1 i_0_0_136 (.A(n_0_0_101), .B1(n_0_0_109), .B2(n_0_0_148), .ZN(
      n_0_0_100));
   NAND2_X1 i_0_0_137 (.A1(n_0_0_148), .A2(n_0_0_102), .ZN(n_0_0_101));
   INV_X1 i_0_0_138 (.A(n_0_0_103), .ZN(n_0_0_102));
   XNOR2_X1 i_0_0_139 (.A(dividend[4]), .B(n_0_0_104), .ZN(n_0_0_103));
   NAND2_X1 i_0_0_140 (.A1(n_0_0_146), .A2(dividend[12]), .ZN(n_0_0_104));
   OAI211_X1 i_0_0_141 (.A(n_0_0_108), .B(n_0_0_105), .C1(n_0_0_124), .C2(
      n_0_0_118), .ZN(n_0_92));
   AOI221_X1 i_0_0_128 (.A(n_0_0_106), .B1(n_0_0_311), .B2(n_0_37), .C1(n_0_35), 
      .C2(n_0_0_222), .ZN(n_0_0_105));
   AND4_X1 i_0_0_130 (.A1(dividend[12]), .A2(n_0_0_134), .A3(n_0_0_107), 
      .A4(n_0_0_430), .ZN(n_0_0_106));
   AOI21_X1 i_0_0_131 (.A(n_0_20), .B1(n_0_0_120), .B2(n_0_0_422), .ZN(n_0_0_107));
   OAI221_X1 i_0_0_142 (.A(n_0_0_117), .B1(n_0_0_109), .B2(n_0_0_126), .C1(
      n_0_0_111), .C2(n_0_0_151), .ZN(n_0_0_108));
   XNOR2_X1 i_0_0_143 (.A(dividend[8]), .B(n_0_0_110), .ZN(n_0_0_109));
   NAND2_X1 i_0_0_144 (.A1(n_0_0_143), .A2(dividend[12]), .ZN(n_0_0_110));
   MUX2_X1 i_0_0_145 (.A(n_0_0_114), .B(n_0_0_112), .S(n_0_0_148), .Z(n_0_0_111));
   XNOR2_X1 i_0_0_146 (.A(dividend[6]), .B(n_0_0_113), .ZN(n_0_0_112));
   NAND2_X1 i_0_0_147 (.A1(n_0_0_144), .A2(dividend[12]), .ZN(n_0_0_113));
   XNOR2_X1 i_0_0_148 (.A(dividend[10]), .B(n_0_0_115), .ZN(n_0_0_114));
   OAI21_X1 i_0_0_149 (.A(dividend[12]), .B1(n_0_0_142), .B2(dividend[9]), 
      .ZN(n_0_0_115));
   NAND4_X1 i_0_0_153 (.A1(n_0_0_120), .A2(n_0_0_422), .A3(reset), .A4(n_0_0_122), 
      .ZN(n_0_0_116));
   NOR3_X1 i_0_0_150 (.A1(n_0_0_121), .A2(n_0_0_123), .A3(n_0_0_127), .ZN(
      n_0_0_117));
   NAND3_X1 i_0_0_155 (.A1(reset), .A2(n_0_0_422), .A3(n_0_0_123), .ZN(n_0_0_118));
   NOR2_X1 i_0_0_151 (.A1(n_0_0_122), .A2(n_0_0_121), .ZN(n_0_0_119));
   NAND2_X1 i_0_0_152 (.A1(n_0_0_127), .A2(n_0_0_122), .ZN(n_0_0_120));
   NAND2_X1 i_0_0_154 (.A1(reset), .A2(n_0_0_422), .ZN(n_0_0_121));
   INV_X1 i_0_0_156 (.A(n_0_0_123), .ZN(n_0_0_122));
   XNOR2_X1 i_0_0_157 (.A(divisor[13]), .B(cla1_n_0), .ZN(n_0_0_123));
   AOI211_X1 i_0_0_161 (.A(n_0_0_128), .B(n_0_0_125), .C1(n_0_0_127), .C2(
      n_0_0_132), .ZN(n_0_0_124));
   NOR2_X1 i_0_0_162 (.A1(n_0_0_129), .A2(n_0_0_126), .ZN(n_0_0_125));
   NAND2_X1 i_0_0_158 (.A1(n_0_0_151), .A2(n_0_0_148), .ZN(n_0_0_126));
   NOR2_X1 i_0_0_159 (.A1(n_0_0_150), .A2(n_0_0_148), .ZN(n_0_0_127));
   NOR2_X1 i_0_0_165 (.A1(n_0_0_135), .A2(n_0_0_151), .ZN(n_0_0_128));
   INV_X1 i_0_0_166 (.A(n_0_0_130), .ZN(n_0_0_129));
   XNOR2_X1 i_0_0_160 (.A(dividend[7]), .B(n_0_0_131), .ZN(n_0_0_130));
   OAI21_X1 i_0_0_163 (.A(dividend[12]), .B1(n_0_0_144), .B2(dividend[6]), 
      .ZN(n_0_0_131));
   XNOR2_X1 i_0_0_169 (.A(n_0_0_430), .B(n_0_0_133), .ZN(n_0_0_132));
   NOR2_X1 i_0_0_170 (.A1(n_0_0_134), .A2(n_0_0_431), .ZN(n_0_0_133));
   NOR3_X1 i_0_0_164 (.A1(n_0_0_142), .A2(dividend[9]), .A3(dividend[10]), 
      .ZN(n_0_0_134));
   OAI21_X1 i_0_0_172 (.A(n_0_0_136), .B1(n_0_0_140), .B2(n_0_0_148), .ZN(
      n_0_0_135));
   NAND2_X1 i_0_0_173 (.A1(n_0_0_148), .A2(n_0_0_137), .ZN(n_0_0_136));
   INV_X1 i_0_0_174 (.A(n_0_0_138), .ZN(n_0_0_137));
   XNOR2_X1 i_0_0_167 (.A(dividend[5]), .B(n_0_0_139), .ZN(n_0_0_138));
   NAND2_X1 i_0_0_168 (.A1(n_0_0_145), .A2(dividend[12]), .ZN(n_0_0_139));
   XNOR2_X1 i_0_0_177 (.A(dividend[9]), .B(n_0_0_141), .ZN(n_0_0_140));
   NAND2_X1 i_0_0_178 (.A1(n_0_0_142), .A2(dividend[12]), .ZN(n_0_0_141));
   OR2_X1 i_0_0_171 (.A1(n_0_0_143), .A2(dividend[8]), .ZN(n_0_0_142));
   OR3_X1 i_0_0_175 (.A1(n_0_0_144), .A2(dividend[6]), .A3(dividend[7]), 
      .ZN(n_0_0_143));
   OR2_X1 i_0_0_176 (.A1(n_0_0_145), .A2(dividend[5]), .ZN(n_0_0_144));
   OR2_X1 i_0_0_179 (.A1(n_0_0_146), .A2(dividend[4]), .ZN(n_0_0_145));
   OR3_X1 i_0_0_180 (.A1(n_0_0_147), .A2(dividend[2]), .A3(dividend[3]), 
      .ZN(n_0_0_146));
   OR2_X1 i_0_0_181 (.A1(dividend[1]), .A2(dividend[0]), .ZN(n_0_0_147));
   XNOR2_X1 i_0_0_182 (.A(n_0_0_440), .B(n_0_0_149), .ZN(n_0_0_148));
   OAI21_X1 i_0_0_183 (.A(n_0_0_153), .B1(n_0_0_154), .B2(n_0_0_426), .ZN(
      n_0_0_149));
   INV_X1 i_0_0_184 (.A(n_0_0_151), .ZN(n_0_0_150));
   XNOR2_X1 i_0_0_185 (.A(n_0_0_154), .B(n_0_0_152), .ZN(n_0_0_151));
   XNOR2_X1 i_0_0_186 (.A(divisor[14]), .B(n_0_0_432), .ZN(n_0_0_152));
   NAND2_X1 i_0_0_187 (.A1(n_0_0_432), .A2(divisor[14]), .ZN(n_0_0_153));
   NOR2_X1 i_0_0_188 (.A1(divisor[13]), .A2(cla1_n_0), .ZN(n_0_0_154));
   INV_X1 i_0_0_192 (.A(n_0_0_155), .ZN(n_0_93));
   AOI22_X1 i_0_0_193 (.A1(n_0_34), .A2(n_0_0_222), .B1(n_0_0_156), .B2(
      n_0_0_311), .ZN(n_0_0_155));
   XOR2_X1 i_0_0_194 (.A(n_0_36), .B(negated_second_operand_number[0]), .Z(
      n_0_0_156));
   INV_X1 i_0_0_195 (.A(n_0_0_157), .ZN(n_0_94));
   AOI22_X1 i_0_0_196 (.A1(n_0_0_311), .A2(n_0_0_158), .B1(n_0_0_222), .B2(
      n_0_33), .ZN(n_0_0_157));
   XNOR2_X1 i_0_0_197 (.A(n_0_0_160), .B(n_0_0_159), .ZN(n_0_0_158));
   XNOR2_X1 i_0_0_198 (.A(n_0_35), .B(n_0_0_305), .ZN(n_0_0_159));
   AOI21_X1 i_0_0_199 (.A(n_0_0_161), .B1(second_operand_number[1]), .B2(n_0_21), 
      .ZN(n_0_0_160));
   NOR2_X1 i_0_0_200 (.A1(n_0_0_428), .A2(n_0_21), .ZN(n_0_0_161));
   INV_X1 i_0_0_201 (.A(n_0_0_162), .ZN(n_0_95));
   AOI22_X1 i_0_0_202 (.A1(n_0_0_163), .A2(n_0_0_311), .B1(n_0_32), .B2(
      n_0_0_222), .ZN(n_0_0_162));
   XNOR2_X1 i_0_0_203 (.A(n_0_34), .B(n_0_0_164), .ZN(n_0_0_163));
   AOI21_X1 i_0_0_204 (.A(n_0_0_165), .B1(n_0_0_167), .B2(n_0_21), .ZN(n_0_0_164));
   NOR2_X1 i_0_0_205 (.A1(n_0_21), .A2(n_0_0_166), .ZN(n_0_0_165));
   XNOR2_X1 i_0_0_189 (.A(negated_second_operand_number[2]), .B(n_0_0_302), 
      .ZN(n_0_0_166));
   XOR2_X1 i_0_0_207 (.A(second_operand_number[2]), .B(n_0_0_261), .Z(n_0_0_167));
   OAI21_X1 i_0_0_190 (.A(n_0_0_168), .B1(n_0_0_171), .B2(n_0_0_264), .ZN(n_0_96));
   AOI22_X1 i_0_0_191 (.A1(n_0_0_169), .A2(n_0_0_309), .B1(n_0_31), .B2(
      n_0_0_222), .ZN(n_0_0_168));
   XNOR2_X1 i_0_0_206 (.A(n_0_0_300), .B(n_0_0_170), .ZN(n_0_0_169));
   XNOR2_X1 i_0_0_208 (.A(n_0_33), .B(negated_second_operand_number[3]), 
      .ZN(n_0_0_170));
   XNOR2_X1 i_0_0_209 (.A(n_0_0_259), .B(n_0_0_172), .ZN(n_0_0_171));
   XOR2_X1 i_0_0_210 (.A(n_0_33), .B(second_operand_number[3]), .Z(n_0_0_172));
   OAI21_X1 i_0_0_211 (.A(n_0_0_173), .B1(n_0_0_176), .B2(n_0_0_308), .ZN(n_0_97));
   AOI22_X1 i_0_0_212 (.A1(n_0_0_174), .A2(n_0_0_265), .B1(n_0_30), .B2(
      n_0_0_222), .ZN(n_0_0_173));
   XNOR2_X1 i_0_0_213 (.A(n_0_0_256), .B(n_0_0_175), .ZN(n_0_0_174));
   XOR2_X1 i_0_0_214 (.A(n_0_32), .B(second_operand_number[4]), .Z(n_0_0_175));
   XNOR2_X1 i_0_0_215 (.A(n_0_0_297), .B(n_0_0_177), .ZN(n_0_0_176));
   XNOR2_X1 i_0_0_216 (.A(n_0_32), .B(negated_second_operand_number[4]), 
      .ZN(n_0_0_177));
   OAI21_X1 i_0_0_217 (.A(n_0_0_178), .B1(n_0_0_181), .B2(n_0_0_308), .ZN(n_0_98));
   AOI22_X1 i_0_0_218 (.A1(n_0_0_179), .A2(n_0_0_265), .B1(n_0_29), .B2(
      n_0_0_222), .ZN(n_0_0_178));
   XNOR2_X1 i_0_0_219 (.A(n_0_0_252), .B(n_0_0_180), .ZN(n_0_0_179));
   XNOR2_X1 i_0_0_220 (.A(n_0_31), .B(second_operand_number[5]), .ZN(n_0_0_180));
   XNOR2_X1 i_0_0_221 (.A(n_0_0_293), .B(n_0_0_182), .ZN(n_0_0_181));
   XNOR2_X1 i_0_0_222 (.A(n_0_31), .B(negated_second_operand_number[5]), 
      .ZN(n_0_0_182));
   OAI21_X1 i_0_0_226 (.A(n_0_0_183), .B1(n_0_0_184), .B2(n_0_0_308), .ZN(n_0_99));
   AOI22_X1 i_0_0_227 (.A1(n_0_0_186), .A2(n_0_0_265), .B1(n_0_28), .B2(
      n_0_0_222), .ZN(n_0_0_183));
   XNOR2_X1 i_0_0_228 (.A(n_0_0_291), .B(n_0_0_185), .ZN(n_0_0_184));
   XOR2_X1 i_0_0_229 (.A(n_0_30), .B(negated_second_operand_number[6]), .Z(
      n_0_0_185));
   XNOR2_X1 i_0_0_230 (.A(n_0_0_250), .B(n_0_0_187), .ZN(n_0_0_186));
   XNOR2_X1 i_0_0_231 (.A(n_0_30), .B(second_operand_number[6]), .ZN(n_0_0_187));
   OAI21_X1 i_0_0_232 (.A(n_0_0_188), .B1(n_0_0_189), .B2(n_0_0_264), .ZN(
      n_0_100));
   AOI22_X1 i_0_0_233 (.A1(n_0_0_191), .A2(n_0_0_309), .B1(n_0_27), .B2(
      n_0_0_222), .ZN(n_0_0_188));
   XNOR2_X1 i_0_0_234 (.A(n_0_0_247), .B(n_0_0_190), .ZN(n_0_0_189));
   XNOR2_X1 i_0_0_235 (.A(n_0_29), .B(second_operand_number[7]), .ZN(n_0_0_190));
   XNOR2_X1 i_0_0_236 (.A(n_0_0_288), .B(n_0_0_192), .ZN(n_0_0_191));
   XOR2_X1 i_0_0_237 (.A(n_0_29), .B(negated_second_operand_number[7]), .Z(
      n_0_0_192));
   INV_X1 i_0_0_238 (.A(n_0_0_193), .ZN(n_0_101));
   AOI22_X1 i_0_0_239 (.A1(n_0_0_194), .A2(n_0_0_311), .B1(n_0_26), .B2(
      n_0_0_222), .ZN(n_0_0_193));
   XNOR2_X1 i_0_0_240 (.A(n_0_28), .B(n_0_0_195), .ZN(n_0_0_194));
   AOI21_X1 i_0_0_241 (.A(n_0_0_196), .B1(n_0_0_198), .B2(n_0_21), .ZN(n_0_0_195));
   NOR2_X1 i_0_0_242 (.A1(n_0_21), .A2(n_0_0_197), .ZN(n_0_0_196));
   XNOR2_X1 i_0_0_243 (.A(negated_second_operand_number[8]), .B(n_0_0_285), 
      .ZN(n_0_0_197));
   XOR2_X1 i_0_0_244 (.A(second_operand_number[8]), .B(n_0_0_244), .Z(n_0_0_198));
   OAI21_X1 i_0_0_245 (.A(n_0_0_199), .B1(n_0_0_202), .B2(n_0_0_308), .ZN(
      n_0_102));
   AOI22_X1 i_0_0_246 (.A1(n_0_0_200), .A2(n_0_0_265), .B1(n_0_25), .B2(
      n_0_0_222), .ZN(n_0_0_199));
   XNOR2_X1 i_0_0_247 (.A(n_0_0_241), .B(n_0_0_201), .ZN(n_0_0_200));
   XOR2_X1 i_0_0_248 (.A(n_0_27), .B(second_operand_number[9]), .Z(n_0_0_201));
   XNOR2_X1 i_0_0_249 (.A(n_0_0_282), .B(n_0_0_203), .ZN(n_0_0_202));
   XNOR2_X1 i_0_0_250 (.A(n_0_27), .B(negated_second_operand_number[9]), 
      .ZN(n_0_0_203));
   OAI21_X1 i_0_0_251 (.A(n_0_0_204), .B1(n_0_0_207), .B2(n_0_0_264), .ZN(
      n_0_103));
   AOI22_X1 i_0_0_252 (.A1(n_0_0_205), .A2(n_0_0_309), .B1(n_0_24), .B2(
      n_0_0_222), .ZN(n_0_0_204));
   XNOR2_X1 i_0_0_253 (.A(n_0_0_278), .B(n_0_0_206), .ZN(n_0_0_205));
   XNOR2_X1 i_0_0_254 (.A(n_0_26), .B(negated_second_operand_number[10]), 
      .ZN(n_0_0_206));
   XNOR2_X1 i_0_0_255 (.A(n_0_0_238), .B(n_0_0_208), .ZN(n_0_0_207));
   XOR2_X1 i_0_0_256 (.A(n_0_26), .B(second_operand_number[10]), .Z(n_0_0_208));
   OAI21_X1 i_0_0_257 (.A(n_0_0_209), .B1(n_0_0_212), .B2(n_0_0_264), .ZN(
      n_0_104));
   AOI22_X1 i_0_0_258 (.A1(n_0_0_210), .A2(n_0_0_309), .B1(n_0_23), .B2(
      n_0_0_222), .ZN(n_0_0_209));
   XNOR2_X1 i_0_0_259 (.A(n_0_0_276), .B(n_0_0_211), .ZN(n_0_0_210));
   XNOR2_X1 i_0_0_260 (.A(n_0_25), .B(negated_second_operand_number[11]), 
      .ZN(n_0_0_211));
   XNOR2_X1 i_0_0_261 (.A(n_0_0_235), .B(n_0_0_213), .ZN(n_0_0_212));
   XNOR2_X1 i_0_0_262 (.A(n_0_25), .B(second_operand_number[11]), .ZN(n_0_0_213));
   INV_X1 i_0_0_263 (.A(n_0_0_214), .ZN(n_0_105));
   AOI222_X1 i_0_0_264 (.A1(n_0_0_309), .A2(n_0_0_217), .B1(n_0_0_215), .B2(
      n_0_0_265), .C1(n_0_0_222), .C2(n_0_22), .ZN(n_0_0_214));
   XNOR2_X1 i_0_0_223 (.A(n_0_0_233), .B(n_0_0_216), .ZN(n_0_0_215));
   XOR2_X1 i_0_0_224 (.A(n_0_24), .B(second_operand_number[12]), .Z(n_0_0_216));
   XNOR2_X1 i_0_0_225 (.A(n_0_0_272), .B(n_0_0_218), .ZN(n_0_0_217));
   XOR2_X1 i_0_0_265 (.A(n_0_24), .B(negated_second_operand_number[12]), 
      .Z(n_0_0_218));
   OAI21_X1 i_0_0_266 (.A(n_0_0_219), .B1(n_0_0_220), .B2(n_0_0_264), .ZN(
      n_0_106));
   AOI22_X1 i_0_0_267 (.A1(n_0_0_223), .A2(n_0_0_309), .B1(n_0_21), .B2(
      n_0_0_222), .ZN(n_0_0_219));
   XNOR2_X1 i_0_0_268 (.A(n_0_0_230), .B(n_0_0_221), .ZN(n_0_0_220));
   XOR2_X1 i_0_0_269 (.A(n_0_23), .B(second_operand_number[13]), .Z(n_0_0_221));
   NOR2_X1 i_0_0_270 (.A1(n_0_60), .A2(ready), .ZN(n_0_0_222));
   XNOR2_X1 i_0_0_271 (.A(n_0_0_270), .B(n_0_0_224), .ZN(n_0_0_223));
   XNOR2_X1 i_0_0_272 (.A(n_0_23), .B(negated_second_operand_number[13]), 
      .ZN(n_0_0_224));
   OAI22_X1 i_0_0_276 (.A1(n_0_0_225), .A2(n_0_0_264), .B1(n_0_0_266), .B2(
      n_0_0_308), .ZN(n_0_107));
   XNOR2_X1 i_0_0_273 (.A(n_0_0_227), .B(n_0_0_226), .ZN(n_0_0_225));
   XNOR2_X1 i_0_0_274 (.A(n_0_22), .B(second_operand_number[14]), .ZN(n_0_0_226));
   OAI21_X1 i_0_0_275 (.A(n_0_0_228), .B1(second_operand_number[13]), .B2(n_0_23), 
      .ZN(n_0_0_227));
   INV_X1 i_0_0_277 (.A(n_0_0_229), .ZN(n_0_0_228));
   AOI21_X1 i_0_0_278 (.A(n_0_0_230), .B1(second_operand_number[13]), .B2(n_0_23), 
      .ZN(n_0_0_229));
   OAI21_X1 i_0_0_279 (.A(n_0_0_232), .B1(n_0_0_233), .B2(n_0_0_231), .ZN(
      n_0_0_230));
   NOR2_X1 i_0_0_280 (.A1(n_0_24), .A2(second_operand_number[12]), .ZN(n_0_0_231));
   NAND2_X1 i_0_0_281 (.A1(n_0_24), .A2(second_operand_number[12]), .ZN(
      n_0_0_232));
   OAI21_X1 i_0_0_282 (.A(n_0_0_234), .B1(second_operand_number[11]), .B2(n_0_25), 
      .ZN(n_0_0_233));
   NAND2_X1 i_0_0_283 (.A1(n_0_0_235), .A2(n_0_0_263), .ZN(n_0_0_234));
   OAI21_X1 i_0_0_284 (.A(n_0_0_236), .B1(n_0_0_238), .B2(n_0_26), .ZN(n_0_0_235));
   INV_X1 i_0_0_285 (.A(n_0_0_237), .ZN(n_0_0_236));
   AOI21_X1 i_0_0_286 (.A(second_operand_number[10]), .B1(n_0_0_238), .B2(n_0_26), 
      .ZN(n_0_0_237));
   AOI21_X1 i_0_0_287 (.A(n_0_0_239), .B1(n_0_0_240), .B2(n_0_0_241), .ZN(
      n_0_0_238));
   NOR2_X1 i_0_0_288 (.A1(n_0_27), .A2(second_operand_number[9]), .ZN(n_0_0_239));
   NAND2_X1 i_0_0_289 (.A1(n_0_27), .A2(second_operand_number[9]), .ZN(n_0_0_240));
   OAI21_X1 i_0_0_290 (.A(n_0_0_242), .B1(second_operand_number[8]), .B2(n_0_28), 
      .ZN(n_0_0_241));
   INV_X1 i_0_0_291 (.A(n_0_0_243), .ZN(n_0_0_242));
   AOI21_X1 i_0_0_292 (.A(n_0_0_244), .B1(second_operand_number[8]), .B2(n_0_28), 
      .ZN(n_0_0_243));
   OAI21_X1 i_0_0_293 (.A(n_0_0_246), .B1(n_0_0_247), .B2(n_0_0_245), .ZN(
      n_0_0_244));
   NOR2_X1 i_0_0_294 (.A1(n_0_29), .A2(second_operand_number[7]), .ZN(n_0_0_245));
   NAND2_X1 i_0_0_295 (.A1(n_0_29), .A2(second_operand_number[7]), .ZN(n_0_0_246));
   OAI21_X1 i_0_0_296 (.A(n_0_0_248), .B1(second_operand_number[6]), .B2(n_0_30), 
      .ZN(n_0_0_247));
   INV_X1 i_0_0_297 (.A(n_0_0_249), .ZN(n_0_0_248));
   AOI21_X1 i_0_0_298 (.A(n_0_0_250), .B1(second_operand_number[6]), .B2(n_0_30), 
      .ZN(n_0_0_249));
   NAND2_X1 i_0_0_302 (.A1(n_0_0_255), .A2(n_0_0_251), .ZN(n_0_0_250));
   OAI21_X1 i_0_0_303 (.A(n_0_0_252), .B1(second_operand_number[5]), .B2(n_0_31), 
      .ZN(n_0_0_251));
   OAI21_X1 i_0_0_299 (.A(n_0_0_254), .B1(n_0_0_256), .B2(n_0_0_253), .ZN(
      n_0_0_252));
   NOR2_X1 i_0_0_300 (.A1(n_0_32), .A2(second_operand_number[4]), .ZN(n_0_0_253));
   NAND2_X1 i_0_0_301 (.A1(n_0_32), .A2(second_operand_number[4]), .ZN(n_0_0_254));
   NAND2_X1 i_0_0_307 (.A1(n_0_31), .A2(second_operand_number[5]), .ZN(n_0_0_255));
   OAI21_X1 i_0_0_304 (.A(n_0_0_257), .B1(second_operand_number[3]), .B2(n_0_33), 
      .ZN(n_0_0_256));
   INV_X1 i_0_0_305 (.A(n_0_0_258), .ZN(n_0_0_257));
   AOI21_X1 i_0_0_306 (.A(n_0_0_259), .B1(second_operand_number[3]), .B2(n_0_33), 
      .ZN(n_0_0_258));
   NAND2_X1 i_0_0_308 (.A1(n_0_0_262), .A2(n_0_0_260), .ZN(n_0_0_259));
   OAI21_X1 i_0_0_309 (.A(n_0_0_261), .B1(second_operand_number[2]), .B2(n_0_34), 
      .ZN(n_0_0_260));
   AOI21_X1 i_0_0_310 (.A(n_0_0_304), .B1(n_0_0_303), .B2(n_0_0_429), .ZN(
      n_0_0_261));
   NAND2_X1 i_0_0_311 (.A1(n_0_34), .A2(second_operand_number[2]), .ZN(n_0_0_262));
   NAND2_X1 i_0_0_312 (.A1(n_0_25), .A2(second_operand_number[11]), .ZN(
      n_0_0_263));
   NAND2_X1 i_0_0_313 (.A1(n_0_21), .A2(n_0_0_311), .ZN(n_0_0_264));
   NOR2_X1 i_0_0_314 (.A1(n_0_0_433), .A2(n_0_0_310), .ZN(n_0_0_265));
   XNOR2_X1 i_0_0_318 (.A(n_0_0_307), .B(n_0_0_267), .ZN(n_0_0_266));
   OAI21_X1 i_0_0_315 (.A(n_0_0_268), .B1(n_0_0_270), .B2(
      negated_second_operand_number[13]), .ZN(n_0_0_267));
   INV_X1 i_0_0_316 (.A(n_0_0_269), .ZN(n_0_0_268));
   AOI21_X1 i_0_0_317 (.A(n_0_23), .B1(n_0_0_270), .B2(
      negated_second_operand_number[13]), .ZN(n_0_0_269));
   AOI21_X1 i_0_0_319 (.A(n_0_0_271), .B1(n_0_0_272), .B2(n_0_0_275), .ZN(
      n_0_0_270));
   NOR2_X1 i_0_0_320 (.A1(n_0_24), .A2(negated_second_operand_number[12]), 
      .ZN(n_0_0_271));
   OAI21_X1 i_0_0_321 (.A(n_0_0_273), .B1(n_0_0_276), .B2(
      negated_second_operand_number[11]), .ZN(n_0_0_272));
   INV_X1 i_0_0_322 (.A(n_0_0_274), .ZN(n_0_0_273));
   AOI21_X1 i_0_0_323 (.A(n_0_25), .B1(n_0_0_276), .B2(
      negated_second_operand_number[11]), .ZN(n_0_0_274));
   NAND2_X1 i_0_0_324 (.A1(n_0_24), .A2(negated_second_operand_number[12]), 
      .ZN(n_0_0_275));
   NAND2_X1 i_0_0_325 (.A1(n_0_0_281), .A2(n_0_0_277), .ZN(n_0_0_276));
   OAI21_X1 i_0_0_326 (.A(n_0_0_278), .B1(negated_second_operand_number[10]), 
      .B2(n_0_26), .ZN(n_0_0_277));
   AOI21_X1 i_0_0_327 (.A(n_0_0_279), .B1(n_0_0_280), .B2(n_0_0_282), .ZN(
      n_0_0_278));
   NOR2_X1 i_0_0_328 (.A1(n_0_27), .A2(negated_second_operand_number[9]), 
      .ZN(n_0_0_279));
   NAND2_X1 i_0_0_329 (.A1(n_0_27), .A2(negated_second_operand_number[9]), 
      .ZN(n_0_0_280));
   NAND2_X1 i_0_0_330 (.A1(n_0_26), .A2(negated_second_operand_number[10]), 
      .ZN(n_0_0_281));
   OAI21_X1 i_0_0_331 (.A(n_0_0_283), .B1(negated_second_operand_number[8]), 
      .B2(n_0_28), .ZN(n_0_0_282));
   INV_X1 i_0_0_332 (.A(n_0_0_284), .ZN(n_0_0_283));
   AOI21_X1 i_0_0_333 (.A(n_0_0_285), .B1(negated_second_operand_number[8]), 
      .B2(n_0_28), .ZN(n_0_0_284));
   AOI21_X1 i_0_0_334 (.A(n_0_0_287), .B1(n_0_0_286), .B2(n_0_0_288), .ZN(
      n_0_0_285));
   NAND2_X1 i_0_0_338 (.A1(n_0_29), .A2(negated_second_operand_number[7]), 
      .ZN(n_0_0_286));
   NOR2_X1 i_0_0_339 (.A1(n_0_29), .A2(negated_second_operand_number[7]), 
      .ZN(n_0_0_287));
   OAI21_X1 i_0_0_340 (.A(n_0_0_289), .B1(negated_second_operand_number[6]), 
      .B2(n_0_30), .ZN(n_0_0_288));
   INV_X1 i_0_0_341 (.A(n_0_0_290), .ZN(n_0_0_289));
   AOI21_X1 i_0_0_342 (.A(n_0_0_291), .B1(negated_second_operand_number[6]), 
      .B2(n_0_30), .ZN(n_0_0_290));
   AOI21_X1 i_0_0_343 (.A(n_0_0_292), .B1(n_0_0_293), .B2(n_0_0_296), .ZN(
      n_0_0_291));
   NOR2_X1 i_0_0_344 (.A1(n_0_31), .A2(negated_second_operand_number[5]), 
      .ZN(n_0_0_292));
   OAI21_X1 i_0_0_335 (.A(n_0_0_294), .B1(negated_second_operand_number[4]), 
      .B2(n_0_32), .ZN(n_0_0_293));
   NAND2_X1 i_0_0_336 (.A1(n_0_0_297), .A2(n_0_0_295), .ZN(n_0_0_294));
   NAND2_X1 i_0_0_337 (.A1(n_0_32), .A2(negated_second_operand_number[4]), 
      .ZN(n_0_0_295));
   NAND2_X1 i_0_0_348 (.A1(n_0_31), .A2(negated_second_operand_number[5]), 
      .ZN(n_0_0_296));
   AOI21_X1 i_0_0_345 (.A(n_0_0_298), .B1(negated_second_operand_number[3]), 
      .B2(n_0_33), .ZN(n_0_0_297));
   INV_X1 i_0_0_346 (.A(n_0_0_299), .ZN(n_0_0_298));
   OAI21_X1 i_0_0_347 (.A(n_0_0_300), .B1(negated_second_operand_number[3]), 
      .B2(n_0_33), .ZN(n_0_0_299));
   NAND2_X1 i_0_0_349 (.A1(n_0_0_306), .A2(n_0_0_301), .ZN(n_0_0_300));
   OAI21_X1 i_0_0_350 (.A(n_0_0_302), .B1(negated_second_operand_number[2]), 
      .B2(n_0_34), .ZN(n_0_0_301));
   AOI21_X1 i_0_0_351 (.A(n_0_0_304), .B1(n_0_0_303), .B2(n_0_0_428), .ZN(
      n_0_0_302));
   NAND3_X1 i_0_0_352 (.A1(n_0_35), .A2(n_0_36), .A3(
      negated_second_operand_number[0]), .ZN(n_0_0_303));
   AOI21_X1 i_0_0_353 (.A(n_0_35), .B1(n_0_36), .B2(
      negated_second_operand_number[0]), .ZN(n_0_0_304));
   NAND2_X1 i_0_0_357 (.A1(n_0_36), .A2(negated_second_operand_number[0]), 
      .ZN(n_0_0_305));
   NAND2_X1 i_0_0_354 (.A1(n_0_34), .A2(negated_second_operand_number[2]), 
      .ZN(n_0_0_306));
   XNOR2_X1 i_0_0_359 (.A(n_0_22), .B(negated_second_operand_number[14]), 
      .ZN(n_0_0_307));
   NAND2_X1 i_0_0_355 (.A1(n_0_0_311), .A2(n_0_0_433), .ZN(n_0_0_308));
   NOR2_X1 i_0_0_356 (.A1(n_0_0_310), .A2(n_0_21), .ZN(n_0_0_309));
   INV_X1 i_0_0_358 (.A(n_0_0_311), .ZN(n_0_0_310));
   AND2_X1 i_0_0_360 (.A1(n_0_20), .A2(n_0_0_315), .ZN(n_0_0_311));
   OAI21_X1 i_0_0_364 (.A(n_0_0_312), .B1(n_0_0_442), .B2(ready), .ZN(n_0_108));
   NAND2_X1 i_0_0_365 (.A1(ready), .A2(n_0_0_312), .ZN(n_0_109));
   INV_X1 i_0_0_361 (.A(n_0_0_312), .ZN(n_0_60));
   NOR2_X1 i_0_0_362 (.A1(n_0_0_315), .A2(reset), .ZN(n_0_0_312));
   OAI21_X1 i_0_0_368 (.A(n_0_20), .B1(n_0_0_314), .B2(n_0_0_442), .ZN(n_0_110));
   NOR2_X1 i_0_0_369 (.A1(reset), .A2(n_0_0_313), .ZN(n_0_74));
   OAI21_X1 i_0_0_370 (.A(n_0_20), .B1(n_0_0_314), .B2(n_0_0_313), .ZN(n_0_75));
   NOR4_X1 i_0_0_363 (.A1(n_0_37), .A2(n_0_38), .A3(n_0_39), .A4(n_0_40), 
      .ZN(n_0_0_313));
   OR2_X1 i_0_0_366 (.A1(n_0_0_315), .A2(ready), .ZN(n_0_0_314));
   NAND3_X1 i_0_0_367 (.A1(number_of_bits_in_dividend[1]), .A2(
      number_of_bits_in_dividend[0]), .A3(n_0_0_316), .ZN(n_0_0_315));
   AND3_X1 i_0_0_371 (.A1(number_of_bits_in_dividend[4]), .A2(
      number_of_bits_in_dividend[3]), .A3(number_of_bits_in_dividend[2]), 
      .ZN(n_0_0_316));
   AOI21_X1 i_0_0_372 (.A(n_0_0_441), .B1(n_0_0_337), .B2(divisor[0]), .ZN(n_0_4));
   XNOR2_X1 i_0_0_373 (.A(n_0_116), .B(n_0_0_441), .ZN(n_0_5));
   AND2_X1 i_0_0_374 (.A1(n_0_0_335), .A2(n_0_0_318), .ZN(n_0_7));
   OAI21_X1 i_0_0_375 (.A(n_0_117), .B1(n_0_116), .B2(n_0_0_336), .ZN(n_0_0_318));
   XOR2_X1 i_0_0_381 (.A(n_0_118), .B(n_0_0_335), .Z(n_0_8));
   XNOR2_X1 i_0_0_382 (.A(n_0_119), .B(n_0_0_334), .ZN(n_0_9));
   XNOR2_X1 i_0_0_383 (.A(n_0_120), .B(n_0_0_333), .ZN(n_0_10));
   XOR2_X1 i_0_0_384 (.A(n_0_121), .B(n_0_0_332), .Z(n_0_11));
   XOR2_X1 i_0_0_385 (.A(n_0_122), .B(n_0_0_331), .Z(n_0_12));
   XOR2_X1 i_0_0_386 (.A(n_0_123), .B(n_0_0_330), .Z(n_0_13));
   XOR2_X1 i_0_0_387 (.A(n_0_124), .B(n_0_0_329), .Z(n_0_14));
   XOR2_X1 i_0_0_388 (.A(n_0_125), .B(n_0_0_328), .Z(n_0_15));
   NAND2_X1 i_0_0_377 (.A1(n_0_0_384), .A2(n_0_0_408), .ZN(n_0_0_321));
   NAND2_X1 i_0_0_378 (.A1(n_0_0_389), .A2(n_0_0_388), .ZN(n_0_0_322));
   MUX2_X1 i_0_0_379 (.A(n_0_0_399), .B(n_0_0_402), .S(n_0_0_439), .Z(n_0_0_323));
   NOR2_X1 i_0_0_409 (.A1(n_0_118), .A2(n_0_0_335), .ZN(n_0_0_334));
   NOR2_X1 i_0_0_380 (.A1(n_0_0_388), .A2(n_0_0_357), .ZN(n_0_0_337));
   NAND2_X1 i_0_0_391 (.A1(n_0_0_384), .A2(n_0_0_347), .ZN(n_0_0_342));
   NAND2_X1 i_0_0_395 (.A1(n_0_0_388), .A2(n_0_0_344), .ZN(n_0_0_343));
   NAND2_X1 i_0_0_396 (.A1(n_0_0_384), .A2(n_0_0_350), .ZN(n_0_0_345));
   NAND2_X1 i_0_0_397 (.A1(n_0_0_388), .A2(n_0_0_347), .ZN(n_0_0_346));
   OAI22_X1 i_0_0_398 (.A1(n_0_0_418), .A2(n_0_0_353), .B1(n_0_0_351), .B2(
      n_0_0_361), .ZN(n_0_0_347));
   OAI221_X1 i_0_0_399 (.A(n_0_0_349), .B1(n_0_0_372), .B2(n_0_0_381), .C1(
      n_0_0_352), .C2(n_0_0_385), .ZN(n_0_120));
   NAND2_X1 i_0_0_400 (.A1(n_0_0_388), .A2(n_0_0_350), .ZN(n_0_0_349));
   OAI22_X1 i_0_0_401 (.A1(n_0_0_418), .A2(n_0_0_356), .B1(n_0_0_351), .B2(
      n_0_0_365), .ZN(n_0_0_350));
   MUX2_X1 i_0_0_402 (.A(n_0_0_353), .B(n_0_0_360), .S(n_0_0_439), .Z(n_0_0_352));
   OAI21_X1 i_0_0_403 (.A(n_0_0_354), .B1(n_0_0_407), .B2(divisor[0]), .ZN(
      n_0_0_353));
   NAND2_X1 i_0_0_404 (.A1(n_0_0_407), .A2(n_0_0_369), .ZN(n_0_0_354));
   MUX2_X1 i_0_0_405 (.A(n_0_0_356), .B(n_0_0_364), .S(n_0_0_439), .Z(n_0_0_355));
   MUX2_X1 i_0_0_406 (.A(n_0_0_357), .B(n_0_0_375), .S(n_0_0_407), .Z(n_0_0_356));
   NAND2_X1 i_0_0_407 (.A1(divisor[12]), .A2(divisor[0]), .ZN(n_0_0_358));
   NAND2_X1 i_0_0_408 (.A1(n_0_0_417), .A2(divisor[12]), .ZN(n_0_0_362));
   MUX2_X1 i_0_0_410 (.A(n_0_0_364), .B(n_0_0_374), .S(n_0_0_439), .Z(n_0_0_363));
   MUX2_X1 i_0_0_411 (.A(n_0_0_365), .B(n_0_0_412), .S(n_0_0_407), .Z(n_0_0_364));
   NAND2_X1 i_0_0_412 (.A1(n_0_0_416), .A2(divisor[12]), .ZN(n_0_0_366));
   MUX2_X1 i_0_0_413 (.A(n_0_0_368), .B(n_0_0_380), .S(n_0_0_439), .Z(n_0_0_367));
   OAI21_X1 i_0_0_414 (.A(divisor[12]), .B1(n_0_0_416), .B2(divisor[3]), 
      .ZN(n_0_0_370));
   MUX2_X1 i_0_0_415 (.A(n_0_0_374), .B(n_0_0_401), .S(n_0_0_439), .Z(n_0_0_373));
   MUX2_X1 i_0_0_416 (.A(n_0_0_375), .B(n_0_0_399), .S(n_0_0_407), .Z(n_0_0_374));
   XOR2_X1 i_0_0_417 (.A(divisor[5]), .B(n_0_0_376), .Z(n_0_0_375));
   NAND2_X1 i_0_0_418 (.A1(n_0_0_415), .A2(divisor[12]), .ZN(n_0_0_376));
   INV_X1 i_0_0_419 (.A(n_0_0_379), .ZN(n_0_0_378));
   MUX2_X1 i_0_0_420 (.A(n_0_0_392), .B(n_0_0_380), .S(n_0_0_418), .Z(n_0_0_379));
   MUX2_X1 i_0_0_421 (.A(n_0_0_381), .B(n_0_0_390), .S(n_0_0_407), .Z(n_0_0_380));
   XOR2_X1 i_0_0_422 (.A(divisor[6]), .B(n_0_0_382), .Z(n_0_0_381));
   NAND2_X1 i_0_0_423 (.A1(n_0_0_414), .A2(divisor[12]), .ZN(n_0_0_382));
   INV_X1 i_0_0_424 (.A(n_0_0_383), .ZN(n_0_128));
   INV_X1 i_0_0_425 (.A(n_0_0_385), .ZN(n_0_0_384));
   OAI22_X1 i_0_0_426 (.A1(n_0_0_439), .A2(n_0_0_392), .B1(n_0_0_390), .B2(
      n_0_0_398), .ZN(n_0_0_389));
   XOR2_X1 i_0_0_427 (.A(divisor[10]), .B(n_0_0_391), .Z(n_0_0_390));
   OAI21_X1 i_0_0_428 (.A(divisor[12]), .B1(n_0_0_405), .B2(divisor[9]), 
      .ZN(n_0_0_391));
   MUX2_X1 i_0_0_429 (.A(n_0_0_393), .B(n_0_0_394), .S(n_0_0_408), .Z(n_0_0_392));
   NAND3_X1 i_0_0_430 (.A1(divisor[12]), .A2(n_0_0_404), .A3(n_0_0_436), 
      .ZN(n_0_0_393));
   OAI22_X1 i_0_0_431 (.A1(n_0_0_439), .A2(n_0_0_401), .B1(n_0_0_399), .B2(
      n_0_0_398), .ZN(n_0_0_397));
   NAND2_X1 i_0_0_432 (.A1(n_0_0_439), .A2(n_0_0_408), .ZN(n_0_0_398));
   XOR2_X1 i_0_0_433 (.A(divisor[9]), .B(n_0_0_400), .Z(n_0_0_399));
   NAND2_X1 i_0_0_434 (.A1(n_0_0_405), .A2(divisor[12]), .ZN(n_0_0_400));
   MUX2_X1 i_0_0_435 (.A(n_0_0_412), .B(n_0_0_402), .S(n_0_0_407), .Z(n_0_0_401));
   XNOR2_X1 i_0_0_436 (.A(divisor[11]), .B(n_0_0_403), .ZN(n_0_0_402));
   NOR2_X1 i_0_0_437 (.A1(n_0_0_404), .A2(n_0_0_437), .ZN(n_0_0_403));
   NOR3_X1 i_0_0_438 (.A1(n_0_0_405), .A2(divisor[9]), .A3(divisor[10]), 
      .ZN(n_0_0_404));
   NAND2_X1 i_0_0_439 (.A1(n_0_0_406), .A2(n_0_0_435), .ZN(n_0_0_405));
   XOR2_X1 i_0_0_440 (.A(divisor[7]), .B(n_0_0_413), .Z(n_0_0_412));
   OAI21_X1 i_0_0_441 (.A(divisor[12]), .B1(n_0_0_414), .B2(divisor[6]), 
      .ZN(n_0_0_413));
   NOR2_X1 i_0_0_442 (.A1(n_0_0_432), .A2(divisor[14]), .ZN(n_0_0_426));
   INV_X1 i_0_0_443 (.A(negated_second_operand_number[1]), .ZN(n_0_0_428));
   INV_X1 i_0_0_444 (.A(second_operand_number[1]), .ZN(n_0_0_429));
   INV_X1 i_0_0_445 (.A(dividend[11]), .ZN(n_0_0_430));
   INV_X1 i_0_0_522 (.A(dividend[12]), .ZN(n_0_0_431));
   INV_X1 i_0_0_447 (.A(n_0_21), .ZN(n_0_0_433));
   INV_X1 i_0_0_449 (.A(divisor[8]), .ZN(n_0_0_435));
   INV_X1 i_0_0_450 (.A(divisor[11]), .ZN(n_0_0_436));
   INV_X1 i_0_0_451 (.A(n_0_0_388), .ZN(n_0_0_438));
   INV_X1 i_0_0_452 (.A(n_0_0_411), .ZN(n_0_0_440));
   INV_X1 i_0_0_453 (.A(n_0_0_336), .ZN(n_0_0_441));
   INV_X1 i_0_0_454 (.A(n_0_0_313), .ZN(n_0_0_442));
   INV_X1 i_0_0_455 (.A(n_0_0_396), .ZN(n_0_0_411));
   INV_X1 i_0_0_456 (.A(n_0_0_534), .ZN(n_0_0_351));
   OAI21_X1 i_0_0_457 (.A(n_0_0_519), .B1(n_0_0_365), .B2(n_0_0_535), .ZN(
      n_0_0_344));
   INV_X1 i_0_0_458 (.A(n_0_0_424), .ZN(n_0_0_365));
   INV_X1 i_0_0_376 (.A(n_0_0_460), .ZN(n_0_0_329));
   NAND3_X1 i_0_0_389 (.A1(n_0_0_333), .A2(n_0_0_503), .A3(n_0_0_502), .ZN(
      n_0_0_331));
   NAND2_X1 i_0_0_390 (.A1(n_0_0_333), .A2(n_0_0_503), .ZN(n_0_0_332));
   INV_X1 i_0_0_459 (.A(n_0_0_517), .ZN(n_0_117));
   INV_X1 i_0_0_392 (.A(n_0_0_502), .ZN(n_0_121));
   INV_X1 i_0_0_393 (.A(n_0_0_500), .ZN(n_0_122));
   NAND2_X1 i_0_0_394 (.A1(n_0_0_489), .A2(n_0_0_493), .ZN(n_0_124));
   INV_X1 i_0_0_460 (.A(n_0_0_377), .ZN(n_0_127));
   NOR2_X1 i_0_0_461 (.A1(n_0_0_317), .A2(n_0_0_4), .ZN(n_0_0_3));
   OAI22_X1 i_0_0_462 (.A1(n_0_0_379), .A2(n_0_0_385), .B1(n_0_0_393), .B2(
      n_0_0_372), .ZN(n_0_0_4));
   NOR2_X1 i_0_0_463 (.A1(n_0_0_373), .A2(n_0_0_438), .ZN(n_0_0_317));
   AOI21_X1 i_0_0_464 (.A(n_0_0_320), .B1(n_0_0_325), .B2(n_0_0_339), .ZN(
      n_0_0_319));
   NOR2_X1 i_0_0_465 (.A1(n_0_0_402), .A2(n_0_0_372), .ZN(n_0_0_320));
   NOR2_X1 i_0_0_466 (.A1(n_0_0_390), .A2(n_0_0_372), .ZN(n_0_0_324));
   INV_X1 i_0_0_467 (.A(n_0_0_367), .ZN(n_0_0_325));
   AOI21_X1 i_0_0_468 (.A(n_0_0_327), .B1(n_0_0_338), .B2(n_0_0_339), .ZN(
      n_0_0_326));
   NOR2_X1 i_0_0_469 (.A1(n_0_0_399), .A2(n_0_0_372), .ZN(n_0_0_327));
   INV_X1 i_0_0_470 (.A(n_0_0_359), .ZN(n_0_0_338));
   INV_X1 i_0_0_471 (.A(n_0_0_438), .ZN(n_0_0_339));
   OAI22_X1 i_0_0_472 (.A1(n_0_0_352), .A2(n_0_0_438), .B1(n_0_0_412), .B2(
      n_0_0_372), .ZN(n_0_0_340));
   NOR2_X1 i_0_0_473 (.A1(n_0_0_355), .A2(n_0_0_385), .ZN(n_0_0_341));
   INV_X1 i_0_0_474 (.A(n_0_0_371), .ZN(n_0_0_348));
   OAI21_X1 i_0_0_475 (.A(n_0_0_346), .B1(n_0_0_375), .B2(n_0_0_372), .ZN(
      n_0_0_371));
   INV_X1 i_0_0_476 (.A(n_0_0_397), .ZN(n_0_0_386));
   INV_X1 i_0_0_477 (.A(n_0_0_389), .ZN(n_0_0_387));
   INV_X1 i_0_0_478 (.A(n_0_0_384), .ZN(n_0_0_395));
   INV_X1 i_0_0_479 (.A(n_0_0_542), .ZN(n_0_0_396));
   INV_X1 i_0_0_480 (.A(n_0_0_445), .ZN(n_0_0_406));
   NAND2_X1 i_0_0_481 (.A1(n_0_0_451), .A2(n_0_0_459), .ZN(n_0_0_417));
   INV_X1 i_0_0_482 (.A(n_0_0_407), .ZN(n_0_0_408));
   INV_X1 i_0_0_483 (.A(divisor[12]), .ZN(n_0_0_437));
   AOI21_X1 i_0_0_484 (.A(reset), .B1(n_0_0_5), .B2(n_0_0_410), .ZN(n_0_0_409));
   INV_X1 i_0_0_485 (.A(number_of_bits_in_dividend[4]), .ZN(n_0_0_410));
   INV_X1 i_0_0_486 (.A(n_0_0_357), .ZN(n_0_0_419));
   AOI21_X1 i_0_0_487 (.A(n_0_0_421), .B1(n_0_0_381), .B2(n_0_0_407), .ZN(
      n_0_0_420));
   NOR2_X1 i_0_0_488 (.A1(n_0_0_407), .A2(n_0_0_527), .ZN(n_0_0_421));
   XNOR2_X1 i_0_0_489 (.A(n_0_0_370), .B(divisor[4]), .ZN(n_0_0_423));
   INV_X1 i_0_0_490 (.A(n_0_0_524), .ZN(n_0_0_424));
   INV_X1 i_0_0_491 (.A(n_0_0_420), .ZN(n_0_0_360));
   XNOR2_X1 i_0_0_446 (.A(n_0_0_457), .B(n_0_126), .ZN(n_0_16));
   INV_X1 i_0_0_448 (.A(n_0_0_3), .ZN(n_0_126));
   AOI22_X1 i_0_0_492 (.A1(n_0_0_378), .A2(n_0_0_388), .B1(n_0_0_384), .B2(
      n_0_0_397), .ZN(n_0_0_377));
   OR2_X1 i_0_0_493 (.A1(n_0_0_341), .A2(n_0_0_340), .ZN(n_0_0_425));
   OAI22_X1 i_0_0_494 (.A1(n_0_0_359), .A2(n_0_0_385), .B1(n_0_0_372), .B2(
      n_0_0_394), .ZN(n_0_0_427));
   OAI21_X1 i_0_0_495 (.A(n_0_0_434), .B1(n_0_0_420), .B2(n_0_0_439), .ZN(
      n_0_0_359));
   NAND2_X1 i_0_0_496 (.A1(n_0_0_368), .A2(n_0_0_439), .ZN(n_0_0_434));
   OAI21_X1 i_0_0_497 (.A(n_0_0_443), .B1(n_0_0_423), .B2(n_0_0_407), .ZN(
      n_0_0_368));
   NAND2_X1 i_0_0_498 (.A1(n_0_0_394), .A2(n_0_0_407), .ZN(n_0_0_443));
   XOR2_X1 i_0_0_499 (.A(divisor[8]), .B(n_0_0_444), .Z(n_0_0_394));
   NAND2_X1 i_0_0_500 (.A1(n_0_0_445), .A2(divisor[12]), .ZN(n_0_0_444));
   OR3_X1 i_0_0_501 (.A1(n_0_0_414), .A2(divisor[7]), .A3(divisor[6]), .ZN(
      n_0_0_445));
   OR2_X1 i_0_0_502 (.A1(n_0_0_415), .A2(divisor[5]), .ZN(n_0_0_414));
   NAND3_X1 i_0_0_503 (.A1(n_0_0_446), .A2(n_0_0_449), .A3(n_0_0_448), .ZN(
      n_0_0_415));
   INV_X1 i_0_0_504 (.A(n_0_0_416), .ZN(n_0_0_446));
   NAND3_X1 i_0_0_505 (.A1(n_0_0_447), .A2(n_0_0_451), .A3(n_0_0_459), .ZN(
      n_0_0_416));
   INV_X1 i_0_0_506 (.A(divisor[2]), .ZN(n_0_0_447));
   INV_X1 i_0_0_507 (.A(divisor[3]), .ZN(n_0_0_448));
   INV_X1 i_0_0_510 (.A(divisor[4]), .ZN(n_0_0_449));
   NOR2_X1 i_0_0_513 (.A1(n_0_0_355), .A2(n_0_0_438), .ZN(n_0_0_450));
   INV_X1 i_0_0_514 (.A(n_0_0_423), .ZN(n_0_0_369));
   INV_X1 i_0_0_515 (.A(n_0_0_527), .ZN(n_0_0_361));
   INV_X1 i_0_0_516 (.A(divisor[1]), .ZN(n_0_0_451));
   NAND2_X1 i_0_0_517 (.A1(n_0_0_407), .A2(n_0_0_418), .ZN(n_0_0_452));
   INV_X1 i_0_0_518 (.A(n_0_0_439), .ZN(n_0_0_418));
   INV_X1 i_0_0_519 (.A(n_0_0_535), .ZN(n_0_0_453));
   OAI22_X1 i_0_0_520 (.A1(n_0_0_386), .A2(n_0_0_530), .B1(n_0_0_387), .B2(
      n_0_0_395), .ZN(n_0_0_454));
   NAND2_X1 i_0_0_521 (.A1(n_0_0_456), .A2(n_0_0_558), .ZN(n_0_0_455));
   INV_X1 i_0_0_524 (.A(n_0_0_538), .ZN(n_0_0_456));
   INV_X1 i_0_0_508 (.A(n_0_0_458), .ZN(n_0_0_457));
   NAND2_X1 i_0_0_509 (.A1(n_0_0_469), .A2(n_0_0_476), .ZN(n_0_0_458));
   INV_X1 i_0_0_525 (.A(divisor[0]), .ZN(n_0_0_459));
   INV_X1 i_0_0_511 (.A(n_0_0_461), .ZN(n_0_0_460));
   NAND2_X1 i_0_0_512 (.A1(n_0_0_469), .A2(n_0_0_494), .ZN(n_0_0_461));
   NAND2_X1 i_0_0_526 (.A1(n_0_0_496), .A2(n_0_0_560), .ZN(n_0_0_385));
   OAI21_X1 i_0_0_527 (.A(n_0_0_530), .B1(n_0_0_528), .B2(n_0_0_422), .ZN(
      n_0_0_372));
   NAND2_X1 i_0_0_528 (.A1(n_0_0_463), .A2(n_0_0_462), .ZN(n_0_59));
   OAI21_X1 i_0_0_529 (.A(n_0_0_409), .B1(n_0_0_5), .B2(n_0_0_410), .ZN(
      n_0_0_462));
   INV_X1 i_0_0_530 (.A(reset), .ZN(n_0_20));
   INV_X1 i_0_0_523 (.A(n_0_0_463), .ZN(n_0_113));
   NAND4_X1 i_0_0_531 (.A1(n_0_0_486), .A2(reset), .A3(n_0_0_481), .A4(n_0_0_479), 
      .ZN(n_0_0_463));
   INV_X1 i_0_0_532 (.A(n_0_0_516), .ZN(n_0_114));
   NAND2_X1 i_0_0_533 (.A1(n_0_0_513), .A2(n_0_0_515), .ZN(n_0_115));
   NAND2_X1 i_0_0_534 (.A1(n_0_0_509), .A2(n_0_0_507), .ZN(n_0_118));
   INV_X1 i_0_0_535 (.A(n_0_0_464), .ZN(n_0_17));
   OAI21_X1 i_0_0_536 (.A(n_0_0_468), .B1(n_0_0_465), .B2(n_0_0_377), .ZN(
      n_0_0_464));
   INV_X1 i_0_0_537 (.A(n_0_0_466), .ZN(n_0_0_465));
   NAND3_X1 i_0_0_538 (.A1(n_0_0_469), .A2(n_0_0_3), .A3(n_0_0_476), .ZN(
      n_0_0_466));
   AOI21_X1 i_0_0_539 (.A(n_0_0_467), .B1(n_0_0_468), .B2(n_0_0_454), .ZN(n_0_18));
   INV_X1 i_0_0_540 (.A(n_0_0_473), .ZN(n_0_0_467));
   NAND4_X1 i_0_0_541 (.A1(n_0_0_469), .A2(n_0_0_494), .A3(n_0_0_487), .A4(
      n_0_0_481), .ZN(n_0_0_468));
   INV_X1 i_0_0_542 (.A(n_0_0_330), .ZN(n_0_0_469));
   NAND3_X1 i_0_0_543 (.A1(n_0_0_470), .A2(n_0_0_505), .A3(n_0_0_498), .ZN(
      n_0_0_330));
   INV_X1 i_0_0_544 (.A(n_0_0_335), .ZN(n_0_0_470));
   NAND3_X1 i_0_0_545 (.A1(n_0_0_512), .A2(n_0_0_525), .A3(n_0_0_517), .ZN(
      n_0_0_335));
   INV_X1 i_0_0_546 (.A(n_0_0_471), .ZN(n_0_19));
   NAND2_X1 i_0_0_547 (.A1(n_0_0_478), .A2(n_0_0_472), .ZN(n_0_0_471));
   NAND2_X1 i_0_0_548 (.A1(n_0_0_473), .A2(n_0_129), .ZN(n_0_0_472));
   NAND4_X1 i_0_0_549 (.A1(n_0_0_333), .A2(n_0_0_476), .A3(n_0_0_498), .A4(
      n_0_0_474), .ZN(n_0_0_473));
   INV_X1 i_0_0_550 (.A(n_0_0_475), .ZN(n_0_0_474));
   NAND3_X1 i_0_0_551 (.A1(n_0_0_383), .A2(n_0_0_377), .A3(n_0_0_3), .ZN(
      n_0_0_475));
   INV_X1 i_0_0_552 (.A(n_0_0_454), .ZN(n_0_0_383));
   INV_X1 i_0_0_553 (.A(n_0_0_477), .ZN(n_0_0_476));
   NAND3_X1 i_0_0_554 (.A1(n_0_0_487), .A2(n_0_0_494), .A3(n_0_0_483), .ZN(
      n_0_0_477));
   NAND3_X1 i_0_0_555 (.A1(n_0_0_486), .A2(n_0_0_481), .A3(n_0_0_479), .ZN(
      n_0_0_478));
   INV_X1 i_0_0_556 (.A(n_0_0_480), .ZN(n_0_0_479));
   OR2_X1 i_0_0_557 (.A1(n_0_129), .A2(n_0_0_454), .ZN(n_0_0_480));
   OAI21_X1 i_0_0_558 (.A(n_0_0_322), .B1(n_0_0_321), .B2(n_0_0_323), .ZN(
      n_0_129));
   INV_X1 i_0_0_559 (.A(n_0_0_482), .ZN(n_0_0_481));
   NAND3_X1 i_0_0_560 (.A1(n_0_0_483), .A2(n_0_0_377), .A3(n_0_0_3), .ZN(
      n_0_0_482));
   INV_X1 i_0_0_561 (.A(n_0_125), .ZN(n_0_0_483));
   NAND2_X1 i_0_0_562 (.A1(n_0_0_484), .A2(n_0_0_319), .ZN(n_0_125));
   NAND3_X1 i_0_0_563 (.A1(n_0_0_496), .A2(n_0_0_485), .A3(n_0_0_560), .ZN(
      n_0_0_484));
   INV_X1 i_0_0_564 (.A(n_0_0_373), .ZN(n_0_0_485));
   INV_X1 i_0_0_565 (.A(n_0_0_328), .ZN(n_0_0_486));
   NAND4_X1 i_0_0_566 (.A1(n_0_0_333), .A2(n_0_0_498), .A3(n_0_0_494), .A4(
      n_0_0_487), .ZN(n_0_0_328));
   INV_X1 i_0_0_567 (.A(n_0_0_488), .ZN(n_0_0_487));
   NAND2_X1 i_0_0_568 (.A1(n_0_0_489), .A2(n_0_0_493), .ZN(n_0_0_488));
   INV_X1 i_0_0_569 (.A(n_0_0_490), .ZN(n_0_0_489));
   NAND2_X1 i_0_0_570 (.A1(n_0_0_491), .A2(n_0_0_492), .ZN(n_0_0_490));
   NAND4_X1 i_0_0_571 (.A1(n_0_0_535), .A2(n_0_0_325), .A3(n_0_0_560), .A4(
      n_0_0_550), .ZN(n_0_0_491));
   INV_X1 i_0_0_572 (.A(n_0_0_324), .ZN(n_0_0_492));
   OR2_X1 i_0_0_573 (.A1(n_0_0_363), .A2(n_0_0_438), .ZN(n_0_0_493));
   INV_X1 i_0_0_574 (.A(n_0_123), .ZN(n_0_0_494));
   NAND2_X1 i_0_0_575 (.A1(n_0_0_495), .A2(n_0_0_326), .ZN(n_0_123));
   NAND3_X1 i_0_0_576 (.A1(n_0_0_496), .A2(n_0_0_497), .A3(n_0_0_560), .ZN(
      n_0_0_495));
   NOR2_X1 i_0_0_577 (.A1(n_0_0_528), .A2(n_0_0_422), .ZN(n_0_0_496));
   INV_X1 i_0_0_578 (.A(n_0_0_363), .ZN(n_0_0_497));
   INV_X1 i_0_0_579 (.A(n_0_0_499), .ZN(n_0_0_498));
   NAND3_X1 i_0_0_580 (.A1(n_0_0_500), .A2(n_0_0_503), .A3(n_0_0_502), .ZN(
      n_0_0_499));
   INV_X1 i_0_0_581 (.A(n_0_0_501), .ZN(n_0_0_500));
   OR2_X1 i_0_0_582 (.A1(n_0_0_450), .A2(n_0_0_427), .ZN(n_0_0_501));
   INV_X1 i_0_0_583 (.A(n_0_0_425), .ZN(n_0_0_502));
   INV_X1 i_0_0_584 (.A(n_0_120), .ZN(n_0_0_503));
   INV_X1 i_0_0_585 (.A(n_0_0_504), .ZN(n_0_0_333));
   NAND4_X1 i_0_0_586 (.A1(n_0_0_512), .A2(n_0_0_525), .A3(n_0_0_505), .A4(
      n_0_0_517), .ZN(n_0_0_504));
   INV_X1 i_0_0_587 (.A(n_0_0_506), .ZN(n_0_0_505));
   NAND3_X1 i_0_0_588 (.A1(n_0_0_509), .A2(n_0_0_511), .A3(n_0_0_507), .ZN(
      n_0_0_506));
   INV_X1 i_0_0_589 (.A(n_0_0_508), .ZN(n_0_0_507));
   NAND2_X1 i_0_0_590 (.A1(n_0_0_342), .A2(n_0_0_343), .ZN(n_0_0_508));
   OAI211_X1 i_0_0_591 (.A(n_0_0_510), .B(n_0_0_530), .C1(n_0_0_528), .C2(
      n_0_0_422), .ZN(n_0_0_509));
   INV_X1 i_0_0_592 (.A(n_0_0_369), .ZN(n_0_0_510));
   INV_X1 i_0_0_593 (.A(n_0_119), .ZN(n_0_0_511));
   NAND2_X1 i_0_0_594 (.A1(n_0_0_345), .A2(n_0_0_348), .ZN(n_0_119));
   INV_X1 i_0_0_595 (.A(n_0_0_336), .ZN(n_0_0_512));
   NAND3_X1 i_0_0_596 (.A1(n_0_0_516), .A2(n_0_0_513), .A3(n_0_0_515), .ZN(
      n_0_0_336));
   OAI211_X1 i_0_0_597 (.A(n_0_0_530), .B(n_0_0_514), .C1(n_0_0_528), .C2(
      n_0_0_422), .ZN(n_0_0_513));
   INV_X1 i_0_0_598 (.A(n_0_0_357), .ZN(n_0_0_514));
   XNOR2_X1 i_0_0_599 (.A(n_0_0_358), .B(n_0_0_451), .ZN(n_0_0_357));
   NAND3_X1 i_0_0_600 (.A1(n_0_0_388), .A2(divisor[0]), .A3(n_0_0_453), .ZN(
      n_0_0_515));
   OAI211_X1 i_0_0_601 (.A(divisor[0]), .B(n_0_0_530), .C1(n_0_0_528), .C2(
      n_0_0_422), .ZN(n_0_0_516));
   NAND3_X1 i_0_0_602 (.A1(n_0_0_523), .A2(n_0_0_518), .A3(n_0_0_520), .ZN(
      n_0_0_517));
   NAND4_X1 i_0_0_603 (.A1(n_0_0_535), .A2(n_0_0_560), .A3(n_0_0_550), .A4(
      n_0_0_519), .ZN(n_0_0_518));
   NAND2_X1 i_0_0_604 (.A1(n_0_0_534), .A2(n_0_0_419), .ZN(n_0_0_519));
   NAND3_X1 i_0_0_605 (.A1(n_0_0_521), .A2(n_0_0_388), .A3(n_0_0_533), .ZN(
      n_0_0_520));
   NAND3_X1 i_0_0_606 (.A1(n_0_0_407), .A2(n_0_0_522), .A3(n_0_0_439), .ZN(
      n_0_0_521));
   INV_X1 i_0_0_607 (.A(n_0_0_361), .ZN(n_0_0_522));
   OAI211_X1 i_0_0_608 (.A(n_0_0_530), .B(n_0_0_524), .C1(n_0_0_528), .C2(
      n_0_0_422), .ZN(n_0_0_523));
   XOR2_X1 i_0_0_609 (.A(divisor[3]), .B(n_0_0_366), .Z(n_0_0_524));
   INV_X1 i_0_0_610 (.A(n_0_116), .ZN(n_0_0_525));
   NAND3_X1 i_0_0_611 (.A1(n_0_0_526), .A2(n_0_0_531), .A3(n_0_0_529), .ZN(
      n_0_116));
   OAI211_X1 i_0_0_612 (.A(n_0_0_530), .B(n_0_0_527), .C1(n_0_0_528), .C2(
      n_0_0_422), .ZN(n_0_0_526));
   XNOR2_X1 i_0_0_613 (.A(divisor[2]), .B(n_0_0_362), .ZN(n_0_0_527));
   AOI22_X1 i_0_0_614 (.A1(n_0_0_540), .A2(n_0_0_543), .B1(n_0_0_539), .B2(
      n_0_0_536), .ZN(n_0_0_528));
   INV_X1 i_0_0_615 (.A(n_0_0_550), .ZN(n_0_0_422));
   NAND3_X1 i_0_0_616 (.A1(n_0_0_388), .A2(n_0_0_419), .A3(n_0_0_453), .ZN(
      n_0_0_529));
   INV_X1 i_0_0_617 (.A(n_0_0_530), .ZN(n_0_0_388));
   NAND2_X1 i_0_0_618 (.A1(n_0_0_550), .A2(n_0_0_455), .ZN(n_0_0_530));
   NAND4_X1 i_0_0_619 (.A1(n_0_0_535), .A2(n_0_0_560), .A3(n_0_0_550), .A4(
      n_0_0_532), .ZN(n_0_0_531));
   INV_X1 i_0_0_620 (.A(n_0_0_533), .ZN(n_0_0_532));
   NAND2_X1 i_0_0_621 (.A1(n_0_0_534), .A2(divisor[0]), .ZN(n_0_0_533));
   INV_X1 i_0_0_622 (.A(n_0_0_452), .ZN(n_0_0_534));
   NAND2_X1 i_0_0_623 (.A1(n_0_0_407), .A2(n_0_0_439), .ZN(n_0_0_535));
   NAND2_X1 i_0_0_624 (.A1(n_0_0_536), .A2(n_0_0_539), .ZN(n_0_0_439));
   NAND2_X1 i_0_0_625 (.A1(n_0_0_537), .A2(n_0_0_538), .ZN(n_0_0_536));
   NAND2_X1 i_0_0_626 (.A1(n_0_0_552), .A2(n_0_0_548), .ZN(n_0_0_537));
   INV_X1 i_0_0_627 (.A(n_0_0_545), .ZN(n_0_0_538));
   NAND3_X1 i_0_0_628 (.A1(n_0_0_552), .A2(n_0_0_545), .A3(n_0_0_548), .ZN(
      n_0_0_539));
   NAND2_X1 i_0_0_629 (.A1(n_0_0_540), .A2(n_0_0_543), .ZN(n_0_0_407));
   NAND2_X1 i_0_0_630 (.A1(n_0_0_541), .A2(n_0_0_542), .ZN(n_0_0_540));
   NAND2_X1 i_0_0_631 (.A1(n_0_0_544), .A2(n_0_0_548), .ZN(n_0_0_541));
   INV_X1 i_0_0_632 (.A(n_0_0_549), .ZN(n_0_0_542));
   NAND3_X1 i_0_0_633 (.A1(n_0_0_544), .A2(n_0_0_549), .A3(n_0_0_548), .ZN(
      n_0_0_543));
   NAND2_X1 i_0_0_634 (.A1(n_0_0_552), .A2(n_0_0_545), .ZN(n_0_0_544));
   NAND2_X1 i_0_0_635 (.A1(n_0_0_547), .A2(n_0_0_546), .ZN(n_0_0_545));
   INV_X1 i_0_0_636 (.A(cla0_n_0), .ZN(n_0_0_546));
   INV_X1 i_0_0_637 (.A(dividend[13]), .ZN(n_0_0_547));
   NAND2_X1 i_0_0_638 (.A1(dividend[14]), .A2(cla0_n_1), .ZN(n_0_0_548));
   NAND2_X1 i_0_0_639 (.A1(n_0_0_554), .A2(n_0_0_559), .ZN(n_0_0_549));
   NAND2_X1 i_0_0_640 (.A1(n_0_0_551), .A2(n_0_0_559), .ZN(n_0_0_550));
   NAND3_X1 i_0_0_641 (.A1(n_0_0_557), .A2(n_0_0_554), .A3(n_0_0_552), .ZN(
      n_0_0_551));
   NAND2_X1 i_0_0_642 (.A1(n_0_0_432), .A2(n_0_0_553), .ZN(n_0_0_552));
   INV_X1 i_0_0_643 (.A(cla0_n_1), .ZN(n_0_0_553));
   NAND2_X1 i_0_0_644 (.A1(n_0_0_556), .A2(n_0_0_555), .ZN(n_0_0_554));
   INV_X1 i_0_0_645 (.A(cla0_n_2), .ZN(n_0_0_555));
   INV_X1 i_0_0_646 (.A(dividend[15]), .ZN(n_0_0_556));
   OAI21_X1 i_0_0_647 (.A(n_0_0_558), .B1(n_0_0_432), .B2(divisor[14]), .ZN(
      n_0_0_557));
   NAND2_X1 i_0_0_648 (.A1(dividend[13]), .A2(cla0_n_0), .ZN(n_0_0_558));
   INV_X1 i_0_0_649 (.A(dividend[14]), .ZN(n_0_0_432));
   NAND2_X1 i_0_0_650 (.A1(dividend[15]), .A2(cla0_n_2), .ZN(n_0_0_559));
   INV_X1 i_0_0_651 (.A(n_0_0_455), .ZN(n_0_0_560));
   MUX2_X1 overFlow_reg_enable_mux_0 (.A(overFlow), .B(n_0_74), .S(n_0_75), 
      .Z(n_0_111));
   MUX2_X1 ready_reg_enable_mux_0 (.A(ready), .B(n_0_20), .S(n_0_53), .Z(n_0_112));
endmodule
