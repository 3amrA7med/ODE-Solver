/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 16:04:01 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3831160354 */

module datapath__0_35(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   XNOR2_X1 i_0 (.A(p_0[2]), .B(p_0[1]), .ZN(p_1[2]));
   NAND2_X1 i_1 (.A1(n_3), .A2(n_0), .ZN(p_1[3]));
   OAI21_X1 i_2 (.A(p_0[3]), .B1(p_0[2]), .B2(p_0[1]), .ZN(n_0));
   XNOR2_X1 i_3 (.A(p_0[4]), .B(n_3), .ZN(p_1[4]));
   XOR2_X1 i_4 (.A(p_0[5]), .B(n_2), .Z(p_1[5]));
   XOR2_X1 i_5 (.A(p_0[31]), .B(n_1), .Z(p_1[6]));
   OR2_X1 i_6 (.A1(p_0[31]), .A2(n_1), .ZN(p_1[11]));
   NOR3_X1 i_7 (.A1(n_3), .A2(p_0[4]), .A3(p_0[5]), .ZN(n_1));
   NOR2_X1 i_8 (.A1(n_3), .A2(p_0[4]), .ZN(n_2));
   OR3_X1 i_9 (.A1(p_0[3]), .A2(p_0[2]), .A3(p_0[1]), .ZN(n_3));
endmodule

module datapath__0_39(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   XNOR2_X1 i_0 (.A(p_0[2]), .B(p_0[1]), .ZN(p_1[2]));
   NAND2_X1 i_1 (.A1(n_3), .A2(n_0), .ZN(p_1[3]));
   OAI21_X1 i_2 (.A(p_0[3]), .B1(p_0[2]), .B2(p_0[1]), .ZN(n_0));
   XNOR2_X1 i_3 (.A(p_0[4]), .B(n_3), .ZN(p_1[4]));
   XOR2_X1 i_4 (.A(p_0[5]), .B(n_2), .Z(p_1[5]));
   XOR2_X1 i_5 (.A(p_0[31]), .B(n_1), .Z(p_1[6]));
   OR2_X1 i_6 (.A1(p_0[31]), .A2(n_1), .ZN(p_1[11]));
   NOR3_X1 i_7 (.A1(n_3), .A2(p_0[4]), .A3(p_0[5]), .ZN(n_1));
   NOR2_X1 i_8 (.A1(n_3), .A2(p_0[4]), .ZN(n_2));
   OR3_X1 i_9 (.A1(p_0[3]), .A2(p_0[2]), .A3(p_0[1]), .ZN(n_3));
endmodule

module datapath__1_338(PacketSize, p_0);
   input [5:0]PacketSize;
   output [31:0]p_0;

   HA_X1 i_0 (.A(PacketSize[1]), .B(PacketSize[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_1 (.A(PacketSize[4]), .B(n_3), .CO(n_1), .S(p_0[4]));
   INV_X1 i_2 (.A(n_2), .ZN(p_0[2]));
   AOI21_X1 i_3 (.A(n_4), .B1(PacketSize[2]), .B2(n_0), .ZN(n_2));
   OAI21_X1 i_4 (.A(n_3), .B1(n_6), .B2(n_4), .ZN(p_0[3]));
   NAND2_X1 i_5 (.A1(n_6), .A2(n_4), .ZN(n_3));
   NOR2_X1 i_6 (.A1(PacketSize[2]), .A2(n_0), .ZN(n_4));
   INV_X1 i_7 (.A(n_5), .ZN(p_0[5]));
   AOI21_X1 i_8 (.A(p_0[31]), .B1(PacketSize[5]), .B2(n_1), .ZN(n_5));
   NOR2_X1 i_9 (.A1(PacketSize[5]), .A2(n_1), .ZN(p_0[31]));
   INV_X1 i_10 (.A(PacketSize[3]), .ZN(n_6));
endmodule

module datapath__1_339(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   NOR2_X1 i_0 (.A1(p_0[6]), .A2(p_0[5]), .ZN(n_0));
   INV_X1 i_1 (.A(p_0[4]), .ZN(n_1));
   INV_X1 i_2 (.A(p_0[3]), .ZN(n_2));
   NAND3_X1 i_3 (.A1(n_0), .A2(n_1), .A3(n_2), .ZN(n_3));
   INV_X1 i_4 (.A(p_0[1]), .ZN(n_4));
   INV_X1 i_5 (.A(p_0[0]), .ZN(n_5));
   INV_X1 i_6 (.A(p_0[2]), .ZN(n_6));
   NAND3_X1 i_7 (.A1(n_4), .A2(n_5), .A3(n_6), .ZN(n_7));
   NOR2_X1 i_8 (.A1(n_3), .A2(n_7), .ZN(p_1[0]));
   NAND3_X1 i_9 (.A1(n_4), .A2(n_6), .A3(p_0[0]), .ZN(n_8));
   NOR2_X1 i_10 (.A1(n_3), .A2(n_8), .ZN(p_1[1]));
   NAND3_X1 i_11 (.A1(n_6), .A2(n_5), .A3(p_0[1]), .ZN(n_9));
   NOR2_X1 i_12 (.A1(n_3), .A2(n_9), .ZN(p_1[2]));
   NAND3_X1 i_13 (.A1(n_6), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_10));
   NOR2_X1 i_14 (.A1(n_3), .A2(n_10), .ZN(p_1[3]));
   NAND3_X1 i_15 (.A1(n_4), .A2(n_5), .A3(p_0[2]), .ZN(n_11));
   NOR2_X1 i_16 (.A1(n_3), .A2(n_11), .ZN(p_1[4]));
   NAND3_X1 i_17 (.A1(n_4), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_12));
   NOR2_X1 i_18 (.A1(n_3), .A2(n_12), .ZN(p_1[5]));
   NAND3_X1 i_19 (.A1(n_5), .A2(p_0[1]), .A3(p_0[2]), .ZN(n_13));
   NOR2_X1 i_20 (.A1(n_3), .A2(n_13), .ZN(p_1[6]));
   NAND3_X1 i_21 (.A1(p_0[1]), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_14));
   NOR2_X1 i_22 (.A1(n_3), .A2(n_14), .ZN(p_1[7]));
   NAND3_X1 i_23 (.A1(n_0), .A2(n_1), .A3(p_0[3]), .ZN(n_15));
   NOR2_X1 i_24 (.A1(n_15), .A2(n_7), .ZN(p_1[8]));
   NOR2_X1 i_25 (.A1(n_15), .A2(n_8), .ZN(p_1[9]));
   NOR2_X1 i_26 (.A1(n_15), .A2(n_9), .ZN(p_1[10]));
   NOR2_X1 i_27 (.A1(n_15), .A2(n_10), .ZN(p_1[11]));
   NOR2_X1 i_28 (.A1(n_15), .A2(n_11), .ZN(p_1[12]));
   NOR2_X1 i_29 (.A1(n_15), .A2(n_12), .ZN(p_1[13]));
   NOR2_X1 i_30 (.A1(n_15), .A2(n_13), .ZN(p_1[14]));
   NOR2_X1 i_31 (.A1(n_15), .A2(n_14), .ZN(p_1[15]));
   NAND3_X1 i_32 (.A1(n_0), .A2(p_0[4]), .A3(n_2), .ZN(n_16));
   NOR2_X1 i_33 (.A1(n_16), .A2(n_7), .ZN(p_1[16]));
   NOR2_X1 i_34 (.A1(n_16), .A2(n_8), .ZN(p_1[17]));
   NOR2_X1 i_35 (.A1(n_16), .A2(n_9), .ZN(p_1[18]));
   NOR2_X1 i_36 (.A1(n_16), .A2(n_10), .ZN(p_1[19]));
   NOR2_X1 i_37 (.A1(n_16), .A2(n_11), .ZN(p_1[20]));
   NOR2_X1 i_38 (.A1(n_16), .A2(n_12), .ZN(p_1[21]));
   NOR2_X1 i_39 (.A1(n_16), .A2(n_13), .ZN(p_1[22]));
   NOR2_X1 i_40 (.A1(n_16), .A2(n_14), .ZN(p_1[23]));
   NAND3_X1 i_41 (.A1(n_0), .A2(p_0[4]), .A3(p_0[3]), .ZN(n_17));
   NOR2_X1 i_42 (.A1(n_17), .A2(n_7), .ZN(p_1[24]));
   NOR2_X1 i_43 (.A1(n_17), .A2(n_8), .ZN(p_1[25]));
   NOR2_X1 i_44 (.A1(n_17), .A2(n_9), .ZN(p_1[26]));
   NOR2_X1 i_45 (.A1(n_17), .A2(n_10), .ZN(p_1[27]));
   NOR2_X1 i_46 (.A1(n_17), .A2(n_11), .ZN(p_1[28]));
   NOR2_X1 i_47 (.A1(n_17), .A2(n_12), .ZN(p_1[29]));
   NOR2_X1 i_48 (.A1(n_17), .A2(n_13), .ZN(p_1[30]));
   NOR2_X1 i_49 (.A1(n_17), .A2(n_14), .ZN(p_1[31]));
endmodule

module datapath__1_344(PacketSize, p_0);
   input [5:0]PacketSize;
   output [31:0]p_0;

   HA_X1 i_0 (.A(PacketSize[2]), .B(n_2), .CO(n_0), .S(p_0[2]));
   HA_X1 i_1 (.A(PacketSize[4]), .B(n_3), .CO(n_1), .S(p_0[4]));
   OAI21_X1 i_2 (.A(n_2), .B1(n_7), .B2(n_6), .ZN(p_0[1]));
   NAND2_X1 i_3 (.A1(n_7), .A2(n_6), .ZN(n_2));
   OAI21_X1 i_4 (.A(n_3), .B1(n_8), .B2(n_5), .ZN(p_0[3]));
   NAND2_X1 i_5 (.A1(n_8), .A2(n_5), .ZN(n_3));
   INV_X1 i_6 (.A(n_4), .ZN(p_0[5]));
   AOI21_X1 i_7 (.A(p_0[31]), .B1(PacketSize[5]), .B2(n_1), .ZN(n_4));
   NOR2_X1 i_8 (.A1(PacketSize[5]), .A2(n_1), .ZN(p_0[31]));
   INV_X1 i_9 (.A(n_0), .ZN(n_5));
   INV_X1 i_10 (.A(PacketSize[0]), .ZN(n_6));
   INV_X1 i_11 (.A(PacketSize[1]), .ZN(n_7));
   INV_X1 i_12 (.A(PacketSize[3]), .ZN(n_8));
endmodule

module datapath__1_345(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   NOR2_X1 i_0 (.A1(p_0[6]), .A2(p_0[5]), .ZN(n_0));
   INV_X1 i_1 (.A(p_0[4]), .ZN(n_1));
   INV_X1 i_2 (.A(p_0[3]), .ZN(n_2));
   NAND3_X1 i_3 (.A1(n_0), .A2(n_1), .A3(n_2), .ZN(n_3));
   INV_X1 i_4 (.A(p_0[1]), .ZN(n_4));
   INV_X1 i_5 (.A(p_0[0]), .ZN(n_5));
   INV_X1 i_6 (.A(p_0[2]), .ZN(n_6));
   NAND3_X1 i_7 (.A1(n_4), .A2(n_5), .A3(n_6), .ZN(n_7));
   NOR2_X1 i_8 (.A1(n_3), .A2(n_7), .ZN(p_1[0]));
   NAND3_X1 i_9 (.A1(n_4), .A2(n_6), .A3(p_0[0]), .ZN(n_8));
   NOR2_X1 i_10 (.A1(n_3), .A2(n_8), .ZN(p_1[1]));
   NAND3_X1 i_11 (.A1(n_6), .A2(n_5), .A3(p_0[1]), .ZN(n_9));
   NOR2_X1 i_12 (.A1(n_3), .A2(n_9), .ZN(p_1[2]));
   NAND3_X1 i_13 (.A1(n_6), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_10));
   NOR2_X1 i_14 (.A1(n_3), .A2(n_10), .ZN(p_1[3]));
   NAND3_X1 i_15 (.A1(n_4), .A2(n_5), .A3(p_0[2]), .ZN(n_11));
   NOR2_X1 i_16 (.A1(n_3), .A2(n_11), .ZN(p_1[4]));
   NAND3_X1 i_17 (.A1(n_4), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_12));
   NOR2_X1 i_18 (.A1(n_3), .A2(n_12), .ZN(p_1[5]));
   NAND3_X1 i_19 (.A1(n_5), .A2(p_0[1]), .A3(p_0[2]), .ZN(n_13));
   NOR2_X1 i_20 (.A1(n_3), .A2(n_13), .ZN(p_1[6]));
   NAND3_X1 i_21 (.A1(p_0[1]), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_14));
   NOR2_X1 i_22 (.A1(n_3), .A2(n_14), .ZN(p_1[7]));
   NAND3_X1 i_23 (.A1(n_0), .A2(n_1), .A3(p_0[3]), .ZN(n_15));
   NOR2_X1 i_24 (.A1(n_15), .A2(n_7), .ZN(p_1[8]));
   NOR2_X1 i_25 (.A1(n_15), .A2(n_8), .ZN(p_1[9]));
   NOR2_X1 i_26 (.A1(n_15), .A2(n_9), .ZN(p_1[10]));
   NOR2_X1 i_27 (.A1(n_15), .A2(n_10), .ZN(p_1[11]));
   NOR2_X1 i_28 (.A1(n_15), .A2(n_11), .ZN(p_1[12]));
   NOR2_X1 i_29 (.A1(n_15), .A2(n_12), .ZN(p_1[13]));
   NOR2_X1 i_30 (.A1(n_15), .A2(n_13), .ZN(p_1[14]));
   NOR2_X1 i_31 (.A1(n_15), .A2(n_14), .ZN(p_1[15]));
   NAND3_X1 i_32 (.A1(n_0), .A2(p_0[4]), .A3(n_2), .ZN(n_16));
   NOR2_X1 i_33 (.A1(n_16), .A2(n_7), .ZN(p_1[16]));
   NOR2_X1 i_34 (.A1(n_16), .A2(n_8), .ZN(p_1[17]));
   NOR2_X1 i_35 (.A1(n_16), .A2(n_9), .ZN(p_1[18]));
   NOR2_X1 i_36 (.A1(n_16), .A2(n_10), .ZN(p_1[19]));
   NOR2_X1 i_37 (.A1(n_16), .A2(n_11), .ZN(p_1[20]));
   NOR2_X1 i_38 (.A1(n_16), .A2(n_12), .ZN(p_1[21]));
   NOR2_X1 i_39 (.A1(n_16), .A2(n_13), .ZN(p_1[22]));
   NOR2_X1 i_40 (.A1(n_16), .A2(n_14), .ZN(p_1[23]));
   NAND3_X1 i_41 (.A1(n_0), .A2(p_0[4]), .A3(p_0[3]), .ZN(n_17));
   NOR2_X1 i_42 (.A1(n_17), .A2(n_7), .ZN(p_1[24]));
   NOR2_X1 i_43 (.A1(n_17), .A2(n_8), .ZN(p_1[25]));
   NOR2_X1 i_44 (.A1(n_17), .A2(n_9), .ZN(p_1[26]));
   NOR2_X1 i_45 (.A1(n_17), .A2(n_10), .ZN(p_1[27]));
   NOR2_X1 i_46 (.A1(n_17), .A2(n_11), .ZN(p_1[28]));
   NOR2_X1 i_47 (.A1(n_17), .A2(n_12), .ZN(p_1[29]));
   NOR2_X1 i_48 (.A1(n_17), .A2(n_13), .ZN(p_1[30]));
   NOR2_X1 i_49 (.A1(n_17), .A2(n_14), .ZN(p_1[31]));
endmodule

module datapath__1_347(PacketSize, p_0);
   input [5:0]PacketSize;
   output [31:0]p_0;

   HA_X1 i_0 (.A(PacketSize[2]), .B(PacketSize[1]), .CO(n_0), .S(p_0[2]));
   HA_X1 i_1 (.A(PacketSize[4]), .B(n_2), .CO(n_1), .S(p_0[4]));
   OAI21_X1 i_2 (.A(n_2), .B1(n_5), .B2(n_4), .ZN(p_0[3]));
   NAND2_X1 i_3 (.A1(n_5), .A2(n_4), .ZN(n_2));
   INV_X1 i_4 (.A(n_3), .ZN(p_0[5]));
   AOI21_X1 i_5 (.A(p_0[31]), .B1(PacketSize[5]), .B2(n_1), .ZN(n_3));
   NOR2_X1 i_6 (.A1(PacketSize[5]), .A2(n_1), .ZN(p_0[31]));
   INV_X1 i_7 (.A(n_0), .ZN(n_4));
   INV_X1 i_8 (.A(PacketSize[3]), .ZN(n_5));
endmodule

module datapath__1_348(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   NOR2_X1 i_0 (.A1(p_0[6]), .A2(p_0[5]), .ZN(n_0));
   INV_X1 i_1 (.A(p_0[4]), .ZN(n_1));
   INV_X1 i_2 (.A(p_0[3]), .ZN(n_2));
   NAND3_X1 i_3 (.A1(n_0), .A2(n_1), .A3(n_2), .ZN(n_3));
   INV_X1 i_4 (.A(p_0[1]), .ZN(n_4));
   INV_X1 i_5 (.A(p_0[0]), .ZN(n_5));
   INV_X1 i_6 (.A(p_0[2]), .ZN(n_6));
   NAND3_X1 i_7 (.A1(n_4), .A2(n_5), .A3(n_6), .ZN(n_7));
   NOR2_X1 i_8 (.A1(n_3), .A2(n_7), .ZN(p_1[0]));
   NAND3_X1 i_9 (.A1(n_4), .A2(n_6), .A3(p_0[0]), .ZN(n_8));
   NOR2_X1 i_10 (.A1(n_3), .A2(n_8), .ZN(p_1[1]));
   NAND3_X1 i_11 (.A1(n_6), .A2(n_5), .A3(p_0[1]), .ZN(n_9));
   NOR2_X1 i_12 (.A1(n_3), .A2(n_9), .ZN(p_1[2]));
   NAND3_X1 i_13 (.A1(n_6), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_10));
   NOR2_X1 i_14 (.A1(n_3), .A2(n_10), .ZN(p_1[3]));
   NAND3_X1 i_15 (.A1(n_4), .A2(n_5), .A3(p_0[2]), .ZN(n_11));
   NOR2_X1 i_16 (.A1(n_3), .A2(n_11), .ZN(p_1[4]));
   NAND3_X1 i_17 (.A1(n_4), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_12));
   NOR2_X1 i_18 (.A1(n_3), .A2(n_12), .ZN(p_1[5]));
   NAND3_X1 i_19 (.A1(n_5), .A2(p_0[1]), .A3(p_0[2]), .ZN(n_13));
   NOR2_X1 i_20 (.A1(n_3), .A2(n_13), .ZN(p_1[6]));
   NAND3_X1 i_21 (.A1(p_0[1]), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_14));
   NOR2_X1 i_22 (.A1(n_3), .A2(n_14), .ZN(p_1[7]));
   NAND3_X1 i_23 (.A1(n_0), .A2(n_1), .A3(p_0[3]), .ZN(n_15));
   NOR2_X1 i_24 (.A1(n_15), .A2(n_7), .ZN(p_1[8]));
   NOR2_X1 i_25 (.A1(n_15), .A2(n_8), .ZN(p_1[9]));
   NOR2_X1 i_26 (.A1(n_15), .A2(n_9), .ZN(p_1[10]));
   NOR2_X1 i_27 (.A1(n_15), .A2(n_10), .ZN(p_1[11]));
   NOR2_X1 i_28 (.A1(n_15), .A2(n_11), .ZN(p_1[12]));
   NOR2_X1 i_29 (.A1(n_15), .A2(n_12), .ZN(p_1[13]));
   NOR2_X1 i_30 (.A1(n_15), .A2(n_13), .ZN(p_1[14]));
   NOR2_X1 i_31 (.A1(n_15), .A2(n_14), .ZN(p_1[15]));
   NAND3_X1 i_32 (.A1(n_0), .A2(p_0[4]), .A3(n_2), .ZN(n_16));
   NOR2_X1 i_33 (.A1(n_16), .A2(n_7), .ZN(p_1[16]));
   NOR2_X1 i_34 (.A1(n_16), .A2(n_8), .ZN(p_1[17]));
   NOR2_X1 i_35 (.A1(n_16), .A2(n_9), .ZN(p_1[18]));
   NOR2_X1 i_36 (.A1(n_16), .A2(n_10), .ZN(p_1[19]));
   NOR2_X1 i_37 (.A1(n_16), .A2(n_11), .ZN(p_1[20]));
   NOR2_X1 i_38 (.A1(n_16), .A2(n_12), .ZN(p_1[21]));
   NOR2_X1 i_39 (.A1(n_16), .A2(n_13), .ZN(p_1[22]));
   NOR2_X1 i_40 (.A1(n_16), .A2(n_14), .ZN(p_1[23]));
   NAND3_X1 i_41 (.A1(n_0), .A2(p_0[4]), .A3(p_0[3]), .ZN(n_17));
   NOR2_X1 i_42 (.A1(n_17), .A2(n_7), .ZN(p_1[24]));
   NOR2_X1 i_43 (.A1(n_17), .A2(n_8), .ZN(p_1[25]));
   NOR2_X1 i_44 (.A1(n_17), .A2(n_9), .ZN(p_1[26]));
   NOR2_X1 i_45 (.A1(n_17), .A2(n_10), .ZN(p_1[27]));
   NOR2_X1 i_46 (.A1(n_17), .A2(n_11), .ZN(p_1[28]));
   NOR2_X1 i_47 (.A1(n_17), .A2(n_12), .ZN(p_1[29]));
   NOR2_X1 i_48 (.A1(n_17), .A2(n_13), .ZN(p_1[30]));
   NOR2_X1 i_49 (.A1(n_17), .A2(n_14), .ZN(p_1[31]));
endmodule

module datapath__1_350(PacketSize, p_0);
   input [5:0]PacketSize;
   output [31:0]p_0;

   HA_X1 i_0 (.A(PacketSize[1]), .B(PacketSize[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_1 (.A(PacketSize[2]), .B(n_0), .CO(n_1), .S(p_0[2]));
   HA_X1 i_2 (.A(PacketSize[4]), .B(n_3), .CO(n_2), .S(p_0[4]));
   OAI21_X1 i_3 (.A(n_3), .B1(n_6), .B2(n_5), .ZN(p_0[3]));
   NAND2_X1 i_4 (.A1(n_6), .A2(n_5), .ZN(n_3));
   INV_X1 i_5 (.A(n_4), .ZN(p_0[5]));
   AOI21_X1 i_6 (.A(p_0[31]), .B1(PacketSize[5]), .B2(n_2), .ZN(n_4));
   NOR2_X1 i_7 (.A1(PacketSize[5]), .A2(n_2), .ZN(p_0[31]));
   INV_X1 i_8 (.A(n_1), .ZN(n_5));
   INV_X1 i_9 (.A(PacketSize[3]), .ZN(n_6));
endmodule

module datapath__1_351(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   NOR2_X1 i_0 (.A1(p_0[6]), .A2(p_0[5]), .ZN(n_0));
   INV_X1 i_1 (.A(p_0[4]), .ZN(n_1));
   INV_X1 i_2 (.A(p_0[3]), .ZN(n_2));
   NAND3_X1 i_3 (.A1(n_0), .A2(n_1), .A3(n_2), .ZN(n_3));
   INV_X1 i_4 (.A(p_0[1]), .ZN(n_4));
   INV_X1 i_5 (.A(p_0[0]), .ZN(n_5));
   INV_X1 i_6 (.A(p_0[2]), .ZN(n_6));
   NAND3_X1 i_7 (.A1(n_4), .A2(n_5), .A3(n_6), .ZN(n_7));
   NOR2_X1 i_8 (.A1(n_3), .A2(n_7), .ZN(p_1[0]));
   NAND3_X1 i_9 (.A1(n_4), .A2(n_6), .A3(p_0[0]), .ZN(n_8));
   NOR2_X1 i_10 (.A1(n_3), .A2(n_8), .ZN(p_1[1]));
   NAND3_X1 i_11 (.A1(n_6), .A2(n_5), .A3(p_0[1]), .ZN(n_9));
   NOR2_X1 i_12 (.A1(n_3), .A2(n_9), .ZN(p_1[2]));
   NAND3_X1 i_13 (.A1(n_6), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_10));
   NOR2_X1 i_14 (.A1(n_3), .A2(n_10), .ZN(p_1[3]));
   NAND3_X1 i_15 (.A1(n_4), .A2(n_5), .A3(p_0[2]), .ZN(n_11));
   NOR2_X1 i_16 (.A1(n_3), .A2(n_11), .ZN(p_1[4]));
   NAND3_X1 i_17 (.A1(n_4), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_12));
   NOR2_X1 i_18 (.A1(n_3), .A2(n_12), .ZN(p_1[5]));
   NAND3_X1 i_19 (.A1(n_5), .A2(p_0[1]), .A3(p_0[2]), .ZN(n_13));
   NOR2_X1 i_20 (.A1(n_3), .A2(n_13), .ZN(p_1[6]));
   NAND3_X1 i_21 (.A1(p_0[1]), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_14));
   NOR2_X1 i_22 (.A1(n_3), .A2(n_14), .ZN(p_1[7]));
   NAND3_X1 i_23 (.A1(n_0), .A2(n_1), .A3(p_0[3]), .ZN(n_15));
   NOR2_X1 i_24 (.A1(n_15), .A2(n_7), .ZN(p_1[8]));
   NOR2_X1 i_25 (.A1(n_15), .A2(n_8), .ZN(p_1[9]));
   NOR2_X1 i_26 (.A1(n_15), .A2(n_9), .ZN(p_1[10]));
   NOR2_X1 i_27 (.A1(n_15), .A2(n_10), .ZN(p_1[11]));
   NOR2_X1 i_28 (.A1(n_15), .A2(n_11), .ZN(p_1[12]));
   NOR2_X1 i_29 (.A1(n_15), .A2(n_12), .ZN(p_1[13]));
   NOR2_X1 i_30 (.A1(n_15), .A2(n_13), .ZN(p_1[14]));
   NOR2_X1 i_31 (.A1(n_15), .A2(n_14), .ZN(p_1[15]));
   NAND3_X1 i_32 (.A1(n_0), .A2(p_0[4]), .A3(n_2), .ZN(n_16));
   NOR2_X1 i_33 (.A1(n_16), .A2(n_7), .ZN(p_1[16]));
   NOR2_X1 i_34 (.A1(n_16), .A2(n_8), .ZN(p_1[17]));
   NOR2_X1 i_35 (.A1(n_16), .A2(n_9), .ZN(p_1[18]));
   NOR2_X1 i_36 (.A1(n_16), .A2(n_10), .ZN(p_1[19]));
   NOR2_X1 i_37 (.A1(n_16), .A2(n_11), .ZN(p_1[20]));
   NOR2_X1 i_38 (.A1(n_16), .A2(n_12), .ZN(p_1[21]));
   NOR2_X1 i_39 (.A1(n_16), .A2(n_13), .ZN(p_1[22]));
   NOR2_X1 i_40 (.A1(n_16), .A2(n_14), .ZN(p_1[23]));
   NAND3_X1 i_41 (.A1(n_0), .A2(p_0[4]), .A3(p_0[3]), .ZN(n_17));
   NOR2_X1 i_42 (.A1(n_17), .A2(n_7), .ZN(p_1[24]));
   NOR2_X1 i_43 (.A1(n_17), .A2(n_8), .ZN(p_1[25]));
   NOR2_X1 i_44 (.A1(n_17), .A2(n_9), .ZN(p_1[26]));
   NOR2_X1 i_45 (.A1(n_17), .A2(n_10), .ZN(p_1[27]));
   NOR2_X1 i_46 (.A1(n_17), .A2(n_11), .ZN(p_1[28]));
   NOR2_X1 i_47 (.A1(n_17), .A2(n_12), .ZN(p_1[29]));
   NOR2_X1 i_48 (.A1(n_17), .A2(n_13), .ZN(p_1[30]));
   NOR2_X1 i_49 (.A1(n_17), .A2(n_14), .ZN(p_1[31]));
endmodule

module datapath__1_355(PacketSize, p_0);
   input [5:0]PacketSize;
   output [31:0]p_0;

   HA_X1 i_0 (.A(PacketSize[3]), .B(n_3), .CO(n_0), .S(p_0[3]));
   HA_X1 i_1 (.A(PacketSize[4]), .B(n_0), .CO(n_1), .S(p_0[4]));
   INV_X1 i_2 (.A(n_2), .ZN(p_0[1]));
   AOI21_X1 i_3 (.A(n_4), .B1(PacketSize[1]), .B2(PacketSize[0]), .ZN(n_2));
   OAI21_X1 i_4 (.A(n_3), .B1(n_6), .B2(n_4), .ZN(p_0[2]));
   NAND2_X1 i_5 (.A1(n_6), .A2(n_4), .ZN(n_3));
   NOR2_X1 i_6 (.A1(PacketSize[1]), .A2(PacketSize[0]), .ZN(n_4));
   INV_X1 i_7 (.A(n_5), .ZN(p_0[5]));
   AOI21_X1 i_8 (.A(p_0[31]), .B1(PacketSize[5]), .B2(n_1), .ZN(n_5));
   NOR2_X1 i_9 (.A1(PacketSize[5]), .A2(n_1), .ZN(p_0[31]));
   INV_X1 i_10 (.A(PacketSize[2]), .ZN(n_6));
endmodule

module datapath__1_356(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   NOR2_X1 i_0 (.A1(p_0[6]), .A2(p_0[5]), .ZN(n_0));
   INV_X1 i_1 (.A(p_0[4]), .ZN(n_1));
   INV_X1 i_2 (.A(p_0[3]), .ZN(n_2));
   NAND3_X1 i_3 (.A1(n_0), .A2(n_1), .A3(n_2), .ZN(n_3));
   INV_X1 i_4 (.A(p_0[1]), .ZN(n_4));
   INV_X1 i_5 (.A(p_0[0]), .ZN(n_5));
   INV_X1 i_6 (.A(p_0[2]), .ZN(n_6));
   NAND3_X1 i_7 (.A1(n_4), .A2(n_5), .A3(n_6), .ZN(n_7));
   NOR2_X1 i_8 (.A1(n_3), .A2(n_7), .ZN(p_1[0]));
   NAND3_X1 i_9 (.A1(n_4), .A2(n_6), .A3(p_0[0]), .ZN(n_8));
   NOR2_X1 i_10 (.A1(n_3), .A2(n_8), .ZN(p_1[1]));
   NAND3_X1 i_11 (.A1(n_6), .A2(n_5), .A3(p_0[1]), .ZN(n_9));
   NOR2_X1 i_12 (.A1(n_3), .A2(n_9), .ZN(p_1[2]));
   NAND3_X1 i_13 (.A1(n_6), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_10));
   NOR2_X1 i_14 (.A1(n_3), .A2(n_10), .ZN(p_1[3]));
   NAND3_X1 i_15 (.A1(n_4), .A2(n_5), .A3(p_0[2]), .ZN(n_11));
   NOR2_X1 i_16 (.A1(n_3), .A2(n_11), .ZN(p_1[4]));
   NAND3_X1 i_17 (.A1(n_4), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_12));
   NOR2_X1 i_18 (.A1(n_3), .A2(n_12), .ZN(p_1[5]));
   NAND3_X1 i_19 (.A1(n_5), .A2(p_0[1]), .A3(p_0[2]), .ZN(n_13));
   NOR2_X1 i_20 (.A1(n_3), .A2(n_13), .ZN(p_1[6]));
   NAND3_X1 i_21 (.A1(p_0[1]), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_14));
   NOR2_X1 i_22 (.A1(n_3), .A2(n_14), .ZN(p_1[7]));
   NAND3_X1 i_23 (.A1(n_0), .A2(n_1), .A3(p_0[3]), .ZN(n_15));
   NOR2_X1 i_24 (.A1(n_15), .A2(n_7), .ZN(p_1[8]));
   NOR2_X1 i_25 (.A1(n_15), .A2(n_8), .ZN(p_1[9]));
   NOR2_X1 i_26 (.A1(n_15), .A2(n_9), .ZN(p_1[10]));
   NOR2_X1 i_27 (.A1(n_15), .A2(n_10), .ZN(p_1[11]));
   NOR2_X1 i_28 (.A1(n_15), .A2(n_11), .ZN(p_1[12]));
   NOR2_X1 i_29 (.A1(n_15), .A2(n_12), .ZN(p_1[13]));
   NOR2_X1 i_30 (.A1(n_15), .A2(n_13), .ZN(p_1[14]));
   NOR2_X1 i_31 (.A1(n_15), .A2(n_14), .ZN(p_1[15]));
   NAND3_X1 i_32 (.A1(n_0), .A2(p_0[4]), .A3(n_2), .ZN(n_16));
   NOR2_X1 i_33 (.A1(n_16), .A2(n_7), .ZN(p_1[16]));
   NOR2_X1 i_34 (.A1(n_16), .A2(n_8), .ZN(p_1[17]));
   NOR2_X1 i_35 (.A1(n_16), .A2(n_9), .ZN(p_1[18]));
   NOR2_X1 i_36 (.A1(n_16), .A2(n_10), .ZN(p_1[19]));
   NOR2_X1 i_37 (.A1(n_16), .A2(n_11), .ZN(p_1[20]));
   NOR2_X1 i_38 (.A1(n_16), .A2(n_12), .ZN(p_1[21]));
   NOR2_X1 i_39 (.A1(n_16), .A2(n_13), .ZN(p_1[22]));
   NOR2_X1 i_40 (.A1(n_16), .A2(n_14), .ZN(p_1[23]));
   NAND3_X1 i_41 (.A1(n_0), .A2(p_0[4]), .A3(p_0[3]), .ZN(n_17));
   NOR2_X1 i_42 (.A1(n_17), .A2(n_7), .ZN(p_1[24]));
   NOR2_X1 i_43 (.A1(n_17), .A2(n_8), .ZN(p_1[25]));
   NOR2_X1 i_44 (.A1(n_17), .A2(n_9), .ZN(p_1[26]));
   NOR2_X1 i_45 (.A1(n_17), .A2(n_10), .ZN(p_1[27]));
   NOR2_X1 i_46 (.A1(n_17), .A2(n_11), .ZN(p_1[28]));
   NOR2_X1 i_47 (.A1(n_17), .A2(n_12), .ZN(p_1[29]));
   NOR2_X1 i_48 (.A1(n_17), .A2(n_13), .ZN(p_1[30]));
   NOR2_X1 i_49 (.A1(n_17), .A2(n_14), .ZN(p_1[31]));
endmodule

module datapath__1_361(PacketSize, p_0);
   input [5:0]PacketSize;
   output [31:0]p_0;

   HA_X1 i_0 (.A(PacketSize[1]), .B(PacketSize[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_1 (.A(PacketSize[3]), .B(n_3), .CO(n_1), .S(p_0[3]));
   HA_X1 i_2 (.A(PacketSize[4]), .B(n_1), .CO(n_2), .S(p_0[4]));
   OAI21_X1 i_3 (.A(n_3), .B1(n_6), .B2(n_5), .ZN(p_0[2]));
   NAND2_X1 i_4 (.A1(n_6), .A2(n_5), .ZN(n_3));
   INV_X1 i_5 (.A(n_4), .ZN(p_0[5]));
   AOI21_X1 i_6 (.A(p_0[31]), .B1(PacketSize[5]), .B2(n_2), .ZN(n_4));
   NOR2_X1 i_7 (.A1(PacketSize[5]), .A2(n_2), .ZN(p_0[31]));
   INV_X1 i_8 (.A(n_0), .ZN(n_5));
   INV_X1 i_9 (.A(PacketSize[2]), .ZN(n_6));
endmodule

module datapath__1_362(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   NOR2_X1 i_0 (.A1(p_0[6]), .A2(p_0[5]), .ZN(n_0));
   INV_X1 i_1 (.A(p_0[4]), .ZN(n_1));
   INV_X1 i_2 (.A(p_0[3]), .ZN(n_2));
   NAND3_X1 i_3 (.A1(n_0), .A2(n_1), .A3(n_2), .ZN(n_3));
   INV_X1 i_4 (.A(p_0[1]), .ZN(n_4));
   INV_X1 i_5 (.A(p_0[0]), .ZN(n_5));
   INV_X1 i_6 (.A(p_0[2]), .ZN(n_6));
   NAND3_X1 i_7 (.A1(n_4), .A2(n_5), .A3(n_6), .ZN(n_7));
   NOR2_X1 i_8 (.A1(n_3), .A2(n_7), .ZN(p_1[0]));
   NAND3_X1 i_9 (.A1(n_4), .A2(n_6), .A3(p_0[0]), .ZN(n_8));
   NOR2_X1 i_10 (.A1(n_3), .A2(n_8), .ZN(p_1[1]));
   NAND3_X1 i_11 (.A1(n_6), .A2(n_5), .A3(p_0[1]), .ZN(n_9));
   NOR2_X1 i_12 (.A1(n_3), .A2(n_9), .ZN(p_1[2]));
   NAND3_X1 i_13 (.A1(n_6), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_10));
   NOR2_X1 i_14 (.A1(n_3), .A2(n_10), .ZN(p_1[3]));
   NAND3_X1 i_15 (.A1(n_4), .A2(n_5), .A3(p_0[2]), .ZN(n_11));
   NOR2_X1 i_16 (.A1(n_3), .A2(n_11), .ZN(p_1[4]));
   NAND3_X1 i_17 (.A1(n_4), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_12));
   NOR2_X1 i_18 (.A1(n_3), .A2(n_12), .ZN(p_1[5]));
   NAND3_X1 i_19 (.A1(n_5), .A2(p_0[1]), .A3(p_0[2]), .ZN(n_13));
   NOR2_X1 i_20 (.A1(n_3), .A2(n_13), .ZN(p_1[6]));
   NAND3_X1 i_21 (.A1(p_0[1]), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_14));
   NOR2_X1 i_22 (.A1(n_3), .A2(n_14), .ZN(p_1[7]));
   NAND3_X1 i_23 (.A1(n_0), .A2(n_1), .A3(p_0[3]), .ZN(n_15));
   NOR2_X1 i_24 (.A1(n_15), .A2(n_7), .ZN(p_1[8]));
   NOR2_X1 i_25 (.A1(n_15), .A2(n_8), .ZN(p_1[9]));
   NOR2_X1 i_26 (.A1(n_15), .A2(n_9), .ZN(p_1[10]));
   NOR2_X1 i_27 (.A1(n_15), .A2(n_10), .ZN(p_1[11]));
   NOR2_X1 i_28 (.A1(n_15), .A2(n_11), .ZN(p_1[12]));
   NOR2_X1 i_29 (.A1(n_15), .A2(n_12), .ZN(p_1[13]));
   NOR2_X1 i_30 (.A1(n_15), .A2(n_13), .ZN(p_1[14]));
   NOR2_X1 i_31 (.A1(n_15), .A2(n_14), .ZN(p_1[15]));
   NAND3_X1 i_32 (.A1(n_0), .A2(p_0[4]), .A3(n_2), .ZN(n_16));
   NOR2_X1 i_33 (.A1(n_16), .A2(n_7), .ZN(p_1[16]));
   NOR2_X1 i_34 (.A1(n_16), .A2(n_8), .ZN(p_1[17]));
   NOR2_X1 i_35 (.A1(n_16), .A2(n_9), .ZN(p_1[18]));
   NOR2_X1 i_36 (.A1(n_16), .A2(n_10), .ZN(p_1[19]));
   NOR2_X1 i_37 (.A1(n_16), .A2(n_11), .ZN(p_1[20]));
   NOR2_X1 i_38 (.A1(n_16), .A2(n_12), .ZN(p_1[21]));
   NOR2_X1 i_39 (.A1(n_16), .A2(n_13), .ZN(p_1[22]));
   NOR2_X1 i_40 (.A1(n_16), .A2(n_14), .ZN(p_1[23]));
   NAND3_X1 i_41 (.A1(n_0), .A2(p_0[4]), .A3(p_0[3]), .ZN(n_17));
   NOR2_X1 i_42 (.A1(n_17), .A2(n_7), .ZN(p_1[24]));
   NOR2_X1 i_43 (.A1(n_17), .A2(n_8), .ZN(p_1[25]));
   NOR2_X1 i_44 (.A1(n_17), .A2(n_9), .ZN(p_1[26]));
   NOR2_X1 i_45 (.A1(n_17), .A2(n_10), .ZN(p_1[27]));
   NOR2_X1 i_46 (.A1(n_17), .A2(n_11), .ZN(p_1[28]));
   NOR2_X1 i_47 (.A1(n_17), .A2(n_12), .ZN(p_1[29]));
   NOR2_X1 i_48 (.A1(n_17), .A2(n_13), .ZN(p_1[30]));
   NOR2_X1 i_49 (.A1(n_17), .A2(n_14), .ZN(p_1[31]));
endmodule

module datapath__1_366(PacketSize, p_0);
   input [5:0]PacketSize;
   output [31:0]p_0;

   HA_X1 i_0 (.A(PacketSize[2]), .B(n_3), .CO(n_0), .S(p_0[2]));
   HA_X1 i_1 (.A(PacketSize[3]), .B(n_0), .CO(n_1), .S(p_0[3]));
   HA_X1 i_2 (.A(PacketSize[4]), .B(n_1), .CO(n_2), .S(p_0[4]));
   OAI21_X1 i_3 (.A(n_3), .B1(n_6), .B2(n_5), .ZN(p_0[1]));
   NAND2_X1 i_4 (.A1(n_6), .A2(n_5), .ZN(n_3));
   INV_X1 i_5 (.A(n_4), .ZN(p_0[5]));
   AOI21_X1 i_6 (.A(p_0[31]), .B1(PacketSize[5]), .B2(n_2), .ZN(n_4));
   NOR2_X1 i_7 (.A1(PacketSize[5]), .A2(n_2), .ZN(p_0[31]));
   INV_X1 i_8 (.A(PacketSize[0]), .ZN(n_5));
   INV_X1 i_9 (.A(PacketSize[1]), .ZN(n_6));
endmodule

module datapath__1_367(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   NOR2_X1 i_0 (.A1(p_0[6]), .A2(p_0[5]), .ZN(n_0));
   INV_X1 i_1 (.A(p_0[4]), .ZN(n_1));
   INV_X1 i_2 (.A(p_0[3]), .ZN(n_2));
   NAND3_X1 i_3 (.A1(n_0), .A2(n_1), .A3(n_2), .ZN(n_3));
   INV_X1 i_4 (.A(p_0[1]), .ZN(n_4));
   INV_X1 i_5 (.A(p_0[0]), .ZN(n_5));
   INV_X1 i_6 (.A(p_0[2]), .ZN(n_6));
   NAND3_X1 i_7 (.A1(n_4), .A2(n_5), .A3(n_6), .ZN(n_7));
   NOR2_X1 i_8 (.A1(n_3), .A2(n_7), .ZN(p_1[0]));
   NAND3_X1 i_9 (.A1(n_4), .A2(n_6), .A3(p_0[0]), .ZN(n_8));
   NOR2_X1 i_10 (.A1(n_3), .A2(n_8), .ZN(p_1[1]));
   NAND3_X1 i_11 (.A1(n_6), .A2(n_5), .A3(p_0[1]), .ZN(n_9));
   NOR2_X1 i_12 (.A1(n_3), .A2(n_9), .ZN(p_1[2]));
   NAND3_X1 i_13 (.A1(n_6), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_10));
   NOR2_X1 i_14 (.A1(n_3), .A2(n_10), .ZN(p_1[3]));
   NAND3_X1 i_15 (.A1(n_4), .A2(n_5), .A3(p_0[2]), .ZN(n_11));
   NOR2_X1 i_16 (.A1(n_3), .A2(n_11), .ZN(p_1[4]));
   NAND3_X1 i_17 (.A1(n_4), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_12));
   NOR2_X1 i_18 (.A1(n_3), .A2(n_12), .ZN(p_1[5]));
   NAND3_X1 i_19 (.A1(n_5), .A2(p_0[1]), .A3(p_0[2]), .ZN(n_13));
   NOR2_X1 i_20 (.A1(n_3), .A2(n_13), .ZN(p_1[6]));
   NAND3_X1 i_21 (.A1(p_0[1]), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_14));
   NOR2_X1 i_22 (.A1(n_3), .A2(n_14), .ZN(p_1[7]));
   NAND3_X1 i_23 (.A1(n_0), .A2(n_1), .A3(p_0[3]), .ZN(n_15));
   NOR2_X1 i_24 (.A1(n_15), .A2(n_7), .ZN(p_1[8]));
   NOR2_X1 i_25 (.A1(n_15), .A2(n_8), .ZN(p_1[9]));
   NOR2_X1 i_26 (.A1(n_15), .A2(n_9), .ZN(p_1[10]));
   NOR2_X1 i_27 (.A1(n_15), .A2(n_10), .ZN(p_1[11]));
   NOR2_X1 i_28 (.A1(n_15), .A2(n_11), .ZN(p_1[12]));
   NOR2_X1 i_29 (.A1(n_15), .A2(n_12), .ZN(p_1[13]));
   NOR2_X1 i_30 (.A1(n_15), .A2(n_13), .ZN(p_1[14]));
   NOR2_X1 i_31 (.A1(n_15), .A2(n_14), .ZN(p_1[15]));
   NAND3_X1 i_32 (.A1(n_0), .A2(p_0[4]), .A3(n_2), .ZN(n_16));
   NOR2_X1 i_33 (.A1(n_16), .A2(n_7), .ZN(p_1[16]));
   NOR2_X1 i_34 (.A1(n_16), .A2(n_8), .ZN(p_1[17]));
   NOR2_X1 i_35 (.A1(n_16), .A2(n_9), .ZN(p_1[18]));
   NOR2_X1 i_36 (.A1(n_16), .A2(n_10), .ZN(p_1[19]));
   NOR2_X1 i_37 (.A1(n_16), .A2(n_11), .ZN(p_1[20]));
   NOR2_X1 i_38 (.A1(n_16), .A2(n_12), .ZN(p_1[21]));
   NOR2_X1 i_39 (.A1(n_16), .A2(n_13), .ZN(p_1[22]));
   NOR2_X1 i_40 (.A1(n_16), .A2(n_14), .ZN(p_1[23]));
   NAND3_X1 i_41 (.A1(n_0), .A2(p_0[4]), .A3(p_0[3]), .ZN(n_17));
   NOR2_X1 i_42 (.A1(n_17), .A2(n_7), .ZN(p_1[24]));
   NOR2_X1 i_43 (.A1(n_17), .A2(n_8), .ZN(p_1[25]));
   NOR2_X1 i_44 (.A1(n_17), .A2(n_9), .ZN(p_1[26]));
   NOR2_X1 i_45 (.A1(n_17), .A2(n_10), .ZN(p_1[27]));
   NOR2_X1 i_46 (.A1(n_17), .A2(n_11), .ZN(p_1[28]));
   NOR2_X1 i_47 (.A1(n_17), .A2(n_12), .ZN(p_1[29]));
   NOR2_X1 i_48 (.A1(n_17), .A2(n_13), .ZN(p_1[30]));
   NOR2_X1 i_49 (.A1(n_17), .A2(n_14), .ZN(p_1[31]));
endmodule

module datapath__1_369(PacketSize, p_0);
   input [5:0]PacketSize;
   output [31:0]p_0;

   HA_X1 i_0 (.A(PacketSize[2]), .B(PacketSize[1]), .CO(n_0), .S(p_0[2]));
   HA_X1 i_1 (.A(PacketSize[3]), .B(n_0), .CO(n_1), .S(p_0[3]));
   HA_X1 i_2 (.A(PacketSize[4]), .B(n_1), .CO(n_2), .S(p_0[4]));
   INV_X1 i_3 (.A(n_3), .ZN(p_0[5]));
   AOI21_X1 i_4 (.A(p_0[31]), .B1(PacketSize[5]), .B2(n_2), .ZN(n_3));
   NOR2_X1 i_5 (.A1(PacketSize[5]), .A2(n_2), .ZN(p_0[31]));
endmodule

module datapath__1_370(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   NOR2_X1 i_0 (.A1(p_0[6]), .A2(p_0[5]), .ZN(n_0));
   INV_X1 i_1 (.A(p_0[4]), .ZN(n_1));
   INV_X1 i_2 (.A(p_0[3]), .ZN(n_2));
   NAND3_X1 i_3 (.A1(n_0), .A2(n_1), .A3(n_2), .ZN(n_3));
   INV_X1 i_4 (.A(p_0[1]), .ZN(n_4));
   INV_X1 i_5 (.A(p_0[0]), .ZN(n_5));
   INV_X1 i_6 (.A(p_0[2]), .ZN(n_6));
   NAND3_X1 i_7 (.A1(n_4), .A2(n_5), .A3(n_6), .ZN(n_7));
   NOR2_X1 i_8 (.A1(n_3), .A2(n_7), .ZN(p_1[0]));
   NAND3_X1 i_9 (.A1(n_4), .A2(n_6), .A3(p_0[0]), .ZN(n_8));
   NOR2_X1 i_10 (.A1(n_3), .A2(n_8), .ZN(p_1[1]));
   NAND3_X1 i_11 (.A1(n_6), .A2(n_5), .A3(p_0[1]), .ZN(n_9));
   NOR2_X1 i_12 (.A1(n_3), .A2(n_9), .ZN(p_1[2]));
   NAND3_X1 i_13 (.A1(n_6), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_10));
   NOR2_X1 i_14 (.A1(n_3), .A2(n_10), .ZN(p_1[3]));
   NAND3_X1 i_15 (.A1(n_4), .A2(n_5), .A3(p_0[2]), .ZN(n_11));
   NOR2_X1 i_16 (.A1(n_3), .A2(n_11), .ZN(p_1[4]));
   NAND3_X1 i_17 (.A1(n_4), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_12));
   NOR2_X1 i_18 (.A1(n_3), .A2(n_12), .ZN(p_1[5]));
   NAND3_X1 i_19 (.A1(n_5), .A2(p_0[1]), .A3(p_0[2]), .ZN(n_13));
   NOR2_X1 i_20 (.A1(n_3), .A2(n_13), .ZN(p_1[6]));
   NAND3_X1 i_21 (.A1(p_0[1]), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_14));
   NOR2_X1 i_22 (.A1(n_3), .A2(n_14), .ZN(p_1[7]));
   NAND3_X1 i_23 (.A1(n_0), .A2(n_1), .A3(p_0[3]), .ZN(n_15));
   NOR2_X1 i_24 (.A1(n_15), .A2(n_7), .ZN(p_1[8]));
   NOR2_X1 i_25 (.A1(n_15), .A2(n_8), .ZN(p_1[9]));
   NOR2_X1 i_26 (.A1(n_15), .A2(n_9), .ZN(p_1[10]));
   NOR2_X1 i_27 (.A1(n_15), .A2(n_10), .ZN(p_1[11]));
   NOR2_X1 i_28 (.A1(n_15), .A2(n_11), .ZN(p_1[12]));
   NOR2_X1 i_29 (.A1(n_15), .A2(n_12), .ZN(p_1[13]));
   NOR2_X1 i_30 (.A1(n_15), .A2(n_13), .ZN(p_1[14]));
   NOR2_X1 i_31 (.A1(n_15), .A2(n_14), .ZN(p_1[15]));
   NAND3_X1 i_32 (.A1(n_0), .A2(p_0[4]), .A3(n_2), .ZN(n_16));
   NOR2_X1 i_33 (.A1(n_16), .A2(n_7), .ZN(p_1[16]));
   NOR2_X1 i_34 (.A1(n_16), .A2(n_8), .ZN(p_1[17]));
   NOR2_X1 i_35 (.A1(n_16), .A2(n_9), .ZN(p_1[18]));
   NOR2_X1 i_36 (.A1(n_16), .A2(n_10), .ZN(p_1[19]));
   NOR2_X1 i_37 (.A1(n_16), .A2(n_11), .ZN(p_1[20]));
   NOR2_X1 i_38 (.A1(n_16), .A2(n_12), .ZN(p_1[21]));
   NOR2_X1 i_39 (.A1(n_16), .A2(n_13), .ZN(p_1[22]));
   NOR2_X1 i_40 (.A1(n_16), .A2(n_14), .ZN(p_1[23]));
   NAND3_X1 i_41 (.A1(n_0), .A2(p_0[4]), .A3(p_0[3]), .ZN(n_17));
   NOR2_X1 i_42 (.A1(n_17), .A2(n_7), .ZN(p_1[24]));
   NOR2_X1 i_43 (.A1(n_17), .A2(n_8), .ZN(p_1[25]));
   NOR2_X1 i_44 (.A1(n_17), .A2(n_9), .ZN(p_1[26]));
   NOR2_X1 i_45 (.A1(n_17), .A2(n_10), .ZN(p_1[27]));
   NOR2_X1 i_46 (.A1(n_17), .A2(n_11), .ZN(p_1[28]));
   NOR2_X1 i_47 (.A1(n_17), .A2(n_12), .ZN(p_1[29]));
   NOR2_X1 i_48 (.A1(n_17), .A2(n_13), .ZN(p_1[30]));
   NOR2_X1 i_49 (.A1(n_17), .A2(n_14), .ZN(p_1[31]));
endmodule

module datapath__1_372(PacketSize, p_0);
   input [5:0]PacketSize;
   output [31:0]p_0;

   HA_X1 i_0 (.A(PacketSize[1]), .B(PacketSize[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_1 (.A(PacketSize[2]), .B(n_0), .CO(n_1), .S(p_0[2]));
   HA_X1 i_2 (.A(PacketSize[3]), .B(n_1), .CO(n_2), .S(p_0[3]));
   HA_X1 i_3 (.A(PacketSize[4]), .B(n_2), .CO(n_3), .S(p_0[4]));
   INV_X1 i_4 (.A(n_4), .ZN(p_0[5]));
   AOI21_X1 i_5 (.A(p_0[31]), .B1(PacketSize[5]), .B2(n_3), .ZN(n_4));
   NOR2_X1 i_6 (.A1(PacketSize[5]), .A2(n_3), .ZN(p_0[31]));
endmodule

module datapath__1_373(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   NOR2_X1 i_0 (.A1(p_0[6]), .A2(p_0[5]), .ZN(n_0));
   INV_X1 i_1 (.A(p_0[4]), .ZN(n_1));
   INV_X1 i_2 (.A(p_0[3]), .ZN(n_2));
   NAND3_X1 i_3 (.A1(n_0), .A2(n_1), .A3(n_2), .ZN(n_3));
   INV_X1 i_4 (.A(p_0[1]), .ZN(n_4));
   INV_X1 i_5 (.A(p_0[0]), .ZN(n_5));
   INV_X1 i_6 (.A(p_0[2]), .ZN(n_6));
   NAND3_X1 i_7 (.A1(n_4), .A2(n_5), .A3(n_6), .ZN(n_7));
   NOR2_X1 i_8 (.A1(n_3), .A2(n_7), .ZN(p_1[0]));
   NAND3_X1 i_9 (.A1(n_4), .A2(n_6), .A3(p_0[0]), .ZN(n_8));
   NOR2_X1 i_10 (.A1(n_3), .A2(n_8), .ZN(p_1[1]));
   NAND3_X1 i_11 (.A1(n_6), .A2(n_5), .A3(p_0[1]), .ZN(n_9));
   NOR2_X1 i_12 (.A1(n_3), .A2(n_9), .ZN(p_1[2]));
   NAND3_X1 i_13 (.A1(n_6), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_10));
   NOR2_X1 i_14 (.A1(n_3), .A2(n_10), .ZN(p_1[3]));
   NAND3_X1 i_15 (.A1(n_4), .A2(n_5), .A3(p_0[2]), .ZN(n_11));
   NOR2_X1 i_16 (.A1(n_3), .A2(n_11), .ZN(p_1[4]));
   NAND3_X1 i_17 (.A1(n_4), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_12));
   NOR2_X1 i_18 (.A1(n_3), .A2(n_12), .ZN(p_1[5]));
   NAND3_X1 i_19 (.A1(n_5), .A2(p_0[1]), .A3(p_0[2]), .ZN(n_13));
   NOR2_X1 i_20 (.A1(n_3), .A2(n_13), .ZN(p_1[6]));
   NAND3_X1 i_21 (.A1(p_0[1]), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_14));
   NOR2_X1 i_22 (.A1(n_3), .A2(n_14), .ZN(p_1[7]));
   NAND3_X1 i_23 (.A1(n_0), .A2(n_1), .A3(p_0[3]), .ZN(n_15));
   NOR2_X1 i_24 (.A1(n_15), .A2(n_7), .ZN(p_1[8]));
   NOR2_X1 i_25 (.A1(n_15), .A2(n_8), .ZN(p_1[9]));
   NOR2_X1 i_26 (.A1(n_15), .A2(n_9), .ZN(p_1[10]));
   NOR2_X1 i_27 (.A1(n_15), .A2(n_10), .ZN(p_1[11]));
   NOR2_X1 i_28 (.A1(n_15), .A2(n_11), .ZN(p_1[12]));
   NOR2_X1 i_29 (.A1(n_15), .A2(n_12), .ZN(p_1[13]));
   NOR2_X1 i_30 (.A1(n_15), .A2(n_13), .ZN(p_1[14]));
   NOR2_X1 i_31 (.A1(n_15), .A2(n_14), .ZN(p_1[15]));
   NAND3_X1 i_32 (.A1(n_0), .A2(p_0[4]), .A3(n_2), .ZN(n_16));
   NOR2_X1 i_33 (.A1(n_16), .A2(n_7), .ZN(p_1[16]));
   NOR2_X1 i_34 (.A1(n_16), .A2(n_8), .ZN(p_1[17]));
   NOR2_X1 i_35 (.A1(n_16), .A2(n_9), .ZN(p_1[18]));
   NOR2_X1 i_36 (.A1(n_16), .A2(n_10), .ZN(p_1[19]));
   NOR2_X1 i_37 (.A1(n_16), .A2(n_11), .ZN(p_1[20]));
   NOR2_X1 i_38 (.A1(n_16), .A2(n_12), .ZN(p_1[21]));
   NOR2_X1 i_39 (.A1(n_16), .A2(n_13), .ZN(p_1[22]));
   NOR2_X1 i_40 (.A1(n_16), .A2(n_14), .ZN(p_1[23]));
   NAND3_X1 i_41 (.A1(n_0), .A2(p_0[4]), .A3(p_0[3]), .ZN(n_17));
   NOR2_X1 i_42 (.A1(n_17), .A2(n_7), .ZN(p_1[24]));
   NOR2_X1 i_43 (.A1(n_17), .A2(n_8), .ZN(p_1[25]));
   NOR2_X1 i_44 (.A1(n_17), .A2(n_9), .ZN(p_1[26]));
   NOR2_X1 i_45 (.A1(n_17), .A2(n_10), .ZN(p_1[27]));
   NOR2_X1 i_46 (.A1(n_17), .A2(n_11), .ZN(p_1[28]));
   NOR2_X1 i_47 (.A1(n_17), .A2(n_12), .ZN(p_1[29]));
   NOR2_X1 i_48 (.A1(n_17), .A2(n_13), .ZN(p_1[30]));
   NOR2_X1 i_49 (.A1(n_17), .A2(n_14), .ZN(p_1[31]));
endmodule

module datapath__1_378(PacketSize, p_0);
   input [5:0]PacketSize;
   output [31:0]p_0;

   HA_X1 i_0 (.A(PacketSize[5]), .B(n_4), .CO(n_1), .S(n_0));
   INV_X1 i_1 (.A(n_2), .ZN(p_0[1]));
   AOI21_X1 i_2 (.A(n_7), .B1(PacketSize[1]), .B2(PacketSize[0]), .ZN(n_2));
   OAI21_X1 i_3 (.A(n_6), .B1(n_8), .B2(n_7), .ZN(p_0[2]));
   INV_X1 i_4 (.A(n_3), .ZN(p_0[3]));
   AOI21_X1 i_5 (.A(n_5), .B1(PacketSize[3]), .B2(n_6), .ZN(n_3));
   OAI21_X1 i_6 (.A(n_4), .B1(n_9), .B2(n_5), .ZN(p_0[4]));
   NAND2_X1 i_7 (.A1(n_9), .A2(n_5), .ZN(n_4));
   NOR2_X1 i_8 (.A1(PacketSize[3]), .A2(n_6), .ZN(n_5));
   NAND2_X1 i_9 (.A1(n_8), .A2(n_7), .ZN(n_6));
   NOR2_X1 i_10 (.A1(PacketSize[1]), .A2(PacketSize[0]), .ZN(n_7));
   INV_X1 i_11 (.A(n_1), .ZN(p_0[31]));
   INV_X1 i_12 (.A(PacketSize[2]), .ZN(n_8));
   INV_X1 i_13 (.A(PacketSize[4]), .ZN(n_9));
endmodule

module datapath__1_379(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   INV_X1 i_0 (.A(p_0[1]), .ZN(n_0));
   INV_X1 i_1 (.A(p_0[0]), .ZN(n_1));
   INV_X1 i_2 (.A(p_0[2]), .ZN(n_2));
   NAND3_X1 i_3 (.A1(n_0), .A2(n_1), .A3(n_2), .ZN(n_3));
   INV_X1 i_4 (.A(p_0[4]), .ZN(n_4));
   INV_X1 i_5 (.A(p_0[3]), .ZN(n_5));
   INV_X1 i_6 (.A(p_0[6]), .ZN(n_6));
   NAND3_X1 i_7 (.A1(n_4), .A2(n_5), .A3(n_6), .ZN(n_7));
   NOR2_X1 i_8 (.A1(n_3), .A2(n_7), .ZN(p_1[0]));
   NAND3_X1 i_9 (.A1(n_0), .A2(n_2), .A3(p_0[0]), .ZN(n_8));
   NOR2_X1 i_10 (.A1(n_7), .A2(n_8), .ZN(p_1[1]));
   NAND3_X1 i_11 (.A1(n_2), .A2(n_1), .A3(p_0[1]), .ZN(n_9));
   NOR2_X1 i_12 (.A1(n_7), .A2(n_9), .ZN(p_1[2]));
   NAND3_X1 i_13 (.A1(n_2), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_10));
   NOR2_X1 i_14 (.A1(n_7), .A2(n_10), .ZN(p_1[3]));
   NAND3_X1 i_15 (.A1(n_0), .A2(n_1), .A3(p_0[2]), .ZN(n_11));
   NOR2_X1 i_16 (.A1(n_7), .A2(n_11), .ZN(p_1[4]));
   NAND3_X1 i_17 (.A1(n_0), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_12));
   NOR2_X1 i_18 (.A1(n_7), .A2(n_12), .ZN(p_1[5]));
   NAND3_X1 i_19 (.A1(n_1), .A2(p_0[1]), .A3(p_0[2]), .ZN(n_13));
   NOR2_X1 i_20 (.A1(n_7), .A2(n_13), .ZN(p_1[6]));
   NAND3_X1 i_21 (.A1(p_0[1]), .A2(p_0[0]), .A3(p_0[2]), .ZN(n_14));
   NOR2_X1 i_22 (.A1(n_7), .A2(n_14), .ZN(p_1[7]));
   NAND3_X1 i_23 (.A1(n_4), .A2(n_6), .A3(p_0[3]), .ZN(n_15));
   NOR2_X1 i_24 (.A1(n_3), .A2(n_15), .ZN(p_1[8]));
   NOR2_X1 i_25 (.A1(n_8), .A2(n_15), .ZN(p_1[9]));
   NOR2_X1 i_26 (.A1(n_9), .A2(n_15), .ZN(p_1[10]));
   NOR2_X1 i_27 (.A1(n_15), .A2(n_10), .ZN(p_1[11]));
   NOR2_X1 i_28 (.A1(n_11), .A2(n_15), .ZN(p_1[12]));
   NOR2_X1 i_29 (.A1(n_15), .A2(n_12), .ZN(p_1[13]));
   NOR2_X1 i_30 (.A1(n_15), .A2(n_13), .ZN(p_1[14]));
   NOR2_X1 i_31 (.A1(n_15), .A2(n_14), .ZN(p_1[15]));
   NAND3_X1 i_32 (.A1(n_6), .A2(n_5), .A3(p_0[4]), .ZN(n_16));
   NOR2_X1 i_33 (.A1(n_3), .A2(n_16), .ZN(p_1[16]));
   NOR2_X1 i_34 (.A1(n_8), .A2(n_16), .ZN(p_1[17]));
   NOR2_X1 i_35 (.A1(n_9), .A2(n_16), .ZN(p_1[18]));
   NOR2_X1 i_36 (.A1(n_16), .A2(n_10), .ZN(p_1[19]));
   NOR2_X1 i_37 (.A1(n_11), .A2(n_16), .ZN(p_1[20]));
   NOR2_X1 i_38 (.A1(n_16), .A2(n_12), .ZN(p_1[21]));
   NOR2_X1 i_39 (.A1(n_16), .A2(n_13), .ZN(p_1[22]));
   NOR2_X1 i_40 (.A1(n_16), .A2(n_14), .ZN(p_1[23]));
   NAND3_X1 i_41 (.A1(n_6), .A2(p_0[4]), .A3(p_0[3]), .ZN(n_17));
   NOR2_X1 i_42 (.A1(n_3), .A2(n_17), .ZN(p_1[24]));
   NOR2_X1 i_43 (.A1(n_8), .A2(n_17), .ZN(p_1[25]));
   NOR2_X1 i_44 (.A1(n_9), .A2(n_17), .ZN(p_1[26]));
   NOR2_X1 i_45 (.A1(n_10), .A2(n_17), .ZN(p_1[27]));
   NOR2_X1 i_46 (.A1(n_11), .A2(n_17), .ZN(p_1[28]));
   NOR2_X1 i_47 (.A1(n_12), .A2(n_17), .ZN(p_1[29]));
   NOR2_X1 i_48 (.A1(n_13), .A2(n_17), .ZN(p_1[30]));
   NOR2_X1 i_49 (.A1(n_17), .A2(n_14), .ZN(p_1[31]));
endmodule

module datapath__0_22(PacketSize, p_0);
   input [5:0]PacketSize;
   output [11:0]p_0;

   INV_X1 i_0 (.A(PacketSize[1]), .ZN(p_0[1]));
   INV_X1 i_1 (.A(PacketSize[2]), .ZN(p_0[2]));
   INV_X1 i_2 (.A(PacketSize[3]), .ZN(p_0[3]));
   INV_X1 i_3 (.A(PacketSize[4]), .ZN(p_0[4]));
   INV_X1 i_4 (.A(PacketSize[5]), .ZN(p_0[5]));
   INV_X1 i_5 (.A(PacketSize[0]), .ZN(p_0[6]));
endmodule

module datapath__0_24(p_0, Small_Packet_Indication_Bit_Location, p_1);
   input [11:0]p_0;
   input [5:0]Small_Packet_Indication_Bit_Location;
   output [5:0]p_1;

   OR2_X1 i_0 (.A1(p_0[0]), .A2(Small_Packet_Indication_Bit_Location[0]), 
      .ZN(n_0));
   NAND2_X1 i_1 (.A1(p_0[0]), .A2(Small_Packet_Indication_Bit_Location[0]), 
      .ZN(n_1));
   NAND2_X1 i_2 (.A1(n_0), .A2(n_1), .ZN(n_2));
   XNOR2_X1 i_3 (.A(n_2), .B(p_0[6]), .ZN(p_1[0]));
   NAND2_X1 i_4 (.A1(n_0), .A2(p_0[6]), .ZN(n_3));
   NAND2_X1 i_5 (.A1(n_3), .A2(n_1), .ZN(n_4));
   OR2_X1 i_6 (.A1(p_0[1]), .A2(Small_Packet_Indication_Bit_Location[1]), 
      .ZN(n_5));
   NAND2_X1 i_7 (.A1(p_0[1]), .A2(Small_Packet_Indication_Bit_Location[1]), 
      .ZN(n_6));
   NAND2_X1 i_8 (.A1(n_5), .A2(n_6), .ZN(n_7));
   XNOR2_X1 i_9 (.A(n_4), .B(n_7), .ZN(p_1[1]));
   NOR2_X1 i_10 (.A1(p_0[2]), .A2(Small_Packet_Indication_Bit_Location[2]), 
      .ZN(n_8));
   INV_X1 i_11 (.A(n_8), .ZN(n_9));
   NAND2_X1 i_12 (.A1(p_0[2]), .A2(Small_Packet_Indication_Bit_Location[2]), 
      .ZN(n_10));
   NAND2_X1 i_13 (.A1(n_9), .A2(n_10), .ZN(n_11));
   INV_X1 i_14 (.A(n_6), .ZN(n_12));
   OAI21_X1 i_15 (.A(n_5), .B1(n_4), .B2(n_12), .ZN(n_13));
   XOR2_X1 i_16 (.A(n_11), .B(n_13), .Z(p_1[2]));
   OAI21_X1 i_17 (.A(n_10), .B1(n_13), .B2(n_8), .ZN(n_14));
   OR2_X1 i_18 (.A1(p_0[3]), .A2(Small_Packet_Indication_Bit_Location[3]), 
      .ZN(n_15));
   NAND2_X1 i_19 (.A1(p_0[3]), .A2(Small_Packet_Indication_Bit_Location[3]), 
      .ZN(n_16));
   NAND2_X1 i_20 (.A1(n_15), .A2(n_16), .ZN(n_17));
   XNOR2_X1 i_21 (.A(n_14), .B(n_17), .ZN(p_1[3]));
   NAND2_X1 i_22 (.A1(n_5), .A2(n_9), .ZN(n_18));
   OAI211_X1 i_23 (.A(n_10), .B(n_16), .C1(n_18), .C2(n_3), .ZN(n_19));
   AOI21_X1 i_24 (.A(n_18), .B1(n_1), .B2(n_6), .ZN(n_20));
   OAI21_X1 i_25 (.A(n_15), .B1(n_19), .B2(n_20), .ZN(n_21));
   NAND2_X1 i_26 (.A1(p_0[4]), .A2(Small_Packet_Indication_Bit_Location[4]), 
      .ZN(n_22));
   INV_X1 i_27 (.A(n_22), .ZN(n_23));
   NOR2_X1 i_28 (.A1(p_0[4]), .A2(Small_Packet_Indication_Bit_Location[4]), 
      .ZN(n_24));
   NOR2_X1 i_29 (.A1(n_23), .A2(n_24), .ZN(n_25));
   XNOR2_X1 i_30 (.A(n_21), .B(n_25), .ZN(p_1[4]));
   OAI21_X1 i_31 (.A(n_22), .B1(n_21), .B2(n_24), .ZN(n_26));
   XNOR2_X1 i_32 (.A(p_0[5]), .B(Small_Packet_Indication_Bit_Location[5]), 
      .ZN(n_27));
   XNOR2_X1 i_33 (.A(n_26), .B(n_27), .ZN(p_1[5]));
endmodule

module datapath__0_196(p_0, Data_Size, p_1);
   input [31:0]p_0;
   input [5:0]Data_Size;
   output [31:0]p_1;

   INV_X1 i_0 (.A(n_0), .ZN(p_1[0]));
   OAI21_X1 i_1 (.A(n_70), .B1(p_0[0]), .B2(Data_Size[0]), .ZN(n_0));
   XOR2_X1 i_2 (.A(n_70), .B(n_1), .Z(p_1[1]));
   OAI21_X1 i_3 (.A(n_69), .B1(p_0[1]), .B2(Data_Size[1]), .ZN(n_1));
   XNOR2_X1 i_4 (.A(n_68), .B(n_2), .ZN(p_1[2]));
   OAI21_X1 i_5 (.A(n_72), .B1(p_0[2]), .B2(Data_Size[2]), .ZN(n_2));
   XOR2_X1 i_6 (.A(n_66), .B(n_3), .Z(p_1[3]));
   NOR2_X1 i_7 (.A1(n_74), .A2(n_73), .ZN(n_3));
   XNOR2_X1 i_8 (.A(n_64), .B(n_4), .ZN(p_1[4]));
   OAI21_X1 i_9 (.A(n_62), .B1(p_0[4]), .B2(Data_Size[4]), .ZN(n_4));
   XNOR2_X1 i_10 (.A(n_60), .B(n_5), .ZN(p_1[5]));
   OAI21_X1 i_11 (.A(n_63), .B1(p_0[5]), .B2(Data_Size[5]), .ZN(n_5));
   INV_X1 i_12 (.A(n_6), .ZN(p_1[6]));
   OAI21_X1 i_13 (.A(n_57), .B1(p_0[6]), .B2(n_58), .ZN(n_6));
   INV_X1 i_14 (.A(n_7), .ZN(p_1[7]));
   OAI21_X1 i_15 (.A(n_55), .B1(p_0[7]), .B2(n_56), .ZN(n_7));
   INV_X1 i_16 (.A(n_8), .ZN(p_1[8]));
   OAI21_X1 i_17 (.A(n_13), .B1(n_23), .B2(n_54), .ZN(n_8));
   AOI21_X1 i_18 (.A(n_12), .B1(n_75), .B2(n_13), .ZN(p_1[9]));
   AOI21_X1 i_19 (.A(n_10), .B1(n_76), .B2(n_11), .ZN(p_1[10]));
   NOR2_X1 i_20 (.A1(n_52), .A2(n_9), .ZN(p_1[11]));
   NOR2_X1 i_21 (.A1(p_0[11]), .A2(n_10), .ZN(n_9));
   NOR2_X1 i_22 (.A1(n_76), .A2(n_11), .ZN(n_10));
   INV_X1 i_23 (.A(n_12), .ZN(n_11));
   NOR2_X1 i_24 (.A1(n_75), .A2(n_13), .ZN(n_12));
   NAND2_X1 i_25 (.A1(n_23), .A2(n_54), .ZN(n_13));
   INV_X1 i_26 (.A(n_14), .ZN(p_1[12]));
   OAI21_X1 i_27 (.A(n_21), .B1(p_0[12]), .B2(n_52), .ZN(n_14));
   XNOR2_X1 i_32 (.A(p_0[15]), .B(n_17), .ZN(p_1[15]));
   AOI21_X1 i_38 (.A(n_24), .B1(n_77), .B2(n_50), .ZN(p_1[16]));
   XOR2_X1 i_40 (.A(p_0[18]), .B(n_22), .Z(p_1[18]));
   INV_X1 i_44 (.A(n_25), .ZN(p_1[19]));
   OAI21_X1 i_45 (.A(n_31), .B1(p_0[19]), .B2(n_26), .ZN(n_25));
   NOR4_X1 i_46 (.A1(n_79), .A2(n_78), .A3(n_77), .A4(n_50), .ZN(n_26));
   AOI21_X1 i_47 (.A(n_27), .B1(n_80), .B2(n_31), .ZN(p_1[20]));
   XOR2_X1 i_48 (.A(n_116), .B(n_27), .Z(p_1[21]));
   NOR2_X1 i_49 (.A1(n_80), .A2(n_31), .ZN(n_27));
   INV_X1 i_50 (.A(n_28), .ZN(p_1[22]));
   OAI21_X1 i_51 (.A(n_30), .B1(p_0[22]), .B2(n_29), .ZN(n_28));
   NOR3_X1 i_52 (.A1(n_81), .A2(n_80), .A3(n_31), .ZN(n_29));
   AOI21_X1 i_53 (.A(n_37), .B1(n_82), .B2(n_30), .ZN(p_1[23]));
   OR2_X1 i_54 (.A1(n_48), .A2(n_31), .ZN(n_30));
   OR2_X1 i_55 (.A1(n_50), .A2(n_49), .ZN(n_31));
   XNOR2_X1 i_69 (.A(p_0[29]), .B(n_40), .ZN(p_1[29]));
   INV_X1 i_86 (.A(n_55), .ZN(n_54));
   AOI21_X1 i_100 (.A(n_71), .B1(n_70), .B2(n_69), .ZN(n_68));
   NAND2_X1 i_101 (.A1(p_0[1]), .A2(Data_Size[1]), .ZN(n_69));
   NAND2_X1 i_102 (.A1(p_0[0]), .A2(Data_Size[0]), .ZN(n_70));
   NOR2_X1 i_103 (.A1(p_0[1]), .A2(Data_Size[1]), .ZN(n_71));
   INV_X1 i_111 (.A(p_0[18]), .ZN(n_79));
   INV_X1 i_112 (.A(p_0[20]), .ZN(n_80));
   INV_X1 i_113 (.A(n_116), .ZN(n_81));
   NAND3_X1 i_34 (.A1(n_116), .A2(p_0[22]), .A3(p_0[20]), .ZN(n_48));
   INV_X1 i_35 (.A(p_0[23]), .ZN(n_82));
   INV_X1 i_37 (.A(n_16), .ZN(n_52));
   NAND2_X1 i_56 (.A1(p_0[10]), .A2(n_108), .ZN(n_16));
   INV_X1 i_57 (.A(p_0[10]), .ZN(n_76));
   INV_X1 i_63 (.A(p_0[9]), .ZN(n_75));
   INV_X1 i_65 (.A(n_18), .ZN(p_1[14]));
   NAND2_X1 i_67 (.A1(n_32), .A2(n_17), .ZN(n_18));
   NAND2_X1 i_68 (.A1(n_19), .A2(n_39), .ZN(n_32));
   INV_X1 i_74 (.A(n_117), .ZN(n_39));
   NAND3_X1 i_75 (.A1(n_20), .A2(n_117), .A3(p_0[13]), .ZN(n_17));
   INV_X1 i_83 (.A(p_0[24]), .ZN(n_84));
   INV_X1 i_107 (.A(n_86), .ZN(p_1[28]));
   NAND2_X1 i_108 (.A1(n_40), .A2(n_87), .ZN(n_86));
   NAND2_X1 i_114 (.A1(n_96), .A2(n_88), .ZN(n_87));
   INV_X1 i_115 (.A(p_0[28]), .ZN(n_88));
   NAND2_X1 i_116 (.A1(n_44), .A2(p_0[28]), .ZN(n_40));
   NAND2_X1 i_117 (.A1(n_92), .A2(n_89), .ZN(p_1[31]));
   NAND3_X1 i_118 (.A1(n_44), .A2(n_91), .A3(n_90), .ZN(n_89));
   INV_X1 i_119 (.A(n_93), .ZN(n_90));
   INV_X1 i_121 (.A(p_0[31]), .ZN(n_91));
   OAI21_X1 i_122 (.A(p_0[31]), .B1(n_96), .B2(n_93), .ZN(n_92));
   NAND2_X1 i_123 (.A1(p_0[30]), .A2(n_94), .ZN(n_93));
   INV_X1 i_124 (.A(n_95), .ZN(n_94));
   NAND2_X1 i_125 (.A1(p_0[29]), .A2(p_0[28]), .ZN(n_95));
   NAND2_X1 i_130 (.A1(p_0[25]), .A2(p_0[26]), .ZN(n_100));
   NAND2_X1 i_144 (.A1(p_0[15]), .A2(p_0[12]), .ZN(n_112));
   BUF_X1 rt_shieldBuf__2 (.A(p_0[8]), .Z(n_23));
   INV_X1 i_36 (.A(n_111), .ZN(n_22));
   INV_X1 i_41 (.A(n_119), .ZN(n_77));
   INV_X1 i_42 (.A(n_110), .ZN(n_24));
   BUF_X1 rt_shieldBuf__2__2__0 (.A(p_0[16]), .Z(n_119));
   INV_X1 i_28 (.A(n_143), .ZN(n_106));
   NAND4_X1 i_29 (.A1(p_0[19]), .A2(p_0[18]), .A3(p_0[17]), .A4(p_0[16]), 
      .ZN(n_49));
   NAND2_X1 i_30 (.A1(n_15), .A2(n_63), .ZN(n_58));
   OAI21_X1 i_31 (.A(n_60), .B1(p_0[5]), .B2(Data_Size[5]), .ZN(n_15));
   NAND2_X1 i_33 (.A1(n_127), .A2(n_62), .ZN(n_60));
   NOR2_X1 i_39 (.A1(n_33), .A2(n_74), .ZN(n_64));
   INV_X1 i_43 (.A(n_128), .ZN(n_33));
   INV_X1 i_58 (.A(n_129), .ZN(n_73));
   NOR2_X1 i_59 (.A1(p_0[3]), .A2(Data_Size[3]), .ZN(n_74));
   NAND2_X1 i_60 (.A1(n_67), .A2(n_72), .ZN(n_66));
   NAND4_X1 i_61 (.A1(n_113), .A2(p_0[16]), .A3(p_0[11]), .A4(n_34), .ZN(n_110));
   INV_X1 i_62 (.A(n_35), .ZN(n_34));
   NAND4_X1 i_64 (.A1(n_56), .A2(p_0[8]), .A3(p_0[7]), .A4(n_98), .ZN(n_35));
   INV_X1 i_66 (.A(n_57), .ZN(n_56));
   NAND2_X1 i_70 (.A1(n_126), .A2(n_130), .ZN(n_57));
   INV_X1 i_71 (.A(n_114), .ZN(n_113));
   INV_X1 i_72 (.A(p_0[17]), .ZN(n_78));
   NAND2_X1 i_73 (.A1(n_42), .A2(n_36), .ZN(p_1[26]));
   NAND3_X1 i_76 (.A1(n_37), .A2(n_41), .A3(n_38), .ZN(n_36));
   INV_X1 i_77 (.A(n_43), .ZN(n_38));
   INV_X1 i_78 (.A(p_0[26]), .ZN(n_41));
   OAI21_X1 i_79 (.A(p_0[26]), .B1(n_85), .B2(n_43), .ZN(n_42));
   NAND2_X1 i_80 (.A1(p_0[24]), .A2(p_0[25]), .ZN(n_43));
   INV_X1 i_81 (.A(n_45), .ZN(p_1[30]));
   NAND2_X1 i_82 (.A1(n_61), .A2(n_46), .ZN(n_45));
   NAND2_X1 i_84 (.A1(n_90), .A2(n_44), .ZN(n_46));
   INV_X1 i_85 (.A(n_96), .ZN(n_44));
   NAND4_X1 i_87 (.A1(n_139), .A2(n_53), .A3(n_47), .A4(n_104), .ZN(n_96));
   INV_X1 i_88 (.A(n_51), .ZN(n_47));
   NAND2_X1 i_89 (.A1(p_0[18]), .A2(n_157), .ZN(n_51));
   INV_X1 i_90 (.A(n_59), .ZN(n_53));
   NAND2_X1 i_91 (.A1(p_0[19]), .A2(p_0[22]), .ZN(n_59));
   NAND2_X1 i_92 (.A1(n_65), .A2(n_115), .ZN(n_61));
   NAND4_X1 i_93 (.A1(n_101), .A2(n_107), .A3(n_104), .A4(n_139), .ZN(n_65));
   INV_X1 i_94 (.A(n_97), .ZN(n_83));
   NAND2_X1 i_95 (.A1(n_98), .A2(p_0[8]), .ZN(n_97));
   NOR2_X1 i_96 (.A1(n_112), .A2(n_102), .ZN(n_98));
   NAND2_X1 i_97 (.A1(p_0[10]), .A2(p_0[9]), .ZN(n_102));
   OAI21_X1 i_98 (.A(p_0[6]), .B1(p_0[5]), .B2(Data_Size[5]), .ZN(n_103));
   INV_X1 i_99 (.A(n_105), .ZN(n_104));
   NAND3_X1 i_104 (.A1(p_0[24]), .A2(p_0[27]), .A3(n_99), .ZN(n_105));
   INV_X1 i_105 (.A(n_109), .ZN(n_107));
   NAND2_X1 i_106 (.A1(p_0[29]), .A2(p_0[28]), .ZN(n_109));
   INV_X1 i_109 (.A(p_0[30]), .ZN(n_115));
   BUF_X1 rt_shieldBuf__2__2__1 (.A(p_0[21]), .Z(n_116));
   BUF_X1 rt_shieldBuf__2__2__2 (.A(p_0[14]), .Z(n_117));
   INV_X1 i_110 (.A(n_118), .ZN(n_108));
   NAND2_X1 i_120 (.A1(n_123), .A2(n_121), .ZN(n_118));
   NAND2_X1 i_126 (.A1(n_20), .A2(p_0[13]), .ZN(n_19));
   INV_X1 i_127 (.A(n_120), .ZN(p_1[13]));
   XNOR2_X1 i_128 (.A(n_20), .B(p_0[13]), .ZN(n_120));
   INV_X1 i_129 (.A(n_21), .ZN(n_20));
   NAND4_X1 i_131 (.A1(n_123), .A2(p_0[12]), .A3(p_0[10]), .A4(n_121), .ZN(n_21));
   INV_X1 i_132 (.A(n_122), .ZN(n_121));
   NAND2_X1 i_133 (.A1(p_0[9]), .A2(p_0[8]), .ZN(n_122));
   INV_X1 i_134 (.A(n_124), .ZN(n_123));
   NAND2_X1 i_135 (.A1(p_0[11]), .A2(n_125), .ZN(n_124));
   INV_X1 i_136 (.A(n_55), .ZN(n_125));
   NAND3_X1 i_137 (.A1(n_126), .A2(p_0[7]), .A3(n_130), .ZN(n_55));
   NAND3_X1 i_138 (.A1(n_127), .A2(n_62), .A3(n_63), .ZN(n_126));
   NAND2_X1 i_139 (.A1(p_0[5]), .A2(Data_Size[5]), .ZN(n_63));
   NAND2_X1 i_140 (.A1(p_0[4]), .A2(Data_Size[4]), .ZN(n_62));
   OAI221_X1 i_141 (.A(n_128), .B1(p_0[4]), .B2(Data_Size[4]), .C1(p_0[3]), 
      .C2(Data_Size[3]), .ZN(n_127));
   NAND3_X1 i_142 (.A1(n_129), .A2(n_67), .A3(n_72), .ZN(n_128));
   NAND2_X1 i_143 (.A1(p_0[2]), .A2(Data_Size[2]), .ZN(n_72));
   OAI21_X1 i_145 (.A(n_68), .B1(p_0[2]), .B2(Data_Size[2]), .ZN(n_67));
   NAND2_X1 i_146 (.A1(p_0[3]), .A2(Data_Size[3]), .ZN(n_129));
   INV_X1 i_147 (.A(n_103), .ZN(n_130));
   NAND2_X1 i_148 (.A1(n_133), .A2(n_131), .ZN(p_1[27]));
   NAND4_X1 i_149 (.A1(n_135), .A2(n_101), .A3(n_132), .A4(n_136), .ZN(n_131));
   INV_X1 i_150 (.A(p_0[27]), .ZN(n_132));
   NAND2_X1 i_151 (.A1(n_134), .A2(p_0[27]), .ZN(n_133));
   NAND3_X1 i_152 (.A1(n_135), .A2(n_136), .A3(n_101), .ZN(n_134));
   INV_X1 i_153 (.A(n_50), .ZN(n_135));
   NAND2_X1 i_154 (.A1(n_113), .A2(n_106), .ZN(n_50));
   INV_X1 i_155 (.A(n_137), .ZN(n_136));
   NAND2_X1 i_156 (.A1(p_0[24]), .A2(n_99), .ZN(n_137));
   INV_X1 i_157 (.A(n_100), .ZN(n_99));
   INV_X1 i_158 (.A(n_138), .ZN(n_101));
   NAND3_X1 i_159 (.A1(n_165), .A2(p_0[18]), .A3(n_157), .ZN(n_138));
   INV_X1 i_160 (.A(n_140), .ZN(n_139));
   NAND2_X1 i_161 (.A1(n_142), .A2(n_144), .ZN(n_140));
   INV_X1 i_162 (.A(n_85), .ZN(n_37));
   NAND2_X1 i_163 (.A1(n_149), .A2(n_153), .ZN(n_85));
   AOI21_X1 i_164 (.A(n_141), .B1(n_110), .B2(n_78), .ZN(p_1[17]));
   INV_X1 i_165 (.A(n_111), .ZN(n_141));
   NAND4_X1 i_166 (.A1(n_142), .A2(n_144), .A3(p_0[17]), .A4(n_119), .ZN(n_111));
   INV_X1 i_167 (.A(n_143), .ZN(n_142));
   NAND2_X1 i_168 (.A1(n_123), .A2(n_83), .ZN(n_143));
   INV_X1 i_169 (.A(n_114), .ZN(n_144));
   NAND2_X1 i_170 (.A1(p_0[13]), .A2(p_0[14]), .ZN(n_114));
   NOR2_X1 i_171 (.A1(n_145), .A2(n_151), .ZN(p_1[24]));
   AOI21_X1 i_172 (.A(n_146), .B1(n_149), .B2(n_153), .ZN(n_145));
   INV_X1 i_173 (.A(n_84), .ZN(n_146));
   INV_X1 i_174 (.A(n_147), .ZN(p_1[25]));
   OAI21_X1 i_175 (.A(n_148), .B1(n_151), .B2(p_0[25]), .ZN(n_147));
   NAND3_X1 i_176 (.A1(n_149), .A2(n_38), .A3(n_153), .ZN(n_148));
   INV_X1 i_177 (.A(n_150), .ZN(n_149));
   NAND3_X1 i_178 (.A1(n_163), .A2(p_0[22]), .A3(p_0[19]), .ZN(n_150));
   INV_X1 i_179 (.A(n_152), .ZN(n_151));
   NAND4_X1 i_180 (.A1(n_165), .A2(n_153), .A3(p_0[24]), .A4(n_163), .ZN(n_152));
   INV_X1 i_181 (.A(n_154), .ZN(n_153));
   NAND3_X1 i_182 (.A1(n_157), .A2(n_123), .A3(n_155), .ZN(n_154));
   INV_X1 i_183 (.A(n_156), .ZN(n_155));
   NAND2_X1 i_184 (.A1(p_0[14]), .A2(n_83), .ZN(n_156));
   INV_X1 i_185 (.A(n_158), .ZN(n_157));
   NAND3_X1 i_186 (.A1(n_161), .A2(p_0[23]), .A3(n_159), .ZN(n_158));
   INV_X1 i_187 (.A(n_160), .ZN(n_159));
   NAND2_X1 i_188 (.A1(p_0[20]), .A2(p_0[17]), .ZN(n_160));
   INV_X1 i_189 (.A(n_162), .ZN(n_161));
   NAND2_X1 i_190 (.A1(p_0[21]), .A2(p_0[16]), .ZN(n_162));
   INV_X1 i_191 (.A(n_164), .ZN(n_163));
   NAND2_X1 i_192 (.A1(p_0[18]), .A2(p_0[13]), .ZN(n_164));
   INV_X1 i_193 (.A(n_166), .ZN(n_165));
   NAND2_X1 i_194 (.A1(p_0[19]), .A2(p_0[22]), .ZN(n_166));
endmodule

module datapath__0_197(Data_Size, p_0);
   input [31:0]Data_Size;
   output [31:0]p_0;

   XNOR2_X1 i_1 (.A(Data_Size[7]), .B(Data_Size[6]), .ZN(p_0[7]));
   OR2_X1 i_2 (.A1(Data_Size[7]), .A2(Data_Size[6]), .ZN(n_0));
   XNOR2_X1 i_3 (.A(Data_Size[8]), .B(n_0), .ZN(p_0[8]));
   OR2_X1 i_4 (.A1(Data_Size[8]), .A2(n_0), .ZN(n_1));
   XNOR2_X1 i_5 (.A(Data_Size[9]), .B(n_1), .ZN(p_0[9]));
   OR2_X1 i_6 (.A1(Data_Size[9]), .A2(n_1), .ZN(n_2));
   XNOR2_X1 i_7 (.A(Data_Size[10]), .B(n_2), .ZN(p_0[10]));
   OR2_X1 i_8 (.A1(Data_Size[10]), .A2(n_2), .ZN(n_3));
   XNOR2_X1 i_9 (.A(Data_Size[11]), .B(n_3), .ZN(p_0[11]));
   OR2_X1 i_10 (.A1(Data_Size[11]), .A2(n_3), .ZN(n_4));
   XNOR2_X1 i_11 (.A(Data_Size[12]), .B(n_4), .ZN(p_0[12]));
   OR2_X1 i_12 (.A1(Data_Size[12]), .A2(n_4), .ZN(n_5));
   XNOR2_X1 i_13 (.A(Data_Size[13]), .B(n_5), .ZN(p_0[13]));
   OR2_X1 i_14 (.A1(Data_Size[13]), .A2(n_5), .ZN(n_6));
   XNOR2_X1 i_15 (.A(Data_Size[14]), .B(n_6), .ZN(p_0[14]));
   OR2_X1 i_16 (.A1(Data_Size[14]), .A2(n_6), .ZN(n_7));
   XNOR2_X1 i_17 (.A(Data_Size[15]), .B(n_7), .ZN(p_0[15]));
   OR2_X1 i_18 (.A1(Data_Size[15]), .A2(n_7), .ZN(n_8));
   XNOR2_X1 i_19 (.A(Data_Size[16]), .B(n_8), .ZN(p_0[16]));
   OR2_X1 i_20 (.A1(Data_Size[16]), .A2(n_8), .ZN(n_9));
   XNOR2_X1 i_21 (.A(Data_Size[17]), .B(n_9), .ZN(p_0[17]));
   OR2_X1 i_22 (.A1(Data_Size[17]), .A2(n_9), .ZN(n_10));
   XNOR2_X1 i_23 (.A(Data_Size[18]), .B(n_10), .ZN(p_0[18]));
   OR2_X1 i_24 (.A1(Data_Size[18]), .A2(n_10), .ZN(n_11));
   XNOR2_X1 i_25 (.A(Data_Size[19]), .B(n_11), .ZN(p_0[19]));
   OR2_X1 i_26 (.A1(Data_Size[19]), .A2(n_11), .ZN(n_12));
   XNOR2_X1 i_27 (.A(Data_Size[20]), .B(n_12), .ZN(p_0[20]));
   OR2_X1 i_28 (.A1(Data_Size[20]), .A2(n_12), .ZN(n_13));
   XNOR2_X1 i_29 (.A(Data_Size[21]), .B(n_13), .ZN(p_0[21]));
   OR2_X1 i_30 (.A1(Data_Size[21]), .A2(n_13), .ZN(n_14));
   XNOR2_X1 i_31 (.A(Data_Size[22]), .B(n_14), .ZN(p_0[22]));
   OR2_X1 i_32 (.A1(Data_Size[22]), .A2(n_14), .ZN(n_15));
   XNOR2_X1 i_33 (.A(Data_Size[23]), .B(n_15), .ZN(p_0[23]));
   OR2_X1 i_34 (.A1(Data_Size[23]), .A2(n_15), .ZN(n_16));
   XNOR2_X1 i_35 (.A(Data_Size[24]), .B(n_16), .ZN(p_0[24]));
   OR2_X1 i_36 (.A1(Data_Size[24]), .A2(n_16), .ZN(n_17));
   XNOR2_X1 i_37 (.A(Data_Size[25]), .B(n_17), .ZN(p_0[25]));
   OR2_X1 i_38 (.A1(Data_Size[25]), .A2(n_17), .ZN(n_18));
   XNOR2_X1 i_39 (.A(Data_Size[26]), .B(n_18), .ZN(p_0[26]));
   OR2_X1 i_40 (.A1(Data_Size[26]), .A2(n_18), .ZN(n_19));
   XNOR2_X1 i_41 (.A(Data_Size[27]), .B(n_19), .ZN(p_0[27]));
   OR2_X1 i_42 (.A1(Data_Size[27]), .A2(n_19), .ZN(n_20));
   XNOR2_X1 i_43 (.A(Data_Size[28]), .B(n_20), .ZN(p_0[28]));
   OR2_X1 i_44 (.A1(Data_Size[28]), .A2(n_20), .ZN(n_21));
   XNOR2_X1 i_45 (.A(Data_Size[29]), .B(n_21), .ZN(p_0[29]));
   OR2_X1 i_46 (.A1(Data_Size[29]), .A2(n_21), .ZN(n_22));
   XNOR2_X1 i_47 (.A(Data_Size[30]), .B(n_22), .ZN(p_0[30]));
   OR2_X1 i_48 (.A1(Data_Size[30]), .A2(n_22), .ZN(n_23));
   XNOR2_X1 i_49 (.A(Data_Size[31]), .B(n_23), .ZN(p_0[31]));
endmodule

module datapath__0_393(p_0, p_1, RowsCount);
   output p_0;
   input [37:0]p_1;
   input [15:0]RowsCount;

   INV_X1 i_4 (.A(p_1[9]), .ZN(n_4));
   NAND2_X1 i_5 (.A1(n_4), .A2(RowsCount[9]), .ZN(n_5));
   INV_X1 i_11 (.A(n_5), .ZN(n_11));
   INV_X1 i_22 (.A(p_1[1]), .ZN(n_22));
   INV_X1 i_23 (.A(p_1[2]), .ZN(n_23));
   AOI22_X1 i_24 (.A1(n_22), .A2(RowsCount[1]), .B1(n_23), .B2(RowsCount[2]), 
      .ZN(n_24));
   INV_X1 i_25 (.A(RowsCount[3]), .ZN(n_25));
   INV_X1 i_26 (.A(RowsCount[2]), .ZN(n_26));
   AOI221_X1 i_27 (.A(n_24), .B1(p_1[3]), .B2(n_25), .C1(p_1[2]), .C2(n_26), 
      .ZN(n_27));
   INV_X1 i_28 (.A(RowsCount[4]), .ZN(n_28));
   OAI22_X1 i_29 (.A1(n_25), .A2(p_1[3]), .B1(n_28), .B2(p_1[4]), .ZN(n_29));
   INV_X1 i_30 (.A(p_1[4]), .ZN(n_30));
   INV_X1 i_31 (.A(p_1[5]), .ZN(n_31));
   INV_X1 i_38 (.A(RowsCount[12]), .ZN(n_38));
   NAND2_X1 i_39 (.A1(n_38), .A2(p_1[12]), .ZN(n_39));
   OAI21_X1 i_40 (.A(n_39), .B1(n_38), .B2(p_1[12]), .ZN(n_40));
   INV_X1 i_41 (.A(RowsCount[11]), .ZN(n_41));
   NAND2_X1 i_42 (.A1(n_41), .A2(p_1[11]), .ZN(n_42));
   OAI21_X1 i_44 (.A(n_42), .B1(n_41), .B2(p_1[11]), .ZN(n_44));
   NOR3_X1 i_47 (.A1(n_39), .A2(RowsCount[13]), .A3(RowsCount[14]), .ZN(n_47));
   OAI22_X1 i_48 (.A1(n_40), .A2(n_42), .B1(n_44), .B2(n_1), .ZN(n_48));
   OAI21_X1 i_0 (.A(n_73), .B1(n_6), .B2(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(n_3), .B1(n_2), .B2(n_12), .ZN(n_0));
   INV_X1 i_2 (.A(n_48), .ZN(n_2));
   INV_X1 i_3 (.A(n_47), .ZN(n_3));
   INV_X1 i_6 (.A(n_7), .ZN(n_6));
   NAND2_X1 i_7 (.A1(n_17), .A2(n_8), .ZN(n_7));
   INV_X1 i_8 (.A(n_9), .ZN(n_8));
   NAND2_X1 i_9 (.A1(n_16), .A2(n_10), .ZN(n_9));
   INV_X1 i_10 (.A(n_12), .ZN(n_10));
   OAI21_X1 i_12 (.A(n_13), .B1(n_14), .B2(n_15), .ZN(n_12));
   AOI21_X1 i_13 (.A(RowsCount[14]), .B1(n_39), .B2(RowsCount[13]), .ZN(n_13));
   INV_X1 i_14 (.A(n_42), .ZN(n_14));
   INV_X1 i_15 (.A(n_40), .ZN(n_15));
   NAND2_X1 i_16 (.A1(n_44), .A2(n_1), .ZN(n_16));
   NAND3_X1 i_17 (.A1(n_20), .A2(n_49), .A3(n_18), .ZN(n_17));
   NAND4_X1 i_18 (.A1(n_19), .A2(n_5), .A3(n_1), .A4(n_66), .ZN(n_18));
   OAI21_X1 i_19 (.A(n_71), .B1(RowsCount[9]), .B2(n_4), .ZN(n_19));
   NAND4_X1 i_20 (.A1(n_21), .A2(n_59), .A3(n_43), .A4(n_69), .ZN(n_20));
   INV_X1 i_21 (.A(n_32), .ZN(n_21));
   NAND4_X1 i_32 (.A1(n_33), .A2(n_63), .A3(n_54), .A4(n_36), .ZN(n_32));
   AOI21_X1 i_33 (.A(n_34), .B1(p_1[6]), .B2(n_58), .ZN(n_33));
   INV_X1 i_34 (.A(n_35), .ZN(n_34));
   NAND2_X1 i_35 (.A1(n_31), .A2(RowsCount[5]), .ZN(n_35));
   NAND2_X1 i_36 (.A1(n_37), .A2(RowsCount[6]), .ZN(n_36));
   INV_X1 i_37 (.A(p_1[6]), .ZN(n_37));
   OAI21_X1 i_43 (.A(n_45), .B1(n_29), .B2(n_27), .ZN(n_43));
   INV_X1 i_45 (.A(n_46), .ZN(n_45));
   OAI22_X1 i_46 (.A1(n_30), .A2(RowsCount[4]), .B1(RowsCount[5]), .B2(n_31), 
      .ZN(n_46));
   NAND3_X1 i_49 (.A1(n_59), .A2(n_50), .A3(n_69), .ZN(n_49));
   NAND2_X1 i_50 (.A1(n_53), .A2(n_51), .ZN(n_50));
   NAND3_X1 i_51 (.A1(n_52), .A2(n_71), .A3(n_61), .ZN(n_51));
   INV_X1 i_52 (.A(n_63), .ZN(n_52));
   NAND3_X1 i_53 (.A1(n_56), .A2(n_54), .A3(n_63), .ZN(n_53));
   NAND2_X1 i_54 (.A1(n_55), .A2(RowsCount[7]), .ZN(n_54));
   INV_X1 i_55 (.A(p_1[7]), .ZN(n_55));
   INV_X1 i_56 (.A(n_57), .ZN(n_56));
   NAND2_X1 i_57 (.A1(p_1[6]), .A2(n_58), .ZN(n_57));
   INV_X1 i_58 (.A(RowsCount[6]), .ZN(n_58));
   AOI21_X1 i_59 (.A(n_65), .B1(n_60), .B2(n_63), .ZN(n_59));
   NAND2_X1 i_60 (.A1(n_61), .A2(n_71), .ZN(n_60));
   NAND2_X1 i_61 (.A1(n_62), .A2(RowsCount[8]), .ZN(n_61));
   INV_X1 i_62 (.A(p_1[8]), .ZN(n_62));
   NAND2_X1 i_63 (.A1(p_1[7]), .A2(n_64), .ZN(n_63));
   INV_X1 i_64 (.A(RowsCount[7]), .ZN(n_64));
   AOI21_X1 i_65 (.A(n_70), .B1(n_66), .B2(n_1), .ZN(n_65));
   NAND2_X1 i_66 (.A1(n_67), .A2(RowsCount[10]), .ZN(n_66));
   INV_X1 i_67 (.A(p_1[10]), .ZN(n_67));
   NAND2_X1 i_68 (.A1(p_1[10]), .A2(n_68), .ZN(n_1));
   INV_X1 i_69 (.A(RowsCount[10]), .ZN(n_68));
   OAI21_X1 i_70 (.A(n_71), .B1(n_11), .B2(n_70), .ZN(n_69));
   NOR2_X1 i_71 (.A1(n_4), .A2(RowsCount[9]), .ZN(n_70));
   NAND2_X1 i_72 (.A1(p_1[8]), .A2(n_72), .ZN(n_71));
   INV_X1 i_73 (.A(RowsCount[8]), .ZN(n_72));
   INV_X1 i_74 (.A(RowsCount[15]), .ZN(n_73));
endmodule

module datapath(PacketSize, p_0);
   input [5:0]PacketSize;
   output [31:0]p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0[1]));
   AOI21_X1 i_1 (.A(n_11), .B1(PacketSize[1]), .B2(PacketSize[0]), .ZN(n_0));
   NAND2_X1 i_2 (.A1(n_1), .A2(n_14), .ZN(p_0[3]));
   NAND2_X1 i_3 (.A1(n_7), .A2(PacketSize[3]), .ZN(n_1));
   NAND2_X1 i_4 (.A1(n_2), .A2(n_3), .ZN(p_0[5]));
   OAI21_X1 i_5 (.A(PacketSize[5]), .B1(n_14), .B2(PacketSize[4]), .ZN(n_2));
   INV_X1 i_6 (.A(n_3), .ZN(p_0[31]));
   NAND3_X1 i_7 (.A1(n_5), .A2(n_4), .A3(n_12), .ZN(n_3));
   INV_X1 i_8 (.A(PacketSize[5]), .ZN(n_4));
   INV_X1 i_9 (.A(n_14), .ZN(n_5));
   NAND2_X1 i_10 (.A1(n_7), .A2(n_6), .ZN(p_0[2]));
   OAI21_X1 i_11 (.A(PacketSize[2]), .B1(PacketSize[0]), .B2(PacketSize[1]), 
      .ZN(n_6));
   NAND2_X1 i_12 (.A1(n_11), .A2(n_17), .ZN(n_7));
   NAND2_X1 i_13 (.A1(n_13), .A2(n_8), .ZN(p_0[4]));
   NAND3_X1 i_14 (.A1(n_11), .A2(n_9), .A3(n_12), .ZN(n_8));
   INV_X1 i_15 (.A(n_10), .ZN(n_9));
   NAND2_X1 i_16 (.A1(n_17), .A2(n_18), .ZN(n_10));
   NOR2_X1 i_17 (.A1(PacketSize[0]), .A2(PacketSize[1]), .ZN(n_11));
   INV_X1 i_18 (.A(PacketSize[4]), .ZN(n_12));
   NAND2_X1 i_19 (.A1(n_14), .A2(PacketSize[4]), .ZN(n_13));
   NAND4_X1 i_20 (.A1(n_15), .A2(n_17), .A3(n_18), .A4(n_16), .ZN(n_14));
   INV_X1 i_21 (.A(PacketSize[0]), .ZN(n_15));
   INV_X1 i_22 (.A(PacketSize[1]), .ZN(n_16));
   INV_X1 i_23 (.A(PacketSize[2]), .ZN(n_17));
   INV_X1 i_24 (.A(PacketSize[3]), .ZN(n_18));
endmodule

module datapath__2_420(p_0, Small_Packet_Indication_Bit_Location, p_1);
   input [31:0]p_0;
   input [5:0]Small_Packet_Indication_Bit_Location;
   output p_1;

   INV_X1 i_0 (.A(n_0), .ZN(p_1));
   NAND4_X1 i_1 (.A1(n_11), .A2(n_18), .A3(n_6), .A4(n_1), .ZN(n_0));
   NAND2_X1 i_2 (.A1(n_3), .A2(n_2), .ZN(n_1));
   NAND2_X1 i_3 (.A1(p_0[1]), .A2(Small_Packet_Indication_Bit_Location[1]), 
      .ZN(n_2));
   NAND2_X1 i_4 (.A1(n_5), .A2(n_4), .ZN(n_3));
   INV_X1 i_5 (.A(Small_Packet_Indication_Bit_Location[1]), .ZN(n_4));
   INV_X1 i_6 (.A(p_0[1]), .ZN(n_5));
   NAND2_X1 i_7 (.A1(n_8), .A2(n_7), .ZN(n_6));
   NAND2_X1 i_8 (.A1(p_0[5]), .A2(Small_Packet_Indication_Bit_Location[5]), 
      .ZN(n_7));
   NAND2_X1 i_9 (.A1(n_10), .A2(n_9), .ZN(n_8));
   INV_X1 i_10 (.A(Small_Packet_Indication_Bit_Location[5]), .ZN(n_9));
   INV_X1 i_11 (.A(p_0[5]), .ZN(n_10));
   NOR2_X1 i_12 (.A1(n_12), .A2(n_15), .ZN(n_11));
   OAI21_X1 i_13 (.A(n_13), .B1(p_0[3]), .B2(n_21), .ZN(n_12));
   NAND2_X1 i_14 (.A1(n_14), .A2(Small_Packet_Indication_Bit_Location[2]), 
      .ZN(n_13));
   INV_X1 i_15 (.A(p_0[2]), .ZN(n_14));
   OAI21_X1 i_16 (.A(n_16), .B1(p_0[4]), .B2(n_25), .ZN(n_15));
   NOR2_X1 i_17 (.A1(p_0[6]), .A2(n_17), .ZN(n_16));
   XOR2_X1 i_18 (.A(Small_Packet_Indication_Bit_Location[0]), .B(p_0[0]), 
      .Z(n_17));
   INV_X1 i_19 (.A(n_19), .ZN(n_18));
   NAND3_X1 i_20 (.A1(n_24), .A2(n_20), .A3(n_22), .ZN(n_19));
   NAND2_X1 i_21 (.A1(p_0[3]), .A2(n_21), .ZN(n_20));
   INV_X1 i_22 (.A(Small_Packet_Indication_Bit_Location[3]), .ZN(n_21));
   NAND2_X1 i_23 (.A1(p_0[2]), .A2(n_23), .ZN(n_22));
   INV_X1 i_24 (.A(Small_Packet_Indication_Bit_Location[2]), .ZN(n_23));
   NAND2_X1 i_25 (.A1(p_0[4]), .A2(n_25), .ZN(n_24));
   INV_X1 i_26 (.A(Small_Packet_Indication_Bit_Location[4]), .ZN(n_25));
endmodule

module datapath__2_568(p_0, p_1);
   input [11:0]p_0;
   output [12:0]p_1;

   INV_X1 i_0 (.A(p_0[0]), .ZN(p_1[0]));
   NAND2_X1 i_1 (.A1(p_0[1]), .A2(p_0[0]), .ZN(n_0));
   INV_X1 i_2 (.A(n_0), .ZN(n_1));
   NAND3_X1 i_3 (.A1(p_0[2]), .A2(p_0[0]), .A3(p_0[1]), .ZN(n_2));
   INV_X1 i_4 (.A(p_0[2]), .ZN(n_3));
   NAND2_X1 i_5 (.A1(p_0[0]), .A2(p_0[1]), .ZN(n_4));
   NOR2_X1 i_6 (.A1(n_3), .A2(n_4), .ZN(n_5));
   NAND2_X1 i_7 (.A1(p_0[3]), .A2(n_5), .ZN(n_6));
   NAND2_X1 i_8 (.A1(n_34), .A2(p_0[4]), .ZN(n_7));
   INV_X1 i_9 (.A(n_7), .ZN(n_8));
   NAND2_X1 i_10 (.A1(p_0[5]), .A2(p_0[4]), .ZN(n_9));
   INV_X1 i_11 (.A(n_9), .ZN(n_10));
   NAND2_X1 i_12 (.A1(n_10), .A2(n_34), .ZN(n_11));
   INV_X1 i_13 (.A(n_11), .ZN(n_12));
   NAND3_X1 i_14 (.A1(p_0[5]), .A2(p_0[6]), .A3(p_0[4]), .ZN(n_13));
   NOR2_X1 i_15 (.A1(n_6), .A2(n_13), .ZN(n_14));
   NAND4_X1 i_16 (.A1(p_0[7]), .A2(p_0[5]), .A3(p_0[6]), .A4(p_0[4]), .ZN(n_15));
   INV_X1 i_17 (.A(n_15), .ZN(n_16));
   NAND2_X1 i_18 (.A1(n_36), .A2(p_0[8]), .ZN(n_17));
   INV_X1 i_19 (.A(n_17), .ZN(n_18));
   NAND2_X1 i_20 (.A1(p_0[8]), .A2(p_0[9]), .ZN(n_19));
   INV_X1 i_21 (.A(n_19), .ZN(n_20));
   NAND2_X1 i_22 (.A1(n_36), .A2(n_20), .ZN(n_21));
   INV_X1 i_23 (.A(n_21), .ZN(n_22));
   NAND2_X1 i_24 (.A1(p_0[10]), .A2(p_0[9]), .ZN(n_23));
   INV_X1 i_25 (.A(n_23), .ZN(n_24));
   NAND2_X1 i_26 (.A1(p_0[8]), .A2(n_24), .ZN(n_25));
   INV_X1 i_27 (.A(n_25), .ZN(n_26));
   NAND2_X1 i_28 (.A1(n_36), .A2(n_26), .ZN(n_27));
   INV_X1 i_29 (.A(n_27), .ZN(n_28));
   INV_X1 i_30 (.A(p_0[10]), .ZN(n_29));
   NAND2_X1 i_31 (.A1(p_0[9]), .A2(p_0[11]), .ZN(n_30));
   NOR2_X1 i_32 (.A1(n_29), .A2(n_30), .ZN(n_31));
   NAND2_X1 i_33 (.A1(p_0[8]), .A2(n_31), .ZN(n_32));
   INV_X1 i_34 (.A(n_32), .ZN(n_33));
   INV_X1 i_35 (.A(n_6), .ZN(n_34));
   NAND2_X1 i_36 (.A1(n_16), .A2(n_34), .ZN(n_35));
   INV_X1 i_37 (.A(n_35), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_36), .A2(n_33), .ZN(n_37));
   INV_X1 i_39 (.A(n_37), .ZN(p_1[12]));
   INV_X1 i_40 (.A(p_0[1]), .ZN(n_38));
   XNOR2_X1 i_41 (.A(p_0[0]), .B(n_38), .ZN(p_1[1]));
   XNOR2_X1 i_42 (.A(n_1), .B(n_3), .ZN(p_1[2]));
   XNOR2_X1 i_43 (.A(p_0[3]), .B(n_2), .ZN(p_1[3]));
   INV_X1 i_44 (.A(p_0[4]), .ZN(n_39));
   XNOR2_X1 i_45 (.A(n_34), .B(n_39), .ZN(p_1[4]));
   INV_X1 i_46 (.A(p_0[5]), .ZN(n_40));
   XNOR2_X1 i_47 (.A(n_8), .B(n_40), .ZN(p_1[5]));
   INV_X1 i_48 (.A(p_0[6]), .ZN(n_41));
   XNOR2_X1 i_49 (.A(n_12), .B(n_41), .ZN(p_1[6]));
   INV_X1 i_50 (.A(p_0[7]), .ZN(n_42));
   XNOR2_X1 i_51 (.A(n_14), .B(n_42), .ZN(p_1[7]));
   INV_X1 i_52 (.A(p_0[8]), .ZN(n_43));
   XNOR2_X1 i_53 (.A(n_36), .B(n_43), .ZN(p_1[8]));
   INV_X1 i_54 (.A(p_0[9]), .ZN(n_44));
   XNOR2_X1 i_55 (.A(n_18), .B(n_44), .ZN(p_1[9]));
   XNOR2_X1 i_56 (.A(n_22), .B(n_29), .ZN(p_1[10]));
   INV_X1 i_57 (.A(p_0[11]), .ZN(n_45));
   XNOR2_X1 i_58 (.A(n_28), .B(n_45), .ZN(p_1[11]));
endmodule

module datapath__2_569(p_0, RowsCount, p_1);
   input [12:0]p_0;
   input [15:0]RowsCount;
   output p_1;

   NOR3_X1 i_0 (.A1(RowsCount[14]), .A2(RowsCount[13]), .A3(RowsCount[15]), 
      .ZN(n_0));
   XNOR2_X1 i_1 (.A(p_0[9]), .B(RowsCount[9]), .ZN(n_1));
   XNOR2_X1 i_2 (.A(p_0[10]), .B(RowsCount[10]), .ZN(n_2));
   XNOR2_X1 i_3 (.A(p_0[12]), .B(RowsCount[12]), .ZN(n_3));
   XNOR2_X1 i_4 (.A(p_0[0]), .B(RowsCount[0]), .ZN(n_4));
   XNOR2_X1 i_5 (.A(p_0[1]), .B(RowsCount[1]), .ZN(n_5));
   XNOR2_X1 i_6 (.A(p_0[5]), .B(RowsCount[5]), .ZN(n_6));
   XNOR2_X1 i_7 (.A(p_0[4]), .B(RowsCount[4]), .ZN(n_7));
   INV_X1 i_8 (.A(n_8), .ZN(p_1));
   NAND4_X1 i_9 (.A1(n_30), .A2(n_24), .A3(n_36), .A4(n_9), .ZN(n_8));
   INV_X1 i_10 (.A(n_10), .ZN(n_9));
   NAND2_X1 i_11 (.A1(n_11), .A2(n_3), .ZN(n_10));
   NOR2_X1 i_12 (.A1(n_22), .A2(n_12), .ZN(n_11));
   NAND3_X1 i_13 (.A1(n_13), .A2(n_6), .A3(n_7), .ZN(n_12));
   INV_X1 i_14 (.A(n_14), .ZN(n_13));
   NAND4_X1 i_15 (.A1(n_20), .A2(n_19), .A3(n_17), .A4(n_15), .ZN(n_14));
   INV_X1 i_16 (.A(n_16), .ZN(n_15));
   NAND3_X1 i_17 (.A1(n_5), .A2(n_0), .A3(n_4), .ZN(n_16));
   INV_X1 i_18 (.A(n_18), .ZN(n_17));
   XOR2_X1 i_19 (.A(RowsCount[2]), .B(p_0[2]), .Z(n_18));
   NAND2_X1 i_20 (.A1(n_21), .A2(RowsCount[3]), .ZN(n_19));
   OR2_X1 i_21 (.A1(n_21), .A2(RowsCount[3]), .ZN(n_20));
   INV_X1 i_22 (.A(p_0[3]), .ZN(n_21));
   XNOR2_X1 i_23 (.A(p_0[6]), .B(n_23), .ZN(n_22));
   INV_X1 i_24 (.A(RowsCount[6]), .ZN(n_23));
   INV_X1 i_25 (.A(n_25), .ZN(n_24));
   NAND2_X1 i_26 (.A1(n_26), .A2(n_28), .ZN(n_25));
   NAND2_X1 i_27 (.A1(n_27), .A2(RowsCount[11]), .ZN(n_26));
   INV_X1 i_28 (.A(p_0[11]), .ZN(n_27));
   NAND2_X1 i_29 (.A1(p_0[11]), .A2(n_29), .ZN(n_28));
   INV_X1 i_30 (.A(RowsCount[11]), .ZN(n_29));
   INV_X1 i_31 (.A(n_31), .ZN(n_30));
   NAND4_X1 i_32 (.A1(n_2), .A2(n_1), .A3(n_34), .A4(n_32), .ZN(n_31));
   NAND2_X1 i_33 (.A1(n_33), .A2(RowsCount[8]), .ZN(n_32));
   INV_X1 i_34 (.A(p_0[8]), .ZN(n_33));
   NAND2_X1 i_35 (.A1(p_0[8]), .A2(n_35), .ZN(n_34));
   INV_X1 i_36 (.A(RowsCount[8]), .ZN(n_35));
   INV_X1 i_37 (.A(n_37), .ZN(n_36));
   NAND2_X1 i_38 (.A1(n_38), .A2(n_40), .ZN(n_37));
   NAND2_X1 i_39 (.A1(n_39), .A2(RowsCount[7]), .ZN(n_38));
   INV_X1 i_40 (.A(p_0[7]), .ZN(n_39));
   NAND2_X1 i_41 (.A1(p_0[7]), .A2(n_41), .ZN(n_40));
   INV_X1 i_42 (.A(RowsCount[7]), .ZN(n_41));
endmodule

module TFlipFlop__4_17(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   AOI211_X1 i_0_0 (.A(n_0_0), .B(RST), .C1(Q), .C2(T), .ZN(n_0));
   NOR2_X1 i_0_1 (.A1(Q), .A2(T), .ZN(n_0_0));
endmodule

module TFlipFlop__4_22(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_27(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_32(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_37(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_42(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_47(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_52(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_57(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_62(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_67(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_72(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_77(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_82(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop__4_87(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module TFlipFlop(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module Counter__parameterized0(value, Enable, CLK, RST);
   output [15:0]value;
   input Enable;
   input CLK;
   input RST;

   wire inputs;

   TFlipFlop__4_17 firstBit (.T(Enable), .CLK(CLK), .RST(RST), .Enable(), 
      .Q(value[0]));
   TFlipFlop__4_22 genblk1_1_counterBits (.T(inputs), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[1]));
   TFlipFlop__4_27 genblk1_2_counterBits (.T(n_0), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[2]));
   TFlipFlop__4_32 genblk1_3_counterBits (.T(n_1), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[3]));
   TFlipFlop__4_37 genblk1_4_counterBits (.T(n_2), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[4]));
   TFlipFlop__4_42 genblk1_5_counterBits (.T(n_3), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[5]));
   TFlipFlop__4_47 genblk1_6_counterBits (.T(n_4), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[6]));
   TFlipFlop__4_52 genblk1_7_counterBits (.T(n_5), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[7]));
   TFlipFlop__4_57 genblk1_8_counterBits (.T(n_6), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[8]));
   TFlipFlop__4_62 genblk1_9_counterBits (.T(n_7), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[9]));
   TFlipFlop__4_67 genblk1_10_counterBits (.T(n_8), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[10]));
   TFlipFlop__4_72 genblk1_11_counterBits (.T(n_9), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[11]));
   TFlipFlop__4_77 genblk1_12_counterBits (.T(n_10), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[12]));
   TFlipFlop__4_82 genblk1_13_counterBits (.T(n_11), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[13]));
   TFlipFlop__4_87 genblk1_14_counterBits (.T(n_12), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[14]));
   TFlipFlop genblk1_15_counterBits (.T(n_13), .CLK(CLK), .RST(RST), .Enable(
      Enable), .Q(value[15]));
   AND2_X1 i_0_0 (.A1(Enable), .A2(value[0]), .ZN(inputs));
   AND2_X1 i_0_1 (.A1(inputs), .A2(value[1]), .ZN(n_0));
   AND2_X1 i_0_2 (.A1(n_0), .A2(value[2]), .ZN(n_1));
   AND2_X1 i_0_3 (.A1(n_1), .A2(value[3]), .ZN(n_2));
   AND2_X1 i_0_4 (.A1(n_2), .A2(value[4]), .ZN(n_3));
   AND2_X1 i_0_5 (.A1(n_3), .A2(value[5]), .ZN(n_4));
   AND2_X1 i_0_6 (.A1(n_4), .A2(value[6]), .ZN(n_5));
   AND2_X1 i_0_7 (.A1(n_5), .A2(value[7]), .ZN(n_6));
   AND2_X1 i_0_8 (.A1(n_6), .A2(value[8]), .ZN(n_7));
   AND2_X1 i_0_9 (.A1(n_7), .A2(value[9]), .ZN(n_8));
   AND2_X1 i_0_10 (.A1(n_8), .A2(value[10]), .ZN(n_9));
   AND2_X1 i_0_11 (.A1(n_9), .A2(value[11]), .ZN(n_10));
   AND2_X1 i_0_12 (.A1(n_10), .A2(value[12]), .ZN(n_11));
   AND2_X1 i_0_13 (.A1(n_11), .A2(value[13]), .ZN(n_12));
   AND2_X1 i_0_14 (.A1(n_12), .A2(value[14]), .ZN(n_13));
endmodule

module DFlipFlop__4_2(D, CLK, RST, Enable, Q);
   input D;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   AOI211_X1 i_0_0 (.A(RST), .B(n_0_0), .C1(n_0_1), .C2(Enable), .ZN(n_0));
   NOR2_X1 i_0_1 (.A1(Q), .A2(Enable), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(D), .ZN(n_0_1));
endmodule

module TFlipFlop__4_7(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   AOI211_X1 i_0_0 (.A(n_0_0), .B(RST), .C1(Q), .C2(T), .ZN(n_0));
   NOR2_X1 i_0_1 (.A1(Q), .A2(T), .ZN(n_0_0));
endmodule

module TFlipFlop__4_12(T, CLK, RST, Enable, Q);
   input T;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   NOR2_X1 i_0_0 (.A1(n_0_0), .A2(RST), .ZN(n_0));
   XOR2_X1 i_0_1 (.A(Q), .B(n_0_1), .Z(n_0_0));
   NAND2_X1 i_0_2 (.A1(Enable), .A2(T), .ZN(n_0_1));
endmodule

module Counter(value, Enable, CLK, RST);
   output [1:0]value;
   input Enable;
   input CLK;
   input RST;

   wire inputs;

   TFlipFlop__4_7 firstBit (.T(Enable), .CLK(CLK), .RST(RST), .Enable(), 
      .Q(value[0]));
   TFlipFlop__4_12 genblk1_1_counterBits (.T(inputs), .CLK(CLK), .RST(RST), 
      .Enable(Enable), .Q(value[1]));
   AND2_X1 i_0_0 (.A1(Enable), .A2(value[0]), .ZN(inputs));
endmodule

module DFlipFlop(D, CLK, RST, Enable, Q);
   input D;
   input CLK;
   input RST;
   input Enable;
   output Q;

   wire n_0_0;
   wire n_0_1;

   DFF_X1 Q_reg (.D(n_0), .CK(CLK), .Q(Q), .QN());
   AOI211_X1 i_0_0 (.A(RST), .B(n_0_0), .C1(n_0_1), .C2(Enable), .ZN(n_0));
   NOR2_X1 i_0_1 (.A1(Q), .A2(Enable), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(D), .ZN(n_0_1));
endmodule

module Decoder_Receiver(RST, CLK, CPU_Bus, Loading_Enable, Done_Loading, 
      Done_Processing_Current_Packet, Done_Element, RAM_Address, RAM_Data);
   input RST;
   input CLK;
   input [31:0]CPU_Bus;
   input Loading_Enable;
   output Done_Loading;
   output Done_Processing_Current_Packet;
   output Done_Element;
   output [12:0]RAM_Address;
   output [63:0]RAM_Data;

   wire n_257_0;
   wire n_257_1;
   wire n_257_2;
   wire n_257_3;
   wire n_257_4;
   wire n_257_5;
   wire n_257_6;
   wire n_257_7;
   wire n_257_8;
   wire n_257_9;
   wire n_257_10;
   wire n_257_11;
   wire n_257_0_0;
   wire n_257_0_1;
   wire n_257_0_2;
   wire n_257_0_3;
   wire n_257_0_4;
   wire n_257_0_5;
   wire n_257_0_6;
   wire n_257_0_7;
   wire n_257_0_8;
   wire n_257_0_9;
   wire n_257_0_10;
   wire n_257_0_11;
   wire n_257_0_12;
   wire n_257_0_13;
   wire n_257_0_14;
   wire n_257_0_15;
   wire n_257_0_16;
   wire n_257_0_17;
   wire n_257_0_18;
   wire n_257_0_19;
   wire n_257_0_20;
   wire n_257_0_21;
   wire n_257_0_22;
   wire n_257_0_23;
   wire n_257_0_24;
   wire n_257_0_25;
   wire n_257_0_26;
   wire n_257_0_27;
   wire n_257_0_28;
   wire n_257_0_29;
   wire n_257_0_30;
   wire n_257_0_31;
   wire n_257_0_32;
   wire n_257_0_33;
   wire n_257_0_34;
   wire n_257_0_35;
   wire n_257_0_36;
   wire n_257_0_37;
   wire n_257_0_38;
   wire n_257_0_39;
   wire n_257_0_40;
   wire n_257_0_41;
   wire n_257_0_42;
   wire n_257_0_43;
   wire n_257_0_44;
   wire n_257_0_45;
   wire n_257_0_46;
   wire n_257_0_47;
   wire n_257_0_48;
   wire n_257_0_49;
   wire n_257_0_50;
   wire n_257_0_51;
   wire n_257_0_52;
   wire n_257_0_53;
   wire n_257_0_54;
   wire n_257_0_55;
   wire n_257_0_56;
   wire n_257_0_57;
   wire n_257_0_58;
   wire n_257_0_59;
   wire n_257_0_60;
   wire n_257_0_61;
   wire n_257_0_62;
   wire n_257_0_63;
   wire n_257_0_64;
   wire n_257_0_65;
   wire n_257_0_66;
   wire n_257_0_67;
   wire n_257_0_68;
   wire n_257_0_69;
   wire n_257_0_70;
   wire n_257_0_71;
   wire n_257_0_72;
   wire n_257_0_73;
   wire n_257_0_74;
   wire n_257_0_75;
   wire n_257_0_76;
   wire n_257_0_77;
   wire n_257_0_78;
   wire n_257_0_79;
   wire n_257_0_80;
   wire n_257_0_81;
   wire n_257_0_82;
   wire n_257_0_83;
   wire n_257_0_84;
   wire n_257_0_85;
   wire n_257_0_86;
   wire n_257_0_87;
   wire n_257_0_88;
   wire n_257_0_89;
   wire n_257_0_90;
   wire n_257_0_91;
   wire n_257_0_92;
   wire n_257_0_93;
   wire n_257_0_94;
   wire n_257_0_95;
   wire n_257_0_96;
   wire n_257_0_97;
   wire n_257_0_98;
   wire n_257_0_99;
   wire n_257_0_100;
   wire n_257_0_101;
   wire n_257_0_102;
   wire n_257_0_103;
   wire n_257_0_104;
   wire n_257_0_105;
   wire n_257_0_106;
   wire n_257_0_107;
   wire n_257_0_108;
   wire n_257_0_109;
   wire n_257_0_110;
   wire n_257_0_111;
   wire n_257_0_112;
   wire n_257_0_113;
   wire n_257_0_114;
   wire n_257_0_115;
   wire n_257_0_116;
   wire n_257_0_117;
   wire n_257_0_118;
   wire n_257_0_119;
   wire n_257_0_120;
   wire n_257_0_121;
   wire n_257_0_122;
   wire n_257_0_123;
   wire n_257_0_124;
   wire n_257_0_125;
   wire n_257_0_126;
   wire n_257_12;
   wire n_257_13;
   wire n_257_1_0;
   wire n_257_1_1;
   wire n_257_1_2;
   wire n_257_1_3;
   wire n_257_1_4;
   wire n_257_1_5;
   wire n_257_1_6;
   wire n_257_1_7;
   wire n_257_1_8;
   wire n_257_1_9;
   wire n_257_1_10;
   wire n_257_1_11;
   wire n_257_1_12;
   wire n_257_1_13;
   wire n_257_1_14;
   wire n_257_1_15;
   wire n_257_1_16;
   wire n_257_1_17;
   wire n_257_1_18;
   wire n_257_1_19;
   wire n_257_1_20;
   wire n_257_1_21;
   wire n_257_1_22;
   wire n_257_1_23;
   wire n_257_1_24;
   wire n_257_1_25;
   wire n_257_1_26;
   wire n_257_1_27;
   wire n_257_1_28;
   wire n_257_1_29;
   wire n_257_1_30;
   wire n_257_1_31;
   wire n_257_1_32;
   wire n_257_1_33;
   wire n_257_1_34;
   wire n_257_1_35;
   wire n_257_1_36;
   wire n_257_1_37;
   wire n_257_1_38;
   wire n_257_1_39;
   wire n_257_1_40;
   wire n_257_1_41;
   wire n_257_1_42;
   wire n_257_1_43;
   wire n_257_1_44;
   wire n_257_1_45;
   wire n_257_1_46;
   wire n_257_1_47;
   wire n_257_1_48;
   wire n_257_1_49;
   wire n_257_1_50;
   wire n_257_1_51;
   wire n_257_1_52;
   wire n_257_1_53;
   wire n_257_1_54;
   wire n_257_1_55;
   wire n_257_1_56;
   wire n_257_1_57;
   wire n_257_1_58;
   wire n_257_1_59;
   wire n_257_1_60;
   wire n_257_1_61;
   wire n_257_1_62;
   wire n_257_1_63;
   wire n_257_1_64;
   wire n_257_1_65;
   wire n_257_1_66;
   wire n_257_1_67;
   wire n_257_1_68;
   wire n_257_1_69;
   wire n_257_1_70;
   wire n_257_1_71;
   wire n_257_1_72;
   wire n_257_1_73;
   wire n_257_1_74;
   wire n_257_1_75;
   wire n_257_1_76;
   wire n_257_1_77;
   wire n_257_1_78;
   wire n_257_1_79;
   wire n_257_1_80;
   wire n_257_1_81;
   wire n_257_1_82;
   wire n_257_1_83;
   wire n_257_1_84;
   wire n_257_1_85;
   wire n_257_1_86;
   wire n_257_1_87;
   wire n_257_1_88;
   wire n_257_1_89;
   wire n_257_1_90;
   wire n_257_1_91;
   wire n_257_1_92;
   wire n_257_1_93;
   wire n_257_1_94;
   wire n_257_1_95;
   wire n_257_1_96;
   wire n_257_1_97;
   wire n_257_2_0;
   wire n_257_2_1;
   wire n_257_2_2;
   wire n_257_2_3;
   wire n_257_2_4;
   wire n_257_2_5;
   wire n_257_2_6;
   wire n_257_2_7;
   wire n_257_2_8;
   wire n_257_2_9;
   wire n_257_2_10;
   wire n_257_2_11;
   wire n_257_2_12;
   wire n_257_2_13;
   wire n_257_2_14;
   wire n_257_2_15;
   wire n_257_2_16;
   wire n_257_2_17;
   wire n_257_2_18;
   wire n_257_2_19;
   wire n_257_2_20;
   wire n_257_2_21;
   wire n_257_2_22;
   wire n_257_2_23;
   wire n_257_2_24;
   wire n_257_2_25;
   wire n_257_2_26;
   wire n_257_2_27;
   wire n_257_2_28;
   wire n_257_2_29;
   wire n_257_2_30;
   wire n_257_2_31;
   wire n_257_2_32;
   wire n_257_2_33;
   wire n_257_2_34;
   wire n_257_2_35;
   wire n_257_2_36;
   wire n_257_2_37;
   wire n_257_2_38;
   wire n_257_2_39;
   wire n_257_2_40;
   wire n_257_2_41;
   wire n_257_2_42;
   wire n_257_2_43;
   wire n_257_2_44;
   wire n_257_2_45;
   wire n_257_2_46;
   wire n_257_2_47;
   wire n_257_2_48;
   wire n_257_2_49;
   wire n_257_2_50;
   wire n_257_2_51;
   wire n_257_2_52;
   wire n_257_2_53;
   wire n_257_2_54;
   wire n_257_2_55;
   wire n_257_2_56;
   wire n_257_2_57;
   wire n_257_2_58;
   wire n_257_2_59;
   wire n_257_2_60;
   wire n_257_2_61;
   wire n_257_2_62;
   wire n_257_2_63;
   wire n_257_2_64;
   wire n_257_2_65;
   wire n_257_2_66;
   wire n_257_2_67;
   wire n_257_2_68;
   wire n_257_2_69;
   wire n_257_2_70;
   wire n_257_2_71;
   wire n_257_2_72;
   wire n_257_2_73;
   wire n_257_2_74;
   wire n_257_2_75;
   wire n_257_2_76;
   wire n_257_2_77;
   wire n_257_2_78;
   wire n_257_2_79;
   wire n_257_2_80;
   wire n_257_2_81;
   wire n_257_2_82;
   wire n_257_2_83;
   wire n_257_2_84;
   wire n_257_2_85;
   wire n_257_2_86;
   wire n_257_2_87;
   wire n_257_2_88;
   wire n_257_2_89;
   wire n_257_2_90;
   wire n_257_2_91;
   wire n_257_2_92;
   wire n_257_2_93;
   wire n_257_2_94;
   wire n_257_2_95;
   wire n_257_2_96;
   wire n_257_2_97;
   wire n_257_2_98;
   wire n_257_2_99;
   wire n_257_2_100;
   wire n_257_2_101;
   wire n_257_2_102;
   wire n_257_2_103;
   wire n_257_2_104;
   wire n_257_2_105;
   wire n_257_2_106;
   wire n_257_2_107;
   wire n_257_2_108;
   wire n_257_2_109;
   wire n_257_2_110;
   wire n_257_2_111;
   wire n_257_2_112;
   wire n_257_2_113;
   wire n_257_2_114;
   wire n_257_2_115;
   wire n_257_2_116;
   wire n_257_2_117;
   wire n_257_2_118;
   wire n_257_2_119;
   wire n_257_2_120;
   wire n_257_2_121;
   wire n_257_2_122;
   wire n_257_2_123;
   wire n_257_2_124;
   wire n_257_2_125;
   wire n_257_2_126;
   wire n_257_14;
   wire n_257_15;
   wire n_257_4_0;
   wire n_257_4_1;
   wire n_257_4_2;
   wire n_257_4_3;
   wire n_257_4_4;
   wire n_257_4_5;
   wire n_257_4_6;
   wire n_257_4_7;
   wire n_257_4_8;
   wire n_257_4_9;
   wire n_257_4_10;
   wire n_257_4_11;
   wire n_257_4_12;
   wire n_257_4_13;
   wire n_257_4_14;
   wire n_257_4_15;
   wire n_257_4_16;
   wire n_257_4_17;
   wire n_257_4_18;
   wire n_257_4_19;
   wire n_257_4_20;
   wire n_257_4_21;
   wire n_257_4_22;
   wire n_257_4_23;
   wire n_257_4_24;
   wire n_257_4_25;
   wire n_257_4_26;
   wire n_257_4_27;
   wire n_257_4_28;
   wire n_257_4_29;
   wire n_257_4_30;
   wire n_257_4_31;
   wire n_257_4_32;
   wire n_257_4_33;
   wire n_257_4_34;
   wire n_257_4_35;
   wire n_257_4_36;
   wire n_257_4_37;
   wire n_257_4_38;
   wire n_257_4_39;
   wire n_257_4_40;
   wire n_257_4_41;
   wire n_257_4_42;
   wire n_257_4_43;
   wire n_257_4_44;
   wire n_257_4_45;
   wire n_257_4_46;
   wire n_257_4_47;
   wire n_257_4_48;
   wire n_257_4_49;
   wire n_257_4_50;
   wire n_257_4_51;
   wire n_257_4_52;
   wire n_257_4_53;
   wire n_257_4_54;
   wire n_257_4_55;
   wire n_257_4_56;
   wire n_257_4_57;
   wire n_257_4_58;
   wire n_257_4_59;
   wire n_257_4_60;
   wire n_257_4_61;
   wire n_257_4_62;
   wire n_257_4_63;
   wire n_257_4_64;
   wire n_257_4_65;
   wire n_257_4_66;
   wire n_257_4_67;
   wire n_257_4_68;
   wire n_257_4_69;
   wire n_257_4_70;
   wire n_257_4_71;
   wire n_257_4_72;
   wire n_257_4_73;
   wire n_257_4_74;
   wire n_257_4_75;
   wire n_257_4_76;
   wire n_257_4_77;
   wire n_257_4_78;
   wire n_257_4_79;
   wire n_257_4_80;
   wire n_257_4_81;
   wire n_257_4_82;
   wire n_257_4_83;
   wire n_257_4_84;
   wire n_257_4_85;
   wire n_257_4_86;
   wire n_257_4_87;
   wire n_257_4_88;
   wire n_257_4_89;
   wire n_257_4_90;
   wire n_257_4_91;
   wire n_257_4_92;
   wire n_257_4_93;
   wire n_257_4_94;
   wire n_257_4_95;
   wire n_257_4_96;
   wire n_257_4_97;
   wire n_257_4_98;
   wire n_257_16;
   wire n_257_5_0;
   wire n_257_5_1;
   wire n_257_5_2;
   wire n_257_5_3;
   wire n_257_5_4;
   wire n_257_5_5;
   wire n_257_5_6;
   wire n_257_5_7;
   wire n_257_5_8;
   wire n_257_5_9;
   wire n_257_5_10;
   wire n_257_5_11;
   wire n_257_5_12;
   wire n_257_5_13;
   wire n_257_5_14;
   wire n_257_5_15;
   wire n_257_5_16;
   wire n_257_5_17;
   wire n_257_5_18;
   wire n_257_5_19;
   wire n_257_5_20;
   wire n_257_5_21;
   wire n_257_5_22;
   wire n_257_5_23;
   wire n_257_5_24;
   wire n_257_5_25;
   wire n_257_5_26;
   wire n_257_5_27;
   wire n_257_5_28;
   wire n_257_5_29;
   wire n_257_5_30;
   wire n_257_5_31;
   wire n_257_5_32;
   wire n_257_5_33;
   wire n_257_5_34;
   wire n_257_5_35;
   wire n_257_5_36;
   wire n_257_5_37;
   wire n_257_5_38;
   wire n_257_5_39;
   wire n_257_5_40;
   wire n_257_5_41;
   wire n_257_5_42;
   wire n_257_5_43;
   wire n_257_5_44;
   wire n_257_5_45;
   wire n_257_5_46;
   wire n_257_5_47;
   wire n_257_5_48;
   wire n_257_5_49;
   wire n_257_5_50;
   wire n_257_5_51;
   wire n_257_5_52;
   wire n_257_5_53;
   wire n_257_5_54;
   wire n_257_5_55;
   wire n_257_5_56;
   wire n_257_5_57;
   wire n_257_5_58;
   wire n_257_5_59;
   wire n_257_5_60;
   wire n_257_5_61;
   wire n_257_5_62;
   wire n_257_5_63;
   wire n_257_5_64;
   wire n_257_5_65;
   wire n_257_5_66;
   wire n_257_5_67;
   wire n_257_5_68;
   wire n_257_5_69;
   wire n_257_5_70;
   wire n_257_5_71;
   wire n_257_5_72;
   wire n_257_5_73;
   wire n_257_5_74;
   wire n_257_5_75;
   wire n_257_5_76;
   wire n_257_5_77;
   wire n_257_5_78;
   wire n_257_5_79;
   wire n_257_5_80;
   wire n_257_5_81;
   wire n_257_5_82;
   wire n_257_5_83;
   wire n_257_5_84;
   wire n_257_5_85;
   wire n_257_5_86;
   wire n_257_5_87;
   wire n_257_5_88;
   wire n_257_5_89;
   wire n_257_5_90;
   wire n_257_5_91;
   wire n_257_5_92;
   wire n_257_5_93;
   wire n_257_5_94;
   wire n_257_5_95;
   wire n_257_5_96;
   wire n_257_5_97;
   wire n_257_5_98;
   wire n_257_17;
   wire n_257_7_0;
   wire n_257_7_1;
   wire n_257_7_2;
   wire n_257_7_3;
   wire n_257_7_4;
   wire n_257_7_5;
   wire n_257_7_6;
   wire n_257_7_7;
   wire n_257_7_8;
   wire n_257_7_9;
   wire n_257_7_10;
   wire n_257_7_11;
   wire n_257_7_12;
   wire n_257_7_13;
   wire n_257_7_14;
   wire n_257_7_15;
   wire n_257_7_16;
   wire n_257_7_17;
   wire n_257_7_18;
   wire n_257_7_19;
   wire n_257_7_20;
   wire n_257_7_21;
   wire n_257_7_22;
   wire n_257_7_23;
   wire n_257_7_24;
   wire n_257_7_25;
   wire n_257_7_26;
   wire n_257_7_27;
   wire n_257_7_28;
   wire n_257_7_29;
   wire n_257_7_30;
   wire n_257_7_31;
   wire n_257_7_32;
   wire n_257_7_33;
   wire n_257_7_34;
   wire n_257_7_35;
   wire n_257_7_36;
   wire n_257_7_37;
   wire n_257_7_38;
   wire n_257_7_39;
   wire n_257_7_40;
   wire n_257_7_41;
   wire n_257_7_42;
   wire n_257_7_43;
   wire n_257_7_44;
   wire n_257_7_45;
   wire n_257_7_46;
   wire n_257_7_47;
   wire n_257_7_48;
   wire n_257_7_49;
   wire n_257_7_50;
   wire n_257_7_51;
   wire n_257_7_52;
   wire n_257_7_53;
   wire n_257_7_54;
   wire n_257_7_55;
   wire n_257_7_56;
   wire n_257_7_57;
   wire n_257_7_58;
   wire n_257_7_59;
   wire n_257_7_60;
   wire n_257_7_61;
   wire n_257_7_62;
   wire n_257_7_63;
   wire n_257_7_64;
   wire n_257_7_65;
   wire n_257_7_66;
   wire n_257_7_67;
   wire n_257_7_68;
   wire n_257_7_69;
   wire n_257_7_70;
   wire n_257_7_71;
   wire n_257_7_72;
   wire n_257_7_73;
   wire n_257_7_74;
   wire n_257_7_75;
   wire n_257_7_76;
   wire n_257_7_77;
   wire n_257_7_78;
   wire n_257_7_79;
   wire n_257_7_80;
   wire n_257_7_81;
   wire n_257_7_82;
   wire n_257_7_83;
   wire n_257_7_84;
   wire n_257_7_85;
   wire n_257_7_86;
   wire n_257_7_87;
   wire n_257_7_88;
   wire n_257_7_89;
   wire n_257_7_90;
   wire n_257_7_91;
   wire n_257_7_92;
   wire n_257_7_93;
   wire n_257_7_94;
   wire n_257_7_95;
   wire n_257_7_96;
   wire n_257_7_97;
   wire n_257_18;
   wire n_257_8_0;
   wire n_257_8_1;
   wire n_257_8_2;
   wire n_257_8_3;
   wire n_257_8_4;
   wire n_257_8_5;
   wire n_257_8_6;
   wire n_257_8_7;
   wire n_257_8_8;
   wire n_257_8_9;
   wire n_257_8_10;
   wire n_257_8_11;
   wire n_257_8_12;
   wire n_257_8_13;
   wire n_257_8_14;
   wire n_257_8_15;
   wire n_257_8_16;
   wire n_257_8_17;
   wire n_257_8_18;
   wire n_257_8_19;
   wire n_257_8_20;
   wire n_257_8_21;
   wire n_257_8_22;
   wire n_257_8_23;
   wire n_257_8_24;
   wire n_257_8_25;
   wire n_257_8_26;
   wire n_257_8_27;
   wire n_257_8_28;
   wire n_257_8_29;
   wire n_257_8_30;
   wire n_257_8_31;
   wire n_257_8_32;
   wire n_257_8_33;
   wire n_257_8_34;
   wire n_257_8_35;
   wire n_257_8_36;
   wire n_257_8_37;
   wire n_257_8_38;
   wire n_257_8_39;
   wire n_257_8_40;
   wire n_257_8_41;
   wire n_257_8_42;
   wire n_257_8_43;
   wire n_257_8_44;
   wire n_257_8_45;
   wire n_257_8_46;
   wire n_257_8_47;
   wire n_257_8_48;
   wire n_257_8_49;
   wire n_257_8_50;
   wire n_257_8_51;
   wire n_257_8_52;
   wire n_257_8_53;
   wire n_257_8_54;
   wire n_257_8_55;
   wire n_257_8_56;
   wire n_257_8_57;
   wire n_257_8_58;
   wire n_257_8_59;
   wire n_257_8_60;
   wire n_257_8_61;
   wire n_257_8_62;
   wire n_257_8_63;
   wire n_257_8_64;
   wire n_257_8_65;
   wire n_257_8_66;
   wire n_257_8_67;
   wire n_257_8_68;
   wire n_257_8_69;
   wire n_257_8_70;
   wire n_257_8_71;
   wire n_257_8_72;
   wire n_257_8_73;
   wire n_257_8_74;
   wire n_257_8_75;
   wire n_257_8_76;
   wire n_257_8_77;
   wire n_257_8_78;
   wire n_257_8_79;
   wire n_257_8_80;
   wire n_257_8_81;
   wire n_257_8_82;
   wire n_257_8_83;
   wire n_257_8_84;
   wire n_257_8_85;
   wire n_257_8_86;
   wire n_257_8_87;
   wire n_257_8_88;
   wire n_257_8_89;
   wire n_257_8_90;
   wire n_257_8_91;
   wire n_257_8_92;
   wire n_257_8_93;
   wire n_257_8_94;
   wire n_257_8_95;
   wire n_257_8_96;
   wire n_257_8_97;
   wire n_257_19;
   wire n_257_9_0;
   wire n_257_9_1;
   wire n_257_9_2;
   wire n_257_9_3;
   wire n_257_9_4;
   wire n_257_9_5;
   wire n_257_9_6;
   wire n_257_9_7;
   wire n_257_9_8;
   wire n_257_9_9;
   wire n_257_9_10;
   wire n_257_9_11;
   wire n_257_9_12;
   wire n_257_9_13;
   wire n_257_9_14;
   wire n_257_9_15;
   wire n_257_9_16;
   wire n_257_9_17;
   wire n_257_9_18;
   wire n_257_9_19;
   wire n_257_9_20;
   wire n_257_9_21;
   wire n_257_9_22;
   wire n_257_9_23;
   wire n_257_9_24;
   wire n_257_9_25;
   wire n_257_9_26;
   wire n_257_9_27;
   wire n_257_9_28;
   wire n_257_9_29;
   wire n_257_9_30;
   wire n_257_9_31;
   wire n_257_9_32;
   wire n_257_9_33;
   wire n_257_9_34;
   wire n_257_9_35;
   wire n_257_9_36;
   wire n_257_9_37;
   wire n_257_9_38;
   wire n_257_9_39;
   wire n_257_9_40;
   wire n_257_9_41;
   wire n_257_9_42;
   wire n_257_9_43;
   wire n_257_9_44;
   wire n_257_9_45;
   wire n_257_9_46;
   wire n_257_9_47;
   wire n_257_9_48;
   wire n_257_9_49;
   wire n_257_9_50;
   wire n_257_9_51;
   wire n_257_9_52;
   wire n_257_9_53;
   wire n_257_9_54;
   wire n_257_9_55;
   wire n_257_9_56;
   wire n_257_9_57;
   wire n_257_9_58;
   wire n_257_9_59;
   wire n_257_9_60;
   wire n_257_9_61;
   wire n_257_9_62;
   wire n_257_9_63;
   wire n_257_9_64;
   wire n_257_9_65;
   wire n_257_9_66;
   wire n_257_9_67;
   wire n_257_9_68;
   wire n_257_9_69;
   wire n_257_9_70;
   wire n_257_9_71;
   wire n_257_9_72;
   wire n_257_9_73;
   wire n_257_9_74;
   wire n_257_9_75;
   wire n_257_9_76;
   wire n_257_9_77;
   wire n_257_9_78;
   wire n_257_9_79;
   wire n_257_9_80;
   wire n_257_9_81;
   wire n_257_9_82;
   wire n_257_9_83;
   wire n_257_9_84;
   wire n_257_9_85;
   wire n_257_9_86;
   wire n_257_9_87;
   wire n_257_9_88;
   wire n_257_9_89;
   wire n_257_9_90;
   wire n_257_9_91;
   wire n_257_9_92;
   wire n_257_9_93;
   wire n_257_9_94;
   wire n_257_9_95;
   wire n_257_9_96;
   wire n_257_9_97;
   wire n_257_9_98;
   wire n_257_20;
   wire n_257_10_0;
   wire n_257_10_1;
   wire n_257_10_2;
   wire n_257_10_3;
   wire n_257_10_4;
   wire n_257_10_5;
   wire n_257_10_6;
   wire n_257_10_7;
   wire n_257_10_8;
   wire n_257_10_9;
   wire n_257_10_10;
   wire n_257_10_11;
   wire n_257_10_12;
   wire n_257_10_13;
   wire n_257_10_14;
   wire n_257_10_15;
   wire n_257_10_16;
   wire n_257_10_17;
   wire n_257_10_18;
   wire n_257_10_19;
   wire n_257_10_20;
   wire n_257_10_21;
   wire n_257_10_22;
   wire n_257_10_23;
   wire n_257_10_24;
   wire n_257_10_25;
   wire n_257_10_26;
   wire n_257_10_27;
   wire n_257_10_28;
   wire n_257_10_29;
   wire n_257_10_30;
   wire n_257_10_31;
   wire n_257_10_32;
   wire n_257_10_33;
   wire n_257_10_34;
   wire n_257_10_35;
   wire n_257_10_36;
   wire n_257_10_37;
   wire n_257_10_38;
   wire n_257_10_39;
   wire n_257_10_40;
   wire n_257_10_41;
   wire n_257_10_42;
   wire n_257_10_43;
   wire n_257_10_44;
   wire n_257_10_45;
   wire n_257_10_46;
   wire n_257_10_47;
   wire n_257_10_48;
   wire n_257_10_49;
   wire n_257_10_50;
   wire n_257_10_51;
   wire n_257_10_52;
   wire n_257_10_53;
   wire n_257_10_54;
   wire n_257_10_55;
   wire n_257_10_56;
   wire n_257_10_57;
   wire n_257_10_58;
   wire n_257_10_59;
   wire n_257_10_60;
   wire n_257_10_61;
   wire n_257_10_62;
   wire n_257_10_63;
   wire n_257_10_64;
   wire n_257_10_65;
   wire n_257_10_66;
   wire n_257_10_67;
   wire n_257_10_68;
   wire n_257_10_69;
   wire n_257_10_70;
   wire n_257_10_71;
   wire n_257_10_72;
   wire n_257_10_73;
   wire n_257_10_74;
   wire n_257_10_75;
   wire n_257_10_76;
   wire n_257_10_77;
   wire n_257_10_78;
   wire n_257_10_79;
   wire n_257_10_80;
   wire n_257_10_81;
   wire n_257_10_82;
   wire n_257_10_83;
   wire n_257_10_84;
   wire n_257_10_85;
   wire n_257_10_86;
   wire n_257_10_87;
   wire n_257_10_88;
   wire n_257_10_89;
   wire n_257_10_90;
   wire n_257_10_91;
   wire n_257_10_92;
   wire n_257_10_93;
   wire n_257_10_94;
   wire n_257_10_95;
   wire n_257_10_96;
   wire n_257_10_97;
   wire n_257_10_98;
   wire n_257_11_0;
   wire n_257_11_1;
   wire n_257_11_2;
   wire n_257_11_3;
   wire n_257_11_4;
   wire n_257_11_5;
   wire n_257_11_6;
   wire n_257_11_7;
   wire n_257_11_8;
   wire n_257_11_9;
   wire n_257_11_10;
   wire n_257_11_11;
   wire n_257_11_12;
   wire n_257_11_13;
   wire n_257_11_14;
   wire n_257_11_15;
   wire n_257_11_16;
   wire n_257_11_17;
   wire n_257_11_18;
   wire n_257_11_19;
   wire n_257_11_20;
   wire n_257_11_21;
   wire n_257_11_22;
   wire n_257_11_23;
   wire n_257_11_24;
   wire n_257_11_25;
   wire n_257_11_26;
   wire n_257_11_27;
   wire n_257_11_28;
   wire n_257_11_29;
   wire n_257_11_30;
   wire n_257_11_31;
   wire n_257_11_32;
   wire n_257_11_33;
   wire n_257_11_34;
   wire n_257_11_35;
   wire n_257_11_36;
   wire n_257_11_37;
   wire n_257_11_38;
   wire n_257_11_39;
   wire n_257_11_40;
   wire n_257_11_41;
   wire n_257_11_42;
   wire n_257_11_43;
   wire n_257_11_44;
   wire n_257_11_45;
   wire n_257_11_46;
   wire n_257_11_47;
   wire n_257_11_48;
   wire n_257_11_49;
   wire n_257_11_50;
   wire n_257_11_51;
   wire n_257_11_52;
   wire n_257_11_53;
   wire n_257_11_54;
   wire n_257_11_55;
   wire n_257_11_56;
   wire n_257_11_57;
   wire n_257_11_58;
   wire n_257_11_59;
   wire n_257_11_60;
   wire n_257_11_61;
   wire n_257_11_62;
   wire n_257_11_63;
   wire n_257_11_64;
   wire n_257_11_65;
   wire n_257_11_66;
   wire n_257_11_67;
   wire n_257_11_68;
   wire n_257_11_69;
   wire n_257_11_70;
   wire n_257_11_71;
   wire n_257_11_72;
   wire n_257_11_73;
   wire n_257_11_74;
   wire n_257_11_75;
   wire n_257_11_76;
   wire n_257_11_77;
   wire n_257_11_78;
   wire n_257_11_79;
   wire n_257_11_80;
   wire n_257_11_81;
   wire n_257_11_82;
   wire n_257_11_83;
   wire n_257_11_84;
   wire n_257_11_85;
   wire n_257_11_86;
   wire n_257_11_87;
   wire n_257_11_88;
   wire n_257_11_89;
   wire n_257_11_90;
   wire n_257_11_91;
   wire n_257_11_92;
   wire n_257_11_93;
   wire n_257_11_94;
   wire n_257_11_95;
   wire n_257_11_96;
   wire n_257_11_97;
   wire n_257_11_98;
   wire n_257_11_99;
   wire n_257_11_100;
   wire n_257_11_101;
   wire n_257_11_102;
   wire n_257_11_103;
   wire n_257_11_104;
   wire n_257_11_105;
   wire n_257_11_106;
   wire n_257_11_107;
   wire n_257_11_108;
   wire n_257_11_109;
   wire n_257_11_110;
   wire n_257_11_111;
   wire n_257_11_112;
   wire n_257_11_113;
   wire n_257_11_114;
   wire n_257_11_115;
   wire n_257_11_116;
   wire n_257_11_117;
   wire n_257_11_118;
   wire n_257_11_119;
   wire n_257_11_120;
   wire n_257_11_121;
   wire n_257_11_122;
   wire n_257_11_123;
   wire n_257_11_124;
   wire n_257_11_125;
   wire n_257_11_126;
   wire n_257_21;
   wire n_257_22;
   wire n_257_12_0;
   wire n_257_12_1;
   wire n_257_12_2;
   wire n_257_12_3;
   wire n_257_12_4;
   wire n_257_12_5;
   wire n_257_12_6;
   wire n_257_12_7;
   wire n_257_12_8;
   wire n_257_12_9;
   wire n_257_12_10;
   wire n_257_12_11;
   wire n_257_12_12;
   wire n_257_12_13;
   wire n_257_12_14;
   wire n_257_12_15;
   wire n_257_12_16;
   wire n_257_12_17;
   wire n_257_12_18;
   wire n_257_12_19;
   wire n_257_12_20;
   wire n_257_12_21;
   wire n_257_12_22;
   wire n_257_12_23;
   wire n_257_12_24;
   wire n_257_12_25;
   wire n_257_12_26;
   wire n_257_12_27;
   wire n_257_12_28;
   wire n_257_12_29;
   wire n_257_12_30;
   wire n_257_12_31;
   wire n_257_12_32;
   wire n_257_12_33;
   wire n_257_12_34;
   wire n_257_12_35;
   wire n_257_12_36;
   wire n_257_12_37;
   wire n_257_12_38;
   wire n_257_12_39;
   wire n_257_12_40;
   wire n_257_12_41;
   wire n_257_12_42;
   wire n_257_12_43;
   wire n_257_12_44;
   wire n_257_12_45;
   wire n_257_12_46;
   wire n_257_12_47;
   wire n_257_12_48;
   wire n_257_12_49;
   wire n_257_12_50;
   wire n_257_12_51;
   wire n_257_12_52;
   wire n_257_12_53;
   wire n_257_12_54;
   wire n_257_12_55;
   wire n_257_12_56;
   wire n_257_12_57;
   wire n_257_12_58;
   wire n_257_12_59;
   wire n_257_12_60;
   wire n_257_12_61;
   wire n_257_12_62;
   wire n_257_12_63;
   wire n_257_12_64;
   wire n_257_12_65;
   wire n_257_12_66;
   wire n_257_12_67;
   wire n_257_12_68;
   wire n_257_12_69;
   wire n_257_12_70;
   wire n_257_12_71;
   wire n_257_12_72;
   wire n_257_12_73;
   wire n_257_12_74;
   wire n_257_12_75;
   wire n_257_12_76;
   wire n_257_12_77;
   wire n_257_12_78;
   wire n_257_12_79;
   wire n_257_12_80;
   wire n_257_12_81;
   wire n_257_12_82;
   wire n_257_12_83;
   wire n_257_12_84;
   wire n_257_12_85;
   wire n_257_12_86;
   wire n_257_12_87;
   wire n_257_12_88;
   wire n_257_12_89;
   wire n_257_12_90;
   wire n_257_12_91;
   wire n_257_12_92;
   wire n_257_12_93;
   wire n_257_12_94;
   wire n_257_12_95;
   wire n_257_12_96;
   wire n_257_12_97;
   wire n_257_23;
   wire n_257_13_0;
   wire n_257_13_1;
   wire n_257_13_2;
   wire n_257_13_3;
   wire n_257_13_4;
   wire n_257_13_5;
   wire n_257_13_6;
   wire n_257_13_7;
   wire n_257_13_8;
   wire n_257_13_9;
   wire n_257_13_10;
   wire n_257_13_11;
   wire n_257_13_12;
   wire n_257_13_13;
   wire n_257_13_14;
   wire n_257_13_15;
   wire n_257_13_16;
   wire n_257_13_17;
   wire n_257_13_18;
   wire n_257_13_19;
   wire n_257_13_20;
   wire n_257_13_21;
   wire n_257_13_22;
   wire n_257_13_23;
   wire n_257_13_24;
   wire n_257_13_25;
   wire n_257_13_26;
   wire n_257_13_27;
   wire n_257_13_28;
   wire n_257_13_29;
   wire n_257_13_30;
   wire n_257_13_31;
   wire n_257_13_32;
   wire n_257_13_33;
   wire n_257_13_34;
   wire n_257_13_35;
   wire n_257_13_36;
   wire n_257_13_37;
   wire n_257_13_38;
   wire n_257_13_39;
   wire n_257_13_40;
   wire n_257_13_41;
   wire n_257_13_42;
   wire n_257_13_43;
   wire n_257_13_44;
   wire n_257_13_45;
   wire n_257_13_46;
   wire n_257_13_47;
   wire n_257_13_48;
   wire n_257_13_49;
   wire n_257_13_50;
   wire n_257_13_51;
   wire n_257_13_52;
   wire n_257_13_53;
   wire n_257_13_54;
   wire n_257_13_55;
   wire n_257_13_56;
   wire n_257_13_57;
   wire n_257_13_58;
   wire n_257_13_59;
   wire n_257_13_60;
   wire n_257_13_61;
   wire n_257_13_62;
   wire n_257_13_63;
   wire n_257_13_64;
   wire n_257_13_65;
   wire n_257_13_66;
   wire n_257_13_67;
   wire n_257_13_68;
   wire n_257_13_69;
   wire n_257_13_70;
   wire n_257_13_71;
   wire n_257_13_72;
   wire n_257_13_73;
   wire n_257_13_74;
   wire n_257_13_75;
   wire n_257_13_76;
   wire n_257_13_77;
   wire n_257_13_78;
   wire n_257_13_79;
   wire n_257_13_80;
   wire n_257_13_81;
   wire n_257_13_82;
   wire n_257_13_83;
   wire n_257_13_84;
   wire n_257_13_85;
   wire n_257_13_86;
   wire n_257_13_87;
   wire n_257_13_88;
   wire n_257_24;
   wire n_257_14_0;
   wire n_257_14_1;
   wire n_257_14_2;
   wire n_257_14_3;
   wire n_257_14_4;
   wire n_257_14_5;
   wire n_257_14_6;
   wire n_257_14_7;
   wire n_257_14_8;
   wire n_257_14_9;
   wire n_257_14_10;
   wire n_257_14_11;
   wire n_257_14_12;
   wire n_257_14_13;
   wire n_257_14_14;
   wire n_257_14_15;
   wire n_257_14_16;
   wire n_257_14_17;
   wire n_257_14_18;
   wire n_257_14_19;
   wire n_257_14_20;
   wire n_257_14_21;
   wire n_257_14_22;
   wire n_257_14_23;
   wire n_257_14_24;
   wire n_257_14_25;
   wire n_257_14_26;
   wire n_257_14_27;
   wire n_257_14_28;
   wire n_257_14_29;
   wire n_257_14_30;
   wire n_257_14_31;
   wire n_257_14_32;
   wire n_257_14_33;
   wire n_257_14_34;
   wire n_257_14_35;
   wire n_257_14_36;
   wire n_257_14_37;
   wire n_257_14_38;
   wire n_257_14_39;
   wire n_257_14_40;
   wire n_257_14_41;
   wire n_257_14_42;
   wire n_257_14_43;
   wire n_257_14_44;
   wire n_257_14_45;
   wire n_257_14_46;
   wire n_257_14_47;
   wire n_257_14_48;
   wire n_257_14_49;
   wire n_257_14_50;
   wire n_257_14_51;
   wire n_257_14_52;
   wire n_257_14_53;
   wire n_257_14_54;
   wire n_257_14_55;
   wire n_257_14_56;
   wire n_257_14_57;
   wire n_257_14_58;
   wire n_257_14_59;
   wire n_257_14_60;
   wire n_257_14_61;
   wire n_257_14_62;
   wire n_257_14_63;
   wire n_257_14_64;
   wire n_257_14_65;
   wire n_257_14_66;
   wire n_257_14_67;
   wire n_257_14_68;
   wire n_257_14_69;
   wire n_257_14_70;
   wire n_257_14_71;
   wire n_257_14_72;
   wire n_257_14_73;
   wire n_257_14_74;
   wire n_257_14_75;
   wire n_257_14_76;
   wire n_257_14_77;
   wire n_257_14_78;
   wire n_257_14_79;
   wire n_257_14_80;
   wire n_257_14_81;
   wire n_257_14_82;
   wire n_257_14_83;
   wire n_257_14_84;
   wire n_257_14_85;
   wire n_257_14_86;
   wire n_257_14_87;
   wire n_257_14_88;
   wire n_257_14_89;
   wire n_257_14_90;
   wire n_257_14_91;
   wire n_257_14_92;
   wire n_257_14_93;
   wire n_257_14_94;
   wire n_257_14_95;
   wire n_257_14_96;
   wire n_257_14_97;
   wire n_257_14_98;
   wire n_257_15_0;
   wire n_257_15_1;
   wire n_257_15_2;
   wire n_257_15_3;
   wire n_257_15_4;
   wire n_257_15_5;
   wire n_257_15_6;
   wire n_257_15_7;
   wire n_257_15_8;
   wire n_257_15_9;
   wire n_257_15_10;
   wire n_257_15_11;
   wire n_257_15_12;
   wire n_257_15_13;
   wire n_257_15_14;
   wire n_257_15_15;
   wire n_257_15_16;
   wire n_257_15_17;
   wire n_257_15_18;
   wire n_257_15_19;
   wire n_257_15_20;
   wire n_257_15_21;
   wire n_257_15_22;
   wire n_257_15_23;
   wire n_257_15_24;
   wire n_257_15_25;
   wire n_257_15_26;
   wire n_257_15_27;
   wire n_257_15_28;
   wire n_257_15_29;
   wire n_257_15_30;
   wire n_257_15_31;
   wire n_257_15_32;
   wire n_257_15_33;
   wire n_257_15_34;
   wire n_257_15_35;
   wire n_257_15_36;
   wire n_257_15_37;
   wire n_257_15_38;
   wire n_257_15_39;
   wire n_257_15_40;
   wire n_257_15_41;
   wire n_257_15_42;
   wire n_257_15_43;
   wire n_257_15_44;
   wire n_257_15_45;
   wire n_257_15_46;
   wire n_257_15_47;
   wire n_257_15_48;
   wire n_257_15_49;
   wire n_257_15_50;
   wire n_257_15_51;
   wire n_257_15_52;
   wire n_257_15_53;
   wire n_257_15_54;
   wire n_257_15_55;
   wire n_257_15_56;
   wire n_257_15_57;
   wire n_257_15_58;
   wire n_257_15_59;
   wire n_257_15_60;
   wire n_257_15_61;
   wire n_257_15_62;
   wire n_257_15_63;
   wire n_257_15_64;
   wire n_257_15_65;
   wire n_257_15_66;
   wire n_257_15_67;
   wire n_257_15_68;
   wire n_257_15_69;
   wire n_257_15_70;
   wire n_257_15_71;
   wire n_257_15_72;
   wire n_257_15_73;
   wire n_257_15_74;
   wire n_257_15_75;
   wire n_257_15_76;
   wire n_257_15_77;
   wire n_257_15_78;
   wire n_257_15_79;
   wire n_257_15_80;
   wire n_257_15_81;
   wire n_257_15_82;
   wire n_257_15_83;
   wire n_257_15_84;
   wire n_257_15_85;
   wire n_257_15_86;
   wire n_257_15_87;
   wire n_257_15_88;
   wire n_257_15_89;
   wire n_257_15_90;
   wire n_257_15_91;
   wire n_257_15_92;
   wire n_257_15_93;
   wire n_257_15_94;
   wire n_257_15_95;
   wire n_257_15_96;
   wire n_257_15_97;
   wire n_257_15_98;
   wire n_257_15_99;
   wire n_257_15_100;
   wire n_257_15_101;
   wire n_257_15_102;
   wire n_257_15_103;
   wire n_257_15_104;
   wire n_257_15_105;
   wire n_257_15_106;
   wire n_257_15_107;
   wire n_257_15_108;
   wire n_257_15_109;
   wire n_257_15_110;
   wire n_257_15_111;
   wire n_257_15_112;
   wire n_257_15_113;
   wire n_257_15_114;
   wire n_257_15_115;
   wire n_257_15_116;
   wire n_257_15_117;
   wire n_257_15_118;
   wire n_257_15_119;
   wire n_257_15_120;
   wire n_257_15_121;
   wire n_257_15_122;
   wire n_257_15_123;
   wire n_257_15_124;
   wire n_257_15_125;
   wire n_257_15_126;
   wire n_257_25;
   wire n_257_16_0;
   wire n_257_16_1;
   wire n_257_16_2;
   wire n_257_16_3;
   wire n_257_16_4;
   wire n_257_16_5;
   wire n_257_16_6;
   wire n_257_16_7;
   wire n_257_16_8;
   wire n_257_16_9;
   wire n_257_16_10;
   wire n_257_16_11;
   wire n_257_16_12;
   wire n_257_16_13;
   wire n_257_16_14;
   wire n_257_16_15;
   wire n_257_16_16;
   wire n_257_16_17;
   wire n_257_16_18;
   wire n_257_16_19;
   wire n_257_16_20;
   wire n_257_16_21;
   wire n_257_16_22;
   wire n_257_16_23;
   wire n_257_16_24;
   wire n_257_16_25;
   wire n_257_16_26;
   wire n_257_16_27;
   wire n_257_16_28;
   wire n_257_16_29;
   wire n_257_16_30;
   wire n_257_16_31;
   wire n_257_16_32;
   wire n_257_16_33;
   wire n_257_16_34;
   wire n_257_16_35;
   wire n_257_16_36;
   wire n_257_16_37;
   wire n_257_16_38;
   wire n_257_16_39;
   wire n_257_16_40;
   wire n_257_16_41;
   wire n_257_16_42;
   wire n_257_16_43;
   wire n_257_16_44;
   wire n_257_16_45;
   wire n_257_16_46;
   wire n_257_16_47;
   wire n_257_16_48;
   wire n_257_16_49;
   wire n_257_16_50;
   wire n_257_16_51;
   wire n_257_16_52;
   wire n_257_16_53;
   wire n_257_16_54;
   wire n_257_16_55;
   wire n_257_16_56;
   wire n_257_16_57;
   wire n_257_16_58;
   wire n_257_16_59;
   wire n_257_16_60;
   wire n_257_16_61;
   wire n_257_16_62;
   wire n_257_16_63;
   wire n_257_16_64;
   wire n_257_16_65;
   wire n_257_16_66;
   wire n_257_16_67;
   wire n_257_16_68;
   wire n_257_16_69;
   wire n_257_16_70;
   wire n_257_16_71;
   wire n_257_16_72;
   wire n_257_16_73;
   wire n_257_16_74;
   wire n_257_16_75;
   wire n_257_16_76;
   wire n_257_16_77;
   wire n_257_16_78;
   wire n_257_16_79;
   wire n_257_16_80;
   wire n_257_16_81;
   wire n_257_16_82;
   wire n_257_16_83;
   wire n_257_16_84;
   wire n_257_16_85;
   wire n_257_16_86;
   wire n_257_16_87;
   wire n_257_16_88;
   wire n_257_16_89;
   wire n_257_16_90;
   wire n_257_16_91;
   wire n_257_16_92;
   wire n_257_16_93;
   wire n_257_16_94;
   wire n_257_16_95;
   wire n_257_16_96;
   wire n_257_16_97;
   wire n_257_16_98;
   wire n_257_16_99;
   wire n_257_16_100;
   wire n_257_16_101;
   wire n_257_16_102;
   wire n_257_16_103;
   wire n_257_16_104;
   wire n_257_16_105;
   wire n_257_16_106;
   wire n_257_16_107;
   wire n_257_16_108;
   wire n_257_16_109;
   wire n_257_16_110;
   wire n_257_16_111;
   wire n_257_16_112;
   wire n_257_16_113;
   wire n_257_16_114;
   wire n_257_16_115;
   wire n_257_16_116;
   wire n_257_16_117;
   wire n_257_16_118;
   wire n_257_16_119;
   wire n_257_16_120;
   wire n_257_16_121;
   wire n_257_16_122;
   wire n_257_16_123;
   wire n_257_16_124;
   wire n_257_16_125;
   wire n_257_16_126;
   wire n_257_26;
   wire n_257_27;
   wire n_257_17_0;
   wire n_257_17_1;
   wire n_257_17_2;
   wire n_257_17_3;
   wire n_257_17_4;
   wire n_257_17_5;
   wire n_257_17_6;
   wire n_257_17_7;
   wire n_257_17_8;
   wire n_257_17_9;
   wire n_257_17_10;
   wire n_257_17_11;
   wire n_257_17_12;
   wire n_257_17_13;
   wire n_257_17_14;
   wire n_257_17_15;
   wire n_257_17_16;
   wire n_257_17_17;
   wire n_257_17_18;
   wire n_257_17_19;
   wire n_257_17_20;
   wire n_257_17_21;
   wire n_257_17_22;
   wire n_257_17_23;
   wire n_257_17_24;
   wire n_257_17_25;
   wire n_257_17_26;
   wire n_257_17_27;
   wire n_257_17_28;
   wire n_257_17_29;
   wire n_257_17_30;
   wire n_257_17_31;
   wire n_257_17_32;
   wire n_257_17_33;
   wire n_257_17_34;
   wire n_257_17_35;
   wire n_257_17_36;
   wire n_257_17_37;
   wire n_257_17_38;
   wire n_257_17_39;
   wire n_257_17_40;
   wire n_257_17_41;
   wire n_257_17_42;
   wire n_257_17_43;
   wire n_257_17_44;
   wire n_257_17_45;
   wire n_257_17_46;
   wire n_257_17_47;
   wire n_257_17_48;
   wire n_257_17_49;
   wire n_257_17_50;
   wire n_257_17_51;
   wire n_257_17_52;
   wire n_257_17_53;
   wire n_257_17_54;
   wire n_257_17_55;
   wire n_257_17_56;
   wire n_257_17_57;
   wire n_257_17_58;
   wire n_257_17_59;
   wire n_257_17_60;
   wire n_257_17_61;
   wire n_257_17_62;
   wire n_257_17_63;
   wire n_257_17_64;
   wire n_257_17_65;
   wire n_257_17_66;
   wire n_257_17_67;
   wire n_257_17_68;
   wire n_257_17_69;
   wire n_257_17_70;
   wire n_257_17_71;
   wire n_257_17_72;
   wire n_257_17_73;
   wire n_257_17_74;
   wire n_257_17_75;
   wire n_257_17_76;
   wire n_257_17_77;
   wire n_257_17_78;
   wire n_257_17_79;
   wire n_257_17_80;
   wire n_257_17_81;
   wire n_257_17_82;
   wire n_257_17_83;
   wire n_257_17_84;
   wire n_257_17_85;
   wire n_257_17_86;
   wire n_257_17_87;
   wire n_257_17_88;
   wire n_257_17_89;
   wire n_257_17_90;
   wire n_257_17_91;
   wire n_257_17_92;
   wire n_257_17_93;
   wire n_257_17_94;
   wire n_257_17_95;
   wire n_257_17_96;
   wire n_257_17_97;
   wire n_257_17_98;
   wire n_257_28;
   wire n_257_18_0;
   wire n_257_18_1;
   wire n_257_18_2;
   wire n_257_18_3;
   wire n_257_18_4;
   wire n_257_18_5;
   wire n_257_18_6;
   wire n_257_18_7;
   wire n_257_18_8;
   wire n_257_18_9;
   wire n_257_18_10;
   wire n_257_18_11;
   wire n_257_18_12;
   wire n_257_18_13;
   wire n_257_18_14;
   wire n_257_18_15;
   wire n_257_18_16;
   wire n_257_18_17;
   wire n_257_18_18;
   wire n_257_18_19;
   wire n_257_18_20;
   wire n_257_18_21;
   wire n_257_18_22;
   wire n_257_18_23;
   wire n_257_18_24;
   wire n_257_18_25;
   wire n_257_18_26;
   wire n_257_18_27;
   wire n_257_18_28;
   wire n_257_18_29;
   wire n_257_18_30;
   wire n_257_18_31;
   wire n_257_18_32;
   wire n_257_18_33;
   wire n_257_18_34;
   wire n_257_18_35;
   wire n_257_18_36;
   wire n_257_18_37;
   wire n_257_18_38;
   wire n_257_18_39;
   wire n_257_18_40;
   wire n_257_18_41;
   wire n_257_18_42;
   wire n_257_18_43;
   wire n_257_18_44;
   wire n_257_18_45;
   wire n_257_18_46;
   wire n_257_18_47;
   wire n_257_18_48;
   wire n_257_18_49;
   wire n_257_18_50;
   wire n_257_18_51;
   wire n_257_18_52;
   wire n_257_18_53;
   wire n_257_18_54;
   wire n_257_18_55;
   wire n_257_18_56;
   wire n_257_18_57;
   wire n_257_18_58;
   wire n_257_18_59;
   wire n_257_18_60;
   wire n_257_18_61;
   wire n_257_18_62;
   wire n_257_18_63;
   wire n_257_18_64;
   wire n_257_18_65;
   wire n_257_18_66;
   wire n_257_18_67;
   wire n_257_18_68;
   wire n_257_18_69;
   wire n_257_18_70;
   wire n_257_18_71;
   wire n_257_18_72;
   wire n_257_18_73;
   wire n_257_18_74;
   wire n_257_18_75;
   wire n_257_18_76;
   wire n_257_18_77;
   wire n_257_18_78;
   wire n_257_18_79;
   wire n_257_18_80;
   wire n_257_18_81;
   wire n_257_18_82;
   wire n_257_18_83;
   wire n_257_18_84;
   wire n_257_18_85;
   wire n_257_18_86;
   wire n_257_18_87;
   wire n_257_18_88;
   wire n_257_18_89;
   wire n_257_18_90;
   wire n_257_18_91;
   wire n_257_18_92;
   wire n_257_18_93;
   wire n_257_18_94;
   wire n_257_18_95;
   wire n_257_18_96;
   wire n_257_18_97;
   wire n_257_29;
   wire n_257_30;
   wire n_257_31;
   wire n_257_32;
   wire n_257_33;
   wire n_257_34;
   wire n_257_35;
   wire n_257_36;
   wire n_257_37;
   wire n_257_38;
   wire n_257_39;
   wire n_257_40;
   wire n_257_41;
   wire n_257_42;
   wire n_257_43;
   wire n_257_44;
   wire n_257_45;
   wire n_257_46;
   wire n_257_47;
   wire n_257_48;
   wire n_257_49;
   wire n_257_50;
   wire n_257_51;
   wire n_257_52;
   wire n_257_53;
   wire n_257_54;
   wire n_257_55;
   wire n_257_56;
   wire n_257_57;
   wire n_257_58;
   wire n_257_59;
   wire n_257_60;
   wire n_257_61;
   wire n_257_62;
   wire n_257_63;
   wire n_257_64;
   wire n_257_65;
   wire n_257_66;
   wire n_257_67;
   wire n_257_21_0;
   wire n_257_21_1;
   wire n_257_21_2;
   wire n_257_21_3;
   wire n_257_21_4;
   wire n_257_21_5;
   wire n_257_21_6;
   wire n_257_21_7;
   wire n_257_21_8;
   wire n_257_21_9;
   wire n_257_21_10;
   wire n_257_21_11;
   wire n_257_21_12;
   wire n_257_21_13;
   wire n_257_21_14;
   wire n_257_21_15;
   wire n_257_21_16;
   wire n_257_21_17;
   wire n_257_21_18;
   wire n_257_21_19;
   wire n_257_21_20;
   wire n_257_21_21;
   wire n_257_21_22;
   wire n_257_21_23;
   wire n_257_21_24;
   wire n_257_21_25;
   wire n_257_21_26;
   wire n_257_21_27;
   wire n_257_21_28;
   wire n_257_21_29;
   wire n_257_21_30;
   wire n_257_21_31;
   wire n_257_21_32;
   wire n_257_21_33;
   wire n_257_21_34;
   wire n_257_21_35;
   wire n_257_21_36;
   wire n_257_21_37;
   wire n_257_21_38;
   wire n_257_21_39;
   wire n_257_21_40;
   wire n_257_21_41;
   wire n_257_21_42;
   wire n_257_21_43;
   wire n_257_21_44;
   wire n_257_21_45;
   wire n_257_21_46;
   wire n_257_21_47;
   wire n_257_21_48;
   wire n_257_21_49;
   wire n_257_21_50;
   wire n_257_21_51;
   wire n_257_21_52;
   wire n_257_21_53;
   wire n_257_21_54;
   wire n_257_21_55;
   wire n_257_21_56;
   wire n_257_21_57;
   wire n_257_21_58;
   wire n_257_21_59;
   wire n_257_21_60;
   wire n_257_21_61;
   wire n_257_21_62;
   wire n_257_21_63;
   wire n_257_21_64;
   wire n_257_21_65;
   wire n_257_21_66;
   wire n_257_21_67;
   wire n_257_21_68;
   wire n_257_21_69;
   wire n_257_21_70;
   wire n_257_21_71;
   wire n_257_21_72;
   wire n_257_21_73;
   wire n_257_21_74;
   wire n_257_21_75;
   wire n_257_21_76;
   wire n_257_21_77;
   wire n_257_21_78;
   wire n_257_21_79;
   wire n_257_21_80;
   wire n_257_21_81;
   wire n_257_21_82;
   wire n_257_21_83;
   wire n_257_21_84;
   wire n_257_21_85;
   wire n_257_21_86;
   wire n_257_21_87;
   wire n_257_21_88;
   wire n_257_21_89;
   wire n_257_21_90;
   wire n_257_21_91;
   wire n_257_21_92;
   wire n_257_21_93;
   wire n_257_21_94;
   wire n_257_21_95;
   wire n_257_21_96;
   wire n_257_21_97;
   wire n_257_21_98;
   wire n_257_68;
   wire n_257_22_0;
   wire n_257_22_1;
   wire n_257_22_2;
   wire n_257_22_3;
   wire n_257_22_4;
   wire n_257_22_5;
   wire n_257_22_6;
   wire n_257_22_7;
   wire n_257_22_8;
   wire n_257_22_9;
   wire n_257_22_10;
   wire n_257_22_11;
   wire n_257_22_12;
   wire n_257_22_13;
   wire n_257_22_14;
   wire n_257_22_15;
   wire n_257_22_16;
   wire n_257_22_17;
   wire n_257_22_18;
   wire n_257_22_19;
   wire n_257_22_20;
   wire n_257_22_21;
   wire n_257_22_22;
   wire n_257_22_23;
   wire n_257_22_24;
   wire n_257_22_25;
   wire n_257_22_26;
   wire n_257_22_27;
   wire n_257_22_28;
   wire n_257_22_29;
   wire n_257_22_30;
   wire n_257_22_31;
   wire n_257_22_32;
   wire n_257_22_33;
   wire n_257_22_34;
   wire n_257_22_35;
   wire n_257_22_36;
   wire n_257_22_37;
   wire n_257_22_38;
   wire n_257_22_39;
   wire n_257_22_40;
   wire n_257_22_41;
   wire n_257_22_42;
   wire n_257_22_43;
   wire n_257_22_44;
   wire n_257_22_45;
   wire n_257_22_46;
   wire n_257_22_47;
   wire n_257_22_48;
   wire n_257_22_49;
   wire n_257_22_50;
   wire n_257_22_51;
   wire n_257_22_52;
   wire n_257_22_53;
   wire n_257_22_54;
   wire n_257_22_55;
   wire n_257_22_56;
   wire n_257_22_57;
   wire n_257_22_58;
   wire n_257_22_59;
   wire n_257_22_60;
   wire n_257_22_61;
   wire n_257_22_62;
   wire n_257_22_63;
   wire n_257_22_64;
   wire n_257_22_65;
   wire n_257_22_66;
   wire n_257_22_67;
   wire n_257_22_68;
   wire n_257_22_69;
   wire n_257_22_70;
   wire n_257_22_71;
   wire n_257_22_72;
   wire n_257_22_73;
   wire n_257_22_74;
   wire n_257_22_75;
   wire n_257_22_76;
   wire n_257_22_77;
   wire n_257_22_78;
   wire n_257_22_79;
   wire n_257_22_80;
   wire n_257_22_81;
   wire n_257_22_82;
   wire n_257_22_83;
   wire n_257_22_84;
   wire n_257_22_85;
   wire n_257_22_86;
   wire n_257_22_87;
   wire n_257_22_88;
   wire n_257_22_89;
   wire n_257_22_90;
   wire n_257_22_91;
   wire n_257_22_92;
   wire n_257_22_93;
   wire n_257_22_94;
   wire n_257_22_95;
   wire n_257_22_96;
   wire n_257_22_97;
   wire n_257_69;
   wire n_257_70;
   wire n_257_71;
   wire n_257_72;
   wire n_257_73;
   wire n_257_74;
   wire n_257_75;
   wire n_257_76;
   wire n_257_77;
   wire n_257_78;
   wire n_257_79;
   wire n_257_80;
   wire n_257_81;
   wire n_257_82;
   wire n_257_83;
   wire n_257_84;
   wire n_257_85;
   wire n_257_86;
   wire n_257_87;
   wire n_257_88;
   wire n_257_89;
   wire n_257_90;
   wire n_257_91;
   wire n_257_92;
   wire n_257_93;
   wire n_257_94;
   wire n_257_95;
   wire n_257_96;
   wire n_257_97;
   wire n_257_98;
   wire n_257_99;
   wire n_257_100;
   wire n_257_101;
   wire n_257_102;
   wire n_257_103;
   wire n_257_104;
   wire n_257_105;
   wire n_257_106;
   wire n_257_25_0;
   wire n_257_25_1;
   wire n_257_25_2;
   wire n_257_25_3;
   wire n_257_25_4;
   wire n_257_25_5;
   wire n_257_25_6;
   wire n_257_25_7;
   wire n_257_25_8;
   wire n_257_25_9;
   wire n_257_25_10;
   wire n_257_25_11;
   wire n_257_25_12;
   wire n_257_25_13;
   wire n_257_25_14;
   wire n_257_25_15;
   wire n_257_25_16;
   wire n_257_25_17;
   wire n_257_25_18;
   wire n_257_25_19;
   wire n_257_25_20;
   wire n_257_25_21;
   wire n_257_25_22;
   wire n_257_25_23;
   wire n_257_25_24;
   wire n_257_25_25;
   wire n_257_25_26;
   wire n_257_25_27;
   wire n_257_25_28;
   wire n_257_25_29;
   wire n_257_25_30;
   wire n_257_25_31;
   wire n_257_25_32;
   wire n_257_25_33;
   wire n_257_25_34;
   wire n_257_25_35;
   wire n_257_25_36;
   wire n_257_25_37;
   wire n_257_25_38;
   wire n_257_25_39;
   wire n_257_25_40;
   wire n_257_25_41;
   wire n_257_25_42;
   wire n_257_25_43;
   wire n_257_25_44;
   wire n_257_25_45;
   wire n_257_25_46;
   wire n_257_25_47;
   wire n_257_25_48;
   wire n_257_25_49;
   wire n_257_25_50;
   wire n_257_25_51;
   wire n_257_25_52;
   wire n_257_25_53;
   wire n_257_25_54;
   wire n_257_25_55;
   wire n_257_25_56;
   wire n_257_25_57;
   wire n_257_25_58;
   wire n_257_25_59;
   wire n_257_25_60;
   wire n_257_25_61;
   wire n_257_25_62;
   wire n_257_25_63;
   wire n_257_25_64;
   wire n_257_25_65;
   wire n_257_25_66;
   wire n_257_25_67;
   wire n_257_25_68;
   wire n_257_25_69;
   wire n_257_25_70;
   wire n_257_25_71;
   wire n_257_25_72;
   wire n_257_25_73;
   wire n_257_25_74;
   wire n_257_25_75;
   wire n_257_25_76;
   wire n_257_25_77;
   wire n_257_25_78;
   wire n_257_25_79;
   wire n_257_25_80;
   wire n_257_25_81;
   wire n_257_25_82;
   wire n_257_25_83;
   wire n_257_25_84;
   wire n_257_25_85;
   wire n_257_25_86;
   wire n_257_25_87;
   wire n_257_25_88;
   wire n_257_25_89;
   wire n_257_25_90;
   wire n_257_25_91;
   wire n_257_25_92;
   wire n_257_25_93;
   wire n_257_25_94;
   wire n_257_25_95;
   wire n_257_25_96;
   wire n_257_25_97;
   wire n_257_25_98;
   wire n_257_25_99;
   wire n_257_25_100;
   wire n_257_25_101;
   wire n_257_25_102;
   wire n_257_25_103;
   wire n_257_25_104;
   wire n_257_25_105;
   wire n_257_25_106;
   wire n_257_25_107;
   wire n_257_25_108;
   wire n_257_25_109;
   wire n_257_25_110;
   wire n_257_25_111;
   wire n_257_25_112;
   wire n_257_25_113;
   wire n_257_25_114;
   wire n_257_25_115;
   wire n_257_25_116;
   wire n_257_25_117;
   wire n_257_25_118;
   wire n_257_25_119;
   wire n_257_25_120;
   wire n_257_25_121;
   wire n_257_25_122;
   wire n_257_25_123;
   wire n_257_25_124;
   wire n_257_25_125;
   wire n_257_25_126;
   wire n_257_107;
   wire n_257_108;
   wire n_257_109;
   wire n_257_110;
   wire n_257_111;
   wire n_257_112;
   wire n_257_113;
   wire n_257_114;
   wire n_257_115;
   wire n_257_116;
   wire n_257_117;
   wire n_257_118;
   wire n_257_119;
   wire n_257_120;
   wire n_257_121;
   wire n_257_122;
   wire n_257_123;
   wire n_257_124;
   wire n_257_125;
   wire n_257_126;
   wire n_257_127;
   wire n_257_128;
   wire n_257_129;
   wire n_257_130;
   wire n_257_131;
   wire n_257_132;
   wire n_257_133;
   wire n_257_134;
   wire n_257_135;
   wire n_257_136;
   wire n_257_137;
   wire n_257_138;
   wire n_257_139;
   wire n_257_140;
   wire n_257_141;
   wire n_257_142;
   wire n_257_143;
   wire n_257_144;
   wire n_257_28_0;
   wire n_257_28_1;
   wire n_257_28_2;
   wire n_257_28_3;
   wire n_257_28_4;
   wire n_257_28_5;
   wire n_257_28_6;
   wire n_257_28_7;
   wire n_257_28_8;
   wire n_257_28_9;
   wire n_257_28_10;
   wire n_257_28_11;
   wire n_257_28_12;
   wire n_257_28_13;
   wire n_257_28_14;
   wire n_257_28_15;
   wire n_257_28_16;
   wire n_257_28_17;
   wire n_257_28_18;
   wire n_257_28_19;
   wire n_257_28_20;
   wire n_257_28_21;
   wire n_257_28_22;
   wire n_257_28_23;
   wire n_257_28_24;
   wire n_257_28_25;
   wire n_257_28_26;
   wire n_257_28_27;
   wire n_257_28_28;
   wire n_257_28_29;
   wire n_257_28_30;
   wire n_257_28_31;
   wire n_257_28_32;
   wire n_257_28_33;
   wire n_257_28_34;
   wire n_257_28_35;
   wire n_257_28_36;
   wire n_257_28_37;
   wire n_257_28_38;
   wire n_257_28_39;
   wire n_257_28_40;
   wire n_257_28_41;
   wire n_257_28_42;
   wire n_257_28_43;
   wire n_257_28_44;
   wire n_257_28_45;
   wire n_257_28_46;
   wire n_257_28_47;
   wire n_257_28_48;
   wire n_257_28_49;
   wire n_257_28_50;
   wire n_257_28_51;
   wire n_257_28_52;
   wire n_257_28_53;
   wire n_257_28_54;
   wire n_257_28_55;
   wire n_257_28_56;
   wire n_257_28_57;
   wire n_257_28_58;
   wire n_257_28_59;
   wire n_257_28_60;
   wire n_257_28_61;
   wire n_257_28_62;
   wire n_257_28_63;
   wire n_257_28_64;
   wire n_257_28_65;
   wire n_257_28_66;
   wire n_257_28_67;
   wire n_257_28_68;
   wire n_257_28_69;
   wire n_257_28_70;
   wire n_257_28_71;
   wire n_257_28_72;
   wire n_257_28_73;
   wire n_257_28_74;
   wire n_257_28_75;
   wire n_257_28_76;
   wire n_257_28_77;
   wire n_257_28_78;
   wire n_257_28_79;
   wire n_257_28_80;
   wire n_257_28_81;
   wire n_257_28_82;
   wire n_257_28_83;
   wire n_257_28_84;
   wire n_257_28_85;
   wire n_257_28_86;
   wire n_257_28_87;
   wire n_257_28_88;
   wire n_257_28_89;
   wire n_257_28_90;
   wire n_257_28_91;
   wire n_257_28_92;
   wire n_257_28_93;
   wire n_257_28_94;
   wire n_257_28_95;
   wire n_257_28_96;
   wire n_257_28_97;
   wire n_257_28_98;
   wire n_257_28_99;
   wire n_257_28_100;
   wire n_257_28_101;
   wire n_257_28_102;
   wire n_257_28_103;
   wire n_257_28_104;
   wire n_257_28_105;
   wire n_257_28_106;
   wire n_257_28_107;
   wire n_257_28_108;
   wire n_257_28_109;
   wire n_257_28_110;
   wire n_257_28_111;
   wire n_257_28_112;
   wire n_257_28_113;
   wire n_257_28_114;
   wire n_257_28_115;
   wire n_257_28_116;
   wire n_257_28_117;
   wire n_257_28_118;
   wire n_257_28_119;
   wire n_257_28_120;
   wire n_257_28_121;
   wire n_257_28_122;
   wire n_257_28_123;
   wire n_257_28_124;
   wire n_257_28_125;
   wire n_257_28_126;
   wire n_257_145;
   wire n_257_146;
   wire n_257_147;
   wire n_257_148;
   wire n_257_149;
   wire n_257_150;
   wire n_257_151;
   wire n_257_152;
   wire n_257_153;
   wire n_257_154;
   wire n_257_155;
   wire n_257_156;
   wire n_257_157;
   wire n_257_158;
   wire n_257_159;
   wire n_257_160;
   wire n_257_161;
   wire n_257_162;
   wire n_257_163;
   wire n_257_164;
   wire n_257_165;
   wire n_257_166;
   wire n_257_167;
   wire n_257_168;
   wire n_257_169;
   wire n_257_170;
   wire n_257_171;
   wire n_257_172;
   wire n_257_173;
   wire n_257_174;
   wire n_257_175;
   wire n_257_176;
   wire n_257_177;
   wire n_257_178;
   wire n_257_179;
   wire n_257_180;
   wire n_257_181;
   wire n_257_182;
   wire n_257_183;
   wire n_257_184;
   wire n_257_31_0;
   wire n_257_31_1;
   wire n_257_31_2;
   wire n_257_31_3;
   wire n_257_31_4;
   wire n_257_31_5;
   wire n_257_31_6;
   wire n_257_31_7;
   wire n_257_31_8;
   wire n_257_31_9;
   wire n_257_31_10;
   wire n_257_31_11;
   wire n_257_31_12;
   wire n_257_31_13;
   wire n_257_31_14;
   wire n_257_31_15;
   wire n_257_31_16;
   wire n_257_31_17;
   wire n_257_31_18;
   wire n_257_31_19;
   wire n_257_31_20;
   wire n_257_31_21;
   wire n_257_31_22;
   wire n_257_31_23;
   wire n_257_31_24;
   wire n_257_31_25;
   wire n_257_31_26;
   wire n_257_31_27;
   wire n_257_31_28;
   wire n_257_31_29;
   wire n_257_31_30;
   wire n_257_31_31;
   wire n_257_31_32;
   wire n_257_31_33;
   wire n_257_31_34;
   wire n_257_31_35;
   wire n_257_31_36;
   wire n_257_31_37;
   wire n_257_31_38;
   wire n_257_31_39;
   wire n_257_31_40;
   wire n_257_31_41;
   wire n_257_31_42;
   wire n_257_31_43;
   wire n_257_31_44;
   wire n_257_31_45;
   wire n_257_31_46;
   wire n_257_31_47;
   wire n_257_31_48;
   wire n_257_31_49;
   wire n_257_31_50;
   wire n_257_31_51;
   wire n_257_31_52;
   wire n_257_31_53;
   wire n_257_31_54;
   wire n_257_31_55;
   wire n_257_31_56;
   wire n_257_31_57;
   wire n_257_31_58;
   wire n_257_31_59;
   wire n_257_31_60;
   wire n_257_31_61;
   wire n_257_31_62;
   wire n_257_31_63;
   wire n_257_31_64;
   wire n_257_31_65;
   wire n_257_31_66;
   wire n_257_31_67;
   wire n_257_31_68;
   wire n_257_31_69;
   wire n_257_31_70;
   wire n_257_31_71;
   wire n_257_31_72;
   wire n_257_31_73;
   wire n_257_31_74;
   wire n_257_31_75;
   wire n_257_31_76;
   wire n_257_31_77;
   wire n_257_31_78;
   wire n_257_31_79;
   wire n_257_31_80;
   wire n_257_31_81;
   wire n_257_31_82;
   wire n_257_31_83;
   wire n_257_31_84;
   wire n_257_31_85;
   wire n_257_31_86;
   wire n_257_31_87;
   wire n_257_31_88;
   wire n_257_32_0;
   wire n_257_32_1;
   wire n_257_32_2;
   wire n_257_32_3;
   wire n_257_32_4;
   wire n_257_32_5;
   wire n_257_32_6;
   wire n_257_32_7;
   wire n_257_32_8;
   wire n_257_32_9;
   wire n_257_32_10;
   wire n_257_32_11;
   wire n_257_32_12;
   wire n_257_32_13;
   wire n_257_32_14;
   wire n_257_32_15;
   wire n_257_32_16;
   wire n_257_32_17;
   wire n_257_32_18;
   wire n_257_32_19;
   wire n_257_32_20;
   wire n_257_32_21;
   wire n_257_32_22;
   wire n_257_32_23;
   wire n_257_32_24;
   wire n_257_32_25;
   wire n_257_32_26;
   wire n_257_32_27;
   wire n_257_32_28;
   wire n_257_32_29;
   wire n_257_32_30;
   wire n_257_32_31;
   wire n_257_32_32;
   wire n_257_32_33;
   wire n_257_32_34;
   wire n_257_32_35;
   wire n_257_32_36;
   wire n_257_32_37;
   wire n_257_32_38;
   wire n_257_32_39;
   wire n_257_32_40;
   wire n_257_32_41;
   wire n_257_32_42;
   wire n_257_32_43;
   wire n_257_32_44;
   wire n_257_32_45;
   wire n_257_32_46;
   wire n_257_32_47;
   wire n_257_32_48;
   wire n_257_32_49;
   wire n_257_32_50;
   wire n_257_32_51;
   wire n_257_32_52;
   wire n_257_32_53;
   wire n_257_32_54;
   wire n_257_32_55;
   wire n_257_32_56;
   wire n_257_32_57;
   wire n_257_32_58;
   wire n_257_32_59;
   wire n_257_32_60;
   wire n_257_32_61;
   wire n_257_32_62;
   wire n_257_32_63;
   wire n_257_32_64;
   wire n_257_32_65;
   wire n_257_32_66;
   wire n_257_32_67;
   wire n_257_32_68;
   wire n_257_32_69;
   wire n_257_32_70;
   wire n_257_32_71;
   wire n_257_32_72;
   wire n_257_32_73;
   wire n_257_32_74;
   wire n_257_32_75;
   wire n_257_32_76;
   wire n_257_32_77;
   wire n_257_32_78;
   wire n_257_32_79;
   wire n_257_32_80;
   wire n_257_32_81;
   wire n_257_32_82;
   wire n_257_32_83;
   wire n_257_32_84;
   wire n_257_32_85;
   wire n_257_32_86;
   wire n_257_32_87;
   wire n_257_32_88;
   wire n_257_32_89;
   wire n_257_32_90;
   wire n_257_32_91;
   wire n_257_32_92;
   wire n_257_32_93;
   wire n_257_32_94;
   wire n_257_32_95;
   wire n_257_32_96;
   wire n_257_32_97;
   wire n_257_32_98;
   wire n_257_32_99;
   wire n_257_32_100;
   wire n_257_32_101;
   wire n_257_32_102;
   wire n_257_32_103;
   wire n_257_32_104;
   wire n_257_32_105;
   wire n_257_32_106;
   wire n_257_32_107;
   wire n_257_32_108;
   wire n_257_32_109;
   wire n_257_32_110;
   wire n_257_32_111;
   wire n_257_32_112;
   wire n_257_32_113;
   wire n_257_32_114;
   wire n_257_32_115;
   wire n_257_32_116;
   wire n_257_32_117;
   wire n_257_32_118;
   wire n_257_32_119;
   wire n_257_32_120;
   wire n_257_32_121;
   wire n_257_32_122;
   wire n_257_32_123;
   wire n_257_32_124;
   wire n_257_32_125;
   wire n_257_32_126;
   wire n_257_185;
   wire n_257_186;
   wire n_257_187;
   wire n_257_188;
   wire n_257_189;
   wire n_257_190;
   wire n_257_191;
   wire n_257_192;
   wire n_257_193;
   wire n_257_194;
   wire n_257_195;
   wire n_257_196;
   wire n_257_197;
   wire n_257_198;
   wire n_257_199;
   wire n_257_200;
   wire n_257_201;
   wire n_257_202;
   wire n_257_203;
   wire n_257_204;
   wire n_257_205;
   wire n_257_206;
   wire n_257_207;
   wire n_257_208;
   wire n_257_209;
   wire n_257_210;
   wire n_257_211;
   wire n_257_212;
   wire n_257_213;
   wire n_257_214;
   wire n_257_215;
   wire n_257_216;
   wire n_257_217;
   wire n_257_218;
   wire n_257_219;
   wire n_257_220;
   wire n_257_221;
   wire n_257_222;
   wire n_257_223;
   wire n_257_35_0;
   wire n_257_35_1;
   wire n_257_35_2;
   wire n_257_35_3;
   wire n_257_35_4;
   wire n_257_35_5;
   wire n_257_35_6;
   wire n_257_35_7;
   wire n_257_35_8;
   wire n_257_35_9;
   wire n_257_35_10;
   wire n_257_35_11;
   wire n_257_35_12;
   wire n_257_35_13;
   wire n_257_35_14;
   wire n_257_35_15;
   wire n_257_35_16;
   wire n_257_35_17;
   wire n_257_35_18;
   wire n_257_35_19;
   wire n_257_35_20;
   wire n_257_35_21;
   wire n_257_35_22;
   wire n_257_35_23;
   wire n_257_35_24;
   wire n_257_35_25;
   wire n_257_35_26;
   wire n_257_35_27;
   wire n_257_35_28;
   wire n_257_35_29;
   wire n_257_35_30;
   wire n_257_35_31;
   wire n_257_35_32;
   wire n_257_35_33;
   wire n_257_35_34;
   wire n_257_35_35;
   wire n_257_35_36;
   wire n_257_35_37;
   wire n_257_35_38;
   wire n_257_35_39;
   wire n_257_35_40;
   wire n_257_35_41;
   wire n_257_35_42;
   wire n_257_35_43;
   wire n_257_35_44;
   wire n_257_35_45;
   wire n_257_35_46;
   wire n_257_35_47;
   wire n_257_35_48;
   wire n_257_35_49;
   wire n_257_35_50;
   wire n_257_35_51;
   wire n_257_35_52;
   wire n_257_35_53;
   wire n_257_35_54;
   wire n_257_35_55;
   wire n_257_35_56;
   wire n_257_35_57;
   wire n_257_35_58;
   wire n_257_35_59;
   wire n_257_35_60;
   wire n_257_35_61;
   wire n_257_35_62;
   wire n_257_35_63;
   wire n_257_35_64;
   wire n_257_35_65;
   wire n_257_35_66;
   wire n_257_35_67;
   wire n_257_35_68;
   wire n_257_35_69;
   wire n_257_35_70;
   wire n_257_35_71;
   wire n_257_35_72;
   wire n_257_35_73;
   wire n_257_35_74;
   wire n_257_35_75;
   wire n_257_35_76;
   wire n_257_35_77;
   wire n_257_35_78;
   wire n_257_35_79;
   wire n_257_35_80;
   wire n_257_35_81;
   wire n_257_35_82;
   wire n_257_35_83;
   wire n_257_35_84;
   wire n_257_35_85;
   wire n_257_35_86;
   wire n_257_35_87;
   wire n_257_35_88;
   wire n_257_35_89;
   wire n_257_35_90;
   wire n_257_35_91;
   wire n_257_35_92;
   wire n_257_35_93;
   wire n_257_35_94;
   wire n_257_35_95;
   wire n_257_35_96;
   wire n_257_35_97;
   wire n_257_35_98;
   wire n_257_35_99;
   wire n_257_35_100;
   wire n_257_35_101;
   wire n_257_35_102;
   wire n_257_35_103;
   wire n_257_35_104;
   wire n_257_35_105;
   wire n_257_35_106;
   wire n_257_35_107;
   wire n_257_35_108;
   wire n_257_35_109;
   wire n_257_35_110;
   wire n_257_35_111;
   wire n_257_35_112;
   wire n_257_35_113;
   wire n_257_35_114;
   wire n_257_35_115;
   wire n_257_35_116;
   wire n_257_35_117;
   wire n_257_35_118;
   wire n_257_35_119;
   wire n_257_35_120;
   wire n_257_35_121;
   wire n_257_35_122;
   wire n_257_35_123;
   wire n_257_35_124;
   wire n_257_35_125;
   wire n_257_35_126;
   wire n_257_224;
   wire n_257_36_0;
   wire n_257_36_1;
   wire n_257_36_2;
   wire n_257_36_3;
   wire n_257_36_4;
   wire n_257_36_5;
   wire n_257_36_6;
   wire n_257_36_7;
   wire n_257_36_8;
   wire n_257_36_9;
   wire n_257_36_10;
   wire n_257_36_11;
   wire n_257_36_12;
   wire n_257_36_13;
   wire n_257_36_14;
   wire n_257_36_15;
   wire n_257_36_16;
   wire n_257_36_17;
   wire n_257_36_18;
   wire n_257_36_19;
   wire n_257_36_20;
   wire n_257_36_21;
   wire n_257_36_22;
   wire n_257_36_23;
   wire n_257_36_24;
   wire n_257_36_25;
   wire n_257_36_26;
   wire n_257_36_27;
   wire n_257_36_28;
   wire n_257_36_29;
   wire n_257_36_30;
   wire n_257_36_31;
   wire n_257_36_32;
   wire n_257_36_33;
   wire n_257_36_34;
   wire n_257_36_35;
   wire n_257_36_36;
   wire n_257_36_37;
   wire n_257_36_38;
   wire n_257_36_39;
   wire n_257_36_40;
   wire n_257_36_41;
   wire n_257_36_42;
   wire n_257_36_43;
   wire n_257_36_44;
   wire n_257_36_45;
   wire n_257_36_46;
   wire n_257_36_47;
   wire n_257_36_48;
   wire n_257_36_49;
   wire n_257_36_50;
   wire n_257_36_51;
   wire n_257_36_52;
   wire n_257_36_53;
   wire n_257_36_54;
   wire n_257_36_55;
   wire n_257_36_56;
   wire n_257_36_57;
   wire n_257_36_58;
   wire n_257_36_59;
   wire n_257_36_60;
   wire n_257_36_61;
   wire n_257_36_62;
   wire n_257_36_63;
   wire n_257_36_64;
   wire n_257_36_65;
   wire n_257_36_66;
   wire n_257_36_67;
   wire n_257_36_68;
   wire n_257_36_69;
   wire n_257_36_70;
   wire n_257_36_71;
   wire n_257_36_72;
   wire n_257_36_73;
   wire n_257_36_74;
   wire n_257_36_75;
   wire n_257_36_76;
   wire n_257_36_77;
   wire n_257_36_78;
   wire n_257_36_79;
   wire n_257_36_80;
   wire n_257_36_81;
   wire n_257_36_82;
   wire n_257_36_83;
   wire n_257_36_84;
   wire n_257_36_85;
   wire n_257_36_86;
   wire n_257_36_87;
   wire n_257_36_88;
   wire n_257_36_89;
   wire n_257_36_90;
   wire n_257_36_91;
   wire n_257_36_92;
   wire n_257_36_93;
   wire n_257_36_94;
   wire n_257_36_95;
   wire n_257_36_96;
   wire n_257_36_97;
   wire n_257_36_98;
   wire n_257_36_99;
   wire n_257_36_100;
   wire n_257_36_101;
   wire n_257_36_102;
   wire n_257_36_103;
   wire n_257_36_104;
   wire n_257_36_105;
   wire n_257_36_106;
   wire n_257_36_107;
   wire n_257_36_108;
   wire n_257_36_109;
   wire n_257_36_110;
   wire n_257_36_111;
   wire n_257_36_112;
   wire n_257_36_113;
   wire n_257_36_114;
   wire n_257_36_115;
   wire n_257_36_116;
   wire n_257_36_117;
   wire n_257_36_118;
   wire n_257_36_119;
   wire n_257_36_120;
   wire n_257_36_121;
   wire n_257_36_122;
   wire n_257_36_123;
   wire n_257_36_124;
   wire n_257_36_125;
   wire n_257_36_126;
   wire n_257_225;
   wire n_257_226;
   wire n_257_227;
   wire n_257_228;
   wire n_257_229;
   wire n_257_230;
   wire n_257_231;
   wire n_257_232;
   wire n_257_233;
   wire n_257_234;
   wire n_257_235;
   wire n_257_236;
   wire n_257_237;
   wire n_257_238;
   wire n_257_239;
   wire n_257_240;
   wire n_257_241;
   wire n_257_242;
   wire n_257_243;
   wire n_257_244;
   wire n_257_245;
   wire n_257_246;
   wire n_257_247;
   wire n_257_248;
   wire n_257_249;
   wire n_257_250;
   wire n_257_251;
   wire n_257_252;
   wire n_257_253;
   wire n_257_254;
   wire n_257_255;
   wire n_257_256;
   wire n_257_257;
   wire n_257_258;
   wire n_257_259;
   wire n_257_260;
   wire n_257_261;
   wire n_257_262;
   wire n_257_263;
   wire n_257_39_0;
   wire n_257_39_1;
   wire n_257_39_2;
   wire n_257_39_3;
   wire n_257_39_4;
   wire n_257_39_5;
   wire n_257_39_6;
   wire n_257_39_7;
   wire n_257_39_8;
   wire n_257_39_9;
   wire n_257_39_10;
   wire n_257_39_11;
   wire n_257_39_12;
   wire n_257_39_13;
   wire n_257_39_14;
   wire n_257_39_15;
   wire n_257_39_16;
   wire n_257_39_17;
   wire n_257_39_18;
   wire n_257_39_19;
   wire n_257_39_20;
   wire n_257_39_21;
   wire n_257_39_22;
   wire n_257_39_23;
   wire n_257_39_24;
   wire n_257_39_25;
   wire n_257_39_26;
   wire n_257_39_27;
   wire n_257_39_28;
   wire n_257_39_29;
   wire n_257_39_30;
   wire n_257_39_31;
   wire n_257_39_32;
   wire n_257_39_33;
   wire n_257_39_34;
   wire n_257_39_35;
   wire n_257_39_36;
   wire n_257_39_37;
   wire n_257_39_38;
   wire n_257_39_39;
   wire n_257_39_40;
   wire n_257_39_41;
   wire n_257_39_42;
   wire n_257_39_43;
   wire n_257_39_44;
   wire n_257_39_45;
   wire n_257_39_46;
   wire n_257_39_47;
   wire n_257_39_48;
   wire n_257_39_49;
   wire n_257_39_50;
   wire n_257_39_51;
   wire n_257_39_52;
   wire n_257_39_53;
   wire n_257_39_54;
   wire n_257_39_55;
   wire n_257_39_56;
   wire n_257_39_57;
   wire n_257_39_58;
   wire n_257_39_59;
   wire n_257_39_60;
   wire n_257_39_61;
   wire n_257_39_62;
   wire n_257_39_63;
   wire n_257_39_64;
   wire n_257_39_65;
   wire n_257_39_66;
   wire n_257_39_67;
   wire n_257_39_68;
   wire n_257_39_69;
   wire n_257_39_70;
   wire n_257_39_71;
   wire n_257_39_72;
   wire n_257_39_73;
   wire n_257_39_74;
   wire n_257_39_75;
   wire n_257_39_76;
   wire n_257_39_77;
   wire n_257_39_78;
   wire n_257_39_79;
   wire n_257_39_80;
   wire n_257_39_81;
   wire n_257_39_82;
   wire n_257_39_83;
   wire n_257_39_84;
   wire n_257_39_85;
   wire n_257_39_86;
   wire n_257_39_87;
   wire n_257_39_88;
   wire n_257_39_89;
   wire n_257_39_90;
   wire n_257_39_91;
   wire n_257_39_92;
   wire n_257_39_93;
   wire n_257_39_94;
   wire n_257_39_95;
   wire n_257_39_96;
   wire n_257_39_97;
   wire n_257_39_98;
   wire n_257_39_99;
   wire n_257_39_100;
   wire n_257_39_101;
   wire n_257_39_102;
   wire n_257_39_103;
   wire n_257_39_104;
   wire n_257_39_105;
   wire n_257_39_106;
   wire n_257_39_107;
   wire n_257_39_108;
   wire n_257_39_109;
   wire n_257_39_110;
   wire n_257_39_111;
   wire n_257_39_112;
   wire n_257_39_113;
   wire n_257_39_114;
   wire n_257_39_115;
   wire n_257_39_116;
   wire n_257_39_117;
   wire n_257_39_118;
   wire n_257_39_119;
   wire n_257_39_120;
   wire n_257_39_121;
   wire n_257_39_122;
   wire n_257_39_123;
   wire n_257_39_124;
   wire n_257_39_125;
   wire n_257_39_126;
   wire n_257_264;
   wire n_257_40_0;
   wire n_257_40_1;
   wire n_257_40_2;
   wire n_257_40_3;
   wire n_257_40_4;
   wire n_257_40_5;
   wire n_257_40_6;
   wire n_257_40_7;
   wire n_257_40_8;
   wire n_257_40_9;
   wire n_257_40_10;
   wire n_257_40_11;
   wire n_257_40_12;
   wire n_257_40_13;
   wire n_257_40_14;
   wire n_257_40_15;
   wire n_257_40_16;
   wire n_257_40_17;
   wire n_257_40_18;
   wire n_257_40_19;
   wire n_257_40_20;
   wire n_257_40_21;
   wire n_257_40_22;
   wire n_257_40_23;
   wire n_257_40_24;
   wire n_257_40_25;
   wire n_257_40_26;
   wire n_257_40_27;
   wire n_257_40_28;
   wire n_257_40_29;
   wire n_257_40_30;
   wire n_257_40_31;
   wire n_257_40_32;
   wire n_257_40_33;
   wire n_257_40_34;
   wire n_257_40_35;
   wire n_257_40_36;
   wire n_257_40_37;
   wire n_257_40_38;
   wire n_257_40_39;
   wire n_257_40_40;
   wire n_257_40_41;
   wire n_257_40_42;
   wire n_257_40_43;
   wire n_257_40_44;
   wire n_257_40_45;
   wire n_257_40_46;
   wire n_257_40_47;
   wire n_257_40_48;
   wire n_257_40_49;
   wire n_257_40_50;
   wire n_257_40_51;
   wire n_257_40_52;
   wire n_257_40_53;
   wire n_257_40_54;
   wire n_257_40_55;
   wire n_257_40_56;
   wire n_257_40_57;
   wire n_257_40_58;
   wire n_257_40_59;
   wire n_257_40_60;
   wire n_257_40_61;
   wire n_257_40_62;
   wire n_257_40_63;
   wire n_257_40_64;
   wire n_257_40_65;
   wire n_257_40_66;
   wire n_257_40_67;
   wire n_257_40_68;
   wire n_257_40_69;
   wire n_257_40_70;
   wire n_257_40_71;
   wire n_257_40_72;
   wire n_257_40_73;
   wire n_257_40_74;
   wire n_257_40_75;
   wire n_257_40_76;
   wire n_257_40_77;
   wire n_257_40_78;
   wire n_257_40_79;
   wire n_257_40_80;
   wire n_257_40_81;
   wire n_257_40_82;
   wire n_257_40_83;
   wire n_257_40_84;
   wire n_257_40_85;
   wire n_257_40_86;
   wire n_257_40_87;
   wire n_257_40_88;
   wire n_257_40_89;
   wire n_257_40_90;
   wire n_257_40_91;
   wire n_257_40_92;
   wire n_257_40_93;
   wire n_257_40_94;
   wire n_257_40_95;
   wire n_257_40_96;
   wire n_257_40_97;
   wire n_257_40_98;
   wire n_257_40_99;
   wire n_257_40_100;
   wire n_257_40_101;
   wire n_257_40_102;
   wire n_257_40_103;
   wire n_257_40_104;
   wire n_257_40_105;
   wire n_257_40_106;
   wire n_257_40_107;
   wire n_257_40_108;
   wire n_257_40_109;
   wire n_257_40_110;
   wire n_257_40_111;
   wire n_257_40_112;
   wire n_257_40_113;
   wire n_257_40_114;
   wire n_257_40_115;
   wire n_257_40_116;
   wire n_257_40_117;
   wire n_257_40_118;
   wire n_257_40_119;
   wire n_257_40_120;
   wire n_257_40_121;
   wire n_257_40_122;
   wire n_257_40_123;
   wire n_257_40_124;
   wire n_257_40_125;
   wire n_257_40_126;
   wire n_257_265;
   wire n_257_266;
   wire n_257_267;
   wire n_257_268;
   wire n_257_269;
   wire n_257_270;
   wire n_257_271;
   wire n_257_272;
   wire n_257_273;
   wire n_257_274;
   wire n_257_275;
   wire n_257_276;
   wire n_257_277;
   wire n_257_278;
   wire n_257_279;
   wire n_257_280;
   wire n_257_281;
   wire n_257_282;
   wire n_257_283;
   wire n_257_284;
   wire n_257_285;
   wire n_257_286;
   wire n_257_287;
   wire n_257_288;
   wire n_257_289;
   wire n_257_290;
   wire n_257_291;
   wire n_257_292;
   wire n_257_293;
   wire n_257_294;
   wire n_257_295;
   wire n_257_296;
   wire n_257_297;
   wire n_257_298;
   wire n_257_299;
   wire n_257_300;
   wire n_257_301;
   wire n_257_302;
   wire n_257_303;
   wire n_257_43_0;
   wire n_257_43_1;
   wire n_257_43_2;
   wire n_257_43_3;
   wire n_257_43_4;
   wire n_257_43_5;
   wire n_257_43_6;
   wire n_257_43_7;
   wire n_257_43_8;
   wire n_257_43_9;
   wire n_257_43_10;
   wire n_257_43_11;
   wire n_257_43_12;
   wire n_257_43_13;
   wire n_257_43_14;
   wire n_257_43_15;
   wire n_257_43_16;
   wire n_257_43_17;
   wire n_257_43_18;
   wire n_257_43_19;
   wire n_257_43_20;
   wire n_257_43_21;
   wire n_257_43_22;
   wire n_257_43_23;
   wire n_257_43_24;
   wire n_257_43_25;
   wire n_257_43_26;
   wire n_257_43_27;
   wire n_257_43_28;
   wire n_257_43_29;
   wire n_257_43_30;
   wire n_257_43_31;
   wire n_257_43_32;
   wire n_257_43_33;
   wire n_257_43_34;
   wire n_257_43_35;
   wire n_257_43_36;
   wire n_257_43_37;
   wire n_257_43_38;
   wire n_257_43_39;
   wire n_257_43_40;
   wire n_257_43_41;
   wire n_257_43_42;
   wire n_257_43_43;
   wire n_257_43_44;
   wire n_257_43_45;
   wire n_257_43_46;
   wire n_257_43_47;
   wire n_257_43_48;
   wire n_257_43_49;
   wire n_257_43_50;
   wire n_257_43_51;
   wire n_257_43_52;
   wire n_257_43_53;
   wire n_257_43_54;
   wire n_257_43_55;
   wire n_257_43_56;
   wire n_257_43_57;
   wire n_257_43_58;
   wire n_257_43_59;
   wire n_257_43_60;
   wire n_257_43_61;
   wire n_257_43_62;
   wire n_257_43_63;
   wire n_257_43_64;
   wire n_257_43_65;
   wire n_257_43_66;
   wire n_257_43_67;
   wire n_257_43_68;
   wire n_257_43_69;
   wire n_257_43_70;
   wire n_257_43_71;
   wire n_257_43_72;
   wire n_257_43_73;
   wire n_257_43_74;
   wire n_257_43_75;
   wire n_257_43_76;
   wire n_257_43_77;
   wire n_257_43_78;
   wire n_257_43_79;
   wire n_257_43_80;
   wire n_257_43_81;
   wire n_257_43_82;
   wire n_257_43_83;
   wire n_257_43_84;
   wire n_257_43_85;
   wire n_257_43_86;
   wire n_257_43_87;
   wire n_257_43_88;
   wire n_257_43_89;
   wire n_257_43_90;
   wire n_257_43_91;
   wire n_257_43_92;
   wire n_257_43_93;
   wire n_257_43_94;
   wire n_257_43_95;
   wire n_257_43_96;
   wire n_257_43_97;
   wire n_257_43_98;
   wire n_257_43_99;
   wire n_257_43_100;
   wire n_257_43_101;
   wire n_257_43_102;
   wire n_257_43_103;
   wire n_257_43_104;
   wire n_257_43_105;
   wire n_257_43_106;
   wire n_257_43_107;
   wire n_257_43_108;
   wire n_257_43_109;
   wire n_257_43_110;
   wire n_257_43_111;
   wire n_257_43_112;
   wire n_257_43_113;
   wire n_257_43_114;
   wire n_257_43_115;
   wire n_257_43_116;
   wire n_257_43_117;
   wire n_257_43_118;
   wire n_257_43_119;
   wire n_257_43_120;
   wire n_257_43_121;
   wire n_257_43_122;
   wire n_257_43_123;
   wire n_257_43_124;
   wire n_257_43_125;
   wire n_257_43_126;
   wire n_257_304;
   wire n_257_305;
   wire n_257_306;
   wire n_257_307;
   wire n_257_308;
   wire n_257_309;
   wire n_257_310;
   wire n_257_311;
   wire n_257_312;
   wire n_257_313;
   wire n_257_314;
   wire n_257_315;
   wire n_257_316;
   wire n_257_317;
   wire n_257_318;
   wire n_257_319;
   wire n_257_320;
   wire n_257_321;
   wire n_257_322;
   wire n_257_323;
   wire n_257_324;
   wire n_257_325;
   wire n_257_326;
   wire n_257_327;
   wire n_257_328;
   wire n_257_329;
   wire n_257_330;
   wire n_257_331;
   wire n_257_332;
   wire n_257_333;
   wire n_257_334;
   wire n_257_335;
   wire n_257_336;
   wire n_257_337;
   wire n_257_338;
   wire n_257_339;
   wire n_257_340;
   wire n_257_341;
   wire n_257_342;
   wire n_257_46_0;
   wire n_257_46_1;
   wire n_257_46_2;
   wire n_257_46_3;
   wire n_257_46_4;
   wire n_257_46_5;
   wire n_257_46_6;
   wire n_257_46_7;
   wire n_257_46_8;
   wire n_257_46_9;
   wire n_257_46_10;
   wire n_257_46_11;
   wire n_257_46_12;
   wire n_257_46_13;
   wire n_257_46_14;
   wire n_257_46_15;
   wire n_257_46_16;
   wire n_257_46_17;
   wire n_257_46_18;
   wire n_257_46_19;
   wire n_257_46_20;
   wire n_257_46_21;
   wire n_257_46_22;
   wire n_257_46_23;
   wire n_257_46_24;
   wire n_257_46_25;
   wire n_257_46_26;
   wire n_257_46_27;
   wire n_257_46_28;
   wire n_257_46_29;
   wire n_257_46_30;
   wire n_257_46_31;
   wire n_257_46_32;
   wire n_257_46_33;
   wire n_257_46_34;
   wire n_257_46_35;
   wire n_257_46_36;
   wire n_257_46_37;
   wire n_257_46_38;
   wire n_257_46_39;
   wire n_257_46_40;
   wire n_257_46_41;
   wire n_257_46_42;
   wire n_257_46_43;
   wire n_257_46_44;
   wire n_257_46_45;
   wire n_257_46_46;
   wire n_257_46_47;
   wire n_257_46_48;
   wire n_257_46_49;
   wire n_257_46_50;
   wire n_257_46_51;
   wire n_257_46_52;
   wire n_257_46_53;
   wire n_257_46_54;
   wire n_257_46_55;
   wire n_257_46_56;
   wire n_257_46_57;
   wire n_257_46_58;
   wire n_257_46_59;
   wire n_257_46_60;
   wire n_257_46_61;
   wire n_257_46_62;
   wire n_257_46_63;
   wire n_257_46_64;
   wire n_257_46_65;
   wire n_257_46_66;
   wire n_257_46_67;
   wire n_257_46_68;
   wire n_257_46_69;
   wire n_257_46_70;
   wire n_257_46_71;
   wire n_257_46_72;
   wire n_257_46_73;
   wire n_257_46_74;
   wire n_257_46_75;
   wire n_257_46_76;
   wire n_257_46_77;
   wire n_257_46_78;
   wire n_257_46_79;
   wire n_257_46_80;
   wire n_257_46_81;
   wire n_257_46_82;
   wire n_257_46_83;
   wire n_257_46_84;
   wire n_257_46_85;
   wire n_257_46_86;
   wire n_257_46_87;
   wire n_257_46_88;
   wire n_257_46_89;
   wire n_257_46_90;
   wire n_257_46_91;
   wire n_257_46_92;
   wire n_257_46_93;
   wire n_257_46_94;
   wire n_257_46_95;
   wire n_257_46_96;
   wire n_257_46_97;
   wire n_257_343;
   wire n_257_344;
   wire n_257_345;
   wire n_257_346;
   wire n_257_347;
   wire n_257_348;
   wire n_257_349;
   wire n_257_350;
   wire n_257_351;
   wire n_257_352;
   wire n_257_353;
   wire n_257_354;
   wire n_257_355;
   wire n_257_356;
   wire n_257_357;
   wire n_257_358;
   wire n_257_359;
   wire n_257_360;
   wire n_257_361;
   wire n_257_362;
   wire n_257_363;
   wire n_257_364;
   wire n_257_365;
   wire n_257_366;
   wire n_257_367;
   wire n_257_368;
   wire n_257_369;
   wire n_257_370;
   wire n_257_371;
   wire n_257_372;
   wire n_257_373;
   wire n_257_374;
   wire n_257_375;
   wire n_257_376;
   wire n_257_377;
   wire n_257_378;
   wire n_257_379;
   wire n_257_380;
   wire n_257_381;
   wire n_257_49_0;
   wire n_257_49_1;
   wire n_257_49_2;
   wire n_257_49_3;
   wire n_257_49_4;
   wire n_257_49_5;
   wire n_257_49_6;
   wire n_257_49_7;
   wire n_257_49_8;
   wire n_257_49_9;
   wire n_257_49_10;
   wire n_257_49_11;
   wire n_257_49_12;
   wire n_257_49_13;
   wire n_257_49_14;
   wire n_257_49_15;
   wire n_257_49_16;
   wire n_257_49_17;
   wire n_257_49_18;
   wire n_257_49_19;
   wire n_257_49_20;
   wire n_257_49_21;
   wire n_257_49_22;
   wire n_257_49_23;
   wire n_257_49_24;
   wire n_257_49_25;
   wire n_257_49_26;
   wire n_257_49_27;
   wire n_257_49_28;
   wire n_257_49_29;
   wire n_257_49_30;
   wire n_257_49_31;
   wire n_257_49_32;
   wire n_257_49_33;
   wire n_257_49_34;
   wire n_257_49_35;
   wire n_257_49_36;
   wire n_257_49_37;
   wire n_257_49_38;
   wire n_257_49_39;
   wire n_257_49_40;
   wire n_257_49_41;
   wire n_257_49_42;
   wire n_257_49_43;
   wire n_257_49_44;
   wire n_257_49_45;
   wire n_257_49_46;
   wire n_257_49_47;
   wire n_257_49_48;
   wire n_257_49_49;
   wire n_257_49_50;
   wire n_257_49_51;
   wire n_257_49_52;
   wire n_257_49_53;
   wire n_257_49_54;
   wire n_257_49_55;
   wire n_257_49_56;
   wire n_257_49_57;
   wire n_257_49_58;
   wire n_257_49_59;
   wire n_257_49_60;
   wire n_257_49_61;
   wire n_257_49_62;
   wire n_257_49_63;
   wire n_257_49_64;
   wire n_257_49_65;
   wire n_257_49_66;
   wire n_257_49_67;
   wire n_257_49_68;
   wire n_257_49_69;
   wire n_257_49_70;
   wire n_257_49_71;
   wire n_257_49_72;
   wire n_257_49_73;
   wire n_257_49_74;
   wire n_257_49_75;
   wire n_257_49_76;
   wire n_257_49_77;
   wire n_257_49_78;
   wire n_257_49_79;
   wire n_257_49_80;
   wire n_257_49_81;
   wire n_257_49_82;
   wire n_257_49_83;
   wire n_257_49_84;
   wire n_257_49_85;
   wire n_257_49_86;
   wire n_257_49_87;
   wire n_257_49_88;
   wire n_257_49_89;
   wire n_257_49_90;
   wire n_257_49_91;
   wire n_257_49_92;
   wire n_257_49_93;
   wire n_257_49_94;
   wire n_257_49_95;
   wire n_257_49_96;
   wire n_257_49_97;
   wire n_257_49_98;
   wire n_257_50_0;
   wire n_257_50_1;
   wire n_257_50_2;
   wire n_257_50_3;
   wire n_257_50_4;
   wire n_257_50_5;
   wire n_257_50_6;
   wire n_257_50_7;
   wire n_257_50_8;
   wire n_257_50_9;
   wire n_257_50_10;
   wire n_257_50_11;
   wire n_257_50_12;
   wire n_257_50_13;
   wire n_257_50_14;
   wire n_257_50_15;
   wire n_257_50_16;
   wire n_257_50_17;
   wire n_257_50_18;
   wire n_257_50_19;
   wire n_257_50_20;
   wire n_257_50_21;
   wire n_257_50_22;
   wire n_257_50_23;
   wire n_257_50_24;
   wire n_257_50_25;
   wire n_257_50_26;
   wire n_257_50_27;
   wire n_257_50_28;
   wire n_257_50_29;
   wire n_257_50_30;
   wire n_257_50_31;
   wire n_257_50_32;
   wire n_257_50_33;
   wire n_257_50_34;
   wire n_257_50_35;
   wire n_257_50_36;
   wire n_257_50_37;
   wire n_257_50_38;
   wire n_257_50_39;
   wire n_257_50_40;
   wire n_257_50_41;
   wire n_257_50_42;
   wire n_257_50_43;
   wire n_257_50_44;
   wire n_257_50_45;
   wire n_257_50_46;
   wire n_257_50_47;
   wire n_257_50_48;
   wire n_257_50_49;
   wire n_257_50_50;
   wire n_257_50_51;
   wire n_257_50_52;
   wire n_257_50_53;
   wire n_257_50_54;
   wire n_257_50_55;
   wire n_257_50_56;
   wire n_257_50_57;
   wire n_257_50_58;
   wire n_257_50_59;
   wire n_257_50_60;
   wire n_257_50_61;
   wire n_257_50_62;
   wire n_257_50_63;
   wire n_257_50_64;
   wire n_257_50_65;
   wire n_257_50_66;
   wire n_257_50_67;
   wire n_257_50_68;
   wire n_257_50_69;
   wire n_257_50_70;
   wire n_257_50_71;
   wire n_257_50_72;
   wire n_257_50_73;
   wire n_257_50_74;
   wire n_257_50_75;
   wire n_257_50_76;
   wire n_257_50_77;
   wire n_257_50_78;
   wire n_257_50_79;
   wire n_257_50_80;
   wire n_257_50_81;
   wire n_257_50_82;
   wire n_257_50_83;
   wire n_257_50_84;
   wire n_257_50_85;
   wire n_257_50_86;
   wire n_257_50_87;
   wire n_257_50_88;
   wire n_257_50_89;
   wire n_257_50_90;
   wire n_257_50_91;
   wire n_257_50_92;
   wire n_257_50_93;
   wire n_257_50_94;
   wire n_257_50_95;
   wire n_257_50_96;
   wire n_257_50_97;
   wire n_257_50_98;
   wire n_257_50_99;
   wire n_257_50_100;
   wire n_257_50_101;
   wire n_257_50_102;
   wire n_257_50_103;
   wire n_257_50_104;
   wire n_257_50_105;
   wire n_257_50_106;
   wire n_257_50_107;
   wire n_257_50_108;
   wire n_257_50_109;
   wire n_257_50_110;
   wire n_257_50_111;
   wire n_257_50_112;
   wire n_257_50_113;
   wire n_257_50_114;
   wire n_257_50_115;
   wire n_257_50_116;
   wire n_257_50_117;
   wire n_257_50_118;
   wire n_257_50_119;
   wire n_257_50_120;
   wire n_257_50_121;
   wire n_257_50_122;
   wire n_257_50_123;
   wire n_257_50_124;
   wire n_257_50_125;
   wire n_257_50_126;
   wire n_257_382;
   wire n_257_383;
   wire n_257_384;
   wire n_257_385;
   wire n_257_386;
   wire n_257_387;
   wire n_257_388;
   wire n_257_389;
   wire n_257_390;
   wire n_257_391;
   wire n_257_392;
   wire n_257_393;
   wire n_257_394;
   wire n_257_395;
   wire n_257_396;
   wire n_257_397;
   wire n_257_398;
   wire n_257_399;
   wire n_257_400;
   wire n_257_401;
   wire n_257_402;
   wire n_257_403;
   wire n_257_404;
   wire n_257_405;
   wire n_257_406;
   wire n_257_407;
   wire n_257_408;
   wire n_257_409;
   wire n_257_410;
   wire n_257_411;
   wire n_257_412;
   wire n_257_413;
   wire n_257_414;
   wire n_257_415;
   wire n_257_416;
   wire n_257_417;
   wire n_257_418;
   wire n_257_419;
   wire n_257_53_0;
   wire n_257_53_1;
   wire n_257_53_2;
   wire n_257_420;
   wire n_257_54_0;
   wire n_257_54_1;
   wire n_257_421;
   wire n_257_422;
   wire n_257_55_0;
   wire n_257_55_1;
   wire n_257_55_2;
   wire n_257_56_0;
   wire n_257_56_1;
   wire n_257_423;
   wire n_257_424;
   wire n_257_57_0;
   wire n_257_57_1;
   wire n_257_57_2;
   wire n_257_58_0;
   wire n_257_58_1;
   wire n_257_425;
   wire n_257_59_0;
   wire n_257_59_1;
   wire n_257_59_2;
   wire n_257_426;
   wire n_257_427;
   wire n_257_60_0;
   wire n_257_61_0;
   wire n_257_61_1;
   wire n_257_61_2;
   wire n_257_428;
   wire n_257_62_0;
   wire n_257_62_1;
   wire n_257_62_2;
   wire n_257_429;
   wire n_257_63_0;
   wire n_257_63_1;
   wire n_257_63_2;
   wire n_257_63_3;
   wire n_257_430;
   wire n_257_64_0;
   wire n_257_64_1;
   wire n_257_431;
   wire n_257_432;
   wire n_257_65_0;
   wire n_257_65_1;
   wire n_257_65_2;
   wire n_257_65_3;
   wire n_257_65_4;
   wire n_257_65_5;
   wire n_257_66_0;
   wire n_257_66_1;
   wire n_257_66_2;
   wire n_257_433;
   wire n_257_67_0;
   wire n_257_67_1;
   wire n_257_67_2;
   wire n_257_67_3;
   wire n_257_67_4;
   wire n_257_67_5;
   wire n_257_67_6;
   wire n_257_67_7;
   wire n_257_67_8;
   wire n_257_67_9;
   wire n_257_67_10;
   wire n_257_67_11;
   wire n_257_67_12;
   wire n_257_67_13;
   wire n_257_67_14;
   wire n_257_67_15;
   wire n_257_67_16;
   wire n_257_67_17;
   wire n_257_67_18;
   wire n_257_67_19;
   wire n_257_67_20;
   wire n_257_67_21;
   wire n_257_67_22;
   wire n_257_67_23;
   wire n_257_67_24;
   wire n_257_67_25;
   wire n_257_67_26;
   wire n_257_67_27;
   wire n_257_67_28;
   wire n_257_67_29;
   wire n_257_67_30;
   wire n_257_67_31;
   wire n_257_67_32;
   wire n_257_67_33;
   wire n_257_67_34;
   wire n_257_67_35;
   wire n_257_67_36;
   wire n_257_67_37;
   wire n_257_67_38;
   wire n_257_67_39;
   wire n_257_67_40;
   wire n_257_67_41;
   wire n_257_67_42;
   wire n_257_67_43;
   wire n_257_67_44;
   wire n_257_67_45;
   wire n_257_67_46;
   wire n_257_67_47;
   wire n_257_67_48;
   wire n_257_67_49;
   wire n_257_67_50;
   wire n_257_67_51;
   wire n_257_67_52;
   wire n_257_67_53;
   wire n_257_67_54;
   wire n_257_67_55;
   wire n_257_67_56;
   wire n_257_67_57;
   wire n_257_67_58;
   wire n_257_67_59;
   wire n_257_67_60;
   wire n_257_67_61;
   wire n_257_67_62;
   wire n_257_67_63;
   wire n_257_67_64;
   wire n_257_67_65;
   wire n_257_67_66;
   wire n_257_67_67;
   wire n_257_67_68;
   wire n_257_67_69;
   wire n_257_67_70;
   wire n_257_67_71;
   wire n_257_67_72;
   wire n_257_67_73;
   wire n_257_67_74;
   wire n_257_67_75;
   wire n_257_67_76;
   wire n_257_67_77;
   wire n_257_67_78;
   wire n_257_67_79;
   wire n_257_67_80;
   wire n_257_67_81;
   wire n_257_67_82;
   wire n_257_67_83;
   wire n_257_67_84;
   wire n_257_67_85;
   wire n_257_67_86;
   wire n_257_67_87;
   wire n_257_67_88;
   wire n_257_67_89;
   wire n_257_67_90;
   wire n_257_67_91;
   wire n_257_67_92;
   wire n_257_67_93;
   wire n_257_67_94;
   wire n_257_67_95;
   wire n_257_67_96;
   wire n_257_67_97;
   wire n_257_67_98;
   wire n_257_67_99;
   wire n_257_67_100;
   wire n_257_67_101;
   wire n_257_67_102;
   wire n_257_67_103;
   wire n_257_67_104;
   wire n_257_67_105;
   wire n_257_67_106;
   wire n_257_67_107;
   wire n_257_67_108;
   wire n_257_67_109;
   wire n_257_67_110;
   wire n_257_67_111;
   wire n_257_67_112;
   wire n_257_67_113;
   wire n_257_67_114;
   wire n_257_67_115;
   wire n_257_67_116;
   wire n_257_67_117;
   wire n_257_67_118;
   wire n_257_67_119;
   wire n_257_67_120;
   wire n_257_67_121;
   wire n_257_67_122;
   wire n_257_67_123;
   wire n_257_67_124;
   wire n_257_67_125;
   wire n_257_67_126;
   wire n_257_434;
   wire n_257_68_0;
   wire n_257_68_1;
   wire n_257_435;
   wire n_257_69_0;
   wire n_257_69_1;
   wire n_257_436;
   wire n_257_70_0;
   wire n_257_70_1;
   wire n_257_437;
   wire n_257_71_0;
   wire n_257_71_1;
   wire n_257_438;
   wire n_257_72_0;
   wire n_257_72_1;
   wire n_257_439;
   wire n_257_73_0;
   wire n_257_73_1;
   wire n_257_440;
   wire n_257_74_0;
   wire n_257_441;
   wire n_257_75_0;
   wire n_257_75_1;
   wire n_257_75_2;
   wire n_257_75_3;
   wire n_257_75_4;
   wire n_257_75_5;
   wire n_257_75_6;
   wire n_257_75_7;
   wire n_257_75_8;
   wire n_257_75_9;
   wire n_257_75_10;
   wire n_257_75_11;
   wire n_257_75_12;
   wire n_257_75_13;
   wire n_257_75_14;
   wire n_257_75_15;
   wire n_257_75_16;
   wire n_257_75_17;
   wire n_257_75_18;
   wire n_257_75_19;
   wire n_257_75_20;
   wire n_257_75_21;
   wire n_257_75_22;
   wire n_257_75_23;
   wire n_257_75_24;
   wire n_257_75_25;
   wire n_257_75_26;
   wire n_257_75_27;
   wire n_257_75_28;
   wire n_257_75_29;
   wire n_257_75_30;
   wire n_257_75_31;
   wire n_257_75_32;
   wire n_257_75_33;
   wire n_257_444;
   wire n_257_449;
   wire n_257_448;
   wire n_257_75_34;
   wire n_257_451;
   wire n_257_75_35;
   wire n_257_450;
   wire n_257_452;
   wire n_257_453;
   wire n_257_454;
   wire n_257_455;
   wire n_257_456;
   wire n_257_457;
   wire n_257_458;
   wire n_257_459;
   wire n_257_75_36;
   wire n_257_460;
   wire n_257_461;
   wire n_257_462;
   wire n_257_463;
   wire n_257_464;
   wire n_257_465;
   wire n_257_466;
   wire n_257_467;
   wire n_257_75_37;
   wire n_257_75_38;
   wire n_257_468;
   wire n_257_469;
   wire n_257_470;
   wire n_257_471;
   wire n_257_472;
   wire n_257_473;
   wire n_257_474;
   wire n_257_475;
   wire n_257_75_39;
   wire n_257_476;
   wire n_257_477;
   wire n_257_478;
   wire n_257_479;
   wire n_257_480;
   wire n_257_481;
   wire n_257_482;
   wire n_257_483;
   wire n_257_75_40;
   wire n_257_75_41;
   wire n_257_75_42;
   wire n_257_485;
   wire n_257_486;
   wire n_257_487;
   wire n_257_488;
   wire n_257_489;
   wire n_257_490;
   wire n_257_491;
   wire n_257_492;
   wire n_257_75_43;
   wire n_257_493;
   wire n_257_494;
   wire n_257_495;
   wire n_257_496;
   wire n_257_497;
   wire n_257_498;
   wire n_257_499;
   wire n_257_500;
   wire n_257_75_44;
   wire n_257_501;
   wire n_257_502;
   wire n_257_503;
   wire n_257_504;
   wire n_257_505;
   wire n_257_506;
   wire n_257_507;
   wire n_257_508;
   wire n_257_75_45;
   wire n_257_509;
   wire n_257_510;
   wire n_257_511;
   wire n_257_512;
   wire n_257_513;
   wire n_257_514;
   wire n_257_515;
   wire n_257_516;
   wire n_257_75_46;
   wire n_257_517;
   wire n_257_518;
   wire n_257_519;
   wire n_257_520;
   wire n_257_521;
   wire n_257_522;
   wire n_257_523;
   wire n_257_524;
   wire n_257_75_47;
   wire n_257_525;
   wire n_257_526;
   wire n_257_527;
   wire n_257_528;
   wire n_257_529;
   wire n_257_530;
   wire n_257_531;
   wire n_257_532;
   wire n_257_75_48;
   wire n_257_75_49;
   wire n_257_533;
   wire n_257_534;
   wire n_257_535;
   wire n_257_536;
   wire n_257_537;
   wire n_257_538;
   wire n_257_539;
   wire n_257_540;
   wire n_257_75_50;
   wire n_257_541;
   wire n_257_542;
   wire n_257_543;
   wire n_257_544;
   wire n_257_545;
   wire n_257_546;
   wire n_257_547;
   wire n_257_548;
   wire n_257_75_51;
   wire n_257_549;
   wire n_257_550;
   wire n_257_551;
   wire n_257_552;
   wire n_257_553;
   wire n_257_554;
   wire n_257_555;
   wire n_257_556;
   wire n_257_75_52;
   wire n_257_557;
   wire n_257_558;
   wire n_257_559;
   wire n_257_560;
   wire n_257_561;
   wire n_257_562;
   wire n_257_563;
   wire n_257_564;
   wire n_257_75_53;
   wire n_257_75_54;
   wire n_257_565;
   wire n_257_566;
   wire n_257_567;
   wire n_257_568;
   wire n_257_569;
   wire n_257_570;
   wire n_257_571;
   wire n_257_572;
   wire n_257_75_55;
   wire n_257_573;
   wire n_257_574;
   wire n_257_575;
   wire n_257_576;
   wire n_257_577;
   wire n_257_578;
   wire n_257_579;
   wire n_257_580;
   wire n_257_75_56;
   wire n_257_75_57;
   wire n_257_581;
   wire n_257_582;
   wire n_257_583;
   wire n_257_584;
   wire n_257_585;
   wire n_257_586;
   wire n_257_587;
   wire n_257_588;
   wire n_257_75_58;
   wire n_257_589;
   wire n_257_590;
   wire n_257_591;
   wire n_257_592;
   wire n_257_593;
   wire n_257_594;
   wire n_257_595;
   wire n_257_596;
   wire n_257_75_59;
   wire n_257_75_60;
   wire n_257_75_61;
   wire n_257_597;
   wire n_257_598;
   wire n_257_599;
   wire n_257_600;
   wire n_257_601;
   wire n_257_602;
   wire n_257_603;
   wire n_257_604;
   wire n_257_75_62;
   wire n_257_605;
   wire n_257_606;
   wire n_257_607;
   wire n_257_608;
   wire n_257_609;
   wire n_257_610;
   wire n_257_611;
   wire n_257_612;
   wire n_257_75_63;
   wire n_257_613;
   wire n_257_614;
   wire n_257_615;
   wire n_257_616;
   wire n_257_617;
   wire n_257_618;
   wire n_257_619;
   wire n_257_620;
   wire n_257_75_64;
   wire n_257_621;
   wire n_257_622;
   wire n_257_623;
   wire n_257_624;
   wire n_257_625;
   wire n_257_626;
   wire n_257_627;
   wire n_257_628;
   wire n_257_75_65;
   wire n_257_75_66;
   wire n_257_75_67;
   wire n_257_75_68;
   wire n_257_629;
   wire n_257_630;
   wire n_257_631;
   wire n_257_632;
   wire n_257_633;
   wire n_257_634;
   wire n_257_635;
   wire n_257_636;
   wire n_257_75_69;
   wire n_257_637;
   wire n_257_638;
   wire n_257_639;
   wire n_257_640;
   wire n_257_641;
   wire n_257_642;
   wire n_257_643;
   wire n_257_644;
   wire n_257_75_70;
   wire n_257_645;
   wire n_257_646;
   wire n_257_647;
   wire n_257_648;
   wire n_257_649;
   wire n_257_650;
   wire n_257_651;
   wire n_257_652;
   wire n_257_75_71;
   wire n_257_653;
   wire n_257_654;
   wire n_257_655;
   wire n_257_656;
   wire n_257_657;
   wire n_257_658;
   wire n_257_659;
   wire n_257_660;
   wire n_257_75_72;
   wire n_257_75_73;
   wire n_257_75_74;
   wire n_257_75_75;
   wire n_257_75_76;
   wire n_257_661;
   wire n_257_662;
   wire n_257_663;
   wire n_257_664;
   wire n_257_665;
   wire n_257_666;
   wire n_257_667;
   wire n_257_668;
   wire n_257_75_77;
   wire n_257_669;
   wire n_257_670;
   wire n_257_671;
   wire n_257_672;
   wire n_257_673;
   wire n_257_674;
   wire n_257_675;
   wire n_257_676;
   wire n_257_75_78;
   wire n_257_677;
   wire n_257_678;
   wire n_257_679;
   wire n_257_680;
   wire n_257_681;
   wire n_257_682;
   wire n_257_683;
   wire n_257_684;
   wire n_257_75_79;
   wire n_257_75_80;
   wire n_257_685;
   wire n_257_686;
   wire n_257_687;
   wire n_257_688;
   wire n_257_689;
   wire n_257_690;
   wire n_257_691;
   wire n_257_692;
   wire n_257_75_81;
   wire n_257_693;
   wire n_257_694;
   wire n_257_695;
   wire n_257_696;
   wire n_257_697;
   wire n_257_698;
   wire n_257_699;
   wire n_257_700;
   wire n_257_75_82;
   wire n_257_75_83;
   wire n_257_75_84;
   wire n_257_75_85;
   wire n_257_701;
   wire n_257_702;
   wire n_257_703;
   wire n_257_704;
   wire n_257_705;
   wire n_257_706;
   wire n_257_707;
   wire n_257_708;
   wire n_257_75_86;
   wire n_257_709;
   wire n_257_710;
   wire n_257_711;
   wire n_257_712;
   wire n_257_713;
   wire n_257_714;
   wire n_257_715;
   wire n_257_716;
   wire n_257_75_87;
   wire n_257_75_88;
   wire n_257_717;
   wire n_257_718;
   wire n_257_719;
   wire n_257_720;
   wire n_257_721;
   wire n_257_722;
   wire n_257_723;
   wire n_257_724;
   wire n_257_75_89;
   wire n_257_725;
   wire n_257_726;
   wire n_257_727;
   wire n_257_728;
   wire n_257_729;
   wire n_257_730;
   wire n_257_731;
   wire n_257_732;
   wire n_257_75_90;
   wire n_257_75_91;
   wire n_257_75_92;
   wire n_257_75_93;
   wire n_257_733;
   wire n_257_734;
   wire n_257_735;
   wire n_257_736;
   wire n_257_737;
   wire n_257_738;
   wire n_257_739;
   wire n_257_740;
   wire n_257_75_94;
   wire n_257_741;
   wire n_257_742;
   wire n_257_743;
   wire n_257_744;
   wire n_257_745;
   wire n_257_746;
   wire n_257_747;
   wire n_257_748;
   wire n_257_75_95;
   wire n_257_75_96;
   wire n_257_749;
   wire n_257_750;
   wire n_257_751;
   wire n_257_752;
   wire n_257_753;
   wire n_257_754;
   wire n_257_755;
   wire n_257_756;
   wire n_257_75_97;
   wire n_257_757;
   wire n_257_758;
   wire n_257_759;
   wire n_257_760;
   wire n_257_761;
   wire n_257_762;
   wire n_257_763;
   wire n_257_764;
   wire n_257_75_98;
   wire n_257_75_99;
   wire n_257_75_100;
   wire n_257_75_101;
   wire n_257_765;
   wire n_257_766;
   wire n_257_767;
   wire n_257_768;
   wire n_257_769;
   wire n_257_770;
   wire n_257_771;
   wire n_257_772;
   wire n_257_75_102;
   wire n_257_773;
   wire n_257_774;
   wire n_257_775;
   wire n_257_776;
   wire n_257_777;
   wire n_257_778;
   wire n_257_779;
   wire n_257_780;
   wire n_257_75_103;
   wire n_257_75_104;
   wire n_257_781;
   wire n_257_782;
   wire n_257_783;
   wire n_257_784;
   wire n_257_785;
   wire n_257_786;
   wire n_257_787;
   wire n_257_788;
   wire n_257_75_105;
   wire n_257_789;
   wire n_257_790;
   wire n_257_791;
   wire n_257_792;
   wire n_257_793;
   wire n_257_794;
   wire n_257_795;
   wire n_257_796;
   wire n_257_75_106;
   wire n_257_75_107;
   wire n_257_75_108;
   wire n_257_75_109;
   wire n_257_797;
   wire n_257_798;
   wire n_257_799;
   wire n_257_800;
   wire n_257_801;
   wire n_257_802;
   wire n_257_803;
   wire n_257_804;
   wire n_257_75_110;
   wire n_257_805;
   wire n_257_806;
   wire n_257_807;
   wire n_257_808;
   wire n_257_809;
   wire n_257_810;
   wire n_257_811;
   wire n_257_812;
   wire n_257_75_111;
   wire n_257_75_112;
   wire n_257_813;
   wire n_257_814;
   wire n_257_815;
   wire n_257_816;
   wire n_257_817;
   wire n_257_818;
   wire n_257_819;
   wire n_257_820;
   wire n_257_75_113;
   wire n_257_821;
   wire n_257_75_114;
   wire n_257_822;
   wire n_257_75_115;
   wire n_257_823;
   wire n_257_75_116;
   wire n_257_824;
   wire n_257_75_117;
   wire n_257_825;
   wire n_257_75_118;
   wire n_257_826;
   wire n_257_75_119;
   wire n_257_827;
   wire n_257_75_120;
   wire n_257_828;
   wire n_257_75_121;
   wire n_257_75_122;
   wire n_257_75_123;
   wire n_257_75_124;
   wire n_257_75_125;
   wire n_257_75_126;
   wire n_257_75_127;
   wire n_257_829;
   wire n_257_830;
   wire n_257_831;
   wire n_257_832;
   wire n_257_833;
   wire n_257_834;
   wire n_257_835;
   wire n_257_836;
   wire n_257_75_128;
   wire n_257_837;
   wire n_257_838;
   wire n_257_839;
   wire n_257_840;
   wire n_257_841;
   wire n_257_842;
   wire n_257_843;
   wire n_257_844;
   wire n_257_75_129;
   wire n_257_75_130;
   wire n_257_845;
   wire n_257_846;
   wire n_257_847;
   wire n_257_848;
   wire n_257_849;
   wire n_257_850;
   wire n_257_851;
   wire n_257_852;
   wire n_257_75_131;
   wire n_257_853;
   wire n_257_854;
   wire n_257_855;
   wire n_257_856;
   wire n_257_857;
   wire n_257_858;
   wire n_257_859;
   wire n_257_860;
   wire n_257_75_132;
   wire n_257_75_133;
   wire n_257_75_134;
   wire n_257_75_135;
   wire n_257_861;
   wire n_257_862;
   wire n_257_863;
   wire n_257_864;
   wire n_257_865;
   wire n_257_866;
   wire n_257_867;
   wire n_257_868;
   wire n_257_75_136;
   wire n_257_869;
   wire n_257_870;
   wire n_257_871;
   wire n_257_872;
   wire n_257_873;
   wire n_257_874;
   wire n_257_875;
   wire n_257_876;
   wire n_257_75_137;
   wire n_257_75_138;
   wire n_257_877;
   wire n_257_878;
   wire n_257_879;
   wire n_257_880;
   wire n_257_881;
   wire n_257_882;
   wire n_257_883;
   wire n_257_884;
   wire n_257_75_139;
   wire n_257_885;
   wire n_257_75_140;
   wire n_257_886;
   wire n_257_75_141;
   wire n_257_887;
   wire n_257_75_142;
   wire n_257_888;
   wire n_257_75_143;
   wire n_257_889;
   wire n_257_75_144;
   wire n_257_890;
   wire n_257_75_145;
   wire n_257_891;
   wire n_257_75_146;
   wire n_257_892;
   wire n_257_75_147;
   wire n_257_75_148;
   wire n_257_75_149;
   wire n_257_75_150;
   wire n_257_75_151;
   wire n_257_75_152;
   wire n_257_893;
   wire n_257_894;
   wire n_257_895;
   wire n_257_896;
   wire n_257_897;
   wire n_257_898;
   wire n_257_75_153;
   wire n_257_899;
   wire n_257_900;
   wire n_257_901;
   wire n_257_902;
   wire n_257_903;
   wire n_257_904;
   wire n_257_905;
   wire n_257_906;
   wire n_257_75_154;
   wire n_257_907;
   wire n_257_908;
   wire n_257_909;
   wire n_257_910;
   wire n_257_911;
   wire n_257_912;
   wire n_257_913;
   wire n_257_914;
   wire n_257_75_155;
   wire n_257_915;
   wire n_257_916;
   wire n_257_917;
   wire n_257_918;
   wire n_257_919;
   wire n_257_920;
   wire n_257_921;
   wire n_257_922;
   wire n_257_75_156;
   wire n_257_923;
   wire n_257_75_157;
   wire n_257_924;
   wire n_257_75_158;
   wire n_257_925;
   wire n_257_75_159;
   wire n_257_926;
   wire n_257_75_160;
   wire n_257_927;
   wire n_257_75_161;
   wire n_257_928;
   wire n_257_75_162;
   wire n_257_929;
   wire n_257_75_163;
   wire n_257_930;
   wire n_257_75_164;
   wire n_257_75_165;
   wire n_257_75_166;
   wire n_257_75_167;
   wire n_257_75_168;
   wire n_257_75_169;
   wire n_257_75_170;
   wire n_257_75_171;
   wire n_257_75_172;
   wire n_257_931;
   wire n_257_932;
   wire n_257_933;
   wire n_257_934;
   wire n_257_935;
   wire n_257_936;
   wire n_257_937;
   wire n_257_938;
   wire n_257_75_173;
   wire n_257_939;
   wire n_257_940;
   wire n_257_941;
   wire n_257_942;
   wire n_257_943;
   wire n_257_944;
   wire n_257_945;
   wire n_257_946;
   wire n_257_75_174;
   wire n_257_947;
   wire n_257_948;
   wire n_257_949;
   wire n_257_950;
   wire n_257_951;
   wire n_257_952;
   wire n_257_953;
   wire n_257_954;
   wire n_257_75_175;
   wire n_257_955;
   wire n_257_75_176;
   wire n_257_956;
   wire n_257_75_177;
   wire n_257_957;
   wire n_257_75_178;
   wire n_257_958;
   wire n_257_75_179;
   wire n_257_959;
   wire n_257_75_180;
   wire n_257_960;
   wire n_257_75_181;
   wire n_257_961;
   wire n_257_75_182;
   wire n_257_962;
   wire n_257_75_183;
   wire n_257_75_184;
   wire n_257_75_185;
   wire n_257_75_186;
   wire n_257_75_187;
   wire n_257_75_188;
   wire n_257_75_189;
   wire n_257_75_190;
   wire n_257_75_191;
   wire n_257_963;
   wire n_257_964;
   wire n_257_965;
   wire n_257_966;
   wire n_257_967;
   wire n_257_968;
   wire n_257_969;
   wire n_257_970;
   wire n_257_75_192;
   wire n_257_971;
   wire n_257_972;
   wire n_257_973;
   wire n_257_974;
   wire n_257_975;
   wire n_257_976;
   wire n_257_977;
   wire n_257_978;
   wire n_257_75_193;
   wire n_257_979;
   wire n_257_980;
   wire n_257_981;
   wire n_257_982;
   wire n_257_983;
   wire n_257_984;
   wire n_257_985;
   wire n_257_986;
   wire n_257_75_194;
   wire n_257_987;
   wire n_257_75_195;
   wire n_257_988;
   wire n_257_75_196;
   wire n_257_989;
   wire n_257_75_197;
   wire n_257_990;
   wire n_257_75_198;
   wire n_257_991;
   wire n_257_75_199;
   wire n_257_75_200;
   wire n_257_992;
   wire n_257_75_201;
   wire n_257_75_202;
   wire n_257_993;
   wire n_257_75_203;
   wire n_257_75_204;
   wire n_257_994;
   wire n_257_75_205;
   wire n_257_75_206;
   wire n_257_75_207;
   wire n_257_75_208;
   wire n_257_75_209;
   wire n_257_75_210;
   wire n_257_75_211;
   wire n_257_75_212;
   wire n_257_75_213;
   wire n_257_75_214;
   wire n_257_75_215;
   wire n_257_75_216;
   wire n_257_995;
   wire n_257_996;
   wire n_257_997;
   wire n_257_998;
   wire n_257_999;
   wire n_257_1000;
   wire n_257_1001;
   wire n_257_1002;
   wire n_257_75_217;
   wire n_257_1003;
   wire n_257_1004;
   wire n_257_1005;
   wire n_257_1006;
   wire n_257_1007;
   wire n_257_1008;
   wire n_257_1009;
   wire n_257_1010;
   wire n_257_75_218;
   wire n_257_1011;
   wire n_257_1012;
   wire n_257_1013;
   wire n_257_1014;
   wire n_257_1015;
   wire n_257_1016;
   wire n_257_1017;
   wire n_257_1018;
   wire n_257_75_219;
   wire n_257_1019;
   wire n_257_75_220;
   wire n_257_1020;
   wire n_257_75_221;
   wire n_257_1021;
   wire n_257_75_222;
   wire n_257_1022;
   wire n_257_75_223;
   wire n_257_1023;
   wire n_257_75_224;
   wire n_257_1024;
   wire n_257_75_225;
   wire n_257_1025;
   wire n_257_75_226;
   wire n_257_1026;
   wire n_257_75_227;
   wire n_257_75_228;
   wire n_257_75_229;
   wire n_257_1027;
   wire n_257_1028;
   wire n_257_1029;
   wire n_257_1030;
   wire n_257_1031;
   wire n_257_1032;
   wire n_257_1033;
   wire n_257_1034;
   wire n_257_75_230;
   wire n_257_1035;
   wire n_257_1036;
   wire n_257_1037;
   wire n_257_1038;
   wire n_257_1039;
   wire n_257_1040;
   wire n_257_1041;
   wire n_257_1042;
   wire n_257_75_231;
   wire n_257_1043;
   wire n_257_1044;
   wire n_257_1045;
   wire n_257_1046;
   wire n_257_1047;
   wire n_257_1048;
   wire n_257_1049;
   wire n_257_1050;
   wire n_257_75_232;
   wire n_257_1051;
   wire n_257_75_233;
   wire n_257_1052;
   wire n_257_75_234;
   wire n_257_1053;
   wire n_257_75_235;
   wire n_257_1054;
   wire n_257_75_236;
   wire n_257_1055;
   wire n_257_75_237;
   wire n_257_1056;
   wire n_257_75_238;
   wire n_257_1057;
   wire n_257_75_239;
   wire n_257_1058;
   wire n_257_75_240;
   wire n_257_75_241;
   wire n_257_75_242;
   wire n_257_1059;
   wire n_257_1060;
   wire n_257_1061;
   wire n_257_1062;
   wire n_257_1063;
   wire n_257_1064;
   wire n_257_1065;
   wire n_257_1066;
   wire n_257_75_243;
   wire n_257_1067;
   wire n_257_1068;
   wire n_257_1069;
   wire n_257_1070;
   wire n_257_1071;
   wire n_257_1072;
   wire n_257_1073;
   wire n_257_1074;
   wire n_257_75_244;
   wire n_257_1075;
   wire n_257_1076;
   wire n_257_1077;
   wire n_257_1078;
   wire n_257_1079;
   wire n_257_1080;
   wire n_257_1081;
   wire n_257_1082;
   wire n_257_75_245;
   wire n_257_1083;
   wire n_257_75_246;
   wire n_257_1084;
   wire n_257_75_247;
   wire n_257_1085;
   wire n_257_75_248;
   wire n_257_1086;
   wire n_257_75_249;
   wire n_257_1087;
   wire n_257_75_250;
   wire n_257_75_251;
   wire n_257_1088;
   wire n_257_75_252;
   wire n_257_75_253;
   wire n_257_1089;
   wire n_257_75_254;
   wire n_257_75_255;
   wire n_257_75_256;
   wire n_257_75_257;
   wire n_257_1090;
   wire n_257_75_258;
   wire n_257_75_259;
   wire n_257_75_260;
   wire n_257_1092;
   wire n_257_75_261;
   wire n_257_1093;
   wire n_257_1094;
   wire n_257_1095;
   wire n_257_75_262;
   wire n_257_75_263;
   wire n_257_75_264;
   wire n_257_75_265;
   wire n_257_75_266;
   wire n_257_75_267;
   wire n_257_75_268;
   wire n_257_75_269;
   wire n_257_75_270;
   wire n_257_75_271;
   wire n_257_75_272;
   wire n_257_75_273;
   wire n_257_75_274;
   wire n_257_75_275;
   wire n_257_75_276;
   wire n_257_75_277;
   wire n_257_75_278;
   wire n_257_75_279;
   wire n_257_75_280;
   wire n_257_75_281;
   wire n_257_75_282;
   wire n_257_75_283;
   wire n_257_75_284;
   wire n_257_75_285;
   wire n_257_75_286;
   wire n_257_75_287;
   wire n_257_75_288;
   wire n_257_75_289;
   wire n_257_75_290;
   wire n_257_75_291;
   wire n_257_75_292;
   wire n_257_75_293;
   wire n_257_75_294;
   wire n_257_75_295;
   wire n_257_1091;
   wire n_257_75_296;
   wire n_257_75_297;
   wire n_257_75_298;
   wire n_257_443;
   wire n_257_75_299;
   wire n_257_445;
   wire n_257_484;
   wire n_257_75_300;
   wire n_257_75_301;
   wire n_257_75_302;
   wire n_257_75_303;
   wire n_257_75_304;
   wire n_257_75_305;
   wire n_257_75_306;
   wire n_257_75_307;
   wire n_257_442;
   wire n_257_446;
   wire n_257_75_308;
   wire n_257_75_309;
   wire n_257_447;
   wire n_257_75_310;
   wire n_257_75_311;
   wire n_257_75_312;
   wire n_257_75_313;
   wire n_257_75_314;
   wire n_257_75_315;
   wire n_257_75_316;
   wire n_257_1096;
   wire n_257_75_317;
   wire n_257_75_318;
   wire n_257_75_319;
   wire n_257_75_320;
   wire n_257_75_321;
   wire n_257_75_322;
   wire n_257_75_323;
   wire n_257_76_0;
   wire n_257_76_1;
   wire n_257_76_2;
   wire n_257_76_3;
   wire n_257_76_4;
   wire n_257_76_5;
   wire n_257_76_6;
   wire n_257_76_7;
   wire n_257_76_8;
   wire n_257_76_9;
   wire n_257_76_10;
   wire n_257_76_11;
   wire n_257_76_12;
   wire n_257_76_13;
   wire n_257_76_14;
   wire n_257_76_15;
   wire n_257_76_16;
   wire n_257_76_17;
   wire n_257_76_18;
   wire n_257_76_19;
   wire n_257_76_20;
   wire n_257_76_21;
   wire n_257_76_22;
   wire n_257_76_23;
   wire n_257_76_24;
   wire n_257_76_25;
   wire n_257_76_26;
   wire n_257_76_27;
   wire n_257_76_28;
   wire n_257_76_29;
   wire n_257_76_30;
   wire n_257_76_31;
   wire n_257_76_32;
   wire n_257_76_33;
   wire n_257_76_34;
   wire n_257_76_35;
   wire n_257_76_36;
   wire n_257_76_37;
   wire n_257_76_38;
   wire n_257_76_39;
   wire n_257_76_40;
   wire n_257_76_41;
   wire n_257_76_42;
   wire n_257_76_43;
   wire n_257_76_44;
   wire n_257_76_45;
   wire n_257_76_46;
   wire n_257_76_47;
   wire n_257_76_48;
   wire n_257_76_49;
   wire n_257_76_50;
   wire n_257_76_51;
   wire n_257_76_52;
   wire n_257_76_53;
   wire n_257_76_54;
   wire n_257_76_55;
   wire n_257_76_56;
   wire n_257_76_57;
   wire n_257_76_58;
   wire n_257_76_59;
   wire n_257_76_60;
   wire n_257_76_61;
   wire n_257_76_62;
   wire n_257_76_63;
   wire n_257_76_64;
   wire n_257_76_65;
   wire n_257_76_66;
   wire n_257_76_67;
   wire n_257_76_68;
   wire n_257_76_69;
   wire n_257_76_70;
   wire n_257_76_71;
   wire n_257_76_72;
   wire n_257_76_73;
   wire n_257_76_74;
   wire n_257_76_75;
   wire n_257_76_76;
   wire n_257_76_77;
   wire n_257_76_78;
   wire n_257_76_79;
   wire n_257_76_80;
   wire n_257_76_81;
   wire n_257_76_82;
   wire n_257_76_83;
   wire n_257_76_84;
   wire n_257_76_85;
   wire n_257_76_86;
   wire n_257_76_87;
   wire n_257_76_88;
   wire n_257_76_89;
   wire n_257_76_90;
   wire n_257_76_91;
   wire n_257_76_92;
   wire n_257_76_93;
   wire n_257_76_94;
   wire n_257_76_95;
   wire n_257_76_96;
   wire n_257_76_97;
   wire n_257_76_98;
   wire n_257_76_99;
   wire n_257_76_100;
   wire n_257_76_101;
   wire n_257_76_102;
   wire n_257_76_103;
   wire n_257_76_104;
   wire n_257_76_105;
   wire n_257_76_106;
   wire n_257_76_107;
   wire n_257_76_108;
   wire n_257_76_109;
   wire n_257_76_110;
   wire n_257_76_111;
   wire n_257_76_112;
   wire n_257_76_113;
   wire n_257_76_114;
   wire n_257_76_115;
   wire n_257_76_116;
   wire n_257_76_117;
   wire n_257_76_118;
   wire n_257_76_119;
   wire n_257_76_120;
   wire n_257_76_121;
   wire n_257_76_122;
   wire n_257_76_123;
   wire n_257_76_124;
   wire n_257_76_125;
   wire n_257_76_126;
   wire n_257_76_127;
   wire n_257_76_128;
   wire n_257_76_129;
   wire n_257_76_130;
   wire n_257_76_131;
   wire n_257_76_132;
   wire n_257_76_133;
   wire n_257_76_134;
   wire n_257_76_135;
   wire n_257_76_136;
   wire n_257_76_137;
   wire n_257_76_138;
   wire n_257_76_139;
   wire n_257_76_140;
   wire n_257_76_141;
   wire n_257_76_142;
   wire n_257_76_143;
   wire n_257_76_144;
   wire n_257_76_145;
   wire n_257_76_146;
   wire n_257_76_147;
   wire n_257_76_148;
   wire n_257_76_149;
   wire n_257_76_150;
   wire n_257_76_151;
   wire n_257_76_152;
   wire n_257_76_153;
   wire n_257_76_154;
   wire n_257_76_155;
   wire n_257_76_156;
   wire n_257_76_157;
   wire n_257_76_158;
   wire n_257_76_159;
   wire n_257_76_160;
   wire n_257_76_161;
   wire n_257_76_162;
   wire n_257_76_163;
   wire n_257_76_164;
   wire n_257_76_165;
   wire n_257_76_166;
   wire n_257_76_167;
   wire n_257_76_168;
   wire n_257_76_169;
   wire n_257_76_170;
   wire n_257_76_171;
   wire n_257_76_172;
   wire n_257_76_173;
   wire n_257_76_174;
   wire n_257_76_175;
   wire n_257_76_176;
   wire n_257_76_177;
   wire n_257_76_178;
   wire n_257_76_179;
   wire n_257_76_180;
   wire n_257_76_181;
   wire n_257_76_182;
   wire n_257_76_183;
   wire n_257_76_184;
   wire n_257_76_185;
   wire n_257_76_186;
   wire n_257_76_187;
   wire n_257_76_188;
   wire n_257_76_189;
   wire n_257_76_190;
   wire n_257_76_191;
   wire n_257_76_192;
   wire n_257_76_193;
   wire n_257_76_194;
   wire n_257_76_195;
   wire n_257_76_196;
   wire n_257_76_197;
   wire n_257_76_198;
   wire n_257_76_199;
   wire n_257_76_200;
   wire n_257_76_201;
   wire n_257_76_202;
   wire n_257_76_203;
   wire n_257_76_204;
   wire n_257_76_205;
   wire n_257_76_206;
   wire n_257_76_207;
   wire n_257_76_208;
   wire n_257_76_209;
   wire n_257_76_210;
   wire n_257_76_211;
   wire n_257_76_212;
   wire n_257_76_213;
   wire n_257_76_214;
   wire n_257_76_215;
   wire n_257_76_216;
   wire n_257_76_217;
   wire n_257_76_218;
   wire n_257_76_219;
   wire n_257_76_220;
   wire n_257_76_221;
   wire n_257_76_222;
   wire n_257_76_223;
   wire n_257_76_224;
   wire n_257_76_225;
   wire n_257_76_226;
   wire n_257_76_227;
   wire n_257_76_228;
   wire n_257_76_229;
   wire n_257_76_230;
   wire n_257_76_231;
   wire n_257_76_232;
   wire n_257_76_233;
   wire n_257_76_234;
   wire n_257_76_235;
   wire n_257_76_236;
   wire n_257_76_237;
   wire n_257_76_238;
   wire n_257_76_239;
   wire n_257_76_240;
   wire n_257_76_241;
   wire n_257_76_242;
   wire n_257_76_243;
   wire n_257_76_244;
   wire n_257_76_245;
   wire n_257_76_246;
   wire n_257_76_247;
   wire n_257_76_248;
   wire n_257_76_249;
   wire n_257_76_250;
   wire n_257_76_251;
   wire n_257_76_252;
   wire n_257_76_253;
   wire n_257_76_254;
   wire n_257_76_255;
   wire n_257_76_256;
   wire n_257_76_257;
   wire n_257_76_258;
   wire n_257_76_259;
   wire n_257_76_260;
   wire n_257_76_261;
   wire n_257_76_262;
   wire n_257_76_263;
   wire n_257_76_264;
   wire n_257_76_265;
   wire n_257_76_266;
   wire n_257_76_267;
   wire n_257_76_268;
   wire n_257_76_269;
   wire n_257_76_270;
   wire n_257_76_271;
   wire n_257_76_272;
   wire n_257_76_273;
   wire n_257_76_274;
   wire n_257_76_275;
   wire n_257_76_276;
   wire n_257_76_277;
   wire n_257_76_278;
   wire n_257_76_279;
   wire n_257_76_280;
   wire n_257_76_281;
   wire n_257_76_282;
   wire n_257_76_283;
   wire n_257_76_284;
   wire n_257_76_285;
   wire n_257_76_286;
   wire n_257_76_287;
   wire n_257_76_288;
   wire n_257_76_289;
   wire n_257_76_290;
   wire n_257_76_291;
   wire n_257_76_292;
   wire n_257_76_293;
   wire n_257_76_294;
   wire n_257_76_295;
   wire n_257_76_296;
   wire n_257_76_297;
   wire n_257_76_298;
   wire n_257_76_299;
   wire n_257_76_300;
   wire n_257_76_301;
   wire n_257_76_302;
   wire n_257_76_303;
   wire n_257_76_304;
   wire n_257_76_305;
   wire n_257_76_306;
   wire n_257_76_307;
   wire n_257_76_308;
   wire n_257_76_309;
   wire n_257_76_310;
   wire n_257_76_311;
   wire n_257_76_312;
   wire n_257_76_313;
   wire n_257_76_314;
   wire n_257_76_315;
   wire n_257_76_316;
   wire n_257_76_317;
   wire n_257_76_318;
   wire n_257_76_319;
   wire n_257_76_320;
   wire n_257_76_321;
   wire n_257_76_322;
   wire n_257_76_323;
   wire n_257_76_324;
   wire n_257_76_325;
   wire n_257_76_326;
   wire n_257_76_327;
   wire n_257_76_328;
   wire n_257_76_329;
   wire n_257_76_330;
   wire n_257_76_331;
   wire n_257_76_332;
   wire n_257_76_333;
   wire n_257_76_334;
   wire n_257_76_335;
   wire n_257_76_336;
   wire n_257_76_337;
   wire n_257_76_338;
   wire n_257_76_339;
   wire n_257_76_340;
   wire n_257_76_341;
   wire n_257_76_342;
   wire n_257_76_343;
   wire n_257_76_344;
   wire n_257_76_345;
   wire n_257_76_346;
   wire n_257_76_347;
   wire n_257_76_348;
   wire n_257_76_349;
   wire n_257_76_350;
   wire n_257_76_351;
   wire n_257_76_352;
   wire n_257_76_353;
   wire n_257_76_354;
   wire n_257_76_355;
   wire n_257_76_356;
   wire n_257_76_357;
   wire n_257_76_358;
   wire n_257_76_359;
   wire n_257_76_360;
   wire n_257_76_361;
   wire n_257_76_362;
   wire n_257_76_363;
   wire n_257_76_364;
   wire n_257_76_365;
   wire n_257_76_366;
   wire n_257_76_367;
   wire n_257_76_368;
   wire n_257_76_369;
   wire n_257_76_370;
   wire n_257_76_371;
   wire n_257_76_372;
   wire n_257_76_373;
   wire n_257_76_374;
   wire n_257_76_375;
   wire n_257_76_376;
   wire n_257_76_377;
   wire n_257_76_378;
   wire n_257_76_379;
   wire n_257_76_380;
   wire n_257_76_381;
   wire n_257_76_382;
   wire n_257_76_383;
   wire n_257_76_384;
   wire n_257_76_385;
   wire n_257_76_386;
   wire n_257_76_387;
   wire n_257_76_388;
   wire n_257_76_389;
   wire n_257_76_390;
   wire n_257_76_391;
   wire n_257_76_392;
   wire n_257_76_393;
   wire n_257_76_394;
   wire n_257_76_395;
   wire n_257_76_396;
   wire n_257_76_397;
   wire n_257_76_398;
   wire n_257_76_399;
   wire n_257_76_400;
   wire n_257_76_401;
   wire n_257_76_402;
   wire n_257_76_403;
   wire n_257_76_404;
   wire n_257_76_405;
   wire n_257_76_406;
   wire n_257_76_407;
   wire n_257_76_408;
   wire n_257_76_409;
   wire n_257_76_410;
   wire n_257_76_411;
   wire n_257_76_412;
   wire n_257_76_413;
   wire n_257_76_414;
   wire n_257_76_415;
   wire n_257_76_416;
   wire n_257_76_417;
   wire n_257_76_418;
   wire n_257_76_419;
   wire n_257_76_420;
   wire n_257_76_421;
   wire n_257_76_422;
   wire n_257_76_423;
   wire n_257_76_424;
   wire n_257_76_425;
   wire n_257_76_426;
   wire n_257_76_427;
   wire n_257_76_428;
   wire n_257_76_429;
   wire n_257_76_430;
   wire n_257_76_431;
   wire n_257_76_432;
   wire n_257_76_433;
   wire n_257_76_434;
   wire n_257_76_435;
   wire n_257_76_436;
   wire n_257_76_437;
   wire n_257_76_438;
   wire n_257_76_439;
   wire n_257_76_440;
   wire n_257_76_441;
   wire n_257_76_442;
   wire n_257_76_443;
   wire n_257_76_444;
   wire n_257_76_445;
   wire n_257_76_446;
   wire n_257_76_447;
   wire n_257_76_448;
   wire n_257_76_449;
   wire n_257_76_450;
   wire n_257_76_451;
   wire n_257_76_452;
   wire n_257_76_453;
   wire n_257_76_454;
   wire n_257_76_455;
   wire n_257_76_456;
   wire n_257_76_457;
   wire n_257_76_458;
   wire n_257_76_459;
   wire n_257_76_460;
   wire n_257_76_461;
   wire n_257_76_462;
   wire n_257_76_463;
   wire n_257_76_464;
   wire n_257_76_465;
   wire n_257_76_466;
   wire n_257_76_467;
   wire n_257_76_468;
   wire n_257_76_469;
   wire n_257_76_470;
   wire n_257_76_471;
   wire n_257_76_472;
   wire n_257_76_473;
   wire n_257_76_474;
   wire n_257_76_475;
   wire n_257_76_476;
   wire n_257_76_477;
   wire n_257_76_478;
   wire n_257_76_479;
   wire n_257_76_480;
   wire n_257_76_481;
   wire n_257_76_482;
   wire n_257_76_483;
   wire n_257_76_484;
   wire n_257_76_485;
   wire n_257_76_486;
   wire n_257_76_487;
   wire n_257_76_488;
   wire n_257_76_489;
   wire n_257_76_490;
   wire n_257_76_491;
   wire n_257_76_492;
   wire n_257_76_493;
   wire n_257_76_494;
   wire n_257_76_495;
   wire n_257_76_496;
   wire n_257_76_497;
   wire n_257_76_498;
   wire n_257_76_499;
   wire n_257_76_500;
   wire n_257_76_501;
   wire n_257_76_502;
   wire n_257_76_503;
   wire n_257_76_504;
   wire n_257_76_505;
   wire n_257_76_506;
   wire n_257_76_507;
   wire n_257_76_508;
   wire n_257_76_509;
   wire n_257_76_510;
   wire n_257_76_511;
   wire n_257_76_512;
   wire n_257_76_513;
   wire n_257_76_514;
   wire n_257_76_515;
   wire n_257_76_516;
   wire n_257_76_517;
   wire n_257_76_518;
   wire n_257_76_519;
   wire n_257_76_520;
   wire n_257_76_521;
   wire n_257_76_522;
   wire n_257_76_523;
   wire n_257_76_524;
   wire n_257_76_525;
   wire n_257_76_526;
   wire n_257_76_527;
   wire n_257_76_528;
   wire n_257_76_529;
   wire n_257_76_530;
   wire n_257_76_531;
   wire n_257_76_532;
   wire n_257_76_533;
   wire n_257_76_534;
   wire n_257_76_535;
   wire n_257_76_536;
   wire n_257_76_537;
   wire n_257_76_538;
   wire n_257_76_539;
   wire n_257_76_540;
   wire n_257_76_541;
   wire n_257_76_542;
   wire n_257_76_543;
   wire n_257_76_544;
   wire n_257_76_545;
   wire n_257_76_546;
   wire n_257_76_547;
   wire n_257_76_548;
   wire n_257_76_549;
   wire n_257_76_550;
   wire n_257_76_551;
   wire n_257_76_552;
   wire n_257_76_553;
   wire n_257_76_554;
   wire n_257_76_555;
   wire n_257_76_556;
   wire n_257_76_557;
   wire n_257_76_558;
   wire n_257_76_559;
   wire n_257_76_560;
   wire n_257_76_561;
   wire n_257_76_562;
   wire n_257_76_563;
   wire n_257_76_564;
   wire n_257_76_565;
   wire n_257_76_566;
   wire n_257_76_567;
   wire n_257_76_568;
   wire n_257_76_569;
   wire n_257_76_570;
   wire n_257_76_571;
   wire n_257_76_572;
   wire n_257_76_573;
   wire n_257_76_574;
   wire n_257_76_575;
   wire n_257_76_576;
   wire n_257_76_577;
   wire n_257_76_578;
   wire n_257_76_579;
   wire n_257_76_580;
   wire n_257_76_581;
   wire n_257_76_582;
   wire n_257_76_583;
   wire n_257_76_584;
   wire n_257_76_585;
   wire n_257_76_586;
   wire n_257_76_587;
   wire n_257_76_588;
   wire n_257_76_589;
   wire n_257_76_590;
   wire n_257_76_591;
   wire n_257_76_592;
   wire n_257_76_593;
   wire n_257_76_594;
   wire n_257_76_595;
   wire n_257_76_596;
   wire n_257_76_597;
   wire n_257_76_598;
   wire n_257_76_599;
   wire n_257_76_600;
   wire n_257_76_601;
   wire n_257_76_602;
   wire n_257_76_603;
   wire n_257_76_604;
   wire n_257_76_605;
   wire n_257_76_606;
   wire n_257_76_607;
   wire n_257_76_608;
   wire n_257_76_609;
   wire n_257_76_610;
   wire n_257_76_611;
   wire n_257_76_612;
   wire n_257_76_613;
   wire n_257_76_614;
   wire n_257_76_615;
   wire n_257_76_616;
   wire n_257_76_617;
   wire n_257_76_618;
   wire n_257_76_619;
   wire n_257_76_620;
   wire n_257_76_621;
   wire n_257_76_622;
   wire n_257_76_623;
   wire n_257_76_624;
   wire n_257_76_625;
   wire n_257_76_626;
   wire n_257_76_627;
   wire n_257_76_628;
   wire n_257_76_629;
   wire n_257_76_630;
   wire n_257_76_631;
   wire n_257_76_632;
   wire n_257_76_633;
   wire n_257_76_634;
   wire n_257_76_635;
   wire n_257_76_636;
   wire n_257_76_637;
   wire n_257_76_638;
   wire n_257_76_639;
   wire n_257_76_640;
   wire n_257_76_641;
   wire n_257_76_642;
   wire n_257_76_643;
   wire n_257_76_644;
   wire n_257_76_645;
   wire n_257_76_646;
   wire n_257_76_647;
   wire n_257_76_648;
   wire n_257_76_649;
   wire n_257_76_650;
   wire n_257_76_651;
   wire n_257_76_652;
   wire n_257_76_653;
   wire n_257_76_654;
   wire n_257_76_655;
   wire n_257_76_656;
   wire n_257_76_657;
   wire n_257_76_658;
   wire n_257_76_659;
   wire n_257_76_660;
   wire n_257_76_661;
   wire n_257_76_662;
   wire n_257_76_663;
   wire n_257_76_664;
   wire n_257_76_665;
   wire n_257_76_666;
   wire n_257_76_667;
   wire n_257_76_668;
   wire n_257_76_669;
   wire n_257_76_670;
   wire n_257_76_671;
   wire n_257_76_672;
   wire n_257_76_673;
   wire n_257_76_674;
   wire n_257_76_675;
   wire n_257_76_676;
   wire n_257_76_677;
   wire n_257_76_678;
   wire n_257_76_679;
   wire n_257_76_680;
   wire n_257_76_681;
   wire n_257_76_682;
   wire n_257_76_683;
   wire n_257_76_684;
   wire n_257_76_685;
   wire n_257_76_686;
   wire n_257_76_687;
   wire n_257_76_688;
   wire n_257_76_689;
   wire n_257_76_690;
   wire n_257_76_691;
   wire n_257_76_692;
   wire n_257_76_693;
   wire n_257_76_694;
   wire n_257_76_695;
   wire n_257_76_696;
   wire n_257_76_697;
   wire n_257_76_698;
   wire n_257_76_699;
   wire n_257_76_700;
   wire n_257_76_701;
   wire n_257_76_702;
   wire n_257_76_703;
   wire n_257_76_704;
   wire n_257_76_705;
   wire n_257_76_706;
   wire n_257_76_707;
   wire n_257_76_708;
   wire n_257_76_709;
   wire n_257_76_710;
   wire n_257_76_711;
   wire n_257_76_712;
   wire n_257_76_713;
   wire n_257_76_714;
   wire n_257_76_715;
   wire n_257_76_716;
   wire n_257_76_717;
   wire n_257_76_718;
   wire n_257_76_719;
   wire n_257_76_720;
   wire n_257_76_721;
   wire n_257_76_722;
   wire n_257_76_723;
   wire n_257_76_724;
   wire n_257_76_725;
   wire n_257_76_726;
   wire n_257_76_727;
   wire n_257_76_728;
   wire n_257_76_729;
   wire n_257_76_730;
   wire n_257_76_731;
   wire n_257_76_732;
   wire n_257_76_733;
   wire n_257_76_734;
   wire n_257_76_735;
   wire n_257_76_736;
   wire n_257_76_737;
   wire n_257_76_738;
   wire n_257_76_739;
   wire n_257_76_740;
   wire n_257_76_741;
   wire n_257_76_742;
   wire n_257_76_743;
   wire n_257_76_744;
   wire n_257_76_745;
   wire n_257_76_746;
   wire n_257_76_747;
   wire n_257_76_748;
   wire n_257_76_749;
   wire n_257_76_750;
   wire n_257_76_751;
   wire n_257_76_752;
   wire n_257_76_753;
   wire n_257_76_754;
   wire n_257_76_755;
   wire n_257_76_756;
   wire n_257_76_757;
   wire n_257_76_758;
   wire n_257_76_759;
   wire n_257_76_760;
   wire n_257_76_761;
   wire n_257_76_762;
   wire n_257_76_763;
   wire n_257_76_764;
   wire n_257_76_765;
   wire n_257_76_766;
   wire n_257_76_767;
   wire n_257_76_768;
   wire n_257_76_769;
   wire n_257_76_770;
   wire n_257_76_771;
   wire n_257_76_772;
   wire n_257_76_773;
   wire n_257_76_774;
   wire n_257_76_775;
   wire n_257_76_776;
   wire n_257_76_777;
   wire n_257_76_778;
   wire n_257_76_779;
   wire n_257_76_780;
   wire n_257_76_781;
   wire n_257_76_782;
   wire n_257_76_783;
   wire n_257_76_784;
   wire n_257_76_785;
   wire n_257_76_786;
   wire n_257_76_787;
   wire n_257_76_788;
   wire n_257_76_789;
   wire n_257_76_790;
   wire n_257_76_791;
   wire n_257_76_792;
   wire n_257_76_793;
   wire n_257_76_794;
   wire n_257_76_795;
   wire n_257_76_796;
   wire n_257_76_797;
   wire n_257_76_798;
   wire n_257_76_799;
   wire n_257_76_800;
   wire n_257_76_801;
   wire n_257_76_802;
   wire n_257_76_803;
   wire n_257_76_804;
   wire n_257_76_805;
   wire n_257_76_806;
   wire n_257_76_807;
   wire n_257_76_808;
   wire n_257_76_809;
   wire n_257_76_810;
   wire n_257_76_811;
   wire n_257_76_812;
   wire n_257_76_813;
   wire n_257_76_814;
   wire n_257_76_815;
   wire n_257_76_816;
   wire n_257_76_817;
   wire n_257_76_818;
   wire n_257_76_819;
   wire n_257_76_820;
   wire n_257_76_821;
   wire n_257_76_822;
   wire n_257_76_823;
   wire n_257_76_824;
   wire n_257_76_825;
   wire n_257_76_826;
   wire n_257_76_827;
   wire n_257_76_828;
   wire n_257_76_829;
   wire n_257_76_830;
   wire n_257_76_831;
   wire n_257_76_832;
   wire n_257_76_833;
   wire n_257_76_834;
   wire n_257_76_835;
   wire n_257_76_836;
   wire n_257_76_837;
   wire n_257_76_838;
   wire n_257_76_839;
   wire n_257_76_840;
   wire n_257_76_841;
   wire n_257_76_842;
   wire n_257_76_843;
   wire n_257_76_844;
   wire n_257_76_845;
   wire n_257_76_846;
   wire n_257_76_847;
   wire n_257_76_848;
   wire n_257_76_849;
   wire n_257_76_850;
   wire n_257_76_851;
   wire n_257_76_852;
   wire n_257_76_853;
   wire n_257_76_854;
   wire n_257_76_855;
   wire n_257_76_856;
   wire n_257_76_857;
   wire n_257_76_858;
   wire n_257_76_859;
   wire n_257_76_860;
   wire n_257_76_861;
   wire n_257_76_862;
   wire n_257_76_863;
   wire n_257_76_864;
   wire n_257_76_865;
   wire n_257_76_866;
   wire n_257_76_867;
   wire n_257_76_868;
   wire n_257_76_869;
   wire n_257_76_870;
   wire n_257_76_871;
   wire n_257_76_872;
   wire n_257_76_873;
   wire n_257_76_874;
   wire n_257_76_875;
   wire n_257_76_876;
   wire n_257_76_877;
   wire n_257_76_878;
   wire n_257_76_879;
   wire n_257_76_880;
   wire n_257_76_881;
   wire n_257_76_882;
   wire n_257_76_883;
   wire n_257_76_884;
   wire n_257_76_885;
   wire n_257_76_886;
   wire n_257_76_887;
   wire n_257_76_888;
   wire n_257_76_889;
   wire n_257_76_890;
   wire n_257_76_891;
   wire n_257_76_892;
   wire n_257_76_893;
   wire n_257_76_894;
   wire n_257_76_895;
   wire n_257_76_896;
   wire n_257_76_897;
   wire n_257_76_898;
   wire n_257_76_899;
   wire n_257_76_900;
   wire n_257_76_901;
   wire n_257_76_902;
   wire n_257_76_903;
   wire n_257_76_904;
   wire n_257_76_905;
   wire n_257_76_906;
   wire n_257_76_907;
   wire n_257_76_908;
   wire n_257_76_909;
   wire n_257_76_910;
   wire n_257_76_911;
   wire n_257_76_912;
   wire n_257_76_913;
   wire n_257_76_914;
   wire n_257_76_915;
   wire n_257_76_916;
   wire n_257_76_917;
   wire n_257_76_918;
   wire n_257_76_919;
   wire n_257_76_920;
   wire n_257_76_921;
   wire n_257_76_922;
   wire n_257_76_923;
   wire n_257_76_924;
   wire n_257_76_925;
   wire n_257_76_926;
   wire n_257_76_927;
   wire n_257_76_928;
   wire n_257_76_929;
   wire n_257_76_930;
   wire n_257_76_931;
   wire n_257_76_932;
   wire n_257_76_933;
   wire n_257_76_934;
   wire n_257_76_935;
   wire n_257_76_936;
   wire n_257_76_937;
   wire n_257_76_938;
   wire n_257_76_939;
   wire n_257_76_940;
   wire n_257_76_941;
   wire n_257_76_942;
   wire n_257_76_943;
   wire n_257_76_944;
   wire n_257_76_945;
   wire n_257_76_946;
   wire n_257_76_947;
   wire n_257_76_948;
   wire n_257_76_949;
   wire n_257_76_950;
   wire n_257_76_951;
   wire n_257_76_952;
   wire n_257_76_953;
   wire n_257_76_954;
   wire n_257_76_955;
   wire n_257_76_956;
   wire n_257_76_957;
   wire n_257_76_958;
   wire n_257_76_959;
   wire n_257_76_960;
   wire n_257_76_961;
   wire n_257_76_962;
   wire n_257_76_963;
   wire n_257_76_964;
   wire n_257_76_965;
   wire n_257_76_966;
   wire n_257_76_967;
   wire n_257_76_968;
   wire n_257_76_969;
   wire n_257_76_970;
   wire n_257_76_971;
   wire n_257_76_972;
   wire n_257_76_973;
   wire n_257_76_974;
   wire n_257_76_975;
   wire n_257_76_976;
   wire n_257_76_977;
   wire n_257_76_978;
   wire n_257_76_979;
   wire n_257_76_980;
   wire n_257_76_981;
   wire n_257_76_982;
   wire n_257_76_983;
   wire n_257_76_984;
   wire n_257_76_985;
   wire n_257_76_986;
   wire n_257_76_987;
   wire n_257_76_988;
   wire n_257_76_989;
   wire n_257_76_990;
   wire n_257_76_991;
   wire n_257_76_992;
   wire n_257_76_993;
   wire n_257_76_994;
   wire n_257_76_995;
   wire n_257_76_996;
   wire n_257_76_997;
   wire n_257_76_998;
   wire n_257_76_999;
   wire n_257_76_1000;
   wire n_257_76_1001;
   wire n_257_76_1002;
   wire n_257_76_1003;
   wire n_257_76_1004;
   wire n_257_76_1005;
   wire n_257_76_1006;
   wire n_257_76_1007;
   wire n_257_76_1008;
   wire n_257_76_1009;
   wire n_257_76_1010;
   wire n_257_76_1011;
   wire n_257_76_1012;
   wire n_257_76_1013;
   wire n_257_76_1014;
   wire n_257_76_1015;
   wire n_257_76_1016;
   wire n_257_76_1017;
   wire n_257_76_1018;
   wire n_257_76_1019;
   wire n_257_76_1020;
   wire n_257_76_1021;
   wire n_257_76_1022;
   wire n_257_76_1023;
   wire n_257_76_1024;
   wire n_257_76_1025;
   wire n_257_76_1026;
   wire n_257_76_1027;
   wire n_257_76_1028;
   wire n_257_76_1029;
   wire n_257_76_1030;
   wire n_257_76_1031;
   wire n_257_76_1032;
   wire n_257_76_1033;
   wire n_257_76_1034;
   wire n_257_76_1035;
   wire n_257_76_1036;
   wire n_257_76_1037;
   wire n_257_76_1038;
   wire n_257_76_1039;
   wire n_257_76_1040;
   wire n_257_76_1041;
   wire n_257_76_1042;
   wire n_257_76_1043;
   wire n_257_76_1044;
   wire n_257_76_1045;
   wire n_257_76_1046;
   wire n_257_76_1047;
   wire n_257_76_1048;
   wire n_257_76_1049;
   wire n_257_76_1050;
   wire n_257_76_1051;
   wire n_257_76_1052;
   wire n_257_76_1053;
   wire n_257_76_1054;
   wire n_257_76_1055;
   wire n_257_76_1056;
   wire n_257_76_1057;
   wire n_257_76_1058;
   wire n_257_76_1059;
   wire n_257_76_1060;
   wire n_257_76_1061;
   wire n_257_76_1062;
   wire n_257_76_1063;
   wire n_257_76_1064;
   wire n_257_76_1065;
   wire n_257_76_1066;
   wire n_257_76_1067;
   wire n_257_76_1068;
   wire n_257_76_1069;
   wire n_257_76_1070;
   wire n_257_76_1071;
   wire n_257_76_1072;
   wire n_257_76_1073;
   wire n_257_76_1074;
   wire n_257_76_1075;
   wire n_257_76_1076;
   wire n_257_76_1077;
   wire n_257_76_1078;
   wire n_257_76_1079;
   wire n_257_76_1080;
   wire n_257_76_1081;
   wire n_257_76_1082;
   wire n_257_76_1083;
   wire n_257_76_1084;
   wire n_257_76_1085;
   wire n_257_76_1086;
   wire n_257_76_1087;
   wire n_257_76_1088;
   wire n_257_76_1089;
   wire n_257_76_1090;
   wire n_257_76_1091;
   wire n_257_76_1092;
   wire n_257_76_1093;
   wire n_257_76_1094;
   wire n_257_76_1095;
   wire n_257_76_1096;
   wire n_257_76_1097;
   wire n_257_76_1098;
   wire n_257_76_1099;
   wire n_257_76_1100;
   wire n_257_76_1101;
   wire n_257_76_1102;
   wire n_257_76_1103;
   wire n_257_76_1104;
   wire n_257_76_1105;
   wire n_257_76_1106;
   wire n_257_76_1107;
   wire n_257_76_1108;
   wire n_257_76_1109;
   wire n_257_76_1110;
   wire n_257_76_1111;
   wire n_257_76_1112;
   wire n_257_76_1113;
   wire n_257_76_1114;
   wire n_257_76_1115;
   wire n_257_76_1116;
   wire n_257_76_1117;
   wire n_257_76_1118;
   wire n_257_76_1119;
   wire n_257_76_1120;
   wire n_257_76_1121;
   wire n_257_76_1122;
   wire n_257_76_1123;
   wire n_257_76_1124;
   wire n_257_76_1125;
   wire n_257_76_1126;
   wire n_257_76_1127;
   wire n_257_76_1128;
   wire n_257_76_1129;
   wire n_257_76_1130;
   wire n_257_76_1131;
   wire n_257_76_1132;
   wire n_257_76_1133;
   wire n_257_76_1134;
   wire n_257_76_1135;
   wire n_257_76_1136;
   wire n_257_76_1137;
   wire n_257_76_1138;
   wire n_257_76_1139;
   wire n_257_76_1140;
   wire n_257_76_1141;
   wire n_257_76_1142;
   wire n_257_76_1143;
   wire n_257_76_1144;
   wire n_257_76_1145;
   wire n_257_76_1146;
   wire n_257_76_1147;
   wire n_257_76_1148;
   wire n_257_76_1149;
   wire n_257_76_1150;
   wire n_257_76_1151;
   wire n_257_76_1152;
   wire n_257_76_1153;
   wire n_257_76_1154;
   wire n_257_76_1155;
   wire n_257_76_1156;
   wire n_257_76_1157;
   wire n_257_76_1158;
   wire n_257_76_1159;
   wire n_257_76_1160;
   wire n_257_76_1161;
   wire n_257_76_1162;
   wire n_257_76_1163;
   wire n_257_76_1164;
   wire n_257_76_1165;
   wire n_257_76_1166;
   wire n_257_76_1167;
   wire n_257_76_1168;
   wire n_257_76_1169;
   wire n_257_76_1170;
   wire n_257_76_1171;
   wire n_257_76_1172;
   wire n_257_76_1173;
   wire n_257_76_1174;
   wire n_257_76_1175;
   wire n_257_76_1176;
   wire n_257_76_1177;
   wire n_257_76_1178;
   wire n_257_76_1179;
   wire n_257_76_1180;
   wire n_257_76_1181;
   wire n_257_76_1182;
   wire n_257_76_1183;
   wire n_257_76_1184;
   wire n_257_76_1185;
   wire n_257_76_1186;
   wire n_257_76_1187;
   wire n_257_76_1188;
   wire n_257_76_1189;
   wire n_257_76_1190;
   wire n_257_76_1191;
   wire n_257_76_1192;
   wire n_257_76_1193;
   wire n_257_76_1194;
   wire n_257_76_1195;
   wire n_257_76_1196;
   wire n_257_76_1197;
   wire n_257_76_1198;
   wire n_257_76_1199;
   wire n_257_76_1200;
   wire n_257_76_1201;
   wire n_257_76_1202;
   wire n_257_76_1203;
   wire n_257_76_1204;
   wire n_257_76_1205;
   wire n_257_76_1206;
   wire n_257_76_1207;
   wire n_257_76_1208;
   wire n_257_76_1209;
   wire n_257_76_1210;
   wire n_257_76_1211;
   wire n_257_76_1212;
   wire n_257_76_1213;
   wire n_257_76_1214;
   wire n_257_76_1215;
   wire n_257_76_1216;
   wire n_257_76_1217;
   wire n_257_76_1218;
   wire n_257_76_1219;
   wire n_257_76_1220;
   wire n_257_76_1221;
   wire n_257_76_1222;
   wire n_257_76_1223;
   wire n_257_76_1224;
   wire n_257_76_1225;
   wire n_257_76_1226;
   wire n_257_76_1227;
   wire n_257_76_1228;
   wire n_257_76_1229;
   wire n_257_76_1230;
   wire n_257_76_1231;
   wire n_257_76_1232;
   wire n_257_76_1233;
   wire n_257_76_1234;
   wire n_257_76_1235;
   wire n_257_76_1236;
   wire n_257_76_1237;
   wire n_257_76_1238;
   wire n_257_76_1239;
   wire n_257_76_1240;
   wire n_257_76_1241;
   wire n_257_76_1242;
   wire n_257_76_1243;
   wire n_257_76_1244;
   wire n_257_76_1245;
   wire n_257_76_1246;
   wire n_257_76_1247;
   wire n_257_76_1248;
   wire n_257_76_1249;
   wire n_257_76_1250;
   wire n_257_76_1251;
   wire n_257_76_1252;
   wire n_257_76_1253;
   wire n_257_76_1254;
   wire n_257_76_1255;
   wire n_257_76_1256;
   wire n_257_76_1257;
   wire n_257_76_1258;
   wire n_257_76_1259;
   wire n_257_76_1260;
   wire n_257_76_1261;
   wire n_257_76_1262;
   wire n_257_76_1263;
   wire n_257_76_1264;
   wire n_257_76_1265;
   wire n_257_76_1266;
   wire n_257_76_1267;
   wire n_257_76_1268;
   wire n_257_76_1269;
   wire n_257_76_1270;
   wire n_257_76_1271;
   wire n_257_76_1272;
   wire n_257_76_1273;
   wire n_257_76_1274;
   wire n_257_76_1275;
   wire n_257_76_1276;
   wire n_257_76_1277;
   wire n_257_76_1278;
   wire n_257_76_1279;
   wire n_257_76_1280;
   wire n_257_76_1281;
   wire n_257_76_1282;
   wire n_257_76_1283;
   wire n_257_76_1284;
   wire n_257_76_1285;
   wire n_257_76_1286;
   wire n_257_76_1287;
   wire n_257_76_1288;
   wire n_257_76_1289;
   wire n_257_76_1290;
   wire n_257_76_1291;
   wire n_257_76_1292;
   wire n_257_76_1293;
   wire n_257_76_1294;
   wire n_257_76_1295;
   wire n_257_76_1296;
   wire n_257_76_1297;
   wire n_257_76_1298;
   wire n_257_76_1299;
   wire n_257_76_1300;
   wire n_257_76_1301;
   wire n_257_76_1302;
   wire n_257_76_1303;
   wire n_257_76_1304;
   wire n_257_76_1305;
   wire n_257_76_1306;
   wire n_257_76_1307;
   wire n_257_76_1308;
   wire n_257_76_1309;
   wire n_257_76_1310;
   wire n_257_76_1311;
   wire n_257_76_1312;
   wire n_257_76_1313;
   wire n_257_76_1314;
   wire n_257_76_1315;
   wire n_257_76_1316;
   wire n_257_76_1317;
   wire n_257_76_1318;
   wire n_257_76_1319;
   wire n_257_76_1320;
   wire n_257_76_1321;
   wire n_257_76_1322;
   wire n_257_76_1323;
   wire n_257_76_1324;
   wire n_257_76_1325;
   wire n_257_76_1326;
   wire n_257_76_1327;
   wire n_257_76_1328;
   wire n_257_76_1329;
   wire n_257_76_1330;
   wire n_257_76_1331;
   wire n_257_76_1332;
   wire n_257_76_1333;
   wire n_257_76_1334;
   wire n_257_76_1335;
   wire n_257_76_1336;
   wire n_257_76_1337;
   wire n_257_76_1338;
   wire n_257_76_1339;
   wire n_257_76_1340;
   wire n_257_76_1341;
   wire n_257_76_1342;
   wire n_257_76_1343;
   wire n_257_76_1344;
   wire n_257_76_1345;
   wire n_257_76_1346;
   wire n_257_76_1347;
   wire n_257_76_1348;
   wire n_257_76_1349;
   wire n_257_76_1350;
   wire n_257_76_1351;
   wire n_257_76_1352;
   wire n_257_76_1353;
   wire n_257_76_1354;
   wire n_257_76_1355;
   wire n_257_76_1356;
   wire n_257_76_1357;
   wire n_257_76_1358;
   wire n_257_76_1359;
   wire n_257_76_1360;
   wire n_257_76_1361;
   wire n_257_76_1362;
   wire n_257_76_1363;
   wire n_257_76_1364;
   wire n_257_76_1365;
   wire n_257_76_1366;
   wire n_257_76_1367;
   wire n_257_76_1368;
   wire n_257_76_1369;
   wire n_257_76_1370;
   wire n_257_76_1371;
   wire n_257_76_1372;
   wire n_257_76_1373;
   wire n_257_76_1374;
   wire n_257_76_1375;
   wire n_257_76_1376;
   wire n_257_76_1377;
   wire n_257_76_1378;
   wire n_257_76_1379;
   wire n_257_76_1380;
   wire n_257_76_1381;
   wire n_257_76_1382;
   wire n_257_76_1383;
   wire n_257_76_1384;
   wire n_257_76_1385;
   wire n_257_76_1386;
   wire n_257_76_1387;
   wire n_257_76_1388;
   wire n_257_76_1389;
   wire n_257_76_1390;
   wire n_257_76_1391;
   wire n_257_76_1392;
   wire n_257_76_1393;
   wire n_257_76_1394;
   wire n_257_76_1395;
   wire n_257_76_1396;
   wire n_257_76_1397;
   wire n_257_76_1398;
   wire n_257_76_1399;
   wire n_257_76_1400;
   wire n_257_76_1401;
   wire n_257_76_1402;
   wire n_257_76_1403;
   wire n_257_76_1404;
   wire n_257_76_1405;
   wire n_257_76_1406;
   wire n_257_76_1407;
   wire n_257_76_1408;
   wire n_257_76_1409;
   wire n_257_76_1410;
   wire n_257_76_1411;
   wire n_257_76_1412;
   wire n_257_76_1413;
   wire n_257_76_1414;
   wire n_257_76_1415;
   wire n_257_76_1416;
   wire n_257_76_1417;
   wire n_257_76_1418;
   wire n_257_76_1419;
   wire n_257_76_1420;
   wire n_257_76_1421;
   wire n_257_76_1422;
   wire n_257_76_1423;
   wire n_257_76_1424;
   wire n_257_76_1425;
   wire n_257_76_1426;
   wire n_257_76_1427;
   wire n_257_76_1428;
   wire n_257_76_1429;
   wire n_257_76_1430;
   wire n_257_76_1431;
   wire n_257_76_1432;
   wire n_257_76_1433;
   wire n_257_76_1434;
   wire n_257_76_1435;
   wire n_257_76_1436;
   wire n_257_76_1437;
   wire n_257_76_1438;
   wire n_257_76_1439;
   wire n_257_76_1440;
   wire n_257_76_1441;
   wire n_257_76_1442;
   wire n_257_76_1443;
   wire n_257_76_1444;
   wire n_257_76_1445;
   wire n_257_76_1446;
   wire n_257_76_1447;
   wire n_257_76_1448;
   wire n_257_76_1449;
   wire n_257_76_1450;
   wire n_257_76_1451;
   wire n_257_76_1452;
   wire n_257_76_1453;
   wire n_257_76_1454;
   wire n_257_76_1455;
   wire n_257_76_1456;
   wire n_257_76_1457;
   wire n_257_76_1458;
   wire n_257_76_1459;
   wire n_257_76_1460;
   wire n_257_76_1461;
   wire n_257_76_1462;
   wire n_257_76_1463;
   wire n_257_76_1464;
   wire n_257_76_1465;
   wire n_257_76_1466;
   wire n_257_76_1467;
   wire n_257_76_1468;
   wire n_257_76_1469;
   wire n_257_76_1470;
   wire n_257_76_1471;
   wire n_257_76_1472;
   wire n_257_76_1473;
   wire n_257_76_1474;
   wire n_257_76_1475;
   wire n_257_76_1476;
   wire n_257_76_1477;
   wire n_257_76_1478;
   wire n_257_76_1479;
   wire n_257_76_1480;
   wire n_257_76_1481;
   wire n_257_76_1482;
   wire n_257_76_1483;
   wire n_257_76_1484;
   wire n_257_76_1485;
   wire n_257_76_1486;
   wire n_257_76_1487;
   wire n_257_76_1488;
   wire n_257_76_1489;
   wire n_257_76_1490;
   wire n_257_76_1491;
   wire n_257_76_1492;
   wire n_257_76_1493;
   wire n_257_76_1494;
   wire n_257_76_1495;
   wire n_257_76_1496;
   wire n_257_76_1497;
   wire n_257_76_1498;
   wire n_257_76_1499;
   wire n_257_76_1500;
   wire n_257_76_1501;
   wire n_257_76_1502;
   wire n_257_76_1503;
   wire n_257_76_1504;
   wire n_257_76_1505;
   wire n_257_76_1506;
   wire n_257_76_1507;
   wire n_257_76_1508;
   wire n_257_76_1509;
   wire n_257_76_1510;
   wire n_257_76_1511;
   wire n_257_76_1512;
   wire n_257_76_1513;
   wire n_257_76_1514;
   wire n_257_76_1515;
   wire n_257_76_1516;
   wire n_257_76_1517;
   wire n_257_76_1518;
   wire n_257_76_1519;
   wire n_257_76_1520;
   wire n_257_76_1521;
   wire n_257_76_1522;
   wire n_257_76_1523;
   wire n_257_76_1524;
   wire n_257_76_1525;
   wire n_257_76_1526;
   wire n_257_76_1527;
   wire n_257_76_1528;
   wire n_257_76_1529;
   wire n_257_76_1530;
   wire n_257_76_1531;
   wire n_257_76_1532;
   wire n_257_76_1533;
   wire n_257_76_1534;
   wire n_257_76_1535;
   wire n_257_76_1536;
   wire n_257_76_1537;
   wire n_257_76_1538;
   wire n_257_76_1539;
   wire n_257_76_1540;
   wire n_257_76_1541;
   wire n_257_76_1542;
   wire n_257_76_1543;
   wire n_257_76_1544;
   wire n_257_76_1545;
   wire n_257_76_1546;
   wire n_257_76_1547;
   wire n_257_76_1548;
   wire n_257_76_1549;
   wire n_257_76_1550;
   wire n_257_76_1551;
   wire n_257_76_1552;
   wire n_257_76_1553;
   wire n_257_76_1554;
   wire n_257_76_1555;
   wire n_257_76_1556;
   wire n_257_76_1557;
   wire n_257_76_1558;
   wire n_257_76_1559;
   wire n_257_76_1560;
   wire n_257_76_1561;
   wire n_257_76_1562;
   wire n_257_76_1563;
   wire n_257_76_1564;
   wire n_257_76_1565;
   wire n_257_76_1566;
   wire n_257_76_1567;
   wire n_257_76_1568;
   wire n_257_76_1569;
   wire n_257_76_1570;
   wire n_257_76_1571;
   wire n_257_76_1572;
   wire n_257_76_1573;
   wire n_257_76_1574;
   wire n_257_76_1575;
   wire n_257_76_1576;
   wire n_257_76_1577;
   wire n_257_76_1578;
   wire n_257_76_1579;
   wire n_257_76_1580;
   wire n_257_76_1581;
   wire n_257_76_1582;
   wire n_257_76_1583;
   wire n_257_76_1584;
   wire n_257_76_1585;
   wire n_257_76_1586;
   wire n_257_76_1587;
   wire n_257_76_1588;
   wire n_257_76_1589;
   wire n_257_76_1590;
   wire n_257_76_1591;
   wire n_257_76_1592;
   wire n_257_76_1593;
   wire n_257_76_1594;
   wire n_257_76_1595;
   wire n_257_76_1596;
   wire n_257_76_1597;
   wire n_257_76_1598;
   wire n_257_76_1599;
   wire n_257_76_1600;
   wire n_257_76_1601;
   wire n_257_76_1602;
   wire n_257_76_1603;
   wire n_257_76_1604;
   wire n_257_76_1605;
   wire n_257_76_1606;
   wire n_257_76_1607;
   wire n_257_76_1608;
   wire n_257_76_1609;
   wire n_257_76_1610;
   wire n_257_76_1611;
   wire n_257_76_1612;
   wire n_257_76_1613;
   wire n_257_76_1614;
   wire n_257_76_1615;
   wire n_257_76_1616;
   wire n_257_76_1617;
   wire n_257_76_1618;
   wire n_257_76_1619;
   wire n_257_76_1620;
   wire n_257_76_1621;
   wire n_257_76_1622;
   wire n_257_76_1623;
   wire n_257_76_1624;
   wire n_257_76_1625;
   wire n_257_76_1626;
   wire n_257_76_1627;
   wire n_257_76_1628;
   wire n_257_76_1629;
   wire n_257_76_1630;
   wire n_257_76_1631;
   wire n_257_76_1632;
   wire n_257_76_1633;
   wire n_257_76_1634;
   wire n_257_76_1635;
   wire n_257_76_1636;
   wire n_257_76_1637;
   wire n_257_76_1638;
   wire n_257_76_1639;
   wire n_257_76_1640;
   wire n_257_76_1641;
   wire n_257_76_1642;
   wire n_257_76_1643;
   wire n_257_76_1644;
   wire n_257_76_1645;
   wire n_257_76_1646;
   wire n_257_76_1647;
   wire n_257_76_1648;
   wire n_257_76_1649;
   wire n_257_76_1650;
   wire n_257_76_1651;
   wire n_257_76_1652;
   wire n_257_76_1653;
   wire n_257_76_1654;
   wire n_257_76_1655;
   wire n_257_76_1656;
   wire n_257_76_1657;
   wire n_257_76_1658;
   wire n_257_76_1659;
   wire n_257_76_1660;
   wire n_257_76_1661;
   wire n_257_76_1662;
   wire n_257_76_1663;
   wire n_257_76_1664;
   wire n_257_76_1665;
   wire n_257_76_1666;
   wire n_257_76_1667;
   wire n_257_76_1668;
   wire n_257_76_1669;
   wire n_257_76_1670;
   wire n_257_76_1671;
   wire n_257_76_1672;
   wire n_257_76_1673;
   wire n_257_76_1674;
   wire n_257_76_1675;
   wire n_257_76_1676;
   wire n_257_76_1677;
   wire n_257_76_1678;
   wire n_257_76_1679;
   wire n_257_76_1680;
   wire n_257_76_1681;
   wire n_257_76_1682;
   wire n_257_76_1683;
   wire n_257_76_1684;
   wire n_257_76_1685;
   wire n_257_76_1686;
   wire n_257_76_1687;
   wire n_257_76_1688;
   wire n_257_76_1689;
   wire n_257_76_1690;
   wire n_257_76_1691;
   wire n_257_76_1692;
   wire n_257_76_1693;
   wire n_257_76_1694;
   wire n_257_76_1695;
   wire n_257_76_1696;
   wire n_257_76_1697;
   wire n_257_76_1698;
   wire n_257_76_1699;
   wire n_257_76_1700;
   wire n_257_76_1701;
   wire n_257_76_1702;
   wire n_257_76_1703;
   wire n_257_76_1704;
   wire n_257_76_1705;
   wire n_257_76_1706;
   wire n_257_76_1707;
   wire n_257_76_1708;
   wire n_257_76_1709;
   wire n_257_76_1710;
   wire n_257_76_1711;
   wire n_257_76_1712;
   wire n_257_76_1713;
   wire n_257_76_1714;
   wire n_257_76_1715;
   wire n_257_76_1716;
   wire n_257_76_1717;
   wire n_257_76_1718;
   wire n_257_76_1719;
   wire n_257_76_1720;
   wire n_257_76_1721;
   wire n_257_76_1722;
   wire n_257_76_1723;
   wire n_257_76_1724;
   wire n_257_76_1725;
   wire n_257_76_1726;
   wire n_257_76_1727;
   wire n_257_76_1728;
   wire n_257_76_1729;
   wire n_257_76_1730;
   wire n_257_76_1731;
   wire n_257_76_1732;
   wire n_257_76_1733;
   wire n_257_76_1734;
   wire n_257_76_1735;
   wire n_257_76_1736;
   wire n_257_76_1737;
   wire n_257_76_1738;
   wire n_257_76_1739;
   wire n_257_76_1740;
   wire n_257_76_1741;
   wire n_257_76_1742;
   wire n_257_76_1743;
   wire n_257_76_1744;
   wire n_257_76_1745;
   wire n_257_76_1746;
   wire n_257_76_1747;
   wire n_257_76_1748;
   wire n_257_76_1749;
   wire n_257_76_1750;
   wire n_257_76_1751;
   wire n_257_76_1752;
   wire n_257_76_1753;
   wire n_257_76_1754;
   wire n_257_76_1755;
   wire n_257_76_1756;
   wire n_257_76_1757;
   wire n_257_76_1758;
   wire n_257_76_1759;
   wire n_257_76_1760;
   wire n_257_76_1761;
   wire n_257_76_1762;
   wire n_257_76_1763;
   wire n_257_76_1764;
   wire n_257_76_1765;
   wire n_257_76_1766;
   wire n_257_76_1767;
   wire n_257_76_1768;
   wire n_257_76_1769;
   wire n_257_76_1770;
   wire n_257_76_1771;
   wire n_257_76_1772;
   wire n_257_76_1773;
   wire n_257_76_1774;
   wire n_257_76_1775;
   wire n_257_76_1776;
   wire n_257_76_1777;
   wire n_257_76_1778;
   wire n_257_76_1779;
   wire n_257_76_1780;
   wire n_257_76_1781;
   wire n_257_76_1782;
   wire n_257_76_1783;
   wire n_257_76_1784;
   wire n_257_76_1785;
   wire n_257_76_1786;
   wire n_257_76_1787;
   wire n_257_76_1788;
   wire n_257_76_1789;
   wire n_257_76_1790;
   wire n_257_76_1791;
   wire n_257_76_1792;
   wire n_257_76_1793;
   wire n_257_76_1794;
   wire n_257_76_1795;
   wire n_257_76_1796;
   wire n_257_76_1797;
   wire n_257_76_1798;
   wire n_257_76_1799;
   wire n_257_76_1800;
   wire n_257_76_1801;
   wire n_257_76_1802;
   wire n_257_76_1803;
   wire n_257_76_1804;
   wire n_257_76_1805;
   wire n_257_76_1806;
   wire n_257_76_1807;
   wire n_257_76_1808;
   wire n_257_76_1809;
   wire n_257_76_1810;
   wire n_257_76_1811;
   wire n_257_76_1812;
   wire n_257_76_1813;
   wire n_257_76_1814;
   wire n_257_76_1815;
   wire n_257_76_1816;
   wire n_257_76_1817;
   wire n_257_76_1818;
   wire n_257_76_1819;
   wire n_257_76_1820;
   wire n_257_76_1821;
   wire n_257_76_1822;
   wire n_257_76_1823;
   wire n_257_76_1824;
   wire n_257_76_1825;
   wire n_257_76_1826;
   wire n_257_76_1827;
   wire n_257_76_1828;
   wire n_257_76_1829;
   wire n_257_76_1830;
   wire n_257_76_1831;
   wire n_257_76_1832;
   wire n_257_76_1833;
   wire n_257_76_1834;
   wire n_257_76_1835;
   wire n_257_76_1836;
   wire n_257_76_1837;
   wire n_257_76_1838;
   wire n_257_76_1839;
   wire n_257_76_1840;
   wire n_257_76_1841;
   wire n_257_76_1842;
   wire n_257_76_1843;
   wire n_257_76_1844;
   wire n_257_76_1845;
   wire n_257_76_1846;
   wire n_257_76_1847;
   wire n_257_76_1848;
   wire n_257_76_1849;
   wire n_257_76_1850;
   wire n_257_76_1851;
   wire n_257_76_1852;
   wire n_257_76_1853;
   wire n_257_76_1854;
   wire n_257_76_1855;
   wire n_257_76_1856;
   wire n_257_76_1857;
   wire n_257_76_1858;
   wire n_257_76_1859;
   wire n_257_76_1860;
   wire n_257_76_1861;
   wire n_257_76_1862;
   wire n_257_76_1863;
   wire n_257_76_1864;
   wire n_257_76_1865;
   wire n_257_76_1866;
   wire n_257_76_1867;
   wire n_257_76_1868;
   wire n_257_76_1869;
   wire n_257_76_1870;
   wire n_257_76_1871;
   wire n_257_76_1872;
   wire n_257_76_1873;
   wire n_257_76_1874;
   wire n_257_76_1875;
   wire n_257_76_1876;
   wire n_257_76_1877;
   wire n_257_76_1878;
   wire n_257_76_1879;
   wire n_257_76_1880;
   wire n_257_76_1881;
   wire n_257_76_1882;
   wire n_257_76_1883;
   wire n_257_76_1884;
   wire n_257_76_1885;
   wire n_257_76_1886;
   wire n_257_76_1887;
   wire n_257_76_1888;
   wire n_257_76_1889;
   wire n_257_76_1890;
   wire n_257_76_1891;
   wire n_257_76_1892;
   wire n_257_76_1893;
   wire n_257_76_1894;
   wire n_257_76_1895;
   wire n_257_76_1896;
   wire n_257_76_1897;
   wire n_257_76_1898;
   wire n_257_76_1899;
   wire n_257_76_1900;
   wire n_257_76_1901;
   wire n_257_76_1902;
   wire n_257_76_1903;
   wire n_257_76_1904;
   wire n_257_76_1905;
   wire n_257_76_1906;
   wire n_257_76_1907;
   wire n_257_76_1908;
   wire n_257_76_1909;
   wire n_257_76_1910;
   wire n_257_76_1911;
   wire n_257_76_1912;
   wire n_257_76_1913;
   wire n_257_76_1914;
   wire n_257_76_1915;
   wire n_257_76_1916;
   wire n_257_76_1917;
   wire n_257_76_1918;
   wire n_257_76_1919;
   wire n_257_76_1920;
   wire n_257_76_1921;
   wire n_257_76_1922;
   wire n_257_76_1923;
   wire n_257_76_1924;
   wire n_257_76_1925;
   wire n_257_76_1926;
   wire n_257_76_1927;
   wire n_257_76_1928;
   wire n_257_76_1929;
   wire n_257_76_1930;
   wire n_257_76_1931;
   wire n_257_76_1932;
   wire n_257_76_1933;
   wire n_257_76_1934;
   wire n_257_76_1935;
   wire n_257_76_1936;
   wire n_257_76_1937;
   wire n_257_76_1938;
   wire n_257_76_1939;
   wire n_257_76_1940;
   wire n_257_76_1941;
   wire n_257_76_1942;
   wire n_257_76_1943;
   wire n_257_76_1944;
   wire n_257_76_1945;
   wire n_257_76_1946;
   wire n_257_76_1947;
   wire n_257_76_1948;
   wire n_257_76_1949;
   wire n_257_76_1950;
   wire n_257_76_1951;
   wire n_257_76_1952;
   wire n_257_76_1953;
   wire n_257_76_1954;
   wire n_257_76_1955;
   wire n_257_76_1956;
   wire n_257_76_1957;
   wire n_257_76_1958;
   wire n_257_76_1959;
   wire n_257_76_1960;
   wire n_257_76_1961;
   wire n_257_76_1962;
   wire n_257_76_1963;
   wire n_257_76_1964;
   wire n_257_76_1965;
   wire n_257_76_1966;
   wire n_257_76_1967;
   wire n_257_76_1968;
   wire n_257_76_1969;
   wire n_257_76_1970;
   wire n_257_76_1971;
   wire n_257_76_1972;
   wire n_257_76_1973;
   wire n_257_76_1974;
   wire n_257_76_1975;
   wire n_257_76_1976;
   wire n_257_76_1977;
   wire n_257_76_1978;
   wire n_257_76_1979;
   wire n_257_76_1980;
   wire n_257_76_1981;
   wire n_257_76_1982;
   wire n_257_76_1983;
   wire n_257_76_1984;
   wire n_257_76_1985;
   wire n_257_76_1986;
   wire n_257_76_1987;
   wire n_257_76_1988;
   wire n_257_76_1989;
   wire n_257_76_1990;
   wire n_257_76_1991;
   wire n_257_76_1992;
   wire n_257_76_1993;
   wire n_257_76_1994;
   wire n_257_76_1995;
   wire n_257_76_1996;
   wire n_257_76_1997;
   wire n_257_76_1998;
   wire n_257_76_1999;
   wire n_257_76_2000;
   wire n_257_76_2001;
   wire n_257_76_2002;
   wire n_257_76_2003;
   wire n_257_76_2004;
   wire n_257_76_2005;
   wire n_257_76_2006;
   wire n_257_76_2007;
   wire n_257_76_2008;
   wire n_257_76_2009;
   wire n_257_76_2010;
   wire n_257_76_2011;
   wire n_257_76_2012;
   wire n_257_76_2013;
   wire n_257_76_2014;
   wire n_257_76_2015;
   wire n_257_76_2016;
   wire n_257_76_2017;
   wire n_257_76_2018;
   wire n_257_76_2019;
   wire n_257_76_2020;
   wire n_257_76_2021;
   wire n_257_76_2022;
   wire n_257_76_2023;
   wire n_257_76_2024;
   wire n_257_76_2025;
   wire n_257_76_2026;
   wire n_257_76_2027;
   wire n_257_76_2028;
   wire n_257_76_2029;
   wire n_257_76_2030;
   wire n_257_76_2031;
   wire n_257_76_2032;
   wire n_257_76_2033;
   wire n_257_76_2034;
   wire n_257_76_2035;
   wire n_257_76_2036;
   wire n_257_76_2037;
   wire n_257_76_2038;
   wire n_257_76_2039;
   wire n_257_76_2040;
   wire n_257_76_2041;
   wire n_257_76_2042;
   wire n_257_76_2043;
   wire n_257_76_2044;
   wire n_257_76_2045;
   wire n_257_76_2046;
   wire n_257_76_2047;
   wire n_257_76_2048;
   wire n_257_76_2049;
   wire n_257_76_2050;
   wire n_257_76_2051;
   wire n_257_76_2052;
   wire n_257_76_2053;
   wire n_257_76_2054;
   wire n_257_76_2055;
   wire n_257_76_2056;
   wire n_257_76_2057;
   wire n_257_76_2058;
   wire n_257_76_2059;
   wire n_257_76_2060;
   wire n_257_76_2061;
   wire n_257_76_2062;
   wire n_257_76_2063;
   wire n_257_76_2064;
   wire n_257_76_2065;
   wire n_257_76_2066;
   wire n_257_76_2067;
   wire n_257_76_2068;
   wire n_257_76_2069;
   wire n_257_76_2070;
   wire n_257_76_2071;
   wire n_257_76_2072;
   wire n_257_76_2073;
   wire n_257_76_2074;
   wire n_257_76_2075;
   wire n_257_76_2076;
   wire n_257_76_2077;
   wire n_257_76_2078;
   wire n_257_76_2079;
   wire n_257_76_2080;
   wire n_257_76_2081;
   wire n_257_76_2082;
   wire n_257_76_2083;
   wire n_257_76_2084;
   wire n_257_76_2085;
   wire n_257_76_2086;
   wire n_257_76_2087;
   wire n_257_76_2088;
   wire n_257_76_2089;
   wire n_257_76_2090;
   wire n_257_76_2091;
   wire n_257_76_2092;
   wire n_257_76_2093;
   wire n_257_76_2094;
   wire n_257_76_2095;
   wire n_257_76_2096;
   wire n_257_76_2097;
   wire n_257_76_2098;
   wire n_257_76_2099;
   wire n_257_76_2100;
   wire n_257_76_2101;
   wire n_257_76_2102;
   wire n_257_76_2103;
   wire n_257_76_2104;
   wire n_257_76_2105;
   wire n_257_76_2106;
   wire n_257_76_2107;
   wire n_257_76_2108;
   wire n_257_76_2109;
   wire n_257_76_2110;
   wire n_257_76_2111;
   wire n_257_76_2112;
   wire n_257_76_2113;
   wire n_257_76_2114;
   wire n_257_76_2115;
   wire n_257_76_2116;
   wire n_257_76_2117;
   wire n_257_76_2118;
   wire n_257_76_2119;
   wire n_257_76_2120;
   wire n_257_76_2121;
   wire n_257_76_2122;
   wire n_257_76_2123;
   wire n_257_76_2124;
   wire n_257_76_2125;
   wire n_257_76_2126;
   wire n_257_76_2127;
   wire n_257_76_2128;
   wire n_257_76_2129;
   wire n_257_76_2130;
   wire n_257_76_2131;
   wire n_257_76_2132;
   wire n_257_76_2133;
   wire n_257_76_2134;
   wire n_257_76_2135;
   wire n_257_76_2136;
   wire n_257_76_2137;
   wire n_257_76_2138;
   wire n_257_76_2139;
   wire n_257_76_2140;
   wire n_257_76_2141;
   wire n_257_76_2142;
   wire n_257_76_2143;
   wire n_257_76_2144;
   wire n_257_76_2145;
   wire n_257_76_2146;
   wire n_257_76_2147;
   wire n_257_76_2148;
   wire n_257_76_2149;
   wire n_257_76_2150;
   wire n_257_76_2151;
   wire n_257_76_2152;
   wire n_257_76_2153;
   wire n_257_76_2154;
   wire n_257_76_2155;
   wire n_257_76_2156;
   wire n_257_76_2157;
   wire n_257_76_2158;
   wire n_257_76_2159;
   wire n_257_76_2160;
   wire n_257_76_2161;
   wire n_257_76_2162;
   wire n_257_76_2163;
   wire n_257_76_2164;
   wire n_257_76_2165;
   wire n_257_76_2166;
   wire n_257_76_2167;
   wire n_257_76_2168;
   wire n_257_76_2169;
   wire n_257_76_2170;
   wire n_257_76_2171;
   wire n_257_76_2172;
   wire n_257_76_2173;
   wire n_257_76_2174;
   wire n_257_76_2175;
   wire n_257_76_2176;
   wire n_257_76_2177;
   wire n_257_76_2178;
   wire n_257_76_2179;
   wire n_257_76_2180;
   wire n_257_76_2181;
   wire n_257_76_2182;
   wire n_257_76_2183;
   wire n_257_76_2184;
   wire n_257_76_2185;
   wire n_257_76_2186;
   wire n_257_76_2187;
   wire n_257_76_2188;
   wire n_257_76_2189;
   wire n_257_76_2190;
   wire n_257_76_2191;
   wire n_257_76_2192;
   wire n_257_76_2193;
   wire n_257_76_2194;
   wire n_257_76_2195;
   wire n_257_76_2196;
   wire n_257_76_2197;
   wire n_257_76_2198;
   wire n_257_76_2199;
   wire n_257_76_2200;
   wire n_257_76_2201;
   wire n_257_76_2202;
   wire n_257_76_2203;
   wire n_257_76_2204;
   wire n_257_76_2205;
   wire n_257_76_2206;
   wire n_257_76_2207;
   wire n_257_76_2208;
   wire n_257_76_2209;
   wire n_257_76_2210;
   wire n_257_76_2211;
   wire n_257_76_2212;
   wire n_257_76_2213;
   wire n_257_76_2214;
   wire n_257_76_2215;
   wire n_257_76_2216;
   wire n_257_76_2217;
   wire n_257_76_2218;
   wire n_257_76_2219;
   wire n_257_76_2220;
   wire n_257_76_2221;
   wire n_257_76_2222;
   wire n_257_76_2223;
   wire n_257_76_2224;
   wire n_257_76_2225;
   wire n_257_76_2226;
   wire n_257_76_2227;
   wire n_257_76_2228;
   wire n_257_76_2229;
   wire n_257_76_2230;
   wire n_257_76_2231;
   wire n_257_76_2232;
   wire n_257_76_2233;
   wire n_257_76_2234;
   wire n_257_76_2235;
   wire n_257_76_2236;
   wire n_257_76_2237;
   wire n_257_76_2238;
   wire n_257_76_2239;
   wire n_257_76_2240;
   wire n_257_76_2241;
   wire n_257_76_2242;
   wire n_257_76_2243;
   wire n_257_76_2244;
   wire n_257_76_2245;
   wire n_257_76_2246;
   wire n_257_76_2247;
   wire n_257_76_2248;
   wire n_257_76_2249;
   wire n_257_76_2250;
   wire n_257_76_2251;
   wire n_257_76_2252;
   wire n_257_76_2253;
   wire n_257_76_2254;
   wire n_257_76_2255;
   wire n_257_76_2256;
   wire n_257_76_2257;
   wire n_257_76_2258;
   wire n_257_76_2259;
   wire n_257_76_2260;
   wire n_257_76_2261;
   wire n_257_76_2262;
   wire n_257_76_2263;
   wire n_257_76_2264;
   wire n_257_76_2265;
   wire n_257_76_2266;
   wire n_257_76_2267;
   wire n_257_76_2268;
   wire n_257_76_2269;
   wire n_257_76_2270;
   wire n_257_76_2271;
   wire n_257_76_2272;
   wire n_257_76_2273;
   wire n_257_76_2274;
   wire n_257_76_2275;
   wire n_257_76_2276;
   wire n_257_76_2277;
   wire n_257_76_2278;
   wire n_257_76_2279;
   wire n_257_76_2280;
   wire n_257_76_2281;
   wire n_257_76_2282;
   wire n_257_76_2283;
   wire n_257_76_2284;
   wire n_257_76_2285;
   wire n_257_76_2286;
   wire n_257_76_2287;
   wire n_257_76_2288;
   wire n_257_76_2289;
   wire n_257_76_2290;
   wire n_257_76_2291;
   wire n_257_76_2292;
   wire n_257_76_2293;
   wire n_257_76_2294;
   wire n_257_76_2295;
   wire n_257_76_2296;
   wire n_257_76_2297;
   wire n_257_76_2298;
   wire n_257_76_2299;
   wire n_257_76_2300;
   wire n_257_76_2301;
   wire n_257_76_2302;
   wire n_257_76_2303;
   wire n_257_76_2304;
   wire n_257_76_2305;
   wire n_257_76_2306;
   wire n_257_76_2307;
   wire n_257_76_2308;
   wire n_257_76_2309;
   wire n_257_76_2310;
   wire n_257_76_2311;
   wire n_257_76_2312;
   wire n_257_76_2313;
   wire n_257_76_2314;
   wire n_257_76_2315;
   wire n_257_76_2316;
   wire n_257_76_2317;
   wire n_257_76_2318;
   wire n_257_76_2319;
   wire n_257_76_2320;
   wire n_257_76_2321;
   wire n_257_76_2322;
   wire n_257_76_2323;
   wire n_257_76_2324;
   wire n_257_76_2325;
   wire n_257_76_2326;
   wire n_257_76_2327;
   wire n_257_76_2328;
   wire n_257_76_2329;
   wire n_257_76_2330;
   wire n_257_76_2331;
   wire n_257_76_2332;
   wire n_257_76_2333;
   wire n_257_76_2334;
   wire n_257_76_2335;
   wire n_257_76_2336;
   wire n_257_76_2337;
   wire n_257_76_2338;
   wire n_257_76_2339;
   wire n_257_76_2340;
   wire n_257_76_2341;
   wire n_257_76_2342;
   wire n_257_76_2343;
   wire n_257_76_2344;
   wire n_257_76_2345;
   wire n_257_76_2346;
   wire n_257_76_2347;
   wire n_257_76_2348;
   wire n_257_76_2349;
   wire n_257_76_2350;
   wire n_257_76_2351;
   wire n_257_76_2352;
   wire n_257_76_2353;
   wire n_257_76_2354;
   wire n_257_76_2355;
   wire n_257_76_2356;
   wire n_257_76_2357;
   wire n_257_76_2358;
   wire n_257_76_2359;
   wire n_257_76_2360;
   wire n_257_76_2361;
   wire n_257_76_2362;
   wire n_257_76_2363;
   wire n_257_76_2364;
   wire n_257_76_2365;
   wire n_257_76_2366;
   wire n_257_76_2367;
   wire n_257_76_2368;
   wire n_257_76_2369;
   wire n_257_76_2370;
   wire n_257_76_2371;
   wire n_257_76_2372;
   wire n_257_76_2373;
   wire n_257_76_2374;
   wire n_257_76_2375;
   wire n_257_76_2376;
   wire n_257_76_2377;
   wire n_257_76_2378;
   wire n_257_76_2379;
   wire n_257_76_2380;
   wire n_257_76_2381;
   wire n_257_76_2382;
   wire n_257_76_2383;
   wire n_257_76_2384;
   wire n_257_76_2385;
   wire n_257_76_2386;
   wire n_257_76_2387;
   wire n_257_76_2388;
   wire n_257_76_2389;
   wire n_257_76_2390;
   wire n_257_76_2391;
   wire n_257_76_2392;
   wire n_257_76_2393;
   wire n_257_76_2394;
   wire n_257_76_2395;
   wire n_257_76_2396;
   wire n_257_76_2397;
   wire n_257_76_2398;
   wire n_257_76_2399;
   wire n_257_76_2400;
   wire n_257_76_2401;
   wire n_257_76_2402;
   wire n_257_76_2403;
   wire n_257_76_2404;
   wire n_257_76_2405;
   wire n_257_76_2406;
   wire n_257_76_2407;
   wire n_257_76_2408;
   wire n_257_76_2409;
   wire n_257_76_2410;
   wire n_257_76_2411;
   wire n_257_76_2412;
   wire n_257_76_2413;
   wire n_257_76_2414;
   wire n_257_76_2415;
   wire n_257_76_2416;
   wire n_257_76_2417;
   wire n_257_76_2418;
   wire n_257_76_2419;
   wire n_257_76_2420;
   wire n_257_76_2421;
   wire n_257_76_2422;
   wire n_257_76_2423;
   wire n_257_76_2424;
   wire n_257_76_2425;
   wire n_257_76_2426;
   wire n_257_76_2427;
   wire n_257_76_2428;
   wire n_257_76_2429;
   wire n_257_76_2430;
   wire n_257_76_2431;
   wire n_257_76_2432;
   wire n_257_76_2433;
   wire n_257_76_2434;
   wire n_257_76_2435;
   wire n_257_76_2436;
   wire n_257_76_2437;
   wire n_257_76_2438;
   wire n_257_76_2439;
   wire n_257_76_2440;
   wire n_257_76_2441;
   wire n_257_76_2442;
   wire n_257_76_2443;
   wire n_257_76_2444;
   wire n_257_76_2445;
   wire n_257_76_2446;
   wire n_257_76_2447;
   wire n_257_76_2448;
   wire n_257_76_2449;
   wire n_257_76_2450;
   wire n_257_76_2451;
   wire n_257_76_2452;
   wire n_257_76_2453;
   wire n_257_76_2454;
   wire n_257_76_2455;
   wire n_257_76_2456;
   wire n_257_76_2457;
   wire n_257_76_2458;
   wire n_257_76_2459;
   wire n_257_76_2460;
   wire n_257_76_2461;
   wire n_257_76_2462;
   wire n_257_76_2463;
   wire n_257_76_2464;
   wire n_257_76_2465;
   wire n_257_76_2466;
   wire n_257_76_2467;
   wire n_257_76_2468;
   wire n_257_76_2469;
   wire n_257_76_2470;
   wire n_257_76_2471;
   wire n_257_76_2472;
   wire n_257_76_2473;
   wire n_257_76_2474;
   wire n_257_76_2475;
   wire n_257_76_2476;
   wire n_257_76_2477;
   wire n_257_76_2478;
   wire n_257_76_2479;
   wire n_257_76_2480;
   wire n_257_76_2481;
   wire n_257_76_2482;
   wire n_257_76_2483;
   wire n_257_76_2484;
   wire n_257_76_2485;
   wire n_257_76_2486;
   wire n_257_76_2487;
   wire n_257_76_2488;
   wire n_257_76_2489;
   wire n_257_76_2490;
   wire n_257_76_2491;
   wire n_257_76_2492;
   wire n_257_76_2493;
   wire n_257_76_2494;
   wire n_257_76_2495;
   wire n_257_76_2496;
   wire n_257_76_2497;
   wire n_257_76_2498;
   wire n_257_76_2499;
   wire n_257_76_2500;
   wire n_257_76_2501;
   wire n_257_76_2502;
   wire n_257_76_2503;
   wire n_257_76_2504;
   wire n_257_76_2505;
   wire n_257_76_2506;
   wire n_257_76_2507;
   wire n_257_76_2508;
   wire n_257_76_2509;
   wire n_257_76_2510;
   wire n_257_76_2511;
   wire n_257_76_2512;
   wire n_257_76_2513;
   wire n_257_76_2514;
   wire n_257_76_2515;
   wire n_257_76_2516;
   wire n_257_76_2517;
   wire n_257_76_2518;
   wire n_257_76_2519;
   wire n_257_76_2520;
   wire n_257_76_2521;
   wire n_257_76_2522;
   wire n_257_76_2523;
   wire n_257_76_2524;
   wire n_257_76_2525;
   wire n_257_76_2526;
   wire n_257_76_2527;
   wire n_257_76_2528;
   wire n_257_76_2529;
   wire n_257_76_2530;
   wire n_257_76_2531;
   wire n_257_76_2532;
   wire n_257_76_2533;
   wire n_257_76_2534;
   wire n_257_76_2535;
   wire n_257_76_2536;
   wire n_257_76_2537;
   wire n_257_76_2538;
   wire n_257_76_2539;
   wire n_257_76_2540;
   wire n_257_76_2541;
   wire n_257_76_2542;
   wire n_257_76_2543;
   wire n_257_76_2544;
   wire n_257_76_2545;
   wire n_257_76_2546;
   wire n_257_76_2547;
   wire n_257_76_2548;
   wire n_257_76_2549;
   wire n_257_76_2550;
   wire n_257_76_2551;
   wire n_257_76_2552;
   wire n_257_76_2553;
   wire n_257_76_2554;
   wire n_257_76_2555;
   wire n_257_76_2556;
   wire n_257_76_2557;
   wire n_257_76_2558;
   wire n_257_76_2559;
   wire n_257_76_2560;
   wire n_257_76_2561;
   wire n_257_76_2562;
   wire n_257_76_2563;
   wire n_257_76_2564;
   wire n_257_76_2565;
   wire n_257_76_2566;
   wire n_257_76_2567;
   wire n_257_76_2568;
   wire n_257_76_2569;
   wire n_257_76_2570;
   wire n_257_76_2571;
   wire n_257_76_2572;
   wire n_257_76_2573;
   wire n_257_76_2574;
   wire n_257_76_2575;
   wire n_257_76_2576;
   wire n_257_76_2577;
   wire n_257_76_2578;
   wire n_257_76_2579;
   wire n_257_76_2580;
   wire n_257_76_2581;
   wire n_257_76_2582;
   wire n_257_76_2583;
   wire n_257_76_2584;
   wire n_257_76_2585;
   wire n_257_76_2586;
   wire n_257_76_2587;
   wire n_257_76_2588;
   wire n_257_76_2589;
   wire n_257_76_2590;
   wire n_257_76_2591;
   wire n_257_76_2592;
   wire n_257_76_2593;
   wire n_257_76_2594;
   wire n_257_76_2595;
   wire n_257_76_2596;
   wire n_257_76_2597;
   wire n_257_76_2598;
   wire n_257_76_2599;
   wire n_257_76_2600;
   wire n_257_76_2601;
   wire n_257_76_2602;
   wire n_257_76_2603;
   wire n_257_76_2604;
   wire n_257_76_2605;
   wire n_257_76_2606;
   wire n_257_76_2607;
   wire n_257_76_2608;
   wire n_257_76_2609;
   wire n_257_76_2610;
   wire n_257_76_2611;
   wire n_257_76_2612;
   wire n_257_76_2613;
   wire n_257_76_2614;
   wire n_257_76_2615;
   wire n_257_76_2616;
   wire n_257_76_2617;
   wire n_257_76_2618;
   wire n_257_76_2619;
   wire n_257_76_2620;
   wire n_257_76_2621;
   wire n_257_76_2622;
   wire n_257_76_2623;
   wire n_257_76_2624;
   wire n_257_76_2625;
   wire n_257_76_2626;
   wire n_257_76_2627;
   wire n_257_76_2628;
   wire n_257_76_2629;
   wire n_257_76_2630;
   wire n_257_76_2631;
   wire n_257_76_2632;
   wire n_257_76_2633;
   wire n_257_76_2634;
   wire n_257_76_2635;
   wire n_257_76_2636;
   wire n_257_76_2637;
   wire n_257_76_2638;
   wire n_257_76_2639;
   wire n_257_76_2640;
   wire n_257_76_2641;
   wire n_257_76_2642;
   wire n_257_76_2643;
   wire n_257_76_2644;
   wire n_257_76_2645;
   wire n_257_76_2646;
   wire n_257_76_2647;
   wire n_257_76_2648;
   wire n_257_76_2649;
   wire n_257_76_2650;
   wire n_257_76_2651;
   wire n_257_76_2652;
   wire n_257_76_2653;
   wire n_257_76_2654;
   wire n_257_76_2655;
   wire n_257_76_2656;
   wire n_257_76_2657;
   wire n_257_76_2658;
   wire n_257_76_2659;
   wire n_257_76_2660;
   wire n_257_76_2661;
   wire n_257_76_2662;
   wire n_257_76_2663;
   wire n_257_76_2664;
   wire n_257_76_2665;
   wire n_257_76_2666;
   wire n_257_76_2667;
   wire n_257_76_2668;
   wire n_257_76_2669;
   wire n_257_76_2670;
   wire n_257_76_2671;
   wire n_257_76_2672;
   wire n_257_76_2673;
   wire n_257_76_2674;
   wire n_257_76_2675;
   wire n_257_76_2676;
   wire n_257_76_2677;
   wire n_257_76_2678;
   wire n_257_76_2679;
   wire n_257_76_2680;
   wire n_257_76_2681;
   wire n_257_76_2682;
   wire n_257_76_2683;
   wire n_257_76_2684;
   wire n_257_76_2685;
   wire n_257_76_2686;
   wire n_257_76_2687;
   wire n_257_76_2688;
   wire n_257_76_2689;
   wire n_257_76_2690;
   wire n_257_76_2691;
   wire n_257_76_2692;
   wire n_257_76_2693;
   wire n_257_76_2694;
   wire n_257_76_2695;
   wire n_257_76_2696;
   wire n_257_76_2697;
   wire n_257_76_2698;
   wire n_257_76_2699;
   wire n_257_76_2700;
   wire n_257_76_2701;
   wire n_257_76_2702;
   wire n_257_76_2703;
   wire n_257_76_2704;
   wire n_257_76_2705;
   wire n_257_76_2706;
   wire n_257_76_2707;
   wire n_257_76_2708;
   wire n_257_76_2709;
   wire n_257_76_2710;
   wire n_257_76_2711;
   wire n_257_76_2712;
   wire n_257_76_2713;
   wire n_257_76_2714;
   wire n_257_76_2715;
   wire n_257_76_2716;
   wire n_257_76_2717;
   wire n_257_76_2718;
   wire n_257_76_2719;
   wire n_257_76_2720;
   wire n_257_76_2721;
   wire n_257_76_2722;
   wire n_257_76_2723;
   wire n_257_76_2724;
   wire n_257_76_2725;
   wire n_257_76_2726;
   wire n_257_76_2727;
   wire n_257_76_2728;
   wire n_257_76_2729;
   wire n_257_76_2730;
   wire n_257_76_2731;
   wire n_257_76_2732;
   wire n_257_76_2733;
   wire n_257_76_2734;
   wire n_257_76_2735;
   wire n_257_76_2736;
   wire n_257_76_2737;
   wire n_257_76_2738;
   wire n_257_76_2739;
   wire n_257_76_2740;
   wire n_257_76_2741;
   wire n_257_76_2742;
   wire n_257_76_2743;
   wire n_257_76_2744;
   wire n_257_76_2745;
   wire n_257_76_2746;
   wire n_257_76_2747;
   wire n_257_76_2748;
   wire n_257_76_2749;
   wire n_257_76_2750;
   wire n_257_76_2751;
   wire n_257_76_2752;
   wire n_257_76_2753;
   wire n_257_76_2754;
   wire n_257_76_2755;
   wire n_257_76_2756;
   wire n_257_76_2757;
   wire n_257_76_2758;
   wire n_257_76_2759;
   wire n_257_76_2760;
   wire n_257_76_2761;
   wire n_257_76_2762;
   wire n_257_76_2763;
   wire n_257_76_2764;
   wire n_257_76_2765;
   wire n_257_76_2766;
   wire n_257_76_2767;
   wire n_257_76_2768;
   wire n_257_76_2769;
   wire n_257_76_2770;
   wire n_257_76_2771;
   wire n_257_76_2772;
   wire n_257_76_2773;
   wire n_257_76_2774;
   wire n_257_76_2775;
   wire n_257_76_2776;
   wire n_257_76_2777;
   wire n_257_76_2778;
   wire n_257_76_2779;
   wire n_257_76_2780;
   wire n_257_76_2781;
   wire n_257_76_2782;
   wire n_257_76_2783;
   wire n_257_76_2784;
   wire n_257_76_2785;
   wire n_257_76_2786;
   wire n_257_76_2787;
   wire n_257_76_2788;
   wire n_257_76_2789;
   wire n_257_76_2790;
   wire n_257_76_2791;
   wire n_257_76_2792;
   wire n_257_76_2793;
   wire n_257_76_2794;
   wire n_257_76_2795;
   wire n_257_76_2796;
   wire n_257_76_2797;
   wire n_257_76_2798;
   wire n_257_76_2799;
   wire n_257_76_2800;
   wire n_257_76_2801;
   wire n_257_76_2802;
   wire n_257_76_2803;
   wire n_257_76_2804;
   wire n_257_76_2805;
   wire n_257_76_2806;
   wire n_257_76_2807;
   wire n_257_76_2808;
   wire n_257_76_2809;
   wire n_257_76_2810;
   wire n_257_76_2811;
   wire n_257_76_2812;
   wire n_257_76_2813;
   wire n_257_76_2814;
   wire n_257_76_2815;
   wire n_257_76_2816;
   wire n_257_76_2817;
   wire n_257_76_2818;
   wire n_257_76_2819;
   wire n_257_76_2820;
   wire n_257_76_2821;
   wire n_257_76_2822;
   wire n_257_76_2823;
   wire n_257_76_2824;
   wire n_257_76_2825;
   wire n_257_76_2826;
   wire n_257_76_2827;
   wire n_257_76_2828;
   wire n_257_76_2829;
   wire n_257_76_2830;
   wire n_257_76_2831;
   wire n_257_76_2832;
   wire n_257_76_2833;
   wire n_257_76_2834;
   wire n_257_76_2835;
   wire n_257_76_2836;
   wire n_257_76_2837;
   wire n_257_76_2838;
   wire n_257_76_2839;
   wire n_257_76_2840;
   wire n_257_76_2841;
   wire n_257_76_2842;
   wire n_257_76_2843;
   wire n_257_76_2844;
   wire n_257_76_2845;
   wire n_257_76_2846;
   wire n_257_76_2847;
   wire n_257_76_2848;
   wire n_257_76_2849;
   wire n_257_76_2850;
   wire n_257_76_2851;
   wire n_257_76_2852;
   wire n_257_76_2853;
   wire n_257_76_2854;
   wire n_257_76_2855;
   wire n_257_76_2856;
   wire n_257_76_2857;
   wire n_257_76_2858;
   wire n_257_76_2859;
   wire n_257_76_2860;
   wire n_257_76_2861;
   wire n_257_76_2862;
   wire n_257_76_2863;
   wire n_257_76_2864;
   wire n_257_76_2865;
   wire n_257_76_2866;
   wire n_257_76_2867;
   wire n_257_76_2868;
   wire n_257_76_2869;
   wire n_257_76_2870;
   wire n_257_76_2871;
   wire n_257_76_2872;
   wire n_257_76_2873;
   wire n_257_76_2874;
   wire n_257_76_2875;
   wire n_257_76_2876;
   wire n_257_76_2877;
   wire n_257_76_2878;
   wire n_257_76_2879;
   wire n_257_76_2880;
   wire n_257_76_2881;
   wire n_257_76_2882;
   wire n_257_76_2883;
   wire n_257_76_2884;
   wire n_257_76_2885;
   wire n_257_76_2886;
   wire n_257_76_2887;
   wire n_257_76_2888;
   wire n_257_76_2889;
   wire n_257_76_2890;
   wire n_257_76_2891;
   wire n_257_76_2892;
   wire n_257_76_2893;
   wire n_257_76_2894;
   wire n_257_76_2895;
   wire n_257_76_2896;
   wire n_257_76_2897;
   wire n_257_76_2898;
   wire n_257_76_2899;
   wire n_257_76_2900;
   wire n_257_76_2901;
   wire n_257_76_2902;
   wire n_257_76_2903;
   wire n_257_76_2904;
   wire n_257_76_2905;
   wire n_257_76_2906;
   wire n_257_76_2907;
   wire n_257_76_2908;
   wire n_257_76_2909;
   wire n_257_76_2910;
   wire n_257_76_2911;
   wire n_257_76_2912;
   wire n_257_76_2913;
   wire n_257_76_2914;
   wire n_257_76_2915;
   wire n_257_76_2916;
   wire n_257_76_2917;
   wire n_257_76_2918;
   wire n_257_76_2919;
   wire n_257_76_2920;
   wire n_257_76_2921;
   wire n_257_76_2922;
   wire n_257_76_2923;
   wire n_257_76_2924;
   wire n_257_76_2925;
   wire n_257_76_2926;
   wire n_257_76_2927;
   wire n_257_76_2928;
   wire n_257_76_2929;
   wire n_257_76_2930;
   wire n_257_76_2931;
   wire n_257_76_2932;
   wire n_257_76_2933;
   wire n_257_76_2934;
   wire n_257_76_2935;
   wire n_257_76_2936;
   wire n_257_76_2937;
   wire n_257_76_2938;
   wire n_257_76_2939;
   wire n_257_76_2940;
   wire n_257_76_2941;
   wire n_257_76_2942;
   wire n_257_76_2943;
   wire n_257_76_2944;
   wire n_257_76_2945;
   wire n_257_76_2946;
   wire n_257_76_2947;
   wire n_257_76_2948;
   wire n_257_76_2949;
   wire n_257_76_2950;
   wire n_257_76_2951;
   wire n_257_76_2952;
   wire n_257_76_2953;
   wire n_257_76_2954;
   wire n_257_76_2955;
   wire n_257_76_2956;
   wire n_257_76_2957;
   wire n_257_76_2958;
   wire n_257_76_2959;
   wire n_257_76_2960;
   wire n_257_76_2961;
   wire n_257_76_2962;
   wire n_257_76_2963;
   wire n_257_76_2964;
   wire n_257_76_2965;
   wire n_257_76_2966;
   wire n_257_76_2967;
   wire n_257_76_2968;
   wire n_257_76_2969;
   wire n_257_76_2970;
   wire n_257_76_2971;
   wire n_257_76_2972;
   wire n_257_76_2973;
   wire n_257_76_2974;
   wire n_257_76_2975;
   wire n_257_76_2976;
   wire n_257_76_2977;
   wire n_257_76_2978;
   wire n_257_76_2979;
   wire n_257_76_2980;
   wire n_257_76_2981;
   wire n_257_76_2982;
   wire n_257_76_2983;
   wire n_257_76_2984;
   wire n_257_76_2985;
   wire n_257_76_2986;
   wire n_257_76_2987;
   wire n_257_76_2988;
   wire n_257_76_2989;
   wire n_257_76_2990;
   wire n_257_76_2991;
   wire n_257_76_2992;
   wire n_257_76_2993;
   wire n_257_76_2994;
   wire n_257_76_2995;
   wire n_257_76_2996;
   wire n_257_76_2997;
   wire n_257_76_2998;
   wire n_257_76_2999;
   wire n_257_76_3000;
   wire n_257_76_3001;
   wire n_257_76_3002;
   wire n_257_76_3003;
   wire n_257_76_3004;
   wire n_257_76_3005;
   wire n_257_76_3006;
   wire n_257_76_3007;
   wire n_257_76_3008;
   wire n_257_76_3009;
   wire n_257_76_3010;
   wire n_257_76_3011;
   wire n_257_76_3012;
   wire n_257_76_3013;
   wire n_257_76_3014;
   wire n_257_76_3015;
   wire n_257_76_3016;
   wire n_257_76_3017;
   wire n_257_76_3018;
   wire n_257_76_3019;
   wire n_257_76_3020;
   wire n_257_76_3021;
   wire n_257_76_3022;
   wire n_257_76_3023;
   wire n_257_76_3024;
   wire n_257_76_3025;
   wire n_257_76_3026;
   wire n_257_76_3027;
   wire n_257_76_3028;
   wire n_257_76_3029;
   wire n_257_76_3030;
   wire n_257_76_3031;
   wire n_257_76_3032;
   wire n_257_76_3033;
   wire n_257_76_3034;
   wire n_257_76_3035;
   wire n_257_76_3036;
   wire n_257_76_3037;
   wire n_257_76_3038;
   wire n_257_76_3039;
   wire n_257_76_3040;
   wire n_257_76_3041;
   wire n_257_76_3042;
   wire n_257_76_3043;
   wire n_257_76_3044;
   wire n_257_76_3045;
   wire n_257_76_3046;
   wire n_257_76_3047;
   wire n_257_76_3048;
   wire n_257_76_3049;
   wire n_257_76_3050;
   wire n_257_76_3051;
   wire n_257_76_3052;
   wire n_257_76_3053;
   wire n_257_76_3054;
   wire n_257_76_3055;
   wire n_257_76_3056;
   wire n_257_76_3057;
   wire n_257_76_3058;
   wire n_257_76_3059;
   wire n_257_76_3060;
   wire n_257_76_3061;
   wire n_257_76_3062;
   wire n_257_76_3063;
   wire n_257_76_3064;
   wire n_257_76_3065;
   wire n_257_76_3066;
   wire n_257_76_3067;
   wire n_257_76_3068;
   wire n_257_76_3069;
   wire n_257_76_3070;
   wire n_257_76_3071;
   wire n_257_76_3072;
   wire n_257_76_3073;
   wire n_257_76_3074;
   wire n_257_76_3075;
   wire n_257_76_3076;
   wire n_257_76_3077;
   wire n_257_76_3078;
   wire n_257_76_3079;
   wire n_257_76_3080;
   wire n_257_76_3081;
   wire n_257_76_3082;
   wire n_257_76_3083;
   wire n_257_76_3084;
   wire n_257_76_3085;
   wire n_257_76_3086;
   wire n_257_76_3087;
   wire n_257_76_3088;
   wire n_257_76_3089;
   wire n_257_76_3090;
   wire n_257_76_3091;
   wire n_257_76_3092;
   wire n_257_76_3093;
   wire n_257_76_3094;
   wire n_257_76_3095;
   wire n_257_76_3096;
   wire n_257_76_3097;
   wire n_257_76_3098;
   wire n_257_76_3099;
   wire n_257_76_3100;
   wire n_257_76_3101;
   wire n_257_76_3102;
   wire n_257_76_3103;
   wire n_257_76_3104;
   wire n_257_76_3105;
   wire n_257_76_3106;
   wire n_257_76_3107;
   wire n_257_76_3108;
   wire n_257_76_3109;
   wire n_257_76_3110;
   wire n_257_76_3111;
   wire n_257_76_3112;
   wire n_257_76_3113;
   wire n_257_76_3114;
   wire n_257_76_3115;
   wire n_257_76_3116;
   wire n_257_76_3117;
   wire n_257_76_3118;
   wire n_257_76_3119;
   wire n_257_76_3120;
   wire n_257_76_3121;
   wire n_257_76_3122;
   wire n_257_76_3123;
   wire n_257_76_3124;
   wire n_257_76_3125;
   wire n_257_76_3126;
   wire n_257_76_3127;
   wire n_257_76_3128;
   wire n_257_76_3129;
   wire n_257_76_3130;
   wire n_257_76_3131;
   wire n_257_76_3132;
   wire n_257_76_3133;
   wire n_257_76_3134;
   wire n_257_76_3135;
   wire n_257_76_3136;
   wire n_257_76_3137;
   wire n_257_76_3138;
   wire n_257_76_3139;
   wire n_257_76_3140;
   wire n_257_76_3141;
   wire n_257_76_3142;
   wire n_257_76_3143;
   wire n_257_76_3144;
   wire n_257_76_3145;
   wire n_257_76_3146;
   wire n_257_76_3147;
   wire n_257_76_3148;
   wire n_257_76_3149;
   wire n_257_76_3150;
   wire n_257_76_3151;
   wire n_257_76_3152;
   wire n_257_76_3153;
   wire n_257_76_3154;
   wire n_257_76_3155;
   wire n_257_76_3156;
   wire n_257_76_3157;
   wire n_257_76_3158;
   wire n_257_76_3159;
   wire n_257_76_3160;
   wire n_257_76_3161;
   wire n_257_76_3162;
   wire n_257_76_3163;
   wire n_257_76_3164;
   wire n_257_76_3165;
   wire n_257_76_3166;
   wire n_257_76_3167;
   wire n_257_76_3168;
   wire n_257_76_3169;
   wire n_257_76_3170;
   wire n_257_76_3171;
   wire n_257_76_3172;
   wire n_257_76_3173;
   wire n_257_76_3174;
   wire n_257_76_3175;
   wire n_257_76_3176;
   wire n_257_76_3177;
   wire n_257_76_3178;
   wire n_257_76_3179;
   wire n_257_76_3180;
   wire n_257_76_3181;
   wire n_257_76_3182;
   wire n_257_76_3183;
   wire n_257_76_3184;
   wire n_257_76_3185;
   wire n_257_76_3186;
   wire n_257_76_3187;
   wire n_257_76_3188;
   wire n_257_76_3189;
   wire n_257_76_3190;
   wire n_257_76_3191;
   wire n_257_76_3192;
   wire n_257_76_3193;
   wire n_257_76_3194;
   wire n_257_76_3195;
   wire n_257_76_3196;
   wire n_257_76_3197;
   wire n_257_76_3198;
   wire n_257_76_3199;
   wire n_257_76_3200;
   wire n_257_76_3201;
   wire n_257_76_3202;
   wire n_257_76_3203;
   wire n_257_76_3204;
   wire n_257_76_3205;
   wire n_257_76_3206;
   wire n_257_76_3207;
   wire n_257_76_3208;
   wire n_257_76_3209;
   wire n_257_76_3210;
   wire n_257_76_3211;
   wire n_257_76_3212;
   wire n_257_76_3213;
   wire n_257_76_3214;
   wire n_257_76_3215;
   wire n_257_76_3216;
   wire n_257_76_3217;
   wire n_257_76_3218;
   wire n_257_76_3219;
   wire n_257_76_3220;
   wire n_257_76_3221;
   wire n_257_76_3222;
   wire n_257_76_3223;
   wire n_257_76_3224;
   wire n_257_76_3225;
   wire n_257_76_3226;
   wire n_257_76_3227;
   wire n_257_76_3228;
   wire n_257_76_3229;
   wire n_257_76_3230;
   wire n_257_76_3231;
   wire n_257_76_3232;
   wire n_257_76_3233;
   wire n_257_76_3234;
   wire n_257_76_3235;
   wire n_257_76_3236;
   wire n_257_76_3237;
   wire n_257_76_3238;
   wire n_257_76_3239;
   wire n_257_76_3240;
   wire n_257_76_3241;
   wire n_257_76_3242;
   wire n_257_76_3243;
   wire n_257_76_3244;
   wire n_257_76_3245;
   wire n_257_76_3246;
   wire n_257_76_3247;
   wire n_257_76_3248;
   wire n_257_76_3249;
   wire n_257_76_3250;
   wire n_257_76_3251;
   wire n_257_76_3252;
   wire n_257_76_3253;
   wire n_257_76_3254;
   wire n_257_76_3255;
   wire n_257_76_3256;
   wire n_257_76_3257;
   wire n_257_76_3258;
   wire n_257_76_3259;
   wire n_257_76_3260;
   wire n_257_76_3261;
   wire n_257_76_3262;
   wire n_257_76_3263;
   wire n_257_76_3264;
   wire n_257_76_3265;
   wire n_257_76_3266;
   wire n_257_76_3267;
   wire n_257_76_3268;
   wire n_257_76_3269;
   wire n_257_76_3270;
   wire n_257_76_3271;
   wire n_257_76_3272;
   wire n_257_76_3273;
   wire n_257_76_3274;
   wire n_257_76_3275;
   wire n_257_76_3276;
   wire n_257_76_3277;
   wire n_257_76_3278;
   wire n_257_76_3279;
   wire n_257_76_3280;
   wire n_257_76_3281;
   wire n_257_76_3282;
   wire n_257_76_3283;
   wire n_257_76_3284;
   wire n_257_76_3285;
   wire n_257_76_3286;
   wire n_257_76_3287;
   wire n_257_76_3288;
   wire n_257_76_3289;
   wire n_257_76_3290;
   wire n_257_76_3291;
   wire n_257_76_3292;
   wire n_257_76_3293;
   wire n_257_76_3294;
   wire n_257_76_3295;
   wire n_257_76_3296;
   wire n_257_76_3297;
   wire n_257_76_3298;
   wire n_257_76_3299;
   wire n_257_76_3300;
   wire n_257_76_3301;
   wire n_257_76_3302;
   wire n_257_76_3303;
   wire n_257_76_3304;
   wire n_257_76_3305;
   wire n_257_76_3306;
   wire n_257_76_3307;
   wire n_257_76_3308;
   wire n_257_76_3309;
   wire n_257_76_3310;
   wire n_257_76_3311;
   wire n_257_76_3312;
   wire n_257_76_3313;
   wire n_257_76_3314;
   wire n_257_76_3315;
   wire n_257_76_3316;
   wire n_257_76_3317;
   wire n_257_76_3318;
   wire n_257_76_3319;
   wire n_257_76_3320;
   wire n_257_76_3321;
   wire n_257_76_3322;
   wire n_257_76_3323;
   wire n_257_76_3324;
   wire n_257_76_3325;
   wire n_257_76_3326;
   wire n_257_76_3327;
   wire n_257_76_3328;
   wire n_257_76_3329;
   wire n_257_76_3330;
   wire n_257_76_3331;
   wire n_257_76_3332;
   wire n_257_76_3333;
   wire n_257_76_3334;
   wire n_257_76_3335;
   wire n_257_76_3336;
   wire n_257_76_3337;
   wire n_257_76_3338;
   wire n_257_76_3339;
   wire n_257_76_3340;
   wire n_257_76_3341;
   wire n_257_76_3342;
   wire n_257_76_3343;
   wire n_257_76_3344;
   wire n_257_76_3345;
   wire n_257_76_3346;
   wire n_257_76_3347;
   wire n_257_76_3348;
   wire n_257_76_3349;
   wire n_257_76_3350;
   wire n_257_76_3351;
   wire n_257_76_3352;
   wire n_257_76_3353;
   wire n_257_76_3354;
   wire n_257_76_3355;
   wire n_257_76_3356;
   wire n_257_76_3357;
   wire n_257_76_3358;
   wire n_257_76_3359;
   wire n_257_76_3360;
   wire n_257_76_3361;
   wire n_257_76_3362;
   wire n_257_76_3363;
   wire n_257_76_3364;
   wire n_257_76_3365;
   wire n_257_76_3366;
   wire n_257_76_3367;
   wire n_257_76_3368;
   wire n_257_76_3369;
   wire n_257_76_3370;
   wire n_257_76_3371;
   wire n_257_76_3372;
   wire n_257_76_3373;
   wire n_257_76_3374;
   wire n_257_76_3375;
   wire n_257_76_3376;
   wire n_257_76_3377;
   wire n_257_76_3378;
   wire n_257_76_3379;
   wire n_257_76_3380;
   wire n_257_76_3381;
   wire n_257_76_3382;
   wire n_257_76_3383;
   wire n_257_76_3384;
   wire n_257_76_3385;
   wire n_257_76_3386;
   wire n_257_76_3387;
   wire n_257_76_3388;
   wire n_257_76_3389;
   wire n_257_76_3390;
   wire n_257_76_3391;
   wire n_257_76_3392;
   wire n_257_76_3393;
   wire n_257_76_3394;
   wire n_257_76_3395;
   wire n_257_76_3396;
   wire n_257_76_3397;
   wire n_257_76_3398;
   wire n_257_76_3399;
   wire n_257_76_3400;
   wire n_257_76_3401;
   wire n_257_76_3402;
   wire n_257_76_3403;
   wire n_257_76_3404;
   wire n_257_76_3405;
   wire n_257_76_3406;
   wire n_257_76_3407;
   wire n_257_76_3408;
   wire n_257_76_3409;
   wire n_257_76_3410;
   wire n_257_76_3411;
   wire n_257_76_3412;
   wire n_257_76_3413;
   wire n_257_76_3414;
   wire n_257_76_3415;
   wire n_257_76_3416;
   wire n_257_76_3417;
   wire n_257_76_3418;
   wire n_257_76_3419;
   wire n_257_76_3420;
   wire n_257_76_3421;
   wire n_257_76_3422;
   wire n_257_76_3423;
   wire n_257_76_3424;
   wire n_257_76_3425;
   wire n_257_76_3426;
   wire n_257_76_3427;
   wire n_257_76_3428;
   wire n_257_76_3429;
   wire n_257_76_3430;
   wire n_257_76_3431;
   wire n_257_76_3432;
   wire n_257_76_3433;
   wire n_257_76_3434;
   wire n_257_76_3435;
   wire n_257_76_3436;
   wire n_257_76_3437;
   wire n_257_76_3438;
   wire n_257_76_3439;
   wire n_257_76_3440;
   wire n_257_76_3441;
   wire n_257_76_3442;
   wire n_257_76_3443;
   wire n_257_76_3444;
   wire n_257_76_3445;
   wire n_257_76_3446;
   wire n_257_76_3447;
   wire n_257_76_3448;
   wire n_257_76_3449;
   wire n_257_76_3450;
   wire n_257_76_3451;
   wire n_257_76_3452;
   wire n_257_76_3453;
   wire n_257_76_3454;
   wire n_257_76_3455;
   wire n_257_76_3456;
   wire n_257_76_3457;
   wire n_257_76_3458;
   wire n_257_76_3459;
   wire n_257_76_3460;
   wire n_257_76_3461;
   wire n_257_76_3462;
   wire n_257_76_3463;
   wire n_257_76_3464;
   wire n_257_76_3465;
   wire n_257_76_3466;
   wire n_257_76_3467;
   wire n_257_76_3468;
   wire n_257_76_3469;
   wire n_257_76_3470;
   wire n_257_76_3471;
   wire n_257_76_3472;
   wire n_257_76_3473;
   wire n_257_76_3474;
   wire n_257_76_3475;
   wire n_257_76_3476;
   wire n_257_76_3477;
   wire n_257_76_3478;
   wire n_257_76_3479;
   wire n_257_76_3480;
   wire n_257_76_3481;
   wire n_257_76_3482;
   wire n_257_76_3483;
   wire n_257_76_3484;
   wire n_257_76_3485;
   wire n_257_76_3486;
   wire n_257_76_3487;
   wire n_257_76_3488;
   wire n_257_76_3489;
   wire n_257_76_3490;
   wire n_257_76_3491;
   wire n_257_76_3492;
   wire n_257_76_3493;
   wire n_257_76_3494;
   wire n_257_76_3495;
   wire n_257_76_3496;
   wire n_257_76_3497;
   wire n_257_76_3498;
   wire n_257_76_3499;
   wire n_257_76_3500;
   wire n_257_76_3501;
   wire n_257_76_3502;
   wire n_257_76_3503;
   wire n_257_76_3504;
   wire n_257_76_3505;
   wire n_257_76_3506;
   wire n_257_76_3507;
   wire n_257_76_3508;
   wire n_257_76_3509;
   wire n_257_76_3510;
   wire n_257_76_3511;
   wire n_257_76_3512;
   wire n_257_76_3513;
   wire n_257_76_3514;
   wire n_257_76_3515;
   wire n_257_76_3516;
   wire n_257_76_3517;
   wire n_257_76_3518;
   wire n_257_76_3519;
   wire n_257_76_3520;
   wire n_257_76_3521;
   wire n_257_76_3522;
   wire n_257_76_3523;
   wire n_257_76_3524;
   wire n_257_76_3525;
   wire n_257_76_3526;
   wire n_257_76_3527;
   wire n_257_76_3528;
   wire n_257_76_3529;
   wire n_257_76_3530;
   wire n_257_76_3531;
   wire n_257_76_3532;
   wire n_257_76_3533;
   wire n_257_76_3534;
   wire n_257_76_3535;
   wire n_257_76_3536;
   wire n_257_76_3537;
   wire n_257_76_3538;
   wire n_257_76_3539;
   wire n_257_76_3540;
   wire n_257_76_3541;
   wire n_257_76_3542;
   wire n_257_76_3543;
   wire n_257_76_3544;
   wire n_257_76_3545;
   wire n_257_76_3546;
   wire n_257_76_3547;
   wire n_257_76_3548;
   wire n_257_76_3549;
   wire n_257_76_3550;
   wire n_257_76_3551;
   wire n_257_76_3552;
   wire n_257_76_3553;
   wire n_257_76_3554;
   wire n_257_76_3555;
   wire n_257_76_3556;
   wire n_257_76_3557;
   wire n_257_76_3558;
   wire n_257_76_3559;
   wire n_257_76_3560;
   wire n_257_76_3561;
   wire n_257_76_3562;
   wire n_257_76_3563;
   wire n_257_76_3564;
   wire n_257_76_3565;
   wire n_257_76_3566;
   wire n_257_76_3567;
   wire n_257_76_3568;
   wire n_257_76_3569;
   wire n_257_76_3570;
   wire n_257_76_3571;
   wire n_257_76_3572;
   wire n_257_76_3573;
   wire n_257_76_3574;
   wire n_257_76_3575;
   wire n_257_76_3576;
   wire n_257_76_3577;
   wire n_257_76_3578;
   wire n_257_76_3579;
   wire n_257_76_3580;
   wire n_257_76_3581;
   wire n_257_76_3582;
   wire n_257_76_3583;
   wire n_257_76_3584;
   wire n_257_76_3585;
   wire n_257_76_3586;
   wire n_257_76_3587;
   wire n_257_76_3588;
   wire n_257_76_3589;
   wire n_257_76_3590;
   wire n_257_76_3591;
   wire n_257_76_3592;
   wire n_257_76_3593;
   wire n_257_76_3594;
   wire n_257_76_3595;
   wire n_257_76_3596;
   wire n_257_76_3597;
   wire n_257_76_3598;
   wire n_257_76_3599;
   wire n_257_76_3600;
   wire n_257_76_3601;
   wire n_257_76_3602;
   wire n_257_76_3603;
   wire n_257_76_3604;
   wire n_257_76_3605;
   wire n_257_76_3606;
   wire n_257_76_3607;
   wire n_257_76_3608;
   wire n_257_76_3609;
   wire n_257_76_3610;
   wire n_257_76_3611;
   wire n_257_76_3612;
   wire n_257_76_3613;
   wire n_257_76_3614;
   wire n_257_76_3615;
   wire n_257_76_3616;
   wire n_257_76_3617;
   wire n_257_76_3618;
   wire n_257_76_3619;
   wire n_257_76_3620;
   wire n_257_76_3621;
   wire n_257_76_3622;
   wire n_257_76_3623;
   wire n_257_76_3624;
   wire n_257_76_3625;
   wire n_257_76_3626;
   wire n_257_76_3627;
   wire n_257_76_3628;
   wire n_257_76_3629;
   wire n_257_76_3630;
   wire n_257_76_3631;
   wire n_257_76_3632;
   wire n_257_76_3633;
   wire n_257_76_3634;
   wire n_257_76_3635;
   wire n_257_76_3636;
   wire n_257_76_3637;
   wire n_257_76_3638;
   wire n_257_76_3639;
   wire n_257_76_3640;
   wire n_257_76_3641;
   wire n_257_76_3642;
   wire n_257_76_3643;
   wire n_257_76_3644;
   wire n_257_76_3645;
   wire n_257_76_3646;
   wire n_257_76_3647;
   wire n_257_76_3648;
   wire n_257_76_3649;
   wire n_257_76_3650;
   wire n_257_76_3651;
   wire n_257_76_3652;
   wire n_257_76_3653;
   wire n_257_76_3654;
   wire n_257_76_3655;
   wire n_257_76_3656;
   wire n_257_76_3657;
   wire n_257_76_3658;
   wire n_257_76_3659;
   wire n_257_76_3660;
   wire n_257_76_3661;
   wire n_257_76_3662;
   wire n_257_76_3663;
   wire n_257_76_3664;
   wire n_257_76_3665;
   wire n_257_76_3666;
   wire n_257_76_3667;
   wire n_257_76_3668;
   wire n_257_76_3669;
   wire n_257_76_3670;
   wire n_257_76_3671;
   wire n_257_76_3672;
   wire n_257_76_3673;
   wire n_257_76_3674;
   wire n_257_76_3675;
   wire n_257_76_3676;
   wire n_257_76_3677;
   wire n_257_76_3678;
   wire n_257_76_3679;
   wire n_257_76_3680;
   wire n_257_76_3681;
   wire n_257_76_3682;
   wire n_257_76_3683;
   wire n_257_76_3684;
   wire n_257_76_3685;
   wire n_257_76_3686;
   wire n_257_76_3687;
   wire n_257_76_3688;
   wire n_257_76_3689;
   wire n_257_76_3690;
   wire n_257_76_3691;
   wire n_257_76_3692;
   wire n_257_76_3693;
   wire n_257_76_3694;
   wire n_257_76_3695;
   wire n_257_76_3696;
   wire n_257_76_3697;
   wire n_257_76_3698;
   wire n_257_76_3699;
   wire n_257_76_3700;
   wire n_257_76_3701;
   wire n_257_76_3702;
   wire n_257_76_3703;
   wire n_257_76_3704;
   wire n_257_76_3705;
   wire n_257_76_3706;
   wire n_257_76_3707;
   wire n_257_76_3708;
   wire n_257_76_3709;
   wire n_257_76_3710;
   wire n_257_76_3711;
   wire n_257_76_3712;
   wire n_257_76_3713;
   wire n_257_76_3714;
   wire n_257_76_3715;
   wire n_257_76_3716;
   wire n_257_76_3717;
   wire n_257_76_3718;
   wire n_257_76_3719;
   wire n_257_76_3720;
   wire n_257_76_3721;
   wire n_257_76_3722;
   wire n_257_76_3723;
   wire n_257_76_3724;
   wire n_257_76_3725;
   wire n_257_76_3726;
   wire n_257_76_3727;
   wire n_257_76_3728;
   wire n_257_76_3729;
   wire n_257_76_3730;
   wire n_257_76_3731;
   wire n_257_76_3732;
   wire n_257_76_3733;
   wire n_257_76_3734;
   wire n_257_76_3735;
   wire n_257_76_3736;
   wire n_257_76_3737;
   wire n_257_76_3738;
   wire n_257_76_3739;
   wire n_257_76_3740;
   wire n_257_76_3741;
   wire n_257_76_3742;
   wire n_257_76_3743;
   wire n_257_76_3744;
   wire n_257_76_3745;
   wire n_257_76_3746;
   wire n_257_76_3747;
   wire n_257_76_3748;
   wire n_257_76_3749;
   wire n_257_76_3750;
   wire n_257_76_3751;
   wire n_257_76_3752;
   wire n_257_76_3753;
   wire n_257_76_3754;
   wire n_257_76_3755;
   wire n_257_76_3756;
   wire n_257_76_3757;
   wire n_257_76_3758;
   wire n_257_76_3759;
   wire n_257_76_3760;
   wire n_257_76_3761;
   wire n_257_76_3762;
   wire n_257_76_3763;
   wire n_257_76_3764;
   wire n_257_76_3765;
   wire n_257_76_3766;
   wire n_257_76_3767;
   wire n_257_76_3768;
   wire n_257_76_3769;
   wire n_257_76_3770;
   wire n_257_76_3771;
   wire n_257_76_3772;
   wire n_257_76_3773;
   wire n_257_76_3774;
   wire n_257_76_3775;
   wire n_257_76_3776;
   wire n_257_76_3777;
   wire n_257_76_3778;
   wire n_257_76_3779;
   wire n_257_76_3780;
   wire n_257_76_3781;
   wire n_257_76_3782;
   wire n_257_76_3783;
   wire n_257_76_3784;
   wire n_257_76_3785;
   wire n_257_76_3786;
   wire n_257_76_3787;
   wire n_257_76_3788;
   wire n_257_76_3789;
   wire n_257_76_3790;
   wire n_257_76_3791;
   wire n_257_76_3792;
   wire n_257_76_3793;
   wire n_257_76_3794;
   wire n_257_76_3795;
   wire n_257_76_3796;
   wire n_257_76_3797;
   wire n_257_76_3798;
   wire n_257_76_3799;
   wire n_257_76_3800;
   wire n_257_76_3801;
   wire n_257_76_3802;
   wire n_257_76_3803;
   wire n_257_76_3804;
   wire n_257_76_3805;
   wire n_257_76_3806;
   wire n_257_76_3807;
   wire n_257_76_3808;
   wire n_257_76_3809;
   wire n_257_76_3810;
   wire n_257_76_3811;
   wire n_257_76_3812;
   wire n_257_76_3813;
   wire n_257_76_3814;
   wire n_257_76_3815;
   wire n_257_76_3816;
   wire n_257_76_3817;
   wire n_257_76_3818;
   wire n_257_76_3819;
   wire n_257_76_3820;
   wire n_257_76_3821;
   wire n_257_76_3822;
   wire n_257_76_3823;
   wire n_257_76_3824;
   wire n_257_76_3825;
   wire n_257_76_3826;
   wire n_257_76_3827;
   wire n_257_76_3828;
   wire n_257_76_3829;
   wire n_257_76_3830;
   wire n_257_76_3831;
   wire n_257_76_3832;
   wire n_257_76_3833;
   wire n_257_76_3834;
   wire n_257_76_3835;
   wire n_257_76_3836;
   wire n_257_76_3837;
   wire n_257_76_3838;
   wire n_257_76_3839;
   wire n_257_76_3840;
   wire n_257_76_3841;
   wire n_257_76_3842;
   wire n_257_76_3843;
   wire n_257_76_3844;
   wire n_257_76_3845;
   wire n_257_76_3846;
   wire n_257_76_3847;
   wire n_257_76_3848;
   wire n_257_76_3849;
   wire n_257_76_3850;
   wire n_257_76_3851;
   wire n_257_76_3852;
   wire n_257_76_3853;
   wire n_257_76_3854;
   wire n_257_76_3855;
   wire n_257_76_3856;
   wire n_257_76_3857;
   wire n_257_76_3858;
   wire n_257_76_3859;
   wire n_257_76_3860;
   wire n_257_76_3861;
   wire n_257_76_3862;
   wire n_257_76_3863;
   wire n_257_76_3864;
   wire n_257_76_3865;
   wire n_257_76_3866;
   wire n_257_76_3867;
   wire n_257_76_3868;
   wire n_257_76_3869;
   wire n_257_76_3870;
   wire n_257_76_3871;
   wire n_257_76_3872;
   wire n_257_76_3873;
   wire n_257_76_3874;
   wire n_257_76_3875;
   wire n_257_76_3876;
   wire n_257_76_3877;
   wire n_257_76_3878;
   wire n_257_76_3879;
   wire n_257_76_3880;
   wire n_257_76_3881;
   wire n_257_76_3882;
   wire n_257_76_3883;
   wire n_257_76_3884;
   wire n_257_76_3885;
   wire n_257_76_3886;
   wire n_257_76_3887;
   wire n_257_76_3888;
   wire n_257_76_3889;
   wire n_257_76_3890;
   wire n_257_76_3891;
   wire n_257_76_3892;
   wire n_257_76_3893;
   wire n_257_76_3894;
   wire n_257_76_3895;
   wire n_257_76_3896;
   wire n_257_76_3897;
   wire n_257_76_3898;
   wire n_257_76_3899;
   wire n_257_76_3900;
   wire n_257_76_3901;
   wire n_257_76_3902;
   wire n_257_76_3903;
   wire n_257_76_3904;
   wire n_257_76_3905;
   wire n_257_76_3906;
   wire n_257_76_3907;
   wire n_257_76_3908;
   wire n_257_76_3909;
   wire n_257_76_3910;
   wire n_257_76_3911;
   wire n_257_76_3912;
   wire n_257_76_3913;
   wire n_257_76_3914;
   wire n_257_76_3915;
   wire n_257_76_3916;
   wire n_257_76_3917;
   wire n_257_76_3918;
   wire n_257_76_3919;
   wire n_257_76_3920;
   wire n_257_76_3921;
   wire n_257_76_3922;
   wire n_257_76_3923;
   wire n_257_76_3924;
   wire n_257_76_3925;
   wire n_257_76_3926;
   wire n_257_76_3927;
   wire n_257_76_3928;
   wire n_257_76_3929;
   wire n_257_76_3930;
   wire n_257_76_3931;
   wire n_257_76_3932;
   wire n_257_76_3933;
   wire n_257_76_3934;
   wire n_257_76_3935;
   wire n_257_76_3936;
   wire n_257_76_3937;
   wire n_257_76_3938;
   wire n_257_76_3939;
   wire n_257_76_3940;
   wire n_257_76_3941;
   wire n_257_76_3942;
   wire n_257_76_3943;
   wire n_257_76_3944;
   wire n_257_76_3945;
   wire n_257_76_3946;
   wire n_257_76_3947;
   wire n_257_76_3948;
   wire n_257_76_3949;
   wire n_257_76_3950;
   wire n_257_76_3951;
   wire n_257_76_3952;
   wire n_257_76_3953;
   wire n_257_76_3954;
   wire n_257_76_3955;
   wire n_257_76_3956;
   wire n_257_76_3957;
   wire n_257_76_3958;
   wire n_257_76_3959;
   wire n_257_76_3960;
   wire n_257_76_3961;
   wire n_257_76_3962;
   wire n_257_76_3963;
   wire n_257_76_3964;
   wire n_257_76_3965;
   wire n_257_76_3966;
   wire n_257_76_3967;
   wire n_257_76_3968;
   wire n_257_76_3969;
   wire n_257_76_3970;
   wire n_257_76_3971;
   wire n_257_76_3972;
   wire n_257_76_3973;
   wire n_257_76_3974;
   wire n_257_76_3975;
   wire n_257_76_3976;
   wire n_257_76_3977;
   wire n_257_76_3978;
   wire n_257_76_3979;
   wire n_257_76_3980;
   wire n_257_76_3981;
   wire n_257_76_3982;
   wire n_257_76_3983;
   wire n_257_76_3984;
   wire n_257_76_3985;
   wire n_257_76_3986;
   wire n_257_76_3987;
   wire n_257_76_3988;
   wire n_257_76_3989;
   wire n_257_76_3990;
   wire n_257_76_3991;
   wire n_257_76_3992;
   wire n_257_76_3993;
   wire n_257_76_3994;
   wire n_257_76_3995;
   wire n_257_76_3996;
   wire n_257_76_3997;
   wire n_257_76_3998;
   wire n_257_76_3999;
   wire n_257_76_4000;
   wire n_257_76_4001;
   wire n_257_76_4002;
   wire n_257_76_4003;
   wire n_257_76_4004;
   wire n_257_76_4005;
   wire n_257_76_4006;
   wire n_257_76_4007;
   wire n_257_76_4008;
   wire n_257_76_4009;
   wire n_257_76_4010;
   wire n_257_76_4011;
   wire n_257_76_4012;
   wire n_257_76_4013;
   wire n_257_76_4014;
   wire n_257_76_4015;
   wire n_257_76_4016;
   wire n_257_76_4017;
   wire n_257_76_4018;
   wire n_257_76_4019;
   wire n_257_76_4020;
   wire n_257_76_4021;
   wire n_257_76_4022;
   wire n_257_76_4023;
   wire n_257_76_4024;
   wire n_257_76_4025;
   wire n_257_76_4026;
   wire n_257_76_4027;
   wire n_257_76_4028;
   wire n_257_76_4029;
   wire n_257_76_4030;
   wire n_257_76_4031;
   wire n_257_76_4032;
   wire n_257_76_4033;
   wire n_257_76_4034;
   wire n_257_76_4035;
   wire n_257_76_4036;
   wire n_257_76_4037;
   wire n_257_76_4038;
   wire n_257_76_4039;
   wire n_257_76_4040;
   wire n_257_76_4041;
   wire n_257_76_4042;
   wire n_257_76_4043;
   wire n_257_76_4044;
   wire n_257_76_4045;
   wire n_257_76_4046;
   wire n_257_76_4047;
   wire n_257_76_4048;
   wire n_257_76_4049;
   wire n_257_76_4050;
   wire n_257_76_4051;
   wire n_257_76_4052;
   wire n_257_76_4053;
   wire n_257_76_4054;
   wire n_257_76_4055;
   wire n_257_76_4056;
   wire n_257_76_4057;
   wire n_257_76_4058;
   wire n_257_76_4059;
   wire n_257_76_4060;
   wire n_257_76_4061;
   wire n_257_76_4062;
   wire n_257_76_4063;
   wire n_257_76_4064;
   wire n_257_76_4065;
   wire n_257_76_4066;
   wire n_257_76_4067;
   wire n_257_76_4068;
   wire n_257_76_4069;
   wire n_257_76_4070;
   wire n_257_76_4071;
   wire n_257_76_4072;
   wire n_257_76_4073;
   wire n_257_76_4074;
   wire n_257_76_4075;
   wire n_257_76_4076;
   wire n_257_76_4077;
   wire n_257_76_4078;
   wire n_257_76_4079;
   wire n_257_76_4080;
   wire n_257_76_4081;
   wire n_257_76_4082;
   wire n_257_76_4083;
   wire n_257_76_4084;
   wire n_257_76_4085;
   wire n_257_76_4086;
   wire n_257_76_4087;
   wire n_257_76_4088;
   wire n_257_76_4089;
   wire n_257_76_4090;
   wire n_257_76_4091;
   wire n_257_76_4092;
   wire n_257_76_4093;
   wire n_257_76_4094;
   wire n_257_76_4095;
   wire n_257_76_4096;
   wire n_257_76_4097;
   wire n_257_76_4098;
   wire n_257_76_4099;
   wire n_257_76_4100;
   wire n_257_76_4101;
   wire n_257_76_4102;
   wire n_257_76_4103;
   wire n_257_76_4104;
   wire n_257_76_4105;
   wire n_257_76_4106;
   wire n_257_76_4107;
   wire n_257_76_4108;
   wire n_257_76_4109;
   wire n_257_76_4110;
   wire n_257_76_4111;
   wire n_257_76_4112;
   wire n_257_76_4113;
   wire n_257_76_4114;
   wire n_257_76_4115;
   wire n_257_76_4116;
   wire n_257_76_4117;
   wire n_257_76_4118;
   wire n_257_76_4119;
   wire n_257_76_4120;
   wire n_257_76_4121;
   wire n_257_76_4122;
   wire n_257_76_4123;
   wire n_257_76_4124;
   wire n_257_76_4125;
   wire n_257_76_4126;
   wire n_257_76_4127;
   wire n_257_76_4128;
   wire n_257_76_4129;
   wire n_257_76_4130;
   wire n_257_76_4131;
   wire n_257_76_4132;
   wire n_257_76_4133;
   wire n_257_76_4134;
   wire n_257_76_4135;
   wire n_257_76_4136;
   wire n_257_76_4137;
   wire n_257_76_4138;
   wire n_257_76_4139;
   wire n_257_76_4140;
   wire n_257_76_4141;
   wire n_257_76_4142;
   wire n_257_76_4143;
   wire n_257_76_4144;
   wire n_257_76_4145;
   wire n_257_76_4146;
   wire n_257_76_4147;
   wire n_257_76_4148;
   wire n_257_76_4149;
   wire n_257_76_4150;
   wire n_257_76_4151;
   wire n_257_76_4152;
   wire n_257_76_4153;
   wire n_257_76_4154;
   wire n_257_76_4155;
   wire n_257_76_4156;
   wire n_257_76_4157;
   wire n_257_76_4158;
   wire n_257_76_4159;
   wire n_257_76_4160;
   wire n_257_76_4161;
   wire n_257_76_4162;
   wire n_257_76_4163;
   wire n_257_76_4164;
   wire n_257_76_4165;
   wire n_257_76_4166;
   wire n_257_76_4167;
   wire n_257_76_4168;
   wire n_257_76_4169;
   wire n_257_76_4170;
   wire n_257_76_4171;
   wire n_257_76_4172;
   wire n_257_76_4173;
   wire n_257_76_4174;
   wire n_257_76_4175;
   wire n_257_76_4176;
   wire n_257_76_4177;
   wire n_257_76_4178;
   wire n_257_76_4179;
   wire n_257_76_4180;
   wire n_257_76_4181;
   wire n_257_76_4182;
   wire n_257_76_4183;
   wire n_257_76_4184;
   wire n_257_76_4185;
   wire n_257_76_4186;
   wire n_257_76_4187;
   wire n_257_76_4188;
   wire n_257_76_4189;
   wire n_257_76_4190;
   wire n_257_76_4191;
   wire n_257_76_4192;
   wire n_257_76_4193;
   wire n_257_76_4194;
   wire n_257_76_4195;
   wire n_257_76_4196;
   wire n_257_76_4197;
   wire n_257_76_4198;
   wire n_257_76_4199;
   wire n_257_76_4200;
   wire n_257_76_4201;
   wire n_257_76_4202;
   wire n_257_76_4203;
   wire n_257_76_4204;
   wire n_257_76_4205;
   wire n_257_76_4206;
   wire n_257_76_4207;
   wire n_257_76_4208;
   wire n_257_76_4209;
   wire n_257_76_4210;
   wire n_257_76_4211;
   wire n_257_76_4212;
   wire n_257_76_4213;
   wire n_257_76_4214;
   wire n_257_76_4215;
   wire n_257_76_4216;
   wire n_257_76_4217;
   wire n_257_76_4218;
   wire n_257_76_4219;
   wire n_257_76_4220;
   wire n_257_76_4221;
   wire n_257_76_4222;
   wire n_257_76_4223;
   wire n_257_76_4224;
   wire n_257_76_4225;
   wire n_257_76_4226;
   wire n_257_76_4227;
   wire n_257_76_4228;
   wire n_257_76_4229;
   wire n_257_76_4230;
   wire n_257_76_4231;
   wire n_257_76_4232;
   wire n_257_76_4233;
   wire n_257_76_4234;
   wire n_257_76_4235;
   wire n_257_76_4236;
   wire n_257_76_4237;
   wire n_257_76_4238;
   wire n_257_76_4239;
   wire n_257_76_4240;
   wire n_257_76_4241;
   wire n_257_76_4242;
   wire n_257_76_4243;
   wire n_257_76_4244;
   wire n_257_76_4245;
   wire n_257_76_4246;
   wire n_257_76_4247;
   wire n_257_76_4248;
   wire n_257_76_4249;
   wire n_257_76_4250;
   wire n_257_76_4251;
   wire n_257_76_4252;
   wire n_257_76_4253;
   wire n_257_76_4254;
   wire n_257_76_4255;
   wire n_257_76_4256;
   wire n_257_76_4257;
   wire n_257_76_4258;
   wire n_257_76_4259;
   wire n_257_76_4260;
   wire n_257_76_4261;
   wire n_257_76_4262;
   wire n_257_76_4263;
   wire n_257_76_4264;
   wire n_257_76_4265;
   wire n_257_76_4266;
   wire n_257_76_4267;
   wire n_257_76_4268;
   wire n_257_76_4269;
   wire n_257_76_4270;
   wire n_257_76_4271;
   wire n_257_76_4272;
   wire n_257_76_4273;
   wire n_257_76_4274;
   wire n_257_76_4275;
   wire n_257_76_4276;
   wire n_257_76_4277;
   wire n_257_76_4278;
   wire n_257_76_4279;
   wire n_257_76_4280;
   wire n_257_76_4281;
   wire n_257_76_4282;
   wire n_257_76_4283;
   wire n_257_76_4284;
   wire n_257_76_4285;
   wire n_257_76_4286;
   wire n_257_76_4287;
   wire n_257_76_4288;
   wire n_257_76_4289;
   wire n_257_76_4290;
   wire n_257_76_4291;
   wire n_257_76_4292;
   wire n_257_76_4293;
   wire n_257_76_4294;
   wire n_257_76_4295;
   wire n_257_76_4296;
   wire n_257_76_4297;
   wire n_257_76_4298;
   wire n_257_76_4299;
   wire n_257_76_4300;
   wire n_257_76_4301;
   wire n_257_76_4302;
   wire n_257_76_4303;
   wire n_257_76_4304;
   wire n_257_76_4305;
   wire n_257_76_4306;
   wire n_257_76_4307;
   wire n_257_76_4308;
   wire n_257_76_4309;
   wire n_257_76_4310;
   wire n_257_76_4311;
   wire n_257_76_4312;
   wire n_257_76_4313;
   wire n_257_76_4314;
   wire n_257_76_4315;
   wire n_257_76_4316;
   wire n_257_76_4317;
   wire n_257_76_4318;
   wire n_257_76_4319;
   wire n_257_76_4320;
   wire n_257_76_4321;
   wire n_257_76_4322;
   wire n_257_76_4323;
   wire n_257_76_4324;
   wire n_257_76_4325;
   wire n_257_76_4326;
   wire n_257_76_4327;
   wire n_257_76_4328;
   wire n_257_76_4329;
   wire n_257_76_4330;
   wire n_257_76_4331;
   wire n_257_76_4332;
   wire n_257_76_4333;
   wire n_257_76_4334;
   wire n_257_76_4335;
   wire n_257_76_4336;
   wire n_257_76_4337;
   wire n_257_76_4338;
   wire n_257_76_4339;
   wire n_257_76_4340;
   wire n_257_76_4341;
   wire n_257_76_4342;
   wire n_257_76_4343;
   wire n_257_76_4344;
   wire n_257_76_4345;
   wire n_257_76_4346;
   wire n_257_76_4347;
   wire n_257_76_4348;
   wire n_257_76_4349;
   wire n_257_76_4350;
   wire n_257_76_4351;
   wire n_257_76_4352;
   wire n_257_76_4353;
   wire n_257_76_4354;
   wire n_257_76_4355;
   wire n_257_76_4356;
   wire n_257_76_4357;
   wire n_257_76_4358;
   wire n_257_76_4359;
   wire n_257_76_4360;
   wire n_257_76_4361;
   wire n_257_76_4362;
   wire n_257_76_4363;
   wire n_257_76_4364;
   wire n_257_76_4365;
   wire n_257_76_4366;
   wire n_257_76_4367;
   wire n_257_76_4368;
   wire n_257_76_4369;
   wire n_257_76_4370;
   wire n_257_76_4371;
   wire n_257_76_4372;
   wire n_257_76_4373;
   wire n_257_76_4374;
   wire n_257_76_4375;
   wire n_257_76_4376;
   wire n_257_76_4377;
   wire n_257_76_4378;
   wire n_257_76_4379;
   wire n_257_76_4380;
   wire n_257_76_4381;
   wire n_257_76_4382;
   wire n_257_76_4383;
   wire n_257_76_4384;
   wire n_257_76_4385;
   wire n_257_76_4386;
   wire n_257_76_4387;
   wire n_257_76_4388;
   wire n_257_76_4389;
   wire n_257_76_4390;
   wire n_257_76_4391;
   wire n_257_76_4392;
   wire n_257_76_4393;
   wire n_257_76_4394;
   wire n_257_76_4395;
   wire n_257_76_4396;
   wire n_257_76_4397;
   wire n_257_76_4398;
   wire n_257_76_4399;
   wire n_257_76_4400;
   wire n_257_76_4401;
   wire n_257_76_4402;
   wire n_257_76_4403;
   wire n_257_76_4404;
   wire n_257_76_4405;
   wire n_257_76_4406;
   wire n_257_76_4407;
   wire n_257_76_4408;
   wire n_257_76_4409;
   wire n_257_76_4410;
   wire n_257_76_4411;
   wire n_257_76_4412;
   wire n_257_76_4413;
   wire n_257_76_4414;
   wire n_257_76_4415;
   wire n_257_76_4416;
   wire n_257_76_4417;
   wire n_257_76_4418;
   wire n_257_76_4419;
   wire n_257_76_4420;
   wire n_257_76_4421;
   wire n_257_76_4422;
   wire n_257_76_4423;
   wire n_257_76_4424;
   wire n_257_76_4425;
   wire n_257_76_4426;
   wire n_257_76_4427;
   wire n_257_76_4428;
   wire n_257_76_4429;
   wire n_257_76_4430;
   wire n_257_76_4431;
   wire n_257_76_4432;
   wire n_257_76_4433;
   wire n_257_76_4434;
   wire n_257_76_4435;
   wire n_257_76_4436;
   wire n_257_76_4437;
   wire n_257_76_4438;
   wire n_257_76_4439;
   wire n_257_76_4440;
   wire n_257_76_4441;
   wire n_257_76_4442;
   wire n_257_76_4443;
   wire n_257_76_4444;
   wire n_257_76_4445;
   wire n_257_76_4446;
   wire n_257_76_4447;
   wire n_257_76_4448;
   wire n_257_76_4449;
   wire n_257_76_4450;
   wire n_257_76_4451;
   wire n_257_76_4452;
   wire n_257_76_4453;
   wire n_257_76_4454;
   wire n_257_76_4455;
   wire n_257_76_4456;
   wire n_257_76_4457;
   wire n_257_76_4458;
   wire n_257_76_4459;
   wire n_257_76_4460;
   wire n_257_76_4461;
   wire n_257_76_4462;
   wire n_257_76_4463;
   wire n_257_76_4464;
   wire n_257_76_4465;
   wire n_257_76_4466;
   wire n_257_76_4467;
   wire n_257_76_4468;
   wire n_257_76_4469;
   wire n_257_76_4470;
   wire n_257_76_4471;
   wire n_257_76_4472;
   wire n_257_76_4473;
   wire n_257_76_4474;
   wire n_257_76_4475;
   wire n_257_76_4476;
   wire n_257_76_4477;
   wire n_257_76_4478;
   wire n_257_76_4479;
   wire n_257_76_4480;
   wire n_257_76_4481;
   wire n_257_76_4482;
   wire n_257_76_4483;
   wire n_257_76_4484;
   wire n_257_76_4485;
   wire n_257_76_4486;
   wire n_257_76_4487;
   wire n_257_76_4488;
   wire n_257_76_4489;
   wire n_257_76_4490;
   wire n_257_76_4491;
   wire n_257_76_4492;
   wire n_257_76_4493;
   wire n_257_76_4494;
   wire n_257_76_4495;
   wire n_257_76_4496;
   wire n_257_76_4497;
   wire n_257_76_4498;
   wire n_257_76_4499;
   wire n_257_76_4500;
   wire n_257_76_4501;
   wire n_257_76_4502;
   wire n_257_76_4503;
   wire n_257_76_4504;
   wire n_257_76_4505;
   wire n_257_76_4506;
   wire n_257_76_4507;
   wire n_257_76_4508;
   wire n_257_76_4509;
   wire n_257_76_4510;
   wire n_257_76_4511;
   wire n_257_76_4512;
   wire n_257_76_4513;
   wire n_257_76_4514;
   wire n_257_76_4515;
   wire n_257_76_4516;
   wire n_257_76_4517;
   wire n_257_76_4518;
   wire n_257_76_4519;
   wire n_257_76_4520;
   wire n_257_76_4521;
   wire n_257_76_4522;
   wire n_257_76_4523;
   wire n_257_76_4524;
   wire n_257_76_4525;
   wire n_257_76_4526;
   wire n_257_76_4527;
   wire n_257_76_4528;
   wire n_257_76_4529;
   wire n_257_76_4530;
   wire n_257_76_4531;
   wire n_257_76_4532;
   wire n_257_76_4533;
   wire n_257_76_4534;
   wire n_257_76_4535;
   wire n_257_76_4536;
   wire n_257_76_4537;
   wire n_257_76_4538;
   wire n_257_76_4539;
   wire n_257_76_4540;
   wire n_257_76_4541;
   wire n_257_76_4542;
   wire n_257_76_4543;
   wire n_257_76_4544;
   wire n_257_76_4545;
   wire n_257_76_4546;
   wire n_257_76_4547;
   wire n_257_76_4548;
   wire n_257_76_4549;
   wire n_257_76_4550;
   wire n_257_76_4551;
   wire n_257_76_4552;
   wire n_257_76_4553;
   wire n_257_76_4554;
   wire n_257_76_4555;
   wire n_257_76_4556;
   wire n_257_76_4557;
   wire n_257_76_4558;
   wire n_257_76_4559;
   wire n_257_76_4560;
   wire n_257_76_4561;
   wire n_257_76_4562;
   wire n_257_76_4563;
   wire n_257_76_4564;
   wire n_257_76_4565;
   wire n_257_76_4566;
   wire n_257_76_4567;
   wire n_257_76_4568;
   wire n_257_76_4569;
   wire n_257_76_4570;
   wire n_257_76_4571;
   wire n_257_76_4572;
   wire n_257_76_4573;
   wire n_257_76_4574;
   wire n_257_76_4575;
   wire n_257_76_4576;
   wire n_257_76_4577;
   wire n_257_76_4578;
   wire n_257_76_4579;
   wire n_257_76_4580;
   wire n_257_76_4581;
   wire n_257_76_4582;
   wire n_257_76_4583;
   wire n_257_76_4584;
   wire n_257_76_4585;
   wire n_257_76_4586;
   wire n_257_76_4587;
   wire n_257_76_4588;
   wire n_257_76_4589;
   wire n_257_76_4590;
   wire n_257_76_4591;
   wire n_257_76_4592;
   wire n_257_76_4593;
   wire n_257_76_4594;
   wire n_257_76_4595;
   wire n_257_76_4596;
   wire n_257_76_4597;
   wire n_257_76_4598;
   wire n_257_76_4599;
   wire n_257_76_4600;
   wire n_257_76_4601;
   wire n_257_76_4602;
   wire n_257_76_4603;
   wire n_257_76_4604;
   wire n_257_76_4605;
   wire n_257_76_4606;
   wire n_257_76_4607;
   wire n_257_76_4608;
   wire n_257_76_4609;
   wire n_257_76_4610;
   wire n_257_76_4611;
   wire n_257_76_4612;
   wire n_257_76_4613;
   wire n_257_76_4614;
   wire n_257_76_4615;
   wire n_257_76_4616;
   wire n_257_76_4617;
   wire n_257_76_4618;
   wire n_257_76_4619;
   wire n_257_76_4620;
   wire n_257_76_4621;
   wire n_257_76_4622;
   wire n_257_76_4623;
   wire n_257_76_4624;
   wire n_257_76_4625;
   wire n_257_76_4626;
   wire n_257_76_4627;
   wire n_257_76_4628;
   wire n_257_76_4629;
   wire n_257_76_4630;
   wire n_257_76_4631;
   wire n_257_76_4632;
   wire n_257_76_4633;
   wire n_257_76_4634;
   wire n_257_76_4635;
   wire n_257_76_4636;
   wire n_257_76_4637;
   wire n_257_76_4638;
   wire n_257_76_4639;
   wire n_257_76_4640;
   wire n_257_76_4641;
   wire n_257_76_4642;
   wire n_257_76_4643;
   wire n_257_76_4644;
   wire n_257_76_4645;
   wire n_257_76_4646;
   wire n_257_76_4647;
   wire n_257_76_4648;
   wire n_257_76_4649;
   wire n_257_76_4650;
   wire n_257_76_4651;
   wire n_257_76_4652;
   wire n_257_76_4653;
   wire n_257_76_4654;
   wire n_257_76_4655;
   wire n_257_76_4656;
   wire n_257_76_4657;
   wire n_257_76_4658;
   wire n_257_76_4659;
   wire n_257_76_4660;
   wire n_257_76_4661;
   wire n_257_76_4662;
   wire n_257_76_4663;
   wire n_257_76_4664;
   wire n_257_76_4665;
   wire n_257_76_4666;
   wire n_257_76_4667;
   wire n_257_76_4668;
   wire n_257_76_4669;
   wire n_257_76_4670;
   wire n_257_76_4671;
   wire n_257_76_4672;
   wire n_257_76_4673;
   wire n_257_76_4674;
   wire n_257_76_4675;
   wire n_257_76_4676;
   wire n_257_76_4677;
   wire n_257_76_4678;
   wire n_257_76_4679;
   wire n_257_76_4680;
   wire n_257_76_4681;
   wire n_257_76_4682;
   wire n_257_76_4683;
   wire n_257_76_4684;
   wire n_257_76_4685;
   wire n_257_76_4686;
   wire n_257_76_4687;
   wire n_257_76_4688;
   wire n_257_76_4689;
   wire n_257_76_4690;
   wire n_257_76_4691;
   wire n_257_76_4692;
   wire n_257_76_4693;
   wire n_257_76_4694;
   wire n_257_76_4695;
   wire n_257_76_4696;
   wire n_257_76_4697;
   wire n_257_76_4698;
   wire n_257_76_4699;
   wire n_257_76_4700;
   wire n_257_76_4701;
   wire n_257_76_4702;
   wire n_257_76_4703;
   wire n_257_76_4704;
   wire n_257_76_4705;
   wire n_257_76_4706;
   wire n_257_76_4707;
   wire n_257_76_4708;
   wire n_257_76_4709;
   wire n_257_76_4710;
   wire n_257_76_4711;
   wire n_257_76_4712;
   wire n_257_76_4713;
   wire n_257_76_4714;
   wire n_257_76_4715;
   wire n_257_76_4716;
   wire n_257_76_4717;
   wire n_257_76_4718;
   wire n_257_76_4719;
   wire n_257_76_4720;
   wire n_257_76_4721;
   wire n_257_76_4722;
   wire n_257_76_4723;
   wire n_257_76_4724;
   wire n_257_76_4725;
   wire n_257_76_4726;
   wire n_257_76_4727;
   wire n_257_76_4728;
   wire n_257_76_4729;
   wire n_257_76_4730;
   wire n_257_76_4731;
   wire n_257_76_4732;
   wire n_257_76_4733;
   wire n_257_76_4734;
   wire n_257_76_4735;
   wire n_257_76_4736;
   wire n_257_76_4737;
   wire n_257_76_4738;
   wire n_257_76_4739;
   wire n_257_76_4740;
   wire n_257_76_4741;
   wire n_257_76_4742;
   wire n_257_76_4743;
   wire n_257_76_4744;
   wire n_257_76_4745;
   wire n_257_76_4746;
   wire n_257_76_4747;
   wire n_257_76_4748;
   wire n_257_76_4749;
   wire n_257_76_4750;
   wire n_257_76_4751;
   wire n_257_76_4752;
   wire n_257_76_4753;
   wire n_257_76_4754;
   wire n_257_76_4755;
   wire n_257_76_4756;
   wire n_257_76_4757;
   wire n_257_76_4758;
   wire n_257_76_4759;
   wire n_257_76_4760;
   wire n_257_76_4761;
   wire n_257_76_4762;
   wire n_257_76_4763;
   wire n_257_76_4764;
   wire n_257_76_4765;
   wire n_257_76_4766;
   wire n_257_76_4767;
   wire n_257_76_4768;
   wire n_257_76_4769;
   wire n_257_76_4770;
   wire n_257_76_4771;
   wire n_257_76_4772;
   wire n_257_76_4773;
   wire n_257_76_4774;
   wire n_257_76_4775;
   wire n_257_76_4776;
   wire n_257_76_4777;
   wire n_257_76_4778;
   wire n_257_76_4779;
   wire n_257_76_4780;
   wire n_257_76_4781;
   wire n_257_76_4782;
   wire n_257_76_4783;
   wire n_257_76_4784;
   wire n_257_76_4785;
   wire n_257_76_4786;
   wire n_257_76_4787;
   wire n_257_76_4788;
   wire n_257_76_4789;
   wire n_257_76_4790;
   wire n_257_76_4791;
   wire n_257_76_4792;
   wire n_257_76_4793;
   wire n_257_76_4794;
   wire n_257_76_4795;
   wire n_257_76_4796;
   wire n_257_76_4797;
   wire n_257_76_4798;
   wire n_257_76_4799;
   wire n_257_76_4800;
   wire n_257_76_4801;
   wire n_257_76_4802;
   wire n_257_76_4803;
   wire n_257_76_4804;
   wire n_257_76_4805;
   wire n_257_76_4806;
   wire n_257_76_4807;
   wire n_257_76_4808;
   wire n_257_76_4809;
   wire n_257_76_4810;
   wire n_257_76_4811;
   wire n_257_76_4812;
   wire n_257_76_4813;
   wire n_257_76_4814;
   wire n_257_76_4815;
   wire n_257_76_4816;
   wire n_257_76_4817;
   wire n_257_76_4818;
   wire n_257_76_4819;
   wire n_257_76_4820;
   wire n_257_76_4821;
   wire n_257_76_4822;
   wire n_257_76_4823;
   wire n_257_76_4824;
   wire n_257_76_4825;
   wire n_257_76_4826;
   wire n_257_76_4827;
   wire n_257_76_4828;
   wire n_257_76_4829;
   wire n_257_76_4830;
   wire n_257_76_4831;
   wire n_257_76_4832;
   wire n_257_76_4833;
   wire n_257_76_4834;
   wire n_257_76_4835;
   wire n_257_76_4836;
   wire n_257_76_4837;
   wire n_257_76_4838;
   wire n_257_76_4839;
   wire n_257_76_4840;
   wire n_257_76_4841;
   wire n_257_76_4842;
   wire n_257_76_4843;
   wire n_257_76_4844;
   wire n_257_76_4845;
   wire n_257_76_4846;
   wire n_257_76_4847;
   wire n_257_76_4848;
   wire n_257_76_4849;
   wire n_257_76_4850;
   wire n_257_76_4851;
   wire n_257_76_4852;
   wire n_257_76_4853;
   wire n_257_76_4854;
   wire n_257_76_4855;
   wire n_257_76_4856;
   wire n_257_76_4857;
   wire n_257_76_4858;
   wire n_257_76_4859;
   wire n_257_76_4860;
   wire n_257_76_4861;
   wire n_257_76_4862;
   wire n_257_76_4863;
   wire n_257_76_4864;
   wire n_257_76_4865;
   wire n_257_76_4866;
   wire n_257_76_4867;
   wire n_257_76_4868;
   wire n_257_76_4869;
   wire n_257_76_4870;
   wire n_257_76_4871;
   wire n_257_76_4872;
   wire n_257_76_4873;
   wire n_257_76_4874;
   wire n_257_76_4875;
   wire n_257_76_4876;
   wire n_257_76_4877;
   wire n_257_76_4878;
   wire n_257_76_4879;
   wire n_257_76_4880;
   wire n_257_76_4881;
   wire n_257_76_4882;
   wire n_257_76_4883;
   wire n_257_76_4884;
   wire n_257_76_4885;
   wire n_257_76_4886;
   wire n_257_76_4887;
   wire n_257_76_4888;
   wire n_257_76_4889;
   wire n_257_76_4890;
   wire n_257_76_4891;
   wire n_257_76_4892;
   wire n_257_76_4893;
   wire n_257_76_4894;
   wire n_257_76_4895;
   wire n_257_76_4896;
   wire n_257_76_4897;
   wire n_257_76_4898;
   wire n_257_76_4899;
   wire n_257_76_4900;
   wire n_257_76_4901;
   wire n_257_76_4902;
   wire n_257_76_4903;
   wire n_257_76_4904;
   wire n_257_76_4905;
   wire n_257_76_4906;
   wire n_257_76_4907;
   wire n_257_76_4908;
   wire n_257_76_4909;
   wire n_257_76_4910;
   wire n_257_76_4911;
   wire n_257_76_4912;
   wire n_257_76_4913;
   wire n_257_76_4914;
   wire n_257_76_4915;
   wire n_257_76_4916;
   wire n_257_76_4917;
   wire n_257_76_4918;
   wire n_257_76_4919;
   wire n_257_76_4920;
   wire n_257_76_4921;
   wire n_257_76_4922;
   wire n_257_76_4923;
   wire n_257_76_4924;
   wire n_257_76_4925;
   wire n_257_76_4926;
   wire n_257_76_4927;
   wire n_257_76_4928;
   wire n_257_76_4929;
   wire n_257_76_4930;
   wire n_257_76_4931;
   wire n_257_76_4932;
   wire n_257_76_4933;
   wire n_257_76_4934;
   wire n_257_76_4935;
   wire n_257_76_4936;
   wire n_257_76_4937;
   wire n_257_76_4938;
   wire n_257_76_4939;
   wire n_257_76_4940;
   wire n_257_76_4941;
   wire n_257_76_4942;
   wire n_257_76_4943;
   wire n_257_76_4944;
   wire n_257_76_4945;
   wire n_257_76_4946;
   wire n_257_76_4947;
   wire n_257_76_4948;
   wire n_257_76_4949;
   wire n_257_76_4950;
   wire n_257_76_4951;
   wire n_257_76_4952;
   wire n_257_76_4953;
   wire n_257_76_4954;
   wire n_257_76_4955;
   wire n_257_76_4956;
   wire n_257_76_4957;
   wire n_257_76_4958;
   wire n_257_76_4959;
   wire n_257_76_4960;
   wire n_257_76_4961;
   wire n_257_76_4962;
   wire n_257_76_4963;
   wire n_257_76_4964;
   wire n_257_76_4965;
   wire n_257_76_4966;
   wire n_257_76_4967;
   wire n_257_76_4968;
   wire n_257_76_4969;
   wire n_257_76_4970;
   wire n_257_76_4971;
   wire n_257_76_4972;
   wire n_257_76_4973;
   wire n_257_76_4974;
   wire n_257_76_4975;
   wire n_257_76_4976;
   wire n_257_76_4977;
   wire n_257_76_4978;
   wire n_257_76_4979;
   wire n_257_76_4980;
   wire n_257_76_4981;
   wire n_257_76_4982;
   wire n_257_76_4983;
   wire n_257_76_4984;
   wire n_257_76_4985;
   wire n_257_76_4986;
   wire n_257_76_4987;
   wire n_257_76_4988;
   wire n_257_76_4989;
   wire n_257_76_4990;
   wire n_257_76_4991;
   wire n_257_76_4992;
   wire n_257_76_4993;
   wire n_257_76_4994;
   wire n_257_76_4995;
   wire n_257_76_4996;
   wire n_257_76_4997;
   wire n_257_76_4998;
   wire n_257_76_4999;
   wire n_257_76_5000;
   wire n_257_76_5001;
   wire n_257_76_5002;
   wire n_257_76_5003;
   wire n_257_76_5004;
   wire n_257_76_5005;
   wire n_257_76_5006;
   wire n_257_76_5007;
   wire n_257_76_5008;
   wire n_257_76_5009;
   wire n_257_76_5010;
   wire n_257_76_5011;
   wire n_257_76_5012;
   wire n_257_76_5013;
   wire n_257_76_5014;
   wire n_257_76_5015;
   wire n_257_76_5016;
   wire n_257_76_5017;
   wire n_257_76_5018;
   wire n_257_76_5019;
   wire n_257_76_5020;
   wire n_257_76_5021;
   wire n_257_76_5022;
   wire n_257_76_5023;
   wire n_257_76_5024;
   wire n_257_76_5025;
   wire n_257_76_5026;
   wire n_257_76_5027;
   wire n_257_76_5028;
   wire n_257_76_5029;
   wire n_257_76_5030;
   wire n_257_76_5031;
   wire n_257_76_5032;
   wire n_257_76_5033;
   wire n_257_76_5034;
   wire n_257_76_5035;
   wire n_257_76_5036;
   wire n_257_76_5037;
   wire n_257_76_5038;
   wire n_257_76_5039;
   wire n_257_76_5040;
   wire n_257_76_5041;
   wire n_257_76_5042;
   wire n_257_76_5043;
   wire n_257_76_5044;
   wire n_257_76_5045;
   wire n_257_76_5046;
   wire n_257_76_5047;
   wire n_257_76_5048;
   wire n_257_76_5049;
   wire n_257_76_5050;
   wire n_257_76_5051;
   wire n_257_76_5052;
   wire n_257_76_5053;
   wire n_257_76_5054;
   wire n_257_76_5055;
   wire n_257_76_5056;
   wire n_257_76_5057;
   wire n_257_76_5058;
   wire n_257_76_5059;
   wire n_257_76_5060;
   wire n_257_76_5061;
   wire n_257_76_5062;
   wire n_257_76_5063;
   wire n_257_76_5064;
   wire n_257_76_5065;
   wire n_257_76_5066;
   wire n_257_76_5067;
   wire n_257_76_5068;
   wire n_257_76_5069;
   wire n_257_76_5070;
   wire n_257_76_5071;
   wire n_257_76_5072;
   wire n_257_76_5073;
   wire n_257_76_5074;
   wire n_257_76_5075;
   wire n_257_76_5076;
   wire n_257_76_5077;
   wire n_257_76_5078;
   wire n_257_76_5079;
   wire n_257_76_5080;
   wire n_257_76_5081;
   wire n_257_76_5082;
   wire n_257_76_5083;
   wire n_257_76_5084;
   wire n_257_76_5085;
   wire n_257_76_5086;
   wire n_257_76_5087;
   wire n_257_76_5088;
   wire n_257_76_5089;
   wire n_257_76_5090;
   wire n_257_76_5091;
   wire n_257_76_5092;
   wire n_257_76_5093;
   wire n_257_76_5094;
   wire n_257_76_5095;
   wire n_257_76_5096;
   wire n_257_76_5097;
   wire n_257_76_5098;
   wire n_257_76_5099;
   wire n_257_76_5100;
   wire n_257_76_5101;
   wire n_257_76_5102;
   wire n_257_76_5103;
   wire n_257_76_5104;
   wire n_257_76_5105;
   wire n_257_76_5106;
   wire n_257_76_5107;
   wire n_257_76_5108;
   wire n_257_76_5109;
   wire n_257_76_5110;
   wire n_257_76_5111;
   wire n_257_76_5112;
   wire n_257_76_5113;
   wire n_257_76_5114;
   wire n_257_76_5115;
   wire n_257_76_5116;
   wire n_257_76_5117;
   wire n_257_76_5118;
   wire n_257_76_5119;
   wire n_257_76_5120;
   wire n_257_76_5121;
   wire n_257_76_5122;
   wire n_257_76_5123;
   wire n_257_76_5124;
   wire n_257_76_5125;
   wire n_257_76_5126;
   wire n_257_76_5127;
   wire n_257_76_5128;
   wire n_257_76_5129;
   wire n_257_76_5130;
   wire n_257_76_5131;
   wire n_257_76_5132;
   wire n_257_76_5133;
   wire n_257_76_5134;
   wire n_257_76_5135;
   wire n_257_76_5136;
   wire n_257_76_5137;
   wire n_257_76_5138;
   wire n_257_76_5139;
   wire n_257_76_5140;
   wire n_257_76_5141;
   wire n_257_76_5142;
   wire n_257_76_5143;
   wire n_257_76_5144;
   wire n_257_76_5145;
   wire n_257_76_5146;
   wire n_257_76_5147;
   wire n_257_76_5148;
   wire n_257_76_5149;
   wire n_257_76_5150;
   wire n_257_76_5151;
   wire n_257_76_5152;
   wire n_257_76_5153;
   wire n_257_76_5154;
   wire n_257_76_5155;
   wire n_257_76_5156;
   wire n_257_76_5157;
   wire n_257_76_5158;
   wire n_257_76_5159;
   wire n_257_76_5160;
   wire n_257_76_5161;
   wire n_257_76_5162;
   wire n_257_76_5163;
   wire n_257_76_5164;
   wire n_257_76_5165;
   wire n_257_76_5166;
   wire n_257_76_5167;
   wire n_257_76_5168;
   wire n_257_76_5169;
   wire n_257_76_5170;
   wire n_257_76_5171;
   wire n_257_76_5172;
   wire n_257_76_5173;
   wire n_257_76_5174;
   wire n_257_76_5175;
   wire n_257_76_5176;
   wire n_257_76_5177;
   wire n_257_76_5178;
   wire n_257_76_5179;
   wire n_257_76_5180;
   wire n_257_76_5181;
   wire n_257_76_5182;
   wire n_257_76_5183;
   wire n_257_76_5184;
   wire n_257_76_5185;
   wire n_257_76_5186;
   wire n_257_76_5187;
   wire n_257_76_5188;
   wire n_257_76_5189;
   wire n_257_76_5190;
   wire n_257_76_5191;
   wire n_257_76_5192;
   wire n_257_76_5193;
   wire n_257_76_5194;
   wire n_257_76_5195;
   wire n_257_76_5196;
   wire n_257_76_5197;
   wire n_257_76_5198;
   wire n_257_76_5199;
   wire n_257_76_5200;
   wire n_257_76_5201;
   wire n_257_76_5202;
   wire n_257_76_5203;
   wire n_257_76_5204;
   wire n_257_76_5205;
   wire n_257_76_5206;
   wire n_257_76_5207;
   wire n_257_76_5208;
   wire n_257_76_5209;
   wire n_257_76_5210;
   wire n_257_76_5211;
   wire n_257_76_5212;
   wire n_257_76_5213;
   wire n_257_76_5214;
   wire n_257_76_5215;
   wire n_257_76_5216;
   wire n_257_76_5217;
   wire n_257_76_5218;
   wire n_257_76_5219;
   wire n_257_76_5220;
   wire n_257_76_5221;
   wire n_257_76_5222;
   wire n_257_76_5223;
   wire n_257_76_5224;
   wire n_257_76_5225;
   wire n_257_76_5226;
   wire n_257_76_5227;
   wire n_257_76_5228;
   wire n_257_76_5229;
   wire n_257_76_5230;
   wire n_257_76_5231;
   wire n_257_76_5232;
   wire n_257_76_5233;
   wire n_257_76_5234;
   wire n_257_76_5235;
   wire n_257_76_5236;
   wire n_257_76_5237;
   wire n_257_76_5238;
   wire n_257_76_5239;
   wire n_257_76_5240;
   wire n_257_76_5241;
   wire n_257_76_5242;
   wire n_257_76_5243;
   wire n_257_76_5244;
   wire n_257_76_5245;
   wire n_257_76_5246;
   wire n_257_76_5247;
   wire n_257_76_5248;
   wire n_257_76_5249;
   wire n_257_76_5250;
   wire n_257_76_5251;
   wire n_257_76_5252;
   wire n_257_76_5253;
   wire n_257_76_5254;
   wire n_257_76_5255;
   wire n_257_76_5256;
   wire n_257_76_5257;
   wire n_257_76_5258;
   wire n_257_76_5259;
   wire n_257_76_5260;
   wire n_257_76_5261;
   wire n_257_76_5262;
   wire n_257_76_5263;
   wire n_257_76_5264;
   wire n_257_76_5265;
   wire n_257_76_5266;
   wire n_257_76_5267;
   wire n_257_76_5268;
   wire n_257_76_5269;
   wire n_257_76_5270;
   wire n_257_76_5271;
   wire n_257_76_5272;
   wire n_257_76_5273;
   wire n_257_76_5274;
   wire n_257_76_5275;
   wire n_257_76_5276;
   wire n_257_76_5277;
   wire n_257_76_5278;
   wire n_257_76_5279;
   wire n_257_76_5280;
   wire n_257_76_5281;
   wire n_257_76_5282;
   wire n_257_76_5283;
   wire n_257_76_5284;
   wire n_257_76_5285;
   wire n_257_76_5286;
   wire n_257_76_5287;
   wire n_257_76_5288;
   wire n_257_76_5289;
   wire n_257_76_5290;
   wire n_257_76_5291;
   wire n_257_76_5292;
   wire n_257_76_5293;
   wire n_257_76_5294;
   wire n_257_76_5295;
   wire n_257_76_5296;
   wire n_257_76_5297;
   wire n_257_76_5298;
   wire n_257_76_5299;
   wire n_257_76_5300;
   wire n_257_76_5301;
   wire n_257_76_5302;
   wire n_257_76_5303;
   wire n_257_76_5304;
   wire n_257_76_5305;
   wire n_257_76_5306;
   wire n_257_76_5307;
   wire n_257_76_5308;
   wire n_257_76_5309;
   wire n_257_76_5310;
   wire n_257_76_5311;
   wire n_257_76_5312;
   wire n_257_76_5313;
   wire n_257_76_5314;
   wire n_257_76_5315;
   wire n_257_76_5316;
   wire n_257_76_5317;
   wire n_257_76_5318;
   wire n_257_76_5319;
   wire n_257_76_5320;
   wire n_257_76_5321;
   wire n_257_76_5322;
   wire n_257_76_5323;
   wire n_257_76_5324;
   wire n_257_76_5325;
   wire n_257_76_5326;
   wire n_257_76_5327;
   wire n_257_76_5328;
   wire n_257_76_5329;
   wire n_257_76_5330;
   wire n_257_76_5331;
   wire n_257_76_5332;
   wire n_257_76_5333;
   wire n_257_76_5334;
   wire n_257_76_5335;
   wire n_257_76_5336;
   wire n_257_76_5337;
   wire n_257_76_5338;
   wire n_257_76_5339;
   wire n_257_76_5340;
   wire n_257_76_5341;
   wire n_257_76_5342;
   wire n_257_76_5343;
   wire n_257_76_5344;
   wire n_257_76_5345;
   wire n_257_76_5346;
   wire n_257_76_5347;
   wire n_257_76_5348;
   wire n_257_76_5349;
   wire n_257_76_5350;
   wire n_257_76_5351;
   wire n_257_76_5352;
   wire n_257_76_5353;
   wire n_257_76_5354;
   wire n_257_76_5355;
   wire n_257_76_5356;
   wire n_257_76_5357;
   wire n_257_76_5358;
   wire n_257_76_5359;
   wire n_257_76_5360;
   wire n_257_76_5361;
   wire n_257_76_5362;
   wire n_257_76_5363;
   wire n_257_76_5364;
   wire n_257_76_5365;
   wire n_257_76_5366;
   wire n_257_76_5367;
   wire n_257_76_5368;
   wire n_257_76_5369;
   wire n_257_76_5370;
   wire n_257_76_5371;
   wire n_257_76_5372;
   wire n_257_76_5373;
   wire n_257_76_5374;
   wire n_257_76_5375;
   wire n_257_76_5376;
   wire n_257_76_5377;
   wire n_257_76_5378;
   wire n_257_76_5379;
   wire n_257_76_5380;
   wire n_257_76_5381;
   wire n_257_76_5382;
   wire n_257_76_5383;
   wire n_257_76_5384;
   wire n_257_76_5385;
   wire n_257_76_5386;
   wire n_257_76_5387;
   wire n_257_76_5388;
   wire n_257_76_5389;
   wire n_257_76_5390;
   wire n_257_76_5391;
   wire n_257_76_5392;
   wire n_257_76_5393;
   wire n_257_76_5394;
   wire n_257_76_5395;
   wire n_257_76_5396;
   wire n_257_76_5397;
   wire n_257_76_5398;
   wire n_257_76_5399;
   wire n_257_76_5400;
   wire n_257_76_5401;
   wire n_257_76_5402;
   wire n_257_76_5403;
   wire n_257_76_5404;
   wire n_257_76_5405;
   wire n_257_76_5406;
   wire n_257_76_5407;
   wire n_257_76_5408;
   wire n_257_76_5409;
   wire n_257_76_5410;
   wire n_257_76_5411;
   wire n_257_76_5412;
   wire n_257_76_5413;
   wire n_257_76_5414;
   wire n_257_76_5415;
   wire n_257_76_5416;
   wire n_257_76_5417;
   wire n_257_76_5418;
   wire n_257_76_5419;
   wire n_257_76_5420;
   wire n_257_76_5421;
   wire n_257_76_5422;
   wire n_257_76_5423;
   wire n_257_76_5424;
   wire n_257_76_5425;
   wire n_257_76_5426;
   wire n_257_76_5427;
   wire n_257_76_5428;
   wire n_257_76_5429;
   wire n_257_76_5430;
   wire n_257_76_5431;
   wire n_257_76_5432;
   wire n_257_76_5433;
   wire n_257_76_5434;
   wire n_257_76_5435;
   wire n_257_76_5436;
   wire n_257_76_5437;
   wire n_257_76_5438;
   wire n_257_76_5439;
   wire n_257_76_5440;
   wire n_257_76_5441;
   wire n_257_76_5442;
   wire n_257_76_5443;
   wire n_257_76_5444;
   wire n_257_76_5445;
   wire n_257_76_5446;
   wire n_257_76_5447;
   wire n_257_76_5448;
   wire n_257_76_5449;
   wire n_257_76_5450;
   wire n_257_76_5451;
   wire n_257_76_5452;
   wire n_257_76_5453;
   wire n_257_76_5454;
   wire n_257_76_5455;
   wire n_257_76_5456;
   wire n_257_76_5457;
   wire n_257_76_5458;
   wire n_257_76_5459;
   wire n_257_76_5460;
   wire n_257_76_5461;
   wire n_257_76_5462;
   wire n_257_76_5463;
   wire n_257_76_5464;
   wire n_257_76_5465;
   wire n_257_76_5466;
   wire n_257_76_5467;
   wire n_257_76_5468;
   wire n_257_76_5469;
   wire n_257_76_5470;
   wire n_257_76_5471;
   wire n_257_76_5472;
   wire n_257_76_5473;
   wire n_257_76_5474;
   wire n_257_76_5475;
   wire n_257_76_5476;
   wire n_257_76_5477;
   wire n_257_76_5478;
   wire n_257_76_5479;
   wire n_257_76_5480;
   wire n_257_76_5481;
   wire n_257_76_5482;
   wire n_257_76_5483;
   wire n_257_76_5484;
   wire n_257_76_5485;
   wire n_257_76_5486;
   wire n_257_76_5487;
   wire n_257_76_5488;
   wire n_257_76_5489;
   wire n_257_76_5490;
   wire n_257_76_5491;
   wire n_257_76_5492;
   wire n_257_76_5493;
   wire n_257_76_5494;
   wire n_257_76_5495;
   wire n_257_76_5496;
   wire n_257_76_5497;
   wire n_257_76_5498;
   wire n_257_76_5499;
   wire n_257_76_5500;
   wire n_257_76_5501;
   wire n_257_76_5502;
   wire n_257_76_5503;
   wire n_257_76_5504;
   wire n_257_76_5505;
   wire n_257_76_5506;
   wire n_257_76_5507;
   wire n_257_76_5508;
   wire n_257_76_5509;
   wire n_257_76_5510;
   wire n_257_76_5511;
   wire n_257_76_5512;
   wire n_257_76_5513;
   wire n_257_76_5514;
   wire n_257_76_5515;
   wire n_257_76_5516;
   wire n_257_76_5517;
   wire n_257_76_5518;
   wire n_257_76_5519;
   wire n_257_76_5520;
   wire n_257_76_5521;
   wire n_257_76_5522;
   wire n_257_76_5523;
   wire n_257_76_5524;
   wire n_257_76_5525;
   wire n_257_76_5526;
   wire n_257_76_5527;
   wire n_257_76_5528;
   wire n_257_76_5529;
   wire n_257_76_5530;
   wire n_257_76_5531;
   wire n_257_76_5532;
   wire n_257_76_5533;
   wire n_257_76_5534;
   wire n_257_76_5535;
   wire n_257_76_5536;
   wire n_257_76_5537;
   wire n_257_76_5538;
   wire n_257_76_5539;
   wire n_257_76_5540;
   wire n_257_76_5541;
   wire n_257_76_5542;
   wire n_257_76_5543;
   wire n_257_76_5544;
   wire n_257_76_5545;
   wire n_257_76_5546;
   wire n_257_76_5547;
   wire n_257_76_5548;
   wire n_257_76_5549;
   wire n_257_76_5550;
   wire n_257_76_5551;
   wire n_257_76_5552;
   wire n_257_76_5553;
   wire n_257_76_5554;
   wire n_257_76_5555;
   wire n_257_76_5556;
   wire n_257_76_5557;
   wire n_257_76_5558;
   wire n_257_76_5559;
   wire n_257_76_5560;
   wire n_257_76_5561;
   wire n_257_76_5562;
   wire n_257_76_5563;
   wire n_257_76_5564;
   wire n_257_76_5565;
   wire n_257_76_5566;
   wire n_257_76_5567;
   wire n_257_76_5568;
   wire n_257_76_5569;
   wire n_257_76_5570;
   wire n_257_76_5571;
   wire n_257_76_5572;
   wire n_257_76_5573;
   wire n_257_76_5574;
   wire n_257_76_5575;
   wire n_257_76_5576;
   wire n_257_76_5577;
   wire n_257_76_5578;
   wire n_257_76_5579;
   wire n_257_76_5580;
   wire n_257_76_5581;
   wire n_257_76_5582;
   wire n_257_76_5583;
   wire n_257_76_5584;
   wire n_257_76_5585;
   wire n_257_76_5586;
   wire n_257_76_5587;
   wire n_257_76_5588;
   wire n_257_76_5589;
   wire n_257_76_5590;
   wire n_257_76_5591;
   wire n_257_76_5592;
   wire n_257_76_5593;
   wire n_257_76_5594;
   wire n_257_76_5595;
   wire n_257_76_5596;
   wire n_257_76_5597;
   wire n_257_76_5598;
   wire n_257_76_5599;
   wire n_257_76_5600;
   wire n_257_76_5601;
   wire n_257_76_5602;
   wire n_257_76_5603;
   wire n_257_76_5604;
   wire n_257_76_5605;
   wire n_257_76_5606;
   wire n_257_76_5607;
   wire n_257_76_5608;
   wire n_257_76_5609;
   wire n_257_76_5610;
   wire n_257_76_5611;
   wire n_257_76_5612;
   wire n_257_76_5613;
   wire n_257_76_5614;
   wire n_257_76_5615;
   wire n_257_76_5616;
   wire n_257_76_5617;
   wire n_257_76_5618;
   wire n_257_76_5619;
   wire n_257_76_5620;
   wire n_257_76_5621;
   wire n_257_76_5622;
   wire n_257_76_5623;
   wire n_257_76_5624;
   wire n_257_76_5625;
   wire n_257_76_5626;
   wire n_257_76_5627;
   wire n_257_76_5628;
   wire n_257_76_5629;
   wire n_257_76_5630;
   wire n_257_76_5631;
   wire n_257_76_5632;
   wire n_257_76_5633;
   wire n_257_76_5634;
   wire n_257_76_5635;
   wire n_257_76_5636;
   wire n_257_76_5637;
   wire n_257_76_5638;
   wire n_257_76_5639;
   wire n_257_76_5640;
   wire n_257_76_5641;
   wire n_257_76_5642;
   wire n_257_76_5643;
   wire n_257_76_5644;
   wire n_257_76_5645;
   wire n_257_76_5646;
   wire n_257_76_5647;
   wire n_257_76_5648;
   wire n_257_76_5649;
   wire n_257_76_5650;
   wire n_257_76_5651;
   wire n_257_76_5652;
   wire n_257_76_5653;
   wire n_257_76_5654;
   wire n_257_76_5655;
   wire n_257_76_5656;
   wire n_257_76_5657;
   wire n_257_76_5658;
   wire n_257_76_5659;
   wire n_257_76_5660;
   wire n_257_76_5661;
   wire n_257_76_5662;
   wire n_257_76_5663;
   wire n_257_76_5664;
   wire n_257_76_5665;
   wire n_257_76_5666;
   wire n_257_76_5667;
   wire n_257_76_5668;
   wire n_257_76_5669;
   wire n_257_76_5670;
   wire n_257_76_5671;
   wire n_257_76_5672;
   wire n_257_76_5673;
   wire n_257_76_5674;
   wire n_257_76_5675;
   wire n_257_76_5676;
   wire n_257_76_5677;
   wire n_257_76_5678;
   wire n_257_76_5679;
   wire n_257_76_5680;
   wire n_257_76_5681;
   wire n_257_76_5682;
   wire n_257_76_5683;
   wire n_257_76_5684;
   wire n_257_76_5685;
   wire n_257_76_5686;
   wire n_257_76_5687;
   wire n_257_76_5688;
   wire n_257_76_5689;
   wire n_257_76_5690;
   wire n_257_76_5691;
   wire n_257_76_5692;
   wire n_257_76_5693;
   wire n_257_76_5694;
   wire n_257_76_5695;
   wire n_257_76_5696;
   wire n_257_76_5697;
   wire n_257_76_5698;
   wire n_257_76_5699;
   wire n_257_76_5700;
   wire n_257_76_5701;
   wire n_257_76_5702;
   wire n_257_76_5703;
   wire n_257_76_5704;
   wire n_257_76_5705;
   wire n_257_76_5706;
   wire n_257_76_5707;
   wire n_257_76_5708;
   wire n_257_76_5709;
   wire n_257_76_5710;
   wire n_257_76_5711;
   wire n_257_76_5712;
   wire n_257_76_5713;
   wire n_257_76_5714;
   wire n_257_76_5715;
   wire n_257_76_5716;
   wire n_257_76_5717;
   wire n_257_76_5718;
   wire n_257_76_5719;
   wire n_257_76_5720;
   wire n_257_76_5721;
   wire n_257_76_5722;
   wire n_257_76_5723;
   wire n_257_76_5724;
   wire n_257_76_5725;
   wire n_257_76_5726;
   wire n_257_76_5727;
   wire n_257_76_5728;
   wire n_257_76_5729;
   wire n_257_76_5730;
   wire n_257_76_5731;
   wire n_257_76_5732;
   wire n_257_76_5733;
   wire n_257_76_5734;
   wire n_257_76_5735;
   wire n_257_76_5736;
   wire n_257_76_5737;
   wire n_257_76_5738;
   wire n_257_76_5739;
   wire n_257_76_5740;
   wire n_257_76_5741;
   wire n_257_76_5742;
   wire n_257_76_5743;
   wire n_257_76_5744;
   wire n_257_76_5745;
   wire n_257_76_5746;
   wire n_257_76_5747;
   wire n_257_76_5748;
   wire n_257_76_5749;
   wire n_257_76_5750;
   wire n_257_76_5751;
   wire n_257_76_5752;
   wire n_257_76_5753;
   wire n_257_76_5754;
   wire n_257_76_5755;
   wire n_257_76_5756;
   wire n_257_76_5757;
   wire n_257_76_5758;
   wire n_257_76_5759;
   wire n_257_76_5760;
   wire n_257_76_5761;
   wire n_257_76_5762;
   wire n_257_76_5763;
   wire n_257_76_5764;
   wire n_257_76_5765;
   wire n_257_76_5766;
   wire n_257_76_5767;
   wire n_257_76_5768;
   wire n_257_76_5769;
   wire n_257_76_5770;
   wire n_257_76_5771;
   wire n_257_76_5772;
   wire n_257_76_5773;
   wire n_257_76_5774;
   wire n_257_76_5775;
   wire n_257_76_5776;
   wire n_257_76_5777;
   wire n_257_76_5778;
   wire n_257_76_5779;
   wire n_257_76_5780;
   wire n_257_76_5781;
   wire n_257_76_5782;
   wire n_257_76_5783;
   wire n_257_76_5784;
   wire n_257_76_5785;
   wire n_257_76_5786;
   wire n_257_76_5787;
   wire n_257_76_5788;
   wire n_257_76_5789;
   wire n_257_76_5790;
   wire n_257_76_5791;
   wire n_257_76_5792;
   wire n_257_76_5793;
   wire n_257_76_5794;
   wire n_257_76_5795;
   wire n_257_76_5796;
   wire n_257_76_5797;
   wire n_257_76_5798;
   wire n_257_76_5799;
   wire n_257_76_5800;
   wire n_257_76_5801;
   wire n_257_76_5802;
   wire n_257_76_5803;
   wire n_257_76_5804;
   wire n_257_76_5805;
   wire n_257_76_5806;
   wire n_257_76_5807;
   wire n_257_76_5808;
   wire n_257_76_5809;
   wire n_257_76_5810;
   wire n_257_76_5811;
   wire n_257_76_5812;
   wire n_257_76_5813;
   wire n_257_76_5814;
   wire n_257_76_5815;
   wire n_257_76_5816;
   wire n_257_76_5817;
   wire n_257_76_5818;
   wire n_257_76_5819;
   wire n_257_76_5820;
   wire n_257_76_5821;
   wire n_257_76_5822;
   wire n_257_76_5823;
   wire n_257_76_5824;
   wire n_257_76_5825;
   wire n_257_76_5826;
   wire n_257_76_5827;
   wire n_257_76_5828;
   wire n_257_76_5829;
   wire n_257_76_5830;
   wire n_257_76_5831;
   wire n_257_76_5832;
   wire n_257_76_5833;
   wire n_257_76_5834;
   wire n_257_76_5835;
   wire n_257_76_5836;
   wire n_257_76_5837;
   wire n_257_76_5838;
   wire n_257_76_5839;
   wire n_257_76_5840;
   wire n_257_76_5841;
   wire n_257_76_5842;
   wire n_257_76_5843;
   wire n_257_76_5844;
   wire n_257_76_5845;
   wire n_257_76_5846;
   wire n_257_76_5847;
   wire n_257_76_5848;
   wire n_257_76_5849;
   wire n_257_76_5850;
   wire n_257_76_5851;
   wire n_257_76_5852;
   wire n_257_76_5853;
   wire n_257_76_5854;
   wire n_257_76_5855;
   wire n_257_76_5856;
   wire n_257_76_5857;
   wire n_257_76_5858;
   wire n_257_76_5859;
   wire n_257_76_5860;
   wire n_257_76_5861;
   wire n_257_76_5862;
   wire n_257_76_5863;
   wire n_257_76_5864;
   wire n_257_76_5865;
   wire n_257_76_5866;
   wire n_257_76_5867;
   wire n_257_76_5868;
   wire n_257_76_5869;
   wire n_257_76_5870;
   wire n_257_76_5871;
   wire n_257_76_5872;
   wire n_257_76_5873;
   wire n_257_76_5874;
   wire n_257_76_5875;
   wire n_257_76_5876;
   wire n_257_76_5877;
   wire n_257_76_5878;
   wire n_257_76_5879;
   wire n_257_76_5880;
   wire n_257_76_5881;
   wire n_257_76_5882;
   wire n_257_76_5883;
   wire n_257_76_5884;
   wire n_257_76_5885;
   wire n_257_76_5886;
   wire n_257_76_5887;
   wire n_257_76_5888;
   wire n_257_76_5889;
   wire n_257_76_5890;
   wire n_257_76_5891;
   wire n_257_76_5892;
   wire n_257_76_5893;
   wire n_257_76_5894;
   wire n_257_76_5895;
   wire n_257_76_5896;
   wire n_257_76_5897;
   wire n_257_76_5898;
   wire n_257_76_5899;
   wire n_257_76_5900;
   wire n_257_76_5901;
   wire n_257_76_5902;
   wire n_257_76_5903;
   wire n_257_76_5904;
   wire n_257_76_5905;
   wire n_257_76_5906;
   wire n_257_76_5907;
   wire n_257_76_5908;
   wire n_257_76_5909;
   wire n_257_76_5910;
   wire n_257_76_5911;
   wire n_257_76_5912;
   wire n_257_76_5913;
   wire n_257_76_5914;
   wire n_257_76_5915;
   wire n_257_76_5916;
   wire n_257_76_5917;
   wire n_257_76_5918;
   wire n_257_76_5919;
   wire n_257_76_5920;
   wire n_257_76_5921;
   wire n_257_76_5922;
   wire n_257_76_5923;
   wire n_257_76_5924;
   wire n_257_76_5925;
   wire n_257_76_5926;
   wire n_257_76_5927;
   wire n_257_76_5928;
   wire n_257_76_5929;
   wire n_257_76_5930;
   wire n_257_76_5931;
   wire n_257_76_5932;
   wire n_257_76_5933;
   wire n_257_76_5934;
   wire n_257_76_5935;
   wire n_257_76_5936;
   wire n_257_76_5937;
   wire n_257_76_5938;
   wire n_257_76_5939;
   wire n_257_76_5940;
   wire n_257_76_5941;
   wire n_257_76_5942;
   wire n_257_76_5943;
   wire n_257_76_5944;
   wire n_257_76_5945;
   wire n_257_76_5946;
   wire n_257_76_5947;
   wire n_257_76_5948;
   wire n_257_76_5949;
   wire n_257_76_5950;
   wire n_257_76_5951;
   wire n_257_76_5952;
   wire n_257_76_5953;
   wire n_257_76_5954;
   wire n_257_76_5955;
   wire n_257_76_5956;
   wire n_257_76_5957;
   wire n_257_76_5958;
   wire n_257_76_5959;
   wire n_257_76_5960;
   wire n_257_76_5961;
   wire n_257_76_5962;
   wire n_257_76_5963;
   wire n_257_76_5964;
   wire n_257_76_5965;
   wire n_257_76_5966;
   wire n_257_76_5967;
   wire n_257_76_5968;
   wire n_257_76_5969;
   wire n_257_76_5970;
   wire n_257_76_5971;
   wire n_257_76_5972;
   wire n_257_76_5973;
   wire n_257_76_5974;
   wire n_257_76_5975;
   wire n_257_76_5976;
   wire n_257_76_5977;
   wire n_257_76_5978;
   wire n_257_76_5979;
   wire n_257_76_5980;
   wire n_257_76_5981;
   wire n_257_76_5982;
   wire n_257_76_5983;
   wire n_257_76_5984;
   wire n_257_76_5985;
   wire n_257_76_5986;
   wire n_257_76_5987;
   wire n_257_76_5988;
   wire n_257_76_5989;
   wire n_257_76_5990;
   wire n_257_76_5991;
   wire n_257_76_5992;
   wire n_257_76_5993;
   wire n_257_76_5994;
   wire n_257_76_5995;
   wire n_257_76_5996;
   wire n_257_76_5997;
   wire n_257_76_5998;
   wire n_257_76_5999;
   wire n_257_76_6000;
   wire n_257_76_6001;
   wire n_257_76_6002;
   wire n_257_76_6003;
   wire n_257_76_6004;
   wire n_257_76_6005;
   wire n_257_76_6006;
   wire n_257_76_6007;
   wire n_257_76_6008;
   wire n_257_76_6009;
   wire n_257_76_6010;
   wire n_257_76_6011;
   wire n_257_76_6012;
   wire n_257_76_6013;
   wire n_257_76_6014;
   wire n_257_76_6015;
   wire n_257_76_6016;
   wire n_257_76_6017;
   wire n_257_76_6018;
   wire n_257_76_6019;
   wire n_257_76_6020;
   wire n_257_76_6021;
   wire n_257_76_6022;
   wire n_257_76_6023;
   wire n_257_76_6024;
   wire n_257_76_6025;
   wire n_257_76_6026;
   wire n_257_76_6027;
   wire n_257_76_6028;
   wire n_257_76_6029;
   wire n_257_76_6030;
   wire n_257_76_6031;
   wire n_257_76_6032;
   wire n_257_76_6033;
   wire n_257_76_6034;
   wire n_257_76_6035;
   wire n_257_76_6036;
   wire n_257_76_6037;
   wire n_257_76_6038;
   wire n_257_76_6039;
   wire n_257_76_6040;
   wire n_257_76_6041;
   wire n_257_76_6042;
   wire n_257_76_6043;
   wire n_257_76_6044;
   wire n_257_76_6045;
   wire n_257_76_6046;
   wire n_257_76_6047;
   wire n_257_76_6048;
   wire n_257_76_6049;
   wire n_257_76_6050;
   wire n_257_76_6051;
   wire n_257_76_6052;
   wire n_257_76_6053;
   wire n_257_76_6054;
   wire n_257_76_6055;
   wire n_257_76_6056;
   wire n_257_76_6057;
   wire n_257_76_6058;
   wire n_257_76_6059;
   wire n_257_76_6060;
   wire n_257_76_6061;
   wire n_257_76_6062;
   wire n_257_76_6063;
   wire n_257_76_6064;
   wire n_257_76_6065;
   wire n_257_76_6066;
   wire n_257_76_6067;
   wire n_257_76_6068;
   wire n_257_76_6069;
   wire n_257_76_6070;
   wire n_257_76_6071;
   wire n_257_76_6072;
   wire n_257_76_6073;
   wire n_257_76_6074;
   wire n_257_76_6075;
   wire n_257_76_6076;
   wire n_257_76_6077;
   wire n_257_76_6078;
   wire n_257_76_6079;
   wire n_257_76_6080;
   wire n_257_76_6081;
   wire n_257_76_6082;
   wire n_257_76_6083;
   wire n_257_76_6084;
   wire n_257_76_6085;
   wire n_257_76_6086;
   wire n_257_76_6087;
   wire n_257_76_6088;
   wire n_257_76_6089;
   wire n_257_76_6090;
   wire n_257_76_6091;
   wire n_257_76_6092;
   wire n_257_76_6093;
   wire n_257_76_6094;
   wire n_257_76_6095;
   wire n_257_76_6096;
   wire n_257_76_6097;
   wire n_257_76_6098;
   wire n_257_76_6099;
   wire n_257_76_6100;
   wire n_257_76_6101;
   wire n_257_76_6102;
   wire n_257_76_6103;
   wire n_257_76_6104;
   wire n_257_76_6105;
   wire n_257_76_6106;
   wire n_257_76_6107;
   wire n_257_76_6108;
   wire n_257_76_6109;
   wire n_257_76_6110;
   wire n_257_76_6111;
   wire n_257_76_6112;
   wire n_257_76_6113;
   wire n_257_76_6114;
   wire n_257_76_6115;
   wire n_257_76_6116;
   wire n_257_76_6117;
   wire n_257_76_6118;
   wire n_257_76_6119;
   wire n_257_76_6120;
   wire n_257_76_6121;
   wire n_257_76_6122;
   wire n_257_76_6123;
   wire n_257_76_6124;
   wire n_257_76_6125;
   wire n_257_76_6126;
   wire n_257_76_6127;
   wire n_257_76_6128;
   wire n_257_76_6129;
   wire n_257_76_6130;
   wire n_257_76_6131;
   wire n_257_76_6132;
   wire n_257_76_6133;
   wire n_257_76_6134;
   wire n_257_76_6135;
   wire n_257_76_6136;
   wire n_257_76_6137;
   wire n_257_76_6138;
   wire n_257_76_6139;
   wire n_257_76_6140;
   wire n_257_76_6141;
   wire n_257_76_6142;
   wire n_257_76_6143;
   wire n_257_76_6144;
   wire n_257_76_6145;
   wire n_257_76_6146;
   wire n_257_76_6147;
   wire n_257_76_6148;
   wire n_257_76_6149;
   wire n_257_76_6150;
   wire n_257_76_6151;
   wire n_257_76_6152;
   wire n_257_76_6153;
   wire n_257_76_6154;
   wire n_257_76_6155;
   wire n_257_76_6156;
   wire n_257_76_6157;
   wire n_257_76_6158;
   wire n_257_76_6159;
   wire n_257_76_6160;
   wire n_257_76_6161;
   wire n_257_76_6162;
   wire n_257_76_6163;
   wire n_257_76_6164;
   wire n_257_76_6165;
   wire n_257_76_6166;
   wire n_257_76_6167;
   wire n_257_76_6168;
   wire n_257_76_6169;
   wire n_257_76_6170;
   wire n_257_76_6171;
   wire n_257_76_6172;
   wire n_257_76_6173;
   wire n_257_76_6174;
   wire n_257_76_6175;
   wire n_257_76_6176;
   wire n_257_76_6177;
   wire n_257_76_6178;
   wire n_257_76_6179;
   wire n_257_76_6180;
   wire n_257_76_6181;
   wire n_257_76_6182;
   wire n_257_76_6183;
   wire n_257_76_6184;
   wire n_257_76_6185;
   wire n_257_76_6186;
   wire n_257_76_6187;
   wire n_257_76_6188;
   wire n_257_76_6189;
   wire n_257_76_6190;
   wire n_257_76_6191;
   wire n_257_76_6192;
   wire n_257_76_6193;
   wire n_257_76_6194;
   wire n_257_76_6195;
   wire n_257_76_6196;
   wire n_257_76_6197;
   wire n_257_76_6198;
   wire n_257_76_6199;
   wire n_257_76_6200;
   wire n_257_76_6201;
   wire n_257_76_6202;
   wire n_257_76_6203;
   wire n_257_76_6204;
   wire n_257_76_6205;
   wire n_257_76_6206;
   wire n_257_76_6207;
   wire n_257_76_6208;
   wire n_257_76_6209;
   wire n_257_76_6210;
   wire n_257_76_6211;
   wire n_257_76_6212;
   wire n_257_76_6213;
   wire n_257_76_6214;
   wire n_257_76_6215;
   wire n_257_76_6216;
   wire n_257_76_6217;
   wire n_257_76_6218;
   wire n_257_76_6219;
   wire n_257_76_6220;
   wire n_257_76_6221;
   wire n_257_76_6222;
   wire n_257_76_6223;
   wire n_257_76_6224;
   wire n_257_76_6225;
   wire n_257_76_6226;
   wire n_257_76_6227;
   wire n_257_76_6228;
   wire n_257_76_6229;
   wire n_257_76_6230;
   wire n_257_76_6231;
   wire n_257_76_6232;
   wire n_257_76_6233;
   wire n_257_76_6234;
   wire n_257_76_6235;
   wire n_257_76_6236;
   wire n_257_76_6237;
   wire n_257_76_6238;
   wire n_257_76_6239;
   wire n_257_76_6240;
   wire n_257_76_6241;
   wire n_257_76_6242;
   wire n_257_76_6243;
   wire n_257_76_6244;
   wire n_257_76_6245;
   wire n_257_76_6246;
   wire n_257_76_6247;
   wire n_257_76_6248;
   wire n_257_76_6249;
   wire n_257_76_6250;
   wire n_257_76_6251;
   wire n_257_76_6252;
   wire n_257_76_6253;
   wire n_257_76_6254;
   wire n_257_76_6255;
   wire n_257_76_6256;
   wire n_257_76_6257;
   wire n_257_76_6258;
   wire n_257_76_6259;
   wire n_257_76_6260;
   wire n_257_76_6261;
   wire n_257_76_6262;
   wire n_257_76_6263;
   wire n_257_76_6264;
   wire n_257_76_6265;
   wire n_257_76_6266;
   wire n_257_76_6267;
   wire n_257_76_6268;
   wire n_257_76_6269;
   wire n_257_76_6270;
   wire n_257_76_6271;
   wire n_257_76_6272;
   wire n_257_76_6273;
   wire n_257_76_6274;
   wire n_257_76_6275;
   wire n_257_76_6276;
   wire n_257_76_6277;
   wire n_257_76_6278;
   wire n_257_76_6279;
   wire n_257_76_6280;
   wire n_257_76_6281;
   wire n_257_76_6282;
   wire n_257_76_6283;
   wire n_257_76_6284;
   wire n_257_76_6285;
   wire n_257_76_6286;
   wire n_257_76_6287;
   wire n_257_76_6288;
   wire n_257_76_6289;
   wire n_257_76_6290;
   wire n_257_76_6291;
   wire n_257_76_6292;
   wire n_257_76_6293;
   wire n_257_76_6294;
   wire n_257_76_6295;
   wire n_257_76_6296;
   wire n_257_76_6297;
   wire n_257_76_6298;
   wire n_257_76_6299;
   wire n_257_76_6300;
   wire n_257_76_6301;
   wire n_257_76_6302;
   wire n_257_76_6303;
   wire n_257_76_6304;
   wire n_257_76_6305;
   wire n_257_76_6306;
   wire n_257_76_6307;
   wire n_257_76_6308;
   wire n_257_76_6309;
   wire n_257_76_6310;
   wire n_257_76_6311;
   wire n_257_76_6312;
   wire n_257_76_6313;
   wire n_257_76_6314;
   wire n_257_76_6315;
   wire n_257_76_6316;
   wire n_257_76_6317;
   wire n_257_76_6318;
   wire n_257_76_6319;
   wire n_257_76_6320;
   wire n_257_76_6321;
   wire n_257_76_6322;
   wire n_257_76_6323;
   wire n_257_76_6324;
   wire n_257_76_6325;
   wire n_257_76_6326;
   wire n_257_76_6327;
   wire n_257_76_6328;
   wire n_257_76_6329;
   wire n_257_76_6330;
   wire n_257_76_6331;
   wire n_257_76_6332;
   wire n_257_76_6333;
   wire n_257_76_6334;
   wire n_257_76_6335;
   wire n_257_76_6336;
   wire n_257_76_6337;
   wire n_257_76_6338;
   wire n_257_76_6339;
   wire n_257_76_6340;
   wire n_257_76_6341;
   wire n_257_76_6342;
   wire n_257_76_6343;
   wire n_257_76_6344;
   wire n_257_76_6345;
   wire n_257_76_6346;
   wire n_257_76_6347;
   wire n_257_76_6348;
   wire n_257_76_6349;
   wire n_257_76_6350;
   wire n_257_76_6351;
   wire n_257_76_6352;
   wire n_257_76_6353;
   wire n_257_76_6354;
   wire n_257_76_6355;
   wire n_257_76_6356;
   wire n_257_76_6357;
   wire n_257_76_6358;
   wire n_257_76_6359;
   wire n_257_76_6360;
   wire n_257_76_6361;
   wire n_257_76_6362;
   wire n_257_76_6363;
   wire n_257_76_6364;
   wire n_257_76_6365;
   wire n_257_76_6366;
   wire n_257_76_6367;
   wire n_257_76_6368;
   wire n_257_76_6369;
   wire n_257_76_6370;
   wire n_257_76_6371;
   wire n_257_76_6372;
   wire n_257_76_6373;
   wire n_257_76_6374;
   wire n_257_76_6375;
   wire n_257_76_6376;
   wire n_257_76_6377;
   wire n_257_76_6378;
   wire n_257_76_6379;
   wire n_257_76_6380;
   wire n_257_76_6381;
   wire n_257_76_6382;
   wire n_257_76_6383;
   wire n_257_76_6384;
   wire n_257_76_6385;
   wire n_257_76_6386;
   wire n_257_76_6387;
   wire n_257_76_6388;
   wire n_257_76_6389;
   wire n_257_76_6390;
   wire n_257_76_6391;
   wire n_257_76_6392;
   wire n_257_76_6393;
   wire n_257_76_6394;
   wire n_257_76_6395;
   wire n_257_76_6396;
   wire n_257_76_6397;
   wire n_257_76_6398;
   wire n_257_76_6399;
   wire n_257_76_6400;
   wire n_257_76_6401;
   wire n_257_76_6402;
   wire n_257_76_6403;
   wire n_257_76_6404;
   wire n_257_76_6405;
   wire n_257_76_6406;
   wire n_257_76_6407;
   wire n_257_76_6408;
   wire n_257_76_6409;
   wire n_257_76_6410;
   wire n_257_76_6411;
   wire n_257_76_6412;
   wire n_257_76_6413;
   wire n_257_76_6414;
   wire n_257_76_6415;
   wire n_257_76_6416;
   wire n_257_76_6417;
   wire n_257_76_6418;
   wire n_257_76_6419;
   wire n_257_76_6420;
   wire n_257_76_6421;
   wire n_257_76_6422;
   wire n_257_76_6423;
   wire n_257_76_6424;
   wire n_257_76_6425;
   wire n_257_76_6426;
   wire n_257_76_6427;
   wire n_257_76_6428;
   wire n_257_76_6429;
   wire n_257_76_6430;
   wire n_257_76_6431;
   wire n_257_76_6432;
   wire n_257_76_6433;
   wire n_257_76_6434;
   wire n_257_76_6435;
   wire n_257_76_6436;
   wire n_257_76_6437;
   wire n_257_76_6438;
   wire n_257_76_6439;
   wire n_257_76_6440;
   wire n_257_76_6441;
   wire n_257_76_6442;
   wire n_257_76_6443;
   wire n_257_76_6444;
   wire n_257_76_6445;
   wire n_257_76_6446;
   wire n_257_76_6447;
   wire n_257_76_6448;
   wire n_257_76_6449;
   wire n_257_76_6450;
   wire n_257_76_6451;
   wire n_257_76_6452;
   wire n_257_76_6453;
   wire n_257_76_6454;
   wire n_257_76_6455;
   wire n_257_76_6456;
   wire n_257_76_6457;
   wire n_257_76_6458;
   wire n_257_76_6459;
   wire n_257_76_6460;
   wire n_257_76_6461;
   wire n_257_76_6462;
   wire n_257_76_6463;
   wire n_257_76_6464;
   wire n_257_76_6465;
   wire n_257_76_6466;
   wire n_257_76_6467;
   wire n_257_76_6468;
   wire n_257_76_6469;
   wire n_257_76_6470;
   wire n_257_76_6471;
   wire n_257_76_6472;
   wire n_257_76_6473;
   wire n_257_76_6474;
   wire n_257_76_6475;
   wire n_257_76_6476;
   wire n_257_76_6477;
   wire n_257_76_6478;
   wire n_257_76_6479;
   wire n_257_76_6480;
   wire n_257_76_6481;
   wire n_257_76_6482;
   wire n_257_76_6483;
   wire n_257_76_6484;
   wire n_257_76_6485;
   wire n_257_76_6486;
   wire n_257_76_6487;
   wire n_257_76_6488;
   wire n_257_76_6489;
   wire n_257_76_6490;
   wire n_257_76_6491;
   wire n_257_76_6492;
   wire n_257_76_6493;
   wire n_257_76_6494;
   wire n_257_76_6495;
   wire n_257_76_6496;
   wire n_257_76_6497;
   wire n_257_76_6498;
   wire n_257_76_6499;
   wire n_257_76_6500;
   wire n_257_76_6501;
   wire n_257_76_6502;
   wire n_257_76_6503;
   wire n_257_76_6504;
   wire n_257_76_6505;
   wire n_257_76_6506;
   wire n_257_76_6507;
   wire n_257_76_6508;
   wire n_257_76_6509;
   wire n_257_76_6510;
   wire n_257_76_6511;
   wire n_257_76_6512;
   wire n_257_76_6513;
   wire n_257_76_6514;
   wire n_257_76_6515;
   wire n_257_76_6516;
   wire n_257_76_6517;
   wire n_257_76_6518;
   wire n_257_76_6519;
   wire n_257_76_6520;
   wire n_257_76_6521;
   wire n_257_76_6522;
   wire n_257_76_6523;
   wire n_257_76_6524;
   wire n_257_76_6525;
   wire n_257_76_6526;
   wire n_257_76_6527;
   wire n_257_76_6528;
   wire n_257_76_6529;
   wire n_257_76_6530;
   wire n_257_76_6531;
   wire n_257_76_6532;
   wire n_257_76_6533;
   wire n_257_76_6534;
   wire n_257_76_6535;
   wire n_257_76_6536;
   wire n_257_76_6537;
   wire n_257_76_6538;
   wire n_257_76_6539;
   wire n_257_76_6540;
   wire n_257_76_6541;
   wire n_257_76_6542;
   wire n_257_76_6543;
   wire n_257_76_6544;
   wire n_257_76_6545;
   wire n_257_76_6546;
   wire n_257_76_6547;
   wire n_257_76_6548;
   wire n_257_76_6549;
   wire n_257_76_6550;
   wire n_257_76_6551;
   wire n_257_76_6552;
   wire n_257_76_6553;
   wire n_257_76_6554;
   wire n_257_76_6555;
   wire n_257_76_6556;
   wire n_257_76_6557;
   wire n_257_76_6558;
   wire n_257_76_6559;
   wire n_257_76_6560;
   wire n_257_76_6561;
   wire n_257_76_6562;
   wire n_257_76_6563;
   wire n_257_76_6564;
   wire n_257_76_6565;
   wire n_257_76_6566;
   wire n_257_76_6567;
   wire n_257_76_6568;
   wire n_257_76_6569;
   wire n_257_76_6570;
   wire n_257_76_6571;
   wire n_257_76_6572;
   wire n_257_76_6573;
   wire n_257_76_6574;
   wire n_257_76_6575;
   wire n_257_76_6576;
   wire n_257_76_6577;
   wire n_257_76_6578;
   wire n_257_76_6579;
   wire n_257_76_6580;
   wire n_257_76_6581;
   wire n_257_76_6582;
   wire n_257_76_6583;
   wire n_257_76_6584;
   wire n_257_76_6585;
   wire n_257_76_6586;
   wire n_257_76_6587;
   wire n_257_76_6588;
   wire n_257_76_6589;
   wire n_257_76_6590;
   wire n_257_76_6591;
   wire n_257_76_6592;
   wire n_257_76_6593;
   wire n_257_76_6594;
   wire n_257_76_6595;
   wire n_257_76_6596;
   wire n_257_76_6597;
   wire n_257_76_6598;
   wire n_257_76_6599;
   wire n_257_76_6600;
   wire n_257_76_6601;
   wire n_257_76_6602;
   wire n_257_76_6603;
   wire n_257_76_6604;
   wire n_257_76_6605;
   wire n_257_76_6606;
   wire n_257_76_6607;
   wire n_257_76_6608;
   wire n_257_76_6609;
   wire n_257_76_6610;
   wire n_257_76_6611;
   wire n_257_76_6612;
   wire n_257_76_6613;
   wire n_257_76_6614;
   wire n_257_76_6615;
   wire n_257_76_6616;
   wire n_257_76_6617;
   wire n_257_76_6618;
   wire n_257_76_6619;
   wire n_257_76_6620;
   wire n_257_76_6621;
   wire n_257_76_6622;
   wire n_257_76_6623;
   wire n_257_76_6624;
   wire n_257_76_6625;
   wire n_257_76_6626;
   wire n_257_76_6627;
   wire n_257_76_6628;
   wire n_257_76_6629;
   wire n_257_76_6630;
   wire n_257_76_6631;
   wire n_257_76_6632;
   wire n_257_76_6633;
   wire n_257_76_6634;
   wire n_257_76_6635;
   wire n_257_76_6636;
   wire n_257_76_6637;
   wire n_257_76_6638;
   wire n_257_76_6639;
   wire n_257_76_6640;
   wire n_257_76_6641;
   wire n_257_76_6642;
   wire n_257_76_6643;
   wire n_257_76_6644;
   wire n_257_76_6645;
   wire n_257_76_6646;
   wire n_257_76_6647;
   wire n_257_76_6648;
   wire n_257_76_6649;
   wire n_257_76_6650;
   wire n_257_76_6651;
   wire n_257_76_6652;
   wire n_257_76_6653;
   wire n_257_76_6654;
   wire n_257_76_6655;
   wire n_257_76_6656;
   wire n_257_76_6657;
   wire n_257_76_6658;
   wire n_257_76_6659;
   wire n_257_76_6660;
   wire n_257_76_6661;
   wire n_257_76_6662;
   wire n_257_76_6663;
   wire n_257_76_6664;
   wire n_257_76_6665;
   wire n_257_76_6666;
   wire n_257_76_6667;
   wire n_257_76_6668;
   wire n_257_76_6669;
   wire n_257_76_6670;
   wire n_257_76_6671;
   wire n_257_76_6672;
   wire n_257_76_6673;
   wire n_257_76_6674;
   wire n_257_76_6675;
   wire n_257_76_6676;
   wire n_257_76_6677;
   wire n_257_76_6678;
   wire n_257_76_6679;
   wire n_257_76_6680;
   wire n_257_76_6681;
   wire n_257_76_6682;
   wire n_257_76_6683;
   wire n_257_76_6684;
   wire n_257_76_6685;
   wire n_257_76_6686;
   wire n_257_76_6687;
   wire n_257_76_6688;
   wire n_257_76_6689;
   wire n_257_76_6690;
   wire n_257_76_6691;
   wire n_257_76_6692;
   wire n_257_76_6693;
   wire n_257_76_6694;
   wire n_257_76_6695;
   wire n_257_76_6696;
   wire n_257_76_6697;
   wire n_257_76_6698;
   wire n_257_76_6699;
   wire n_257_76_6700;
   wire n_257_76_6701;
   wire n_257_76_6702;
   wire n_257_76_6703;
   wire n_257_76_6704;
   wire n_257_76_6705;
   wire n_257_76_6706;
   wire n_257_76_6707;
   wire n_257_76_6708;
   wire n_257_76_6709;
   wire n_257_76_6710;
   wire n_257_76_6711;
   wire n_257_76_6712;
   wire n_257_76_6713;
   wire n_257_76_6714;
   wire n_257_76_6715;
   wire n_257_76_6716;
   wire n_257_76_6717;
   wire n_257_76_6718;
   wire n_257_76_6719;
   wire n_257_76_6720;
   wire n_257_76_6721;
   wire n_257_76_6722;
   wire n_257_76_6723;
   wire n_257_76_6724;
   wire n_257_76_6725;
   wire n_257_76_6726;
   wire n_257_76_6727;
   wire n_257_76_6728;
   wire n_257_76_6729;
   wire n_257_76_6730;
   wire n_257_76_6731;
   wire n_257_76_6732;
   wire n_257_76_6733;
   wire n_257_76_6734;
   wire n_257_76_6735;
   wire n_257_76_6736;
   wire n_257_76_6737;
   wire n_257_76_6738;
   wire n_257_76_6739;
   wire n_257_76_6740;
   wire n_257_76_6741;
   wire n_257_76_6742;
   wire n_257_76_6743;
   wire n_257_76_6744;
   wire n_257_76_6745;
   wire n_257_76_6746;
   wire n_257_76_6747;
   wire n_257_76_6748;
   wire n_257_76_6749;
   wire n_257_76_6750;
   wire n_257_76_6751;
   wire n_257_76_6752;
   wire n_257_76_6753;
   wire n_257_76_6754;
   wire n_257_76_6755;
   wire n_257_76_6756;
   wire n_257_76_6757;
   wire n_257_76_6758;
   wire n_257_76_6759;
   wire n_257_76_6760;
   wire n_257_76_6761;
   wire n_257_76_6762;
   wire n_257_76_6763;
   wire n_257_76_6764;
   wire n_257_76_6765;
   wire n_257_76_6766;
   wire n_257_76_6767;
   wire n_257_76_6768;
   wire n_257_76_6769;
   wire n_257_76_6770;
   wire n_257_76_6771;
   wire n_257_76_6772;
   wire n_257_76_6773;
   wire n_257_76_6774;
   wire n_257_76_6775;
   wire n_257_76_6776;
   wire n_257_76_6777;
   wire n_257_76_6778;
   wire n_257_76_6779;
   wire n_257_76_6780;
   wire n_257_76_6781;
   wire n_257_76_6782;
   wire n_257_76_6783;
   wire n_257_76_6784;
   wire n_257_76_6785;
   wire n_257_76_6786;
   wire n_257_76_6787;
   wire n_257_76_6788;
   wire n_257_76_6789;
   wire n_257_76_6790;
   wire n_257_76_6791;
   wire n_257_76_6792;
   wire n_257_76_6793;
   wire n_257_76_6794;
   wire n_257_76_6795;
   wire n_257_76_6796;
   wire n_257_76_6797;
   wire n_257_76_6798;
   wire n_257_76_6799;
   wire n_257_76_6800;
   wire n_257_76_6801;
   wire n_257_76_6802;
   wire n_257_76_6803;
   wire n_257_76_6804;
   wire n_257_76_6805;
   wire n_257_76_6806;
   wire n_257_76_6807;
   wire n_257_76_6808;
   wire n_257_76_6809;
   wire n_257_76_6810;
   wire n_257_76_6811;
   wire n_257_76_6812;
   wire n_257_76_6813;
   wire n_257_76_6814;
   wire n_257_76_6815;
   wire n_257_76_6816;
   wire n_257_76_6817;
   wire n_257_76_6818;
   wire n_257_76_6819;
   wire n_257_76_6820;
   wire n_257_76_6821;
   wire n_257_76_6822;
   wire n_257_76_6823;
   wire n_257_76_6824;
   wire n_257_76_6825;
   wire n_257_76_6826;
   wire n_257_76_6827;
   wire n_257_76_6828;
   wire n_257_76_6829;
   wire n_257_76_6830;
   wire n_257_76_6831;
   wire n_257_76_6832;
   wire n_257_76_6833;
   wire n_257_76_6834;
   wire n_257_76_6835;
   wire n_257_76_6836;
   wire n_257_76_6837;
   wire n_257_76_6838;
   wire n_257_76_6839;
   wire n_257_76_6840;
   wire n_257_76_6841;
   wire n_257_76_6842;
   wire n_257_76_6843;
   wire n_257_76_6844;
   wire n_257_76_6845;
   wire n_257_76_6846;
   wire n_257_76_6847;
   wire n_257_76_6848;
   wire n_257_76_6849;
   wire n_257_76_6850;
   wire n_257_76_6851;
   wire n_257_76_6852;
   wire n_257_76_6853;
   wire n_257_76_6854;
   wire n_257_76_6855;
   wire n_257_76_6856;
   wire n_257_76_6857;
   wire n_257_76_6858;
   wire n_257_76_6859;
   wire n_257_76_6860;
   wire n_257_76_6861;
   wire n_257_76_6862;
   wire n_257_76_6863;
   wire n_257_76_6864;
   wire n_257_76_6865;
   wire n_257_76_6866;
   wire n_257_76_6867;
   wire n_257_76_6868;
   wire n_257_76_6869;
   wire n_257_76_6870;
   wire n_257_76_6871;
   wire n_257_76_6872;
   wire n_257_76_6873;
   wire n_257_76_6874;
   wire n_257_76_6875;
   wire n_257_76_6876;
   wire n_257_76_6877;
   wire n_257_76_6878;
   wire n_257_76_6879;
   wire n_257_76_6880;
   wire n_257_76_6881;
   wire n_257_76_6882;
   wire n_257_76_6883;
   wire n_257_76_6884;
   wire n_257_76_6885;
   wire n_257_76_6886;
   wire n_257_76_6887;
   wire n_257_76_6888;
   wire n_257_76_6889;
   wire n_257_76_6890;
   wire n_257_76_6891;
   wire n_257_76_6892;
   wire n_257_76_6893;
   wire n_257_76_6894;
   wire n_257_76_6895;
   wire n_257_76_6896;
   wire n_257_76_6897;
   wire n_257_76_6898;
   wire n_257_76_6899;
   wire n_257_76_6900;
   wire n_257_76_6901;
   wire n_257_76_6902;
   wire n_257_76_6903;
   wire n_257_76_6904;
   wire n_257_76_6905;
   wire n_257_76_6906;
   wire n_257_76_6907;
   wire n_257_76_6908;
   wire n_257_76_6909;
   wire n_257_76_6910;
   wire n_257_76_6911;
   wire n_257_76_6912;
   wire n_257_76_6913;
   wire n_257_76_6914;
   wire n_257_76_6915;
   wire n_257_76_6916;
   wire n_257_76_6917;
   wire n_257_76_6918;
   wire n_257_76_6919;
   wire n_257_76_6920;
   wire n_257_76_6921;
   wire n_257_76_6922;
   wire n_257_76_6923;
   wire n_257_76_6924;
   wire n_257_76_6925;
   wire n_257_76_6926;
   wire n_257_76_6927;
   wire n_257_76_6928;
   wire n_257_76_6929;
   wire n_257_76_6930;
   wire n_257_76_6931;
   wire n_257_76_6932;
   wire n_257_76_6933;
   wire n_257_76_6934;
   wire n_257_76_6935;
   wire n_257_76_6936;
   wire n_257_76_6937;
   wire n_257_76_6938;
   wire n_257_76_6939;
   wire n_257_76_6940;
   wire n_257_76_6941;
   wire n_257_76_6942;
   wire n_257_76_6943;
   wire n_257_76_6944;
   wire n_257_76_6945;
   wire n_257_76_6946;
   wire n_257_76_6947;
   wire n_257_76_6948;
   wire n_257_76_6949;
   wire n_257_76_6950;
   wire n_257_76_6951;
   wire n_257_76_6952;
   wire n_257_76_6953;
   wire n_257_76_6954;
   wire n_257_76_6955;
   wire n_257_76_6956;
   wire n_257_76_6957;
   wire n_257_76_6958;
   wire n_257_76_6959;
   wire n_257_76_6960;
   wire n_257_76_6961;
   wire n_257_76_6962;
   wire n_257_76_6963;
   wire n_257_76_6964;
   wire n_257_76_6965;
   wire n_257_76_6966;
   wire n_257_76_6967;
   wire n_257_76_6968;
   wire n_257_76_6969;
   wire n_257_76_6970;
   wire n_257_76_6971;
   wire n_257_76_6972;
   wire n_257_76_6973;
   wire n_257_76_6974;
   wire n_257_76_6975;
   wire n_257_76_6976;
   wire n_257_76_6977;
   wire n_257_76_6978;
   wire n_257_76_6979;
   wire n_257_76_6980;
   wire n_257_76_6981;
   wire n_257_76_6982;
   wire n_257_76_6983;
   wire n_257_76_6984;
   wire n_257_76_6985;
   wire n_257_76_6986;
   wire n_257_76_6987;
   wire n_257_76_6988;
   wire n_257_76_6989;
   wire n_257_76_6990;
   wire n_257_76_6991;
   wire n_257_76_6992;
   wire n_257_76_6993;
   wire n_257_76_6994;
   wire n_257_76_6995;
   wire n_257_76_6996;
   wire n_257_76_6997;
   wire n_257_76_6998;
   wire n_257_76_6999;
   wire n_257_76_7000;
   wire n_257_76_7001;
   wire n_257_76_7002;
   wire n_257_76_7003;
   wire n_257_76_7004;
   wire n_257_76_7005;
   wire n_257_76_7006;
   wire n_257_76_7007;
   wire n_257_76_7008;
   wire n_257_76_7009;
   wire n_257_76_7010;
   wire n_257_76_7011;
   wire n_257_76_7012;
   wire n_257_76_7013;
   wire n_257_76_7014;
   wire n_257_76_7015;
   wire n_257_76_7016;
   wire n_257_76_7017;
   wire n_257_76_7018;
   wire n_257_76_7019;
   wire n_257_76_7020;
   wire n_257_76_7021;
   wire n_257_76_7022;
   wire n_257_76_7023;
   wire n_257_76_7024;
   wire n_257_76_7025;
   wire n_257_76_7026;
   wire n_257_76_7027;
   wire n_257_76_7028;
   wire n_257_76_7029;
   wire n_257_76_7030;
   wire n_257_76_7031;
   wire n_257_76_7032;
   wire n_257_76_7033;
   wire n_257_76_7034;
   wire n_257_76_7035;
   wire n_257_76_7036;
   wire n_257_76_7037;
   wire n_257_76_7038;
   wire n_257_76_7039;
   wire n_257_76_7040;
   wire n_257_76_7041;
   wire n_257_76_7042;
   wire n_257_76_7043;
   wire n_257_76_7044;
   wire n_257_76_7045;
   wire n_257_76_7046;
   wire n_257_76_7047;
   wire n_257_76_7048;
   wire n_257_76_7049;
   wire n_257_76_7050;
   wire n_257_76_7051;
   wire n_257_76_7052;
   wire n_257_76_7053;
   wire n_257_76_7054;
   wire n_257_76_7055;
   wire n_257_76_7056;
   wire n_257_76_7057;
   wire n_257_76_7058;
   wire n_257_76_7059;
   wire n_257_76_7060;
   wire n_257_76_7061;
   wire n_257_76_7062;
   wire n_257_76_7063;
   wire n_257_76_7064;
   wire n_257_76_7065;
   wire n_257_76_7066;
   wire n_257_76_7067;
   wire n_257_76_7068;
   wire n_257_76_7069;
   wire n_257_76_7070;
   wire n_257_76_7071;
   wire n_257_76_7072;
   wire n_257_76_7073;
   wire n_257_76_7074;
   wire n_257_76_7075;
   wire n_257_76_7076;
   wire n_257_76_7077;
   wire n_257_76_7078;
   wire n_257_76_7079;
   wire n_257_76_7080;
   wire n_257_76_7081;
   wire n_257_76_7082;
   wire n_257_76_7083;
   wire n_257_76_7084;
   wire n_257_76_7085;
   wire n_257_76_7086;
   wire n_257_76_7087;
   wire n_257_76_7088;
   wire n_257_76_7089;
   wire n_257_76_7090;
   wire n_257_76_7091;
   wire n_257_76_7092;
   wire n_257_76_7093;
   wire n_257_76_7094;
   wire n_257_76_7095;
   wire n_257_76_7096;
   wire n_257_76_7097;
   wire n_257_76_7098;
   wire n_257_76_7099;
   wire n_257_76_7100;
   wire n_257_76_7101;
   wire n_257_76_7102;
   wire n_257_76_7103;
   wire n_257_76_7104;
   wire n_257_76_7105;
   wire n_257_76_7106;
   wire n_257_76_7107;
   wire n_257_76_7108;
   wire n_257_76_7109;
   wire n_257_76_7110;
   wire n_257_76_7111;
   wire n_257_76_7112;
   wire n_257_76_7113;
   wire n_257_76_7114;
   wire n_257_76_7115;
   wire n_257_76_7116;
   wire n_257_76_7117;
   wire n_257_76_7118;
   wire n_257_76_7119;
   wire n_257_76_7120;
   wire n_257_76_7121;
   wire n_257_76_7122;
   wire n_257_76_7123;
   wire n_257_76_7124;
   wire n_257_76_7125;
   wire n_257_76_7126;
   wire n_257_76_7127;
   wire n_257_76_7128;
   wire n_257_76_7129;
   wire n_257_76_7130;
   wire n_257_76_7131;
   wire n_257_76_7132;
   wire n_257_76_7133;
   wire n_257_76_7134;
   wire n_257_76_7135;
   wire n_257_76_7136;
   wire n_257_76_7137;
   wire n_257_76_7138;
   wire n_257_76_7139;
   wire n_257_76_7140;
   wire n_257_76_7141;
   wire n_257_76_7142;
   wire n_257_76_7143;
   wire n_257_76_7144;
   wire n_257_76_7145;
   wire n_257_76_7146;
   wire n_257_76_7147;
   wire n_257_76_7148;
   wire n_257_76_7149;
   wire n_257_76_7150;
   wire n_257_76_7151;
   wire n_257_76_7152;
   wire n_257_76_7153;
   wire n_257_76_7154;
   wire n_257_76_7155;
   wire n_257_76_7156;
   wire n_257_76_7157;
   wire n_257_76_7158;
   wire n_257_76_7159;
   wire n_257_76_7160;
   wire n_257_76_7161;
   wire n_257_76_7162;
   wire n_257_76_7163;
   wire n_257_76_7164;
   wire n_257_76_7165;
   wire n_257_76_7166;
   wire n_257_76_7167;
   wire n_257_76_7168;
   wire n_257_76_7169;
   wire n_257_76_7170;
   wire n_257_76_7171;
   wire n_257_76_7172;
   wire n_257_76_7173;
   wire n_257_76_7174;
   wire n_257_76_7175;
   wire n_257_76_7176;
   wire n_257_76_7177;
   wire n_257_76_7178;
   wire n_257_76_7179;
   wire n_257_76_7180;
   wire n_257_76_7181;
   wire n_257_76_7182;
   wire n_257_76_7183;
   wire n_257_76_7184;
   wire n_257_76_7185;
   wire n_257_76_7186;
   wire n_257_76_7187;
   wire n_257_76_7188;
   wire n_257_76_7189;
   wire n_257_76_7190;
   wire n_257_76_7191;
   wire n_257_76_7192;
   wire n_257_76_7193;
   wire n_257_76_7194;
   wire n_257_76_7195;
   wire n_257_76_7196;
   wire n_257_76_7197;
   wire n_257_76_7198;
   wire n_257_76_7199;
   wire n_257_76_7200;
   wire n_257_76_7201;
   wire n_257_76_7202;
   wire n_257_76_7203;
   wire n_257_76_7204;
   wire n_257_76_7205;
   wire n_257_76_7206;
   wire n_257_76_7207;
   wire n_257_76_7208;
   wire n_257_76_7209;
   wire n_257_76_7210;
   wire n_257_76_7211;
   wire n_257_76_7212;
   wire n_257_76_7213;
   wire n_257_76_7214;
   wire n_257_76_7215;
   wire n_257_76_7216;
   wire n_257_76_7217;
   wire n_257_76_7218;
   wire n_257_76_7219;
   wire n_257_76_7220;
   wire n_257_76_7221;
   wire n_257_76_7222;
   wire n_257_76_7223;
   wire n_257_76_7224;
   wire n_257_76_7225;
   wire n_257_76_7226;
   wire n_257_76_7227;
   wire n_257_76_7228;
   wire n_257_76_7229;
   wire n_257_76_7230;
   wire n_257_76_7231;
   wire n_257_76_7232;
   wire n_257_76_7233;
   wire n_257_76_7234;
   wire n_257_76_7235;
   wire n_257_76_7236;
   wire n_257_76_7237;
   wire n_257_76_7238;
   wire n_257_76_7239;
   wire n_257_76_7240;
   wire n_257_76_7241;
   wire n_257_76_7242;
   wire n_257_76_7243;
   wire n_257_76_7244;
   wire n_257_76_7245;
   wire n_257_76_7246;
   wire n_257_76_7247;
   wire n_257_76_7248;
   wire n_257_76_7249;
   wire n_257_76_7250;
   wire n_257_76_7251;
   wire n_257_76_7252;
   wire n_257_76_7253;
   wire n_257_76_7254;
   wire n_257_76_7255;
   wire n_257_76_7256;
   wire n_257_76_7257;
   wire n_257_76_7258;
   wire n_257_76_7259;
   wire n_257_76_7260;
   wire n_257_76_7261;
   wire n_257_76_7262;
   wire n_257_76_7263;
   wire n_257_76_7264;
   wire n_257_76_7265;
   wire n_257_76_7266;
   wire n_257_76_7267;
   wire n_257_76_7268;
   wire n_257_76_7269;
   wire n_257_76_7270;
   wire n_257_76_7271;
   wire n_257_76_7272;
   wire n_257_76_7273;
   wire n_257_76_7274;
   wire n_257_76_7275;
   wire n_257_76_7276;
   wire n_257_76_7277;
   wire n_257_76_7278;
   wire n_257_76_7279;
   wire n_257_76_7280;
   wire n_257_76_7281;
   wire n_257_76_7282;
   wire n_257_76_7283;
   wire n_257_76_7284;
   wire n_257_76_7285;
   wire n_257_76_7286;
   wire n_257_76_7287;
   wire n_257_76_7288;
   wire n_257_76_7289;
   wire n_257_76_7290;
   wire n_257_76_7291;
   wire n_257_76_7292;
   wire n_257_76_7293;
   wire n_257_76_7294;
   wire n_257_76_7295;
   wire n_257_76_7296;
   wire n_257_76_7297;
   wire n_257_76_7298;
   wire n_257_76_7299;
   wire n_257_76_7300;
   wire n_257_76_7301;
   wire n_257_76_7302;
   wire n_257_76_7303;
   wire n_257_76_7304;
   wire n_257_76_7305;
   wire n_257_76_7306;
   wire n_257_76_7307;
   wire n_257_76_7308;
   wire n_257_76_7309;
   wire n_257_76_7310;
   wire n_257_76_7311;
   wire n_257_76_7312;
   wire n_257_76_7313;
   wire n_257_76_7314;
   wire n_257_76_7315;
   wire n_257_76_7316;
   wire n_257_76_7317;
   wire n_257_76_7318;
   wire n_257_76_7319;
   wire n_257_76_7320;
   wire n_257_76_7321;
   wire n_257_76_7322;
   wire n_257_76_7323;
   wire n_257_76_7324;
   wire n_257_76_7325;
   wire n_257_76_7326;
   wire n_257_76_7327;
   wire n_257_76_7328;
   wire n_257_76_7329;
   wire n_257_76_7330;
   wire n_257_76_7331;
   wire n_257_76_7332;
   wire n_257_76_7333;
   wire n_257_76_7334;
   wire n_257_76_7335;
   wire n_257_76_7336;
   wire n_257_76_7337;
   wire n_257_76_7338;
   wire n_257_76_7339;
   wire n_257_76_7340;
   wire n_257_76_7341;
   wire n_257_76_7342;
   wire n_257_76_7343;
   wire n_257_76_7344;
   wire n_257_76_7345;
   wire n_257_76_7346;
   wire n_257_76_7347;
   wire n_257_76_7348;
   wire n_257_76_7349;
   wire n_257_76_7350;
   wire n_257_76_7351;
   wire n_257_76_7352;
   wire n_257_76_7353;
   wire n_257_76_7354;
   wire n_257_76_7355;
   wire n_257_76_7356;
   wire n_257_76_7357;
   wire n_257_76_7358;
   wire n_257_76_7359;
   wire n_257_76_7360;
   wire n_257_76_7361;
   wire n_257_76_7362;
   wire n_257_76_7363;
   wire n_257_76_7364;
   wire n_257_76_7365;
   wire n_257_76_7366;
   wire n_257_76_7367;
   wire n_257_76_7368;
   wire n_257_76_7369;
   wire n_257_76_7370;
   wire n_257_76_7371;
   wire n_257_76_7372;
   wire n_257_76_7373;
   wire n_257_76_7374;
   wire n_257_76_7375;
   wire n_257_76_7376;
   wire n_257_76_7377;
   wire n_257_76_7378;
   wire n_257_76_7379;
   wire n_257_76_7380;
   wire n_257_76_7381;
   wire n_257_76_7382;
   wire n_257_76_7383;
   wire n_257_76_7384;
   wire n_257_76_7385;
   wire n_257_76_7386;
   wire n_257_76_7387;
   wire n_257_76_7388;
   wire n_257_76_7389;
   wire n_257_76_7390;
   wire n_257_76_7391;
   wire n_257_76_7392;
   wire n_257_76_7393;
   wire n_257_76_7394;
   wire n_257_76_7395;
   wire n_257_76_7396;
   wire n_257_76_7397;
   wire n_257_76_7398;
   wire n_257_76_7399;
   wire n_257_76_7400;
   wire n_257_76_7401;
   wire n_257_76_7402;
   wire n_257_76_7403;
   wire n_257_76_7404;
   wire n_257_76_7405;
   wire n_257_76_7406;
   wire n_257_76_7407;
   wire n_257_76_7408;
   wire n_257_76_7409;
   wire n_257_76_7410;
   wire n_257_76_7411;
   wire n_257_76_7412;
   wire n_257_76_7413;
   wire n_257_76_7414;
   wire n_257_76_7415;
   wire n_257_76_7416;
   wire n_257_76_7417;
   wire n_257_76_7418;
   wire n_257_76_7419;
   wire n_257_76_7420;
   wire n_257_76_7421;
   wire n_257_76_7422;
   wire n_257_76_7423;
   wire n_257_76_7424;
   wire n_257_76_7425;
   wire n_257_76_7426;
   wire n_257_76_7427;
   wire n_257_76_7428;
   wire n_257_76_7429;
   wire n_257_76_7430;
   wire n_257_76_7431;
   wire n_257_76_7432;
   wire n_257_76_7433;
   wire n_257_76_7434;
   wire n_257_76_7435;
   wire n_257_76_7436;
   wire n_257_76_7437;
   wire n_257_76_7438;
   wire n_257_76_7439;
   wire n_257_76_7440;
   wire n_257_76_7441;
   wire n_257_76_7442;
   wire n_257_76_7443;
   wire n_257_76_7444;
   wire n_257_76_7445;
   wire n_257_76_7446;
   wire n_257_76_7447;
   wire n_257_76_7448;
   wire n_257_76_7449;
   wire n_257_76_7450;
   wire n_257_76_7451;
   wire n_257_76_7452;
   wire n_257_76_7453;
   wire n_257_76_7454;
   wire n_257_76_7455;
   wire n_257_76_7456;
   wire n_257_76_7457;
   wire n_257_76_7458;
   wire n_257_76_7459;
   wire n_257_76_7460;
   wire n_257_76_7461;
   wire n_257_76_7462;
   wire n_257_76_7463;
   wire n_257_76_7464;
   wire n_257_76_7465;
   wire n_257_76_7466;
   wire n_257_76_7467;
   wire n_257_76_7468;
   wire n_257_76_7469;
   wire n_257_76_7470;
   wire n_257_76_7471;
   wire n_257_76_7472;
   wire n_257_76_7473;
   wire n_257_76_7474;
   wire n_257_76_7475;
   wire n_257_76_7476;
   wire n_257_76_7477;
   wire n_257_76_7478;
   wire n_257_76_7479;
   wire n_257_76_7480;
   wire n_257_76_7481;
   wire n_257_76_7482;
   wire n_257_76_7483;
   wire n_257_76_7484;
   wire n_257_76_7485;
   wire n_257_76_7486;
   wire n_257_76_7487;
   wire n_257_76_7488;
   wire n_257_76_7489;
   wire n_257_76_7490;
   wire n_257_76_7491;
   wire n_257_76_7492;
   wire n_257_76_7493;
   wire n_257_76_7494;
   wire n_257_76_7495;
   wire n_257_76_7496;
   wire n_257_76_7497;
   wire n_257_76_7498;
   wire n_257_76_7499;
   wire n_257_76_7500;
   wire n_257_76_7501;
   wire n_257_76_7502;
   wire n_257_76_7503;
   wire n_257_76_7504;
   wire n_257_76_7505;
   wire n_257_76_7506;
   wire n_257_76_7507;
   wire n_257_76_7508;
   wire n_257_76_7509;
   wire n_257_76_7510;
   wire n_257_76_7511;
   wire n_257_76_7512;
   wire n_257_76_7513;
   wire n_257_76_7514;
   wire n_257_76_7515;
   wire n_257_76_7516;
   wire n_257_76_7517;
   wire n_257_76_7518;
   wire n_257_76_7519;
   wire n_257_76_7520;
   wire n_257_76_7521;
   wire n_257_76_7522;
   wire n_257_76_7523;
   wire n_257_76_7524;
   wire n_257_76_7525;
   wire n_257_76_7526;
   wire n_257_76_7527;
   wire n_257_76_7528;
   wire n_257_76_7529;
   wire n_257_76_7530;
   wire n_257_76_7531;
   wire n_257_76_7532;
   wire n_257_76_7533;
   wire n_257_76_7534;
   wire n_257_76_7535;
   wire n_257_76_7536;
   wire n_257_76_7537;
   wire n_257_76_7538;
   wire n_257_76_7539;
   wire n_257_76_7540;
   wire n_257_76_7541;
   wire n_257_76_7542;
   wire n_257_76_7543;
   wire n_257_76_7544;
   wire n_257_76_7545;
   wire n_257_76_7546;
   wire n_257_76_7547;
   wire n_257_76_7548;
   wire n_257_76_7549;
   wire n_257_76_7550;
   wire n_257_76_7551;
   wire n_257_76_7552;
   wire n_257_76_7553;
   wire n_257_76_7554;
   wire n_257_76_7555;
   wire n_257_76_7556;
   wire n_257_76_7557;
   wire n_257_76_7558;
   wire n_257_76_7559;
   wire n_257_76_7560;
   wire n_257_76_7561;
   wire n_257_76_7562;
   wire n_257_76_7563;
   wire n_257_76_7564;
   wire n_257_76_7565;
   wire n_257_76_7566;
   wire n_257_76_7567;
   wire n_257_76_7568;
   wire n_257_76_7569;
   wire n_257_76_7570;
   wire n_257_76_7571;
   wire n_257_76_7572;
   wire n_257_76_7573;
   wire n_257_76_7574;
   wire n_257_76_7575;
   wire n_257_76_7576;
   wire n_257_76_7577;
   wire n_257_76_7578;
   wire n_257_76_7579;
   wire n_257_76_7580;
   wire n_257_76_7581;
   wire n_257_76_7582;
   wire n_257_76_7583;
   wire n_257_76_7584;
   wire n_257_76_7585;
   wire n_257_76_7586;
   wire n_257_76_7587;
   wire n_257_76_7588;
   wire n_257_76_7589;
   wire n_257_76_7590;
   wire n_257_76_7591;
   wire n_257_76_7592;
   wire n_257_76_7593;
   wire n_257_76_7594;
   wire n_257_76_7595;
   wire n_257_76_7596;
   wire n_257_76_7597;
   wire n_257_76_7598;
   wire n_257_76_7599;
   wire n_257_76_7600;
   wire n_257_76_7601;
   wire n_257_76_7602;
   wire n_257_76_7603;
   wire n_257_76_7604;
   wire n_257_76_7605;
   wire n_257_76_7606;
   wire n_257_76_7607;
   wire n_257_76_7608;
   wire n_257_76_7609;
   wire n_257_76_7610;
   wire n_257_76_7611;
   wire n_257_76_7612;
   wire n_257_76_7613;
   wire n_257_76_7614;
   wire n_257_76_7615;
   wire n_257_76_7616;
   wire n_257_76_7617;
   wire n_257_76_7618;
   wire n_257_76_7619;
   wire n_257_76_7620;
   wire n_257_76_7621;
   wire n_257_76_7622;
   wire n_257_76_7623;
   wire n_257_76_7624;
   wire n_257_76_7625;
   wire n_257_76_7626;
   wire n_257_76_7627;
   wire n_257_76_7628;
   wire n_257_76_7629;
   wire n_257_76_7630;
   wire n_257_76_7631;
   wire n_257_76_7632;
   wire n_257_76_7633;
   wire n_257_76_7634;
   wire n_257_76_7635;
   wire n_257_76_7636;
   wire n_257_76_7637;
   wire n_257_76_7638;
   wire n_257_76_7639;
   wire n_257_76_7640;
   wire n_257_76_7641;
   wire n_257_76_7642;
   wire n_257_76_7643;
   wire n_257_76_7644;
   wire n_257_76_7645;
   wire n_257_76_7646;
   wire n_257_76_7647;
   wire n_257_76_7648;
   wire n_257_76_7649;
   wire n_257_76_7650;
   wire n_257_76_7651;
   wire n_257_76_7652;
   wire n_257_76_7653;
   wire n_257_76_7654;
   wire n_257_76_7655;
   wire n_257_76_7656;
   wire n_257_76_7657;
   wire n_257_76_7658;
   wire n_257_76_7659;
   wire n_257_76_7660;
   wire n_257_76_7661;
   wire n_257_76_7662;
   wire n_257_76_7663;
   wire n_257_76_7664;
   wire n_257_76_7665;
   wire n_257_76_7666;
   wire n_257_76_7667;
   wire n_257_76_7668;
   wire n_257_76_7669;
   wire n_257_76_7670;
   wire n_257_76_7671;
   wire n_257_76_7672;
   wire n_257_76_7673;
   wire n_257_76_7674;
   wire n_257_76_7675;
   wire n_257_76_7676;
   wire n_257_76_7677;
   wire n_257_76_7678;
   wire n_257_76_7679;
   wire n_257_76_7680;
   wire n_257_76_7681;
   wire n_257_76_7682;
   wire n_257_76_7683;
   wire n_257_76_7684;
   wire n_257_76_7685;
   wire n_257_76_7686;
   wire n_257_76_7687;
   wire n_257_76_7688;
   wire n_257_76_7689;
   wire n_257_76_7690;
   wire n_257_76_7691;
   wire n_257_76_7692;
   wire n_257_76_7693;
   wire n_257_76_7694;
   wire n_257_76_7695;
   wire n_257_76_7696;
   wire n_257_76_7697;
   wire n_257_76_7698;
   wire n_257_76_7699;
   wire n_257_76_7700;
   wire n_257_76_7701;
   wire n_257_76_7702;
   wire n_257_76_7703;
   wire n_257_76_7704;
   wire n_257_76_7705;
   wire n_257_76_7706;
   wire n_257_76_7707;
   wire n_257_76_7708;
   wire n_257_76_7709;
   wire n_257_76_7710;
   wire n_257_76_7711;
   wire n_257_76_7712;
   wire n_257_76_7713;
   wire n_257_76_7714;
   wire n_257_76_7715;
   wire n_257_76_7716;
   wire n_257_76_7717;
   wire n_257_76_7718;
   wire n_257_76_7719;
   wire n_257_76_7720;
   wire n_257_76_7721;
   wire n_257_76_7722;
   wire n_257_76_7723;
   wire n_257_76_7724;
   wire n_257_76_7725;
   wire n_257_76_7726;
   wire n_257_76_7727;
   wire n_257_76_7728;
   wire n_257_76_7729;
   wire n_257_76_7730;
   wire n_257_76_7731;
   wire n_257_76_7732;
   wire n_257_76_7733;
   wire n_257_76_7734;
   wire n_257_76_7735;
   wire n_257_76_7736;
   wire n_257_76_7737;
   wire n_257_76_7738;
   wire n_257_76_7739;
   wire n_257_76_7740;
   wire n_257_76_7741;
   wire n_257_76_7742;
   wire n_257_76_7743;
   wire n_257_76_7744;
   wire n_257_76_7745;
   wire n_257_76_7746;
   wire n_257_76_7747;
   wire n_257_76_7748;
   wire n_257_76_7749;
   wire n_257_76_7750;
   wire n_257_76_7751;
   wire n_257_76_7752;
   wire n_257_76_7753;
   wire n_257_76_7754;
   wire n_257_76_7755;
   wire n_257_76_7756;
   wire n_257_76_7757;
   wire n_257_76_7758;
   wire n_257_76_7759;
   wire n_257_76_7760;
   wire n_257_76_7761;
   wire n_257_76_7762;
   wire n_257_76_7763;
   wire n_257_76_7764;
   wire n_257_76_7765;
   wire n_257_76_7766;
   wire n_257_76_7767;
   wire n_257_76_7768;
   wire n_257_76_7769;
   wire n_257_76_7770;
   wire n_257_76_7771;
   wire n_257_76_7772;
   wire n_257_76_7773;
   wire n_257_76_7774;
   wire n_257_76_7775;
   wire n_257_76_7776;
   wire n_257_76_7777;
   wire n_257_76_7778;
   wire n_257_76_7779;
   wire n_257_76_7780;
   wire n_257_76_7781;
   wire n_257_76_7782;
   wire n_257_76_7783;
   wire n_257_76_7784;
   wire n_257_76_7785;
   wire n_257_76_7786;
   wire n_257_76_7787;
   wire n_257_76_7788;
   wire n_257_76_7789;
   wire n_257_76_7790;
   wire n_257_76_7791;
   wire n_257_76_7792;
   wire n_257_76_7793;
   wire n_257_76_7794;
   wire n_257_76_7795;
   wire n_257_76_7796;
   wire n_257_76_7797;
   wire n_257_76_7798;
   wire n_257_76_7799;
   wire n_257_76_7800;
   wire n_257_76_7801;
   wire n_257_76_7802;
   wire n_257_76_7803;
   wire n_257_76_7804;
   wire n_257_76_7805;
   wire n_257_76_7806;
   wire n_257_76_7807;
   wire n_257_76_7808;
   wire n_257_76_7809;
   wire n_257_76_7810;
   wire n_257_76_7811;
   wire n_257_76_7812;
   wire n_257_76_7813;
   wire n_257_76_7814;
   wire n_257_76_7815;
   wire n_257_76_7816;
   wire n_257_76_7817;
   wire n_257_76_7818;
   wire n_257_76_7819;
   wire n_257_76_7820;
   wire n_257_76_7821;
   wire n_257_76_7822;
   wire n_257_76_7823;
   wire n_257_76_7824;
   wire n_257_76_7825;
   wire n_257_76_7826;
   wire n_257_76_7827;
   wire n_257_76_7828;
   wire n_257_76_7829;
   wire n_257_76_7830;
   wire n_257_76_7831;
   wire n_257_76_7832;
   wire n_257_76_7833;
   wire n_257_76_7834;
   wire n_257_76_7835;
   wire n_257_76_7836;
   wire n_257_76_7837;
   wire n_257_76_7838;
   wire n_257_76_7839;
   wire n_257_76_7840;
   wire n_257_76_7841;
   wire n_257_76_7842;
   wire n_257_76_7843;
   wire n_257_76_7844;
   wire n_257_76_7845;
   wire n_257_76_7846;
   wire n_257_76_7847;
   wire n_257_76_7848;
   wire n_257_76_7849;
   wire n_257_76_7850;
   wire n_257_76_7851;
   wire n_257_76_7852;
   wire n_257_76_7853;
   wire n_257_76_7854;
   wire n_257_76_7855;
   wire n_257_76_7856;
   wire n_257_76_7857;
   wire n_257_76_7858;
   wire n_257_76_7859;
   wire n_257_76_7860;
   wire n_257_76_7861;
   wire n_257_76_7862;
   wire n_257_76_7863;
   wire n_257_76_7864;
   wire n_257_76_7865;
   wire n_257_76_7866;
   wire n_257_76_7867;
   wire n_257_76_7868;
   wire n_257_76_7869;
   wire n_257_76_7870;
   wire n_257_76_7871;
   wire n_257_76_7872;
   wire n_257_76_7873;
   wire n_257_76_7874;
   wire n_257_76_7875;
   wire n_257_76_7876;
   wire n_257_76_7877;
   wire n_257_76_7878;
   wire n_257_76_7879;
   wire n_257_76_7880;
   wire n_257_76_7881;
   wire n_257_76_7882;
   wire n_257_76_7883;
   wire n_257_76_7884;
   wire n_257_76_7885;
   wire n_257_76_7886;
   wire n_257_76_7887;
   wire n_257_76_7888;
   wire n_257_76_7889;
   wire n_257_76_7890;
   wire n_257_76_7891;
   wire n_257_76_7892;
   wire n_257_76_7893;
   wire n_257_76_7894;
   wire n_257_76_7895;
   wire n_257_76_7896;
   wire n_257_76_7897;
   wire n_257_76_7898;
   wire n_257_76_7899;
   wire n_257_76_7900;
   wire n_257_76_7901;
   wire n_257_76_7902;
   wire n_257_76_7903;
   wire n_257_76_7904;
   wire n_257_76_7905;
   wire n_257_76_7906;
   wire n_257_76_7907;
   wire n_257_76_7908;
   wire n_257_76_7909;
   wire n_257_76_7910;
   wire n_257_76_7911;
   wire n_257_76_7912;
   wire n_257_76_7913;
   wire n_257_76_7914;
   wire n_257_76_7915;
   wire n_257_76_7916;
   wire n_257_76_7917;
   wire n_257_76_7918;
   wire n_257_76_7919;
   wire n_257_76_7920;
   wire n_257_76_7921;
   wire n_257_76_7922;
   wire n_257_76_7923;
   wire n_257_76_7924;
   wire n_257_76_7925;
   wire n_257_76_7926;
   wire n_257_76_7927;
   wire n_257_76_7928;
   wire n_257_76_7929;
   wire n_257_76_7930;
   wire n_257_76_7931;
   wire n_257_76_7932;
   wire n_257_76_7933;
   wire n_257_76_7934;
   wire n_257_76_7935;
   wire n_257_76_7936;
   wire n_257_76_7937;
   wire n_257_76_7938;
   wire n_257_76_7939;
   wire n_257_76_7940;
   wire n_257_76_7941;
   wire n_257_76_7942;
   wire n_257_76_7943;
   wire n_257_76_7944;
   wire n_257_76_7945;
   wire n_257_76_7946;
   wire n_257_76_7947;
   wire n_257_76_7948;
   wire n_257_76_7949;
   wire n_257_76_7950;
   wire n_257_76_7951;
   wire n_257_76_7952;
   wire n_257_76_7953;
   wire n_257_76_7954;
   wire n_257_76_7955;
   wire n_257_76_7956;
   wire n_257_76_7957;
   wire n_257_76_7958;
   wire n_257_76_7959;
   wire n_257_76_7960;
   wire n_257_76_7961;
   wire n_257_76_7962;
   wire n_257_76_7963;
   wire n_257_76_7964;
   wire n_257_76_7965;
   wire n_257_76_7966;
   wire n_257_76_7967;
   wire n_257_76_7968;
   wire n_257_76_7969;
   wire n_257_76_7970;
   wire n_257_76_7971;
   wire n_257_76_7972;
   wire n_257_76_7973;
   wire n_257_76_7974;
   wire n_257_76_7975;
   wire n_257_76_7976;
   wire n_257_76_7977;
   wire n_257_76_7978;
   wire n_257_76_7979;
   wire n_257_76_7980;
   wire n_257_76_7981;
   wire n_257_76_7982;
   wire n_257_76_7983;
   wire n_257_76_7984;
   wire n_257_76_7985;
   wire n_257_76_7986;
   wire n_257_76_7987;
   wire n_257_76_7988;
   wire n_257_76_7989;
   wire n_257_76_7990;
   wire n_257_76_7991;
   wire n_257_76_7992;
   wire n_257_76_7993;
   wire n_257_76_7994;
   wire n_257_76_7995;
   wire n_257_76_7996;
   wire n_257_76_7997;
   wire n_257_76_7998;
   wire n_257_76_7999;
   wire n_257_76_8000;
   wire n_257_76_8001;
   wire n_257_76_8002;
   wire n_257_76_8003;
   wire n_257_76_8004;
   wire n_257_76_8005;
   wire n_257_76_8006;
   wire n_257_76_8007;
   wire n_257_76_8008;
   wire n_257_76_8009;
   wire n_257_76_8010;
   wire n_257_76_8011;
   wire n_257_76_8012;
   wire n_257_76_8013;
   wire n_257_76_8014;
   wire n_257_76_8015;
   wire n_257_76_8016;
   wire n_257_76_8017;
   wire n_257_76_8018;
   wire n_257_76_8019;
   wire n_257_76_8020;
   wire n_257_76_8021;
   wire n_257_76_8022;
   wire n_257_76_8023;
   wire n_257_76_8024;
   wire n_257_76_8025;
   wire n_257_76_8026;
   wire n_257_76_8027;
   wire n_257_76_8028;
   wire n_257_76_8029;
   wire n_257_76_8030;
   wire n_257_76_8031;
   wire n_257_76_8032;
   wire n_257_76_8033;
   wire n_257_76_8034;
   wire n_257_76_8035;
   wire n_257_76_8036;
   wire n_257_76_8037;
   wire n_257_76_8038;
   wire n_257_76_8039;
   wire n_257_76_8040;
   wire n_257_76_8041;
   wire n_257_76_8042;
   wire n_257_76_8043;
   wire n_257_76_8044;
   wire n_257_76_8045;
   wire n_257_76_8046;
   wire n_257_76_8047;
   wire n_257_76_8048;
   wire n_257_76_8049;
   wire n_257_76_8050;
   wire n_257_76_8051;
   wire n_257_76_8052;
   wire n_257_76_8053;
   wire n_257_76_8054;
   wire n_257_76_8055;
   wire n_257_76_8056;
   wire n_257_76_8057;
   wire n_257_76_8058;
   wire n_257_76_8059;
   wire n_257_76_8060;
   wire n_257_76_8061;
   wire n_257_76_8062;
   wire n_257_76_8063;
   wire n_257_76_8064;
   wire n_257_76_8065;
   wire n_257_76_8066;
   wire n_257_76_8067;
   wire n_257_76_8068;
   wire n_257_76_8069;
   wire n_257_76_8070;
   wire n_257_76_8071;
   wire n_257_76_8072;
   wire n_257_76_8073;
   wire n_257_76_8074;
   wire n_257_76_8075;
   wire n_257_76_8076;
   wire n_257_76_8077;
   wire n_257_76_8078;
   wire n_257_76_8079;
   wire n_257_76_8080;
   wire n_257_76_8081;
   wire n_257_76_8082;
   wire n_257_76_8083;
   wire n_257_76_8084;
   wire n_257_76_8085;
   wire n_257_76_8086;
   wire n_257_76_8087;
   wire n_257_76_8088;
   wire n_257_76_8089;
   wire n_257_76_8090;
   wire n_257_76_8091;
   wire n_257_76_8092;
   wire n_257_76_8093;
   wire n_257_76_8094;
   wire n_257_76_8095;
   wire n_257_76_8096;
   wire n_257_76_8097;
   wire n_257_76_8098;
   wire n_257_76_8099;
   wire n_257_76_8100;
   wire n_257_76_8101;
   wire n_257_76_8102;
   wire n_257_76_8103;
   wire n_257_76_8104;
   wire n_257_76_8105;
   wire n_257_76_8106;
   wire n_257_76_8107;
   wire n_257_76_8108;
   wire n_257_76_8109;
   wire n_257_76_8110;
   wire n_257_76_8111;
   wire n_257_76_8112;
   wire n_257_76_8113;
   wire n_257_76_8114;
   wire n_257_76_8115;
   wire n_257_76_8116;
   wire n_257_76_8117;
   wire n_257_76_8118;
   wire n_257_76_8119;
   wire n_257_76_8120;
   wire n_257_76_8121;
   wire n_257_76_8122;
   wire n_257_76_8123;
   wire n_257_76_8124;
   wire n_257_76_8125;
   wire n_257_76_8126;
   wire n_257_76_8127;
   wire n_257_76_8128;
   wire n_257_76_8129;
   wire n_257_76_8130;
   wire n_257_76_8131;
   wire n_257_76_8132;
   wire n_257_76_8133;
   wire n_257_76_8134;
   wire n_257_76_8135;
   wire n_257_76_8136;
   wire n_257_76_8137;
   wire n_257_76_8138;
   wire n_257_76_8139;
   wire n_257_76_8140;
   wire n_257_76_8141;
   wire n_257_76_8142;
   wire n_257_76_8143;
   wire n_257_76_8144;
   wire n_257_76_8145;
   wire n_257_76_8146;
   wire n_257_76_8147;
   wire n_257_76_8148;
   wire n_257_76_8149;
   wire n_257_76_8150;
   wire n_257_76_8151;
   wire n_257_76_8152;
   wire n_257_76_8153;
   wire n_257_76_8154;
   wire n_257_76_8155;
   wire n_257_76_8156;
   wire n_257_76_8157;
   wire n_257_76_8158;
   wire n_257_76_8159;
   wire n_257_76_8160;
   wire n_257_76_8161;
   wire n_257_76_8162;
   wire n_257_76_8163;
   wire n_257_76_8164;
   wire n_257_76_8165;
   wire n_257_76_8166;
   wire n_257_76_8167;
   wire n_257_76_8168;
   wire n_257_76_8169;
   wire n_257_76_8170;
   wire n_257_76_8171;
   wire n_257_76_8172;
   wire n_257_76_8173;
   wire n_257_76_8174;
   wire n_257_76_8175;
   wire n_257_76_8176;
   wire n_257_76_8177;
   wire n_257_76_8178;
   wire n_257_76_8179;
   wire n_257_76_8180;
   wire n_257_76_8181;
   wire n_257_76_8182;
   wire n_257_76_8183;
   wire n_257_76_8184;
   wire n_257_76_8185;
   wire n_257_76_8186;
   wire n_257_76_8187;
   wire n_257_76_8188;
   wire n_257_76_8189;
   wire n_257_76_8190;
   wire n_257_76_8191;
   wire n_257_76_8192;
   wire n_257_76_8193;
   wire n_257_76_8194;
   wire n_257_76_8195;
   wire n_257_76_8196;
   wire n_257_76_8197;
   wire n_257_76_8198;
   wire n_257_76_8199;
   wire n_257_76_8200;
   wire n_257_76_8201;
   wire n_257_76_8202;
   wire n_257_76_8203;
   wire n_257_76_8204;
   wire n_257_76_8205;
   wire n_257_76_8206;
   wire n_257_76_8207;
   wire n_257_76_8208;
   wire n_257_76_8209;
   wire n_257_76_8210;
   wire n_257_76_8211;
   wire n_257_76_8212;
   wire n_257_76_8213;
   wire n_257_76_8214;
   wire n_257_76_8215;
   wire n_257_76_8216;
   wire n_257_76_8217;
   wire n_257_76_8218;
   wire n_257_76_8219;
   wire n_257_76_8220;
   wire n_257_76_8221;
   wire n_257_76_8222;
   wire n_257_76_8223;
   wire n_257_76_8224;
   wire n_257_76_8225;
   wire n_257_76_8226;
   wire n_257_76_8227;
   wire n_257_76_8228;
   wire n_257_76_8229;
   wire n_257_76_8230;
   wire n_257_76_8231;
   wire n_257_76_8232;
   wire n_257_76_8233;
   wire n_257_76_8234;
   wire n_257_76_8235;
   wire n_257_76_8236;
   wire n_257_76_8237;
   wire n_257_76_8238;
   wire n_257_76_8239;
   wire n_257_76_8240;
   wire n_257_76_8241;
   wire n_257_76_8242;
   wire n_257_76_8243;
   wire n_257_76_8244;
   wire n_257_76_8245;
   wire n_257_76_8246;
   wire n_257_76_8247;
   wire n_257_76_8248;
   wire n_257_76_8249;
   wire n_257_76_8250;
   wire n_257_76_8251;
   wire n_257_76_8252;
   wire n_257_76_8253;
   wire n_257_76_8254;
   wire n_257_76_8255;
   wire n_257_76_8256;
   wire n_257_76_8257;
   wire n_257_76_8258;
   wire n_257_76_8259;
   wire n_257_76_8260;
   wire n_257_76_8261;
   wire n_257_76_8262;
   wire n_257_76_8263;
   wire n_257_76_8264;
   wire n_257_76_8265;
   wire n_257_76_8266;
   wire n_257_76_8267;
   wire n_257_76_8268;
   wire n_257_76_8269;
   wire n_257_76_8270;
   wire n_257_76_8271;
   wire n_257_76_8272;
   wire n_257_76_8273;
   wire n_257_76_8274;
   wire n_257_76_8275;
   wire n_257_76_8276;
   wire n_257_76_8277;
   wire n_257_76_8278;
   wire n_257_76_8279;
   wire n_257_76_8280;
   wire n_257_76_8281;
   wire n_257_76_8282;
   wire n_257_76_8283;
   wire n_257_76_8284;
   wire n_257_76_8285;
   wire n_257_76_8286;
   wire n_257_76_8287;
   wire n_257_76_8288;
   wire n_257_76_8289;
   wire n_257_76_8290;
   wire n_257_76_8291;
   wire n_257_76_8292;
   wire n_257_76_8293;
   wire n_257_76_8294;
   wire n_257_76_8295;
   wire n_257_76_8296;
   wire n_257_76_8297;
   wire n_257_76_8298;
   wire n_257_76_8299;
   wire n_257_76_8300;
   wire n_257_76_8301;
   wire n_257_76_8302;
   wire n_257_76_8303;
   wire n_257_76_8304;
   wire n_257_76_8305;
   wire n_257_76_8306;
   wire n_257_76_8307;
   wire n_257_76_8308;
   wire n_257_76_8309;
   wire n_257_76_8310;
   wire n_257_76_8311;
   wire n_257_76_8312;
   wire n_257_76_8313;
   wire n_257_76_8314;
   wire n_257_76_8315;
   wire n_257_76_8316;
   wire n_257_76_8317;
   wire n_257_76_8318;
   wire n_257_76_8319;
   wire n_257_76_8320;
   wire n_257_76_8321;
   wire n_257_76_8322;
   wire n_257_76_8323;
   wire n_257_76_8324;
   wire n_257_76_8325;
   wire n_257_76_8326;
   wire n_257_76_8327;
   wire n_257_76_8328;
   wire n_257_76_8329;
   wire n_257_76_8330;
   wire n_257_76_8331;
   wire n_257_76_8332;
   wire n_257_76_8333;
   wire n_257_76_8334;
   wire n_257_76_8335;
   wire n_257_76_8336;
   wire n_257_76_8337;
   wire n_257_76_8338;
   wire n_257_76_8339;
   wire n_257_76_8340;
   wire n_257_76_8341;
   wire n_257_76_8342;
   wire n_257_76_8343;
   wire n_257_76_8344;
   wire n_257_76_8345;
   wire n_257_76_8346;
   wire n_257_76_8347;
   wire n_257_76_8348;
   wire n_257_76_8349;
   wire n_257_76_8350;
   wire n_257_76_8351;
   wire n_257_76_8352;
   wire n_257_76_8353;
   wire n_257_76_8354;
   wire n_257_76_8355;
   wire n_257_76_8356;
   wire n_257_76_8357;
   wire n_257_76_8358;
   wire n_257_76_8359;
   wire n_257_76_8360;
   wire n_257_76_8361;
   wire n_257_76_8362;
   wire n_257_76_8363;
   wire n_257_76_8364;
   wire n_257_76_8365;
   wire n_257_76_8366;
   wire n_257_76_8367;
   wire n_257_76_8368;
   wire n_257_76_8369;
   wire n_257_76_8370;
   wire n_257_76_8371;
   wire n_257_76_8372;
   wire n_257_76_8373;
   wire n_257_76_8374;
   wire n_257_76_8375;
   wire n_257_76_8376;
   wire n_257_76_8377;
   wire n_257_76_8378;
   wire n_257_76_8379;
   wire n_257_76_8380;
   wire n_257_76_8381;
   wire n_257_76_8382;
   wire n_257_76_8383;
   wire n_257_76_8384;
   wire n_257_76_8385;
   wire n_257_76_8386;
   wire n_257_76_8387;
   wire n_257_76_8388;
   wire n_257_76_8389;
   wire n_257_76_8390;
   wire n_257_76_8391;
   wire n_257_76_8392;
   wire n_257_76_8393;
   wire n_257_76_8394;
   wire n_257_76_8395;
   wire n_257_76_8396;
   wire n_257_76_8397;
   wire n_257_76_8398;
   wire n_257_76_8399;
   wire n_257_76_8400;
   wire n_257_76_8401;
   wire n_257_76_8402;
   wire n_257_76_8403;
   wire n_257_76_8404;
   wire n_257_76_8405;
   wire n_257_76_8406;
   wire n_257_76_8407;
   wire n_257_76_8408;
   wire n_257_76_8409;
   wire n_257_76_8410;
   wire n_257_76_8411;
   wire n_257_76_8412;
   wire n_257_76_8413;
   wire n_257_76_8414;
   wire n_257_76_8415;
   wire n_257_76_8416;
   wire n_257_76_8417;
   wire n_257_76_8418;
   wire n_257_76_8419;
   wire n_257_76_8420;
   wire n_257_76_8421;
   wire n_257_76_8422;
   wire n_257_76_8423;
   wire n_257_76_8424;
   wire n_257_76_8425;
   wire n_257_76_8426;
   wire n_257_76_8427;
   wire n_257_76_8428;
   wire n_257_76_8429;
   wire n_257_76_8430;
   wire n_257_76_8431;
   wire n_257_76_8432;
   wire n_257_76_8433;
   wire n_257_76_8434;
   wire n_257_76_8435;
   wire n_257_76_8436;
   wire n_257_76_8437;
   wire n_257_76_8438;
   wire n_257_76_8439;
   wire n_257_76_8440;
   wire n_257_76_8441;
   wire n_257_76_8442;
   wire n_257_76_8443;
   wire n_257_76_8444;
   wire n_257_76_8445;
   wire n_257_76_8446;
   wire n_257_76_8447;
   wire n_257_76_8448;
   wire n_257_76_8449;
   wire n_257_76_8450;
   wire n_257_76_8451;
   wire n_257_76_8452;
   wire n_257_76_8453;
   wire n_257_76_8454;
   wire n_257_76_8455;
   wire n_257_76_8456;
   wire n_257_76_8457;
   wire n_257_76_8458;
   wire n_257_76_8459;
   wire n_257_76_8460;
   wire n_257_76_8461;
   wire n_257_76_8462;
   wire n_257_76_8463;
   wire n_257_76_8464;
   wire n_257_76_8465;
   wire n_257_76_8466;
   wire n_257_76_8467;
   wire n_257_76_8468;
   wire n_257_76_8469;
   wire n_257_76_8470;
   wire n_257_76_8471;
   wire n_257_76_8472;
   wire n_257_76_8473;
   wire n_257_76_8474;
   wire n_257_76_8475;
   wire n_257_76_8476;
   wire n_257_76_8477;
   wire n_257_76_8478;
   wire n_257_76_8479;
   wire n_257_76_8480;
   wire n_257_76_8481;
   wire n_257_76_8482;
   wire n_257_76_8483;
   wire n_257_76_8484;
   wire n_257_76_8485;
   wire n_257_76_8486;
   wire n_257_76_8487;
   wire n_257_76_8488;
   wire n_257_76_8489;
   wire n_257_76_8490;
   wire n_257_76_8491;
   wire n_257_76_8492;
   wire n_257_76_8493;
   wire n_257_76_8494;
   wire n_257_76_8495;
   wire n_257_76_8496;
   wire n_257_76_8497;
   wire n_257_76_8498;
   wire n_257_76_8499;
   wire n_257_76_8500;
   wire n_257_76_8501;
   wire n_257_76_8502;
   wire n_257_76_8503;
   wire n_257_76_8504;
   wire n_257_76_8505;
   wire n_257_76_8506;
   wire n_257_76_8507;
   wire n_257_76_8508;
   wire n_257_76_8509;
   wire n_257_76_8510;
   wire n_257_76_8511;
   wire n_257_76_8512;
   wire n_257_76_8513;
   wire n_257_76_8514;
   wire n_257_76_8515;
   wire n_257_76_8516;
   wire n_257_76_8517;
   wire n_257_76_8518;
   wire n_257_76_8519;
   wire n_257_76_8520;
   wire n_257_76_8521;
   wire n_257_76_8522;
   wire n_257_76_8523;
   wire n_257_76_8524;
   wire n_257_76_8525;
   wire n_257_76_8526;
   wire n_257_76_8527;
   wire n_257_76_8528;
   wire n_257_76_8529;
   wire n_257_76_8530;
   wire n_257_76_8531;
   wire n_257_76_8532;
   wire n_257_76_8533;
   wire n_257_76_8534;
   wire n_257_76_8535;
   wire n_257_76_8536;
   wire n_257_76_8537;
   wire n_257_76_8538;
   wire n_257_76_8539;
   wire n_257_76_8540;
   wire n_257_76_8541;
   wire n_257_76_8542;
   wire n_257_76_8543;
   wire n_257_76_8544;
   wire n_257_76_8545;
   wire n_257_76_8546;
   wire n_257_76_8547;
   wire n_257_76_8548;
   wire n_257_76_8549;
   wire n_257_76_8550;
   wire n_257_76_8551;
   wire n_257_76_8552;
   wire n_257_76_8553;
   wire n_257_76_8554;
   wire n_257_76_8555;
   wire n_257_76_8556;
   wire n_257_76_8557;
   wire n_257_76_8558;
   wire n_257_76_8559;
   wire n_257_76_8560;
   wire n_257_76_8561;
   wire n_257_76_8562;
   wire n_257_76_8563;
   wire n_257_76_8564;
   wire n_257_76_8565;
   wire n_257_76_8566;
   wire n_257_76_8567;
   wire n_257_76_8568;
   wire n_257_76_8569;
   wire n_257_76_8570;
   wire n_257_76_8571;
   wire n_257_76_8572;
   wire n_257_76_8573;
   wire n_257_76_8574;
   wire n_257_76_8575;
   wire n_257_76_8576;
   wire n_257_76_8577;
   wire n_257_76_8578;
   wire n_257_76_8579;
   wire n_257_76_8580;
   wire n_257_76_8581;
   wire n_257_76_8582;
   wire n_257_76_8583;
   wire n_257_76_8584;
   wire n_257_76_8585;
   wire n_257_76_8586;
   wire n_257_76_8587;
   wire n_257_76_8588;
   wire n_257_76_8589;
   wire n_257_76_8590;
   wire n_257_76_8591;
   wire n_257_76_8592;
   wire n_257_76_8593;
   wire n_257_76_8594;
   wire n_257_76_8595;
   wire n_257_76_8596;
   wire n_257_76_8597;
   wire n_257_76_8598;
   wire n_257_76_8599;
   wire n_257_76_8600;
   wire n_257_76_8601;
   wire n_257_76_8602;
   wire n_257_76_8603;
   wire n_257_76_8604;
   wire n_257_76_8605;
   wire n_257_76_8606;
   wire n_257_76_8607;
   wire n_257_76_8608;
   wire n_257_76_8609;
   wire n_257_76_8610;
   wire n_257_76_8611;
   wire n_257_76_8612;
   wire n_257_76_8613;
   wire n_257_76_8614;
   wire n_257_76_8615;
   wire n_257_76_8616;
   wire n_257_76_8617;
   wire n_257_76_8618;
   wire n_257_76_8619;
   wire n_257_76_8620;
   wire n_257_76_8621;
   wire n_257_76_8622;
   wire n_257_76_8623;
   wire n_257_76_8624;
   wire n_257_76_8625;
   wire n_257_76_8626;
   wire n_257_76_8627;
   wire n_257_76_8628;
   wire n_257_76_8629;
   wire n_257_76_8630;
   wire n_257_76_8631;
   wire n_257_76_8632;
   wire n_257_76_8633;
   wire n_257_76_8634;
   wire n_257_76_8635;
   wire n_257_76_8636;
   wire n_257_76_8637;
   wire n_257_76_8638;
   wire n_257_76_8639;
   wire n_257_76_8640;
   wire n_257_76_8641;
   wire n_257_76_8642;
   wire n_257_76_8643;
   wire n_257_76_8644;
   wire n_257_76_8645;
   wire n_257_76_8646;
   wire n_257_76_8647;
   wire n_257_76_8648;
   wire n_257_76_8649;
   wire n_257_76_8650;
   wire n_257_76_8651;
   wire n_257_76_8652;
   wire n_257_76_8653;
   wire n_257_76_8654;
   wire n_257_76_8655;
   wire n_257_76_8656;
   wire n_257_76_8657;
   wire n_257_76_8658;
   wire n_257_76_8659;
   wire n_257_76_8660;
   wire n_257_76_8661;
   wire n_257_76_8662;
   wire n_257_76_8663;
   wire n_257_76_8664;
   wire n_257_76_8665;
   wire n_257_76_8666;
   wire n_257_76_8667;
   wire n_257_76_8668;
   wire n_257_76_8669;
   wire n_257_76_8670;
   wire n_257_76_8671;
   wire n_257_76_8672;
   wire n_257_76_8673;
   wire n_257_76_8674;
   wire n_257_76_8675;
   wire n_257_76_8676;
   wire n_257_76_8677;
   wire n_257_76_8678;
   wire n_257_76_8679;
   wire n_257_76_8680;
   wire n_257_76_8681;
   wire n_257_76_8682;
   wire n_257_76_8683;
   wire n_257_76_8684;
   wire n_257_76_8685;
   wire n_257_76_8686;
   wire n_257_76_8687;
   wire n_257_76_8688;
   wire n_257_76_8689;
   wire n_257_76_8690;
   wire n_257_76_8691;
   wire n_257_76_8692;
   wire n_257_76_8693;
   wire n_257_76_8694;
   wire n_257_76_8695;
   wire n_257_76_8696;
   wire n_257_76_8697;
   wire n_257_76_8698;
   wire n_257_76_8699;
   wire n_257_76_8700;
   wire n_257_76_8701;
   wire n_257_76_8702;
   wire n_257_76_8703;
   wire n_257_76_8704;
   wire n_257_76_8705;
   wire n_257_76_8706;
   wire n_257_76_8707;
   wire n_257_76_8708;
   wire n_257_76_8709;
   wire n_257_76_8710;
   wire n_257_76_8711;
   wire n_257_76_8712;
   wire n_257_76_8713;
   wire n_257_76_8714;
   wire n_257_76_8715;
   wire n_257_76_8716;
   wire n_257_76_8717;
   wire n_257_76_8718;
   wire n_257_76_8719;
   wire n_257_76_8720;
   wire n_257_76_8721;
   wire n_257_76_8722;
   wire n_257_76_8723;
   wire n_257_76_8724;
   wire n_257_76_8725;
   wire n_257_76_8726;
   wire n_257_76_8727;
   wire n_257_76_8728;
   wire n_257_76_8729;
   wire n_257_76_8730;
   wire n_257_76_8731;
   wire n_257_76_8732;
   wire n_257_76_8733;
   wire n_257_76_8734;
   wire n_257_76_8735;
   wire n_257_76_8736;
   wire n_257_76_8737;
   wire n_257_76_8738;
   wire n_257_76_8739;
   wire n_257_76_8740;
   wire n_257_76_8741;
   wire n_257_76_8742;
   wire n_257_76_8743;
   wire n_257_76_8744;
   wire n_257_76_8745;
   wire n_257_76_8746;
   wire n_257_76_8747;
   wire n_257_76_8748;
   wire n_257_76_8749;
   wire n_257_76_8750;
   wire n_257_76_8751;
   wire n_257_76_8752;
   wire n_257_76_8753;
   wire n_257_76_8754;
   wire n_257_76_8755;
   wire n_257_76_8756;
   wire n_257_76_8757;
   wire n_257_76_8758;
   wire n_257_76_8759;
   wire n_257_76_8760;
   wire n_257_76_8761;
   wire n_257_76_8762;
   wire n_257_76_8763;
   wire n_257_76_8764;
   wire n_257_76_8765;
   wire n_257_76_8766;
   wire n_257_76_8767;
   wire n_257_76_8768;
   wire n_257_76_8769;
   wire n_257_76_8770;
   wire n_257_76_8771;
   wire n_257_76_8772;
   wire n_257_76_8773;
   wire n_257_76_8774;
   wire n_257_76_8775;
   wire n_257_76_8776;
   wire n_257_76_8777;
   wire n_257_76_8778;
   wire n_257_76_8779;
   wire n_257_76_8780;
   wire n_257_76_8781;
   wire n_257_76_8782;
   wire n_257_76_8783;
   wire n_257_76_8784;
   wire n_257_76_8785;
   wire n_257_76_8786;
   wire n_257_76_8787;
   wire n_257_76_8788;
   wire n_257_76_8789;
   wire n_257_76_8790;
   wire n_257_76_8791;
   wire n_257_76_8792;
   wire n_257_76_8793;
   wire n_257_76_8794;
   wire n_257_76_8795;
   wire n_257_76_8796;
   wire n_257_76_8797;
   wire n_257_76_8798;
   wire n_257_76_8799;
   wire n_257_76_8800;
   wire n_257_76_8801;
   wire n_257_76_8802;
   wire n_257_76_8803;
   wire n_257_76_8804;
   wire n_257_76_8805;
   wire n_257_76_8806;
   wire n_257_76_8807;
   wire n_257_76_8808;
   wire n_257_76_8809;
   wire n_257_76_8810;
   wire n_257_76_8811;
   wire n_257_76_8812;
   wire n_257_76_8813;
   wire n_257_76_8814;
   wire n_257_76_8815;
   wire n_257_76_8816;
   wire n_257_76_8817;
   wire n_257_76_8818;
   wire n_257_76_8819;
   wire n_257_76_8820;
   wire n_257_76_8821;
   wire n_257_76_8822;
   wire n_257_76_8823;
   wire n_257_76_8824;
   wire n_257_76_8825;
   wire n_257_76_8826;
   wire n_257_76_8827;
   wire n_257_76_8828;
   wire n_257_76_8829;
   wire n_257_76_8830;
   wire n_257_76_8831;
   wire n_257_76_8832;
   wire n_257_76_8833;
   wire n_257_76_8834;
   wire n_257_76_8835;
   wire n_257_76_8836;
   wire n_257_76_8837;
   wire n_257_76_8838;
   wire n_257_76_8839;
   wire n_257_76_8840;
   wire n_257_76_8841;
   wire n_257_76_8842;
   wire n_257_76_8843;
   wire n_257_76_8844;
   wire n_257_76_8845;
   wire n_257_76_8846;
   wire n_257_76_8847;
   wire n_257_76_8848;
   wire n_257_76_8849;
   wire n_257_76_8850;
   wire n_257_76_8851;
   wire n_257_76_8852;
   wire n_257_76_8853;
   wire n_257_76_8854;
   wire n_257_76_8855;
   wire n_257_76_8856;
   wire n_257_76_8857;
   wire n_257_76_8858;
   wire n_257_76_8859;
   wire n_257_76_8860;
   wire n_257_76_8861;
   wire n_257_76_8862;
   wire n_257_76_8863;
   wire n_257_76_8864;
   wire n_257_76_8865;
   wire n_257_76_8866;
   wire n_257_76_8867;
   wire n_257_76_8868;
   wire n_257_76_8869;
   wire n_257_76_8870;
   wire n_257_76_8871;
   wire n_257_76_8872;
   wire n_257_76_8873;
   wire n_257_76_8874;
   wire n_257_76_8875;
   wire n_257_76_8876;
   wire n_257_76_8877;
   wire n_257_76_8878;
   wire n_257_76_8879;
   wire n_257_76_8880;
   wire n_257_76_8881;
   wire n_257_76_8882;
   wire n_257_76_8883;
   wire n_257_76_8884;
   wire n_257_76_8885;
   wire n_257_76_8886;
   wire n_257_76_8887;
   wire n_257_76_8888;
   wire n_257_76_8889;
   wire n_257_76_8890;
   wire n_257_76_8891;
   wire n_257_76_8892;
   wire n_257_76_8893;
   wire n_257_76_8894;
   wire n_257_76_8895;
   wire n_257_76_8896;
   wire n_257_76_8897;
   wire n_257_76_8898;
   wire n_257_76_8899;
   wire n_257_76_8900;
   wire n_257_76_8901;
   wire n_257_76_8902;
   wire n_257_76_8903;
   wire n_257_76_8904;
   wire n_257_76_8905;
   wire n_257_76_8906;
   wire n_257_76_8907;
   wire n_257_76_8908;
   wire n_257_76_8909;
   wire n_257_76_8910;
   wire n_257_76_8911;
   wire n_257_76_8912;
   wire n_257_76_8913;
   wire n_257_76_8914;
   wire n_257_76_8915;
   wire n_257_76_8916;
   wire n_257_76_8917;
   wire n_257_76_8918;
   wire n_257_76_8919;
   wire n_257_76_8920;
   wire n_257_76_8921;
   wire n_257_76_8922;
   wire n_257_76_8923;
   wire n_257_76_8924;
   wire n_257_76_8925;
   wire n_257_76_8926;
   wire n_257_76_8927;
   wire n_257_76_8928;
   wire n_257_76_8929;
   wire n_257_76_8930;
   wire n_257_76_8931;
   wire n_257_76_8932;
   wire n_257_76_8933;
   wire n_257_76_8934;
   wire n_257_76_8935;
   wire n_257_76_8936;
   wire n_257_76_8937;
   wire n_257_76_8938;
   wire n_257_76_8939;
   wire n_257_76_8940;
   wire n_257_76_8941;
   wire n_257_76_8942;
   wire n_257_76_8943;
   wire n_257_76_8944;
   wire n_257_76_8945;
   wire n_257_76_8946;
   wire n_257_76_8947;
   wire n_257_76_8948;
   wire n_257_76_8949;
   wire n_257_76_8950;
   wire n_257_76_8951;
   wire n_257_76_8952;
   wire n_257_76_8953;
   wire n_257_76_8954;
   wire n_257_76_8955;
   wire n_257_76_8956;
   wire n_257_76_8957;
   wire n_257_76_8958;
   wire n_257_76_8959;
   wire n_257_76_8960;
   wire n_257_76_8961;
   wire n_257_76_8962;
   wire n_257_76_8963;
   wire n_257_76_8964;
   wire n_257_76_8965;
   wire n_257_76_8966;
   wire n_257_76_8967;
   wire n_257_76_8968;
   wire n_257_76_8969;
   wire n_257_76_8970;
   wire n_257_76_8971;
   wire n_257_76_8972;
   wire n_257_76_8973;
   wire n_257_76_8974;
   wire n_257_76_8975;
   wire n_257_76_8976;
   wire n_257_76_8977;
   wire n_257_76_8978;
   wire n_257_76_8979;
   wire n_257_76_8980;
   wire n_257_76_8981;
   wire n_257_76_8982;
   wire n_257_76_8983;
   wire n_257_76_8984;
   wire n_257_76_8985;
   wire n_257_76_8986;
   wire n_257_76_8987;
   wire n_257_76_8988;
   wire n_257_76_8989;
   wire n_257_76_8990;
   wire n_257_76_8991;
   wire n_257_76_8992;
   wire n_257_76_8993;
   wire n_257_76_8994;
   wire n_257_76_8995;
   wire n_257_76_8996;
   wire n_257_76_8997;
   wire n_257_76_8998;
   wire n_257_76_8999;
   wire n_257_76_9000;
   wire n_257_76_9001;
   wire n_257_76_9002;
   wire n_257_76_9003;
   wire n_257_76_9004;
   wire n_257_76_9005;
   wire n_257_76_9006;
   wire n_257_76_9007;
   wire n_257_76_9008;
   wire n_257_76_9009;
   wire n_257_76_9010;
   wire n_257_76_9011;
   wire n_257_76_9012;
   wire n_257_76_9013;
   wire n_257_76_9014;
   wire n_257_76_9015;
   wire n_257_76_9016;
   wire n_257_76_9017;
   wire n_257_76_9018;
   wire n_257_76_9019;
   wire n_257_76_9020;
   wire n_257_76_9021;
   wire n_257_76_9022;
   wire n_257_76_9023;
   wire n_257_76_9024;
   wire n_257_76_9025;
   wire n_257_76_9026;
   wire n_257_76_9027;
   wire n_257_76_9028;
   wire n_257_76_9029;
   wire n_257_76_9030;
   wire n_257_76_9031;
   wire n_257_76_9032;
   wire n_257_76_9033;
   wire n_257_76_9034;
   wire n_257_76_9035;
   wire n_257_76_9036;
   wire n_257_76_9037;
   wire n_257_76_9038;
   wire n_257_76_9039;
   wire n_257_76_9040;
   wire n_257_76_9041;
   wire n_257_76_9042;
   wire n_257_76_9043;
   wire n_257_76_9044;
   wire n_257_76_9045;
   wire n_257_76_9046;
   wire n_257_76_9047;
   wire n_257_76_9048;
   wire n_257_76_9049;
   wire n_257_76_9050;
   wire n_257_76_9051;
   wire n_257_76_9052;
   wire n_257_76_9053;
   wire n_257_76_9054;
   wire n_257_76_9055;
   wire n_257_76_9056;
   wire n_257_76_9057;
   wire n_257_76_9058;
   wire n_257_76_9059;
   wire n_257_76_9060;
   wire n_257_76_9061;
   wire n_257_76_9062;
   wire n_257_76_9063;
   wire n_257_76_9064;
   wire n_257_76_9065;
   wire n_257_76_9066;
   wire n_257_76_9067;
   wire n_257_76_9068;
   wire n_257_76_9069;
   wire n_257_76_9070;
   wire n_257_76_9071;
   wire n_257_76_9072;
   wire n_257_76_9073;
   wire n_257_76_9074;
   wire n_257_76_9075;
   wire n_257_76_9076;
   wire n_257_76_9077;
   wire n_257_76_9078;
   wire n_257_76_9079;
   wire n_257_76_9080;
   wire n_257_76_9081;
   wire n_257_76_9082;
   wire n_257_76_9083;
   wire n_257_76_9084;
   wire n_257_76_9085;
   wire n_257_76_9086;
   wire n_257_76_9087;
   wire n_257_76_9088;
   wire n_257_76_9089;
   wire n_257_76_9090;
   wire n_257_76_9091;
   wire n_257_76_9092;
   wire n_257_76_9093;
   wire n_257_76_9094;
   wire n_257_76_9095;
   wire n_257_76_9096;
   wire n_257_76_9097;
   wire n_257_76_9098;
   wire n_257_76_9099;
   wire n_257_76_9100;
   wire n_257_76_9101;
   wire n_257_76_9102;
   wire n_257_76_9103;
   wire n_257_76_9104;
   wire n_257_76_9105;
   wire n_257_76_9106;
   wire n_257_76_9107;
   wire n_257_76_9108;
   wire n_257_76_9109;
   wire n_257_76_9110;
   wire n_257_76_9111;
   wire n_257_76_9112;
   wire n_257_76_9113;
   wire n_257_76_9114;
   wire n_257_76_9115;
   wire n_257_76_9116;
   wire n_257_76_9117;
   wire n_257_76_9118;
   wire n_257_76_9119;
   wire n_257_76_9120;
   wire n_257_76_9121;
   wire n_257_76_9122;
   wire n_257_76_9123;
   wire n_257_76_9124;
   wire n_257_76_9125;
   wire n_257_76_9126;
   wire n_257_76_9127;
   wire n_257_76_9128;
   wire n_257_76_9129;
   wire n_257_76_9130;
   wire n_257_76_9131;
   wire n_257_76_9132;
   wire n_257_76_9133;
   wire n_257_76_9134;
   wire n_257_76_9135;
   wire n_257_76_9136;
   wire n_257_76_9137;
   wire n_257_76_9138;
   wire n_257_76_9139;
   wire n_257_76_9140;
   wire n_257_76_9141;
   wire n_257_76_9142;
   wire n_257_76_9143;
   wire n_257_76_9144;
   wire n_257_76_9145;
   wire n_257_76_9146;
   wire n_257_76_9147;
   wire n_257_76_9148;
   wire n_257_76_9149;
   wire n_257_76_9150;
   wire n_257_76_9151;
   wire n_257_76_9152;
   wire n_257_76_9153;
   wire n_257_76_9154;
   wire n_257_76_9155;
   wire n_257_76_9156;
   wire n_257_76_9157;
   wire n_257_76_9158;
   wire n_257_76_9159;
   wire n_257_76_9160;
   wire n_257_76_9161;
   wire n_257_76_9162;
   wire n_257_76_9163;
   wire n_257_76_9164;
   wire n_257_76_9165;
   wire n_257_76_9166;
   wire n_257_76_9167;
   wire n_257_76_9168;
   wire n_257_76_9169;
   wire n_257_76_9170;
   wire n_257_76_9171;
   wire n_257_76_9172;
   wire n_257_76_9173;
   wire n_257_76_9174;
   wire n_257_76_9175;
   wire n_257_76_9176;
   wire n_257_76_9177;
   wire n_257_76_9178;
   wire n_257_76_9179;
   wire n_257_76_9180;
   wire n_257_76_9181;
   wire n_257_76_9182;
   wire n_257_76_9183;
   wire n_257_76_9184;
   wire n_257_76_9185;
   wire n_257_76_9186;
   wire n_257_76_9187;
   wire n_257_76_9188;
   wire n_257_76_9189;
   wire n_257_76_9190;
   wire n_257_76_9191;
   wire n_257_76_9192;
   wire n_257_76_9193;
   wire n_257_76_9194;
   wire n_257_76_9195;
   wire n_257_76_9196;
   wire n_257_76_9197;
   wire n_257_76_9198;
   wire n_257_76_9199;
   wire n_257_76_9200;
   wire n_257_76_9201;
   wire n_257_76_9202;
   wire n_257_76_9203;
   wire n_257_76_9204;
   wire n_257_76_9205;
   wire n_257_76_9206;
   wire n_257_76_9207;
   wire n_257_76_9208;
   wire n_257_76_9209;
   wire n_257_76_9210;
   wire n_257_76_9211;
   wire n_257_76_9212;
   wire n_257_76_9213;
   wire n_257_76_9214;
   wire n_257_76_9215;
   wire n_257_76_9216;
   wire n_257_76_9217;
   wire n_257_76_9218;
   wire n_257_76_9219;
   wire n_257_76_9220;
   wire n_257_76_9221;
   wire n_257_76_9222;
   wire n_257_76_9223;
   wire n_257_76_9224;
   wire n_257_76_9225;
   wire n_257_76_9226;
   wire n_257_76_9227;
   wire n_257_76_9228;
   wire n_257_76_9229;
   wire n_257_76_9230;
   wire n_257_76_9231;
   wire n_257_76_9232;
   wire n_257_76_9233;
   wire n_257_76_9234;
   wire n_257_76_9235;
   wire n_257_76_9236;
   wire n_257_76_9237;
   wire n_257_76_9238;
   wire n_257_76_9239;
   wire n_257_76_9240;
   wire n_257_76_9241;
   wire n_257_76_9242;
   wire n_257_76_9243;
   wire n_257_76_9244;
   wire n_257_76_9245;
   wire n_257_76_9246;
   wire n_257_76_9247;
   wire n_257_76_9248;
   wire n_257_76_9249;
   wire n_257_76_9250;
   wire n_257_76_9251;
   wire n_257_76_9252;
   wire n_257_76_9253;
   wire n_257_76_9254;
   wire n_257_76_9255;
   wire n_257_76_9256;
   wire n_257_76_9257;
   wire n_257_76_9258;
   wire n_257_76_9259;
   wire n_257_76_9260;
   wire n_257_76_9261;
   wire n_257_76_9262;
   wire n_257_76_9263;
   wire n_257_76_9264;
   wire n_257_76_9265;
   wire n_257_76_9266;
   wire n_257_76_9267;
   wire n_257_76_9268;
   wire n_257_76_9269;
   wire n_257_76_9270;
   wire n_257_76_9271;
   wire n_257_76_9272;
   wire n_257_76_9273;
   wire n_257_76_9274;
   wire n_257_76_9275;
   wire n_257_76_9276;
   wire n_257_76_9277;
   wire n_257_76_9278;
   wire n_257_76_9279;
   wire n_257_76_9280;
   wire n_257_76_9281;
   wire n_257_76_9282;
   wire n_257_76_9283;
   wire n_257_76_9284;
   wire n_257_76_9285;
   wire n_257_76_9286;
   wire n_257_76_9287;
   wire n_257_76_9288;
   wire n_257_76_9289;
   wire n_257_76_9290;
   wire n_257_76_9291;
   wire n_257_76_9292;
   wire n_257_76_9293;
   wire n_257_76_9294;
   wire n_257_76_9295;
   wire n_257_76_9296;
   wire n_257_76_9297;
   wire n_257_76_9298;
   wire n_257_76_9299;
   wire n_257_76_9300;
   wire n_257_76_9301;
   wire n_257_76_9302;
   wire n_257_76_9303;
   wire n_257_76_9304;
   wire n_257_76_9305;
   wire n_257_76_9306;
   wire n_257_76_9307;
   wire n_257_76_9308;
   wire n_257_76_9309;
   wire n_257_76_9310;
   wire n_257_76_9311;
   wire n_257_76_9312;
   wire n_257_76_9313;
   wire n_257_76_9314;
   wire n_257_76_9315;
   wire n_257_76_9316;
   wire n_257_76_9317;
   wire n_257_76_9318;
   wire n_257_76_9319;
   wire n_257_76_9320;
   wire n_257_76_9321;
   wire n_257_76_9322;
   wire n_257_76_9323;
   wire n_257_76_9324;
   wire n_257_76_9325;
   wire n_257_76_9326;
   wire n_257_76_9327;
   wire n_257_76_9328;
   wire n_257_76_9329;
   wire n_257_76_9330;
   wire n_257_76_9331;
   wire n_257_76_9332;
   wire n_257_76_9333;
   wire n_257_76_9334;
   wire n_257_76_9335;
   wire n_257_76_9336;
   wire n_257_76_9337;
   wire n_257_76_9338;
   wire n_257_76_9339;
   wire n_257_76_9340;
   wire n_257_76_9341;
   wire n_257_76_9342;
   wire n_257_76_9343;
   wire n_257_76_9344;
   wire n_257_76_9345;
   wire n_257_76_9346;
   wire n_257_76_9347;
   wire n_257_76_9348;
   wire n_257_76_9349;
   wire n_257_76_9350;
   wire n_257_76_9351;
   wire n_257_76_9352;
   wire n_257_76_9353;
   wire n_257_76_9354;
   wire n_257_76_9355;
   wire n_257_76_9356;
   wire n_257_76_9357;
   wire n_257_76_9358;
   wire n_257_76_9359;
   wire n_257_76_9360;
   wire n_257_76_9361;
   wire n_257_76_9362;
   wire n_257_76_9363;
   wire n_257_76_9364;
   wire n_257_76_9365;
   wire n_257_76_9366;
   wire n_257_76_9367;
   wire n_257_76_9368;
   wire n_257_76_9369;
   wire n_257_76_9370;
   wire n_257_76_9371;
   wire n_257_76_9372;
   wire n_257_76_9373;
   wire n_257_76_9374;
   wire n_257_76_9375;
   wire n_257_76_9376;
   wire n_257_76_9377;
   wire n_257_76_9378;
   wire n_257_76_9379;
   wire n_257_76_9380;
   wire n_257_76_9381;
   wire n_257_76_9382;
   wire n_257_76_9383;
   wire n_257_76_9384;
   wire n_257_76_9385;
   wire n_257_76_9386;
   wire n_257_76_9387;
   wire n_257_76_9388;
   wire n_257_76_9389;
   wire n_257_76_9390;
   wire n_257_76_9391;
   wire n_257_76_9392;
   wire n_257_76_9393;
   wire n_257_76_9394;
   wire n_257_76_9395;
   wire n_257_76_9396;
   wire n_257_76_9397;
   wire n_257_76_9398;
   wire n_257_76_9399;
   wire n_257_76_9400;
   wire n_257_76_9401;
   wire n_257_76_9402;
   wire n_257_76_9403;
   wire n_257_76_9404;
   wire n_257_76_9405;
   wire n_257_76_9406;
   wire n_257_76_9407;
   wire n_257_76_9408;
   wire n_257_76_9409;
   wire n_257_76_9410;
   wire n_257_76_9411;
   wire n_257_76_9412;
   wire n_257_76_9413;
   wire n_257_76_9414;
   wire n_257_76_9415;
   wire n_257_76_9416;
   wire n_257_76_9417;
   wire n_257_76_9418;
   wire n_257_76_9419;
   wire n_257_76_9420;
   wire n_257_76_9421;
   wire n_257_76_9422;
   wire n_257_76_9423;
   wire n_257_76_9424;
   wire n_257_76_9425;
   wire n_257_76_9426;
   wire n_257_76_9427;
   wire n_257_76_9428;
   wire n_257_76_9429;
   wire n_257_76_9430;
   wire n_257_76_9431;
   wire n_257_76_9432;
   wire n_257_76_9433;
   wire n_257_76_9434;
   wire n_257_76_9435;
   wire n_257_76_9436;
   wire n_257_76_9437;
   wire n_257_76_9438;
   wire n_257_76_9439;
   wire n_257_76_9440;
   wire n_257_76_9441;
   wire n_257_76_9442;
   wire n_257_76_9443;
   wire n_257_76_9444;
   wire n_257_76_9445;
   wire n_257_76_9446;
   wire n_257_76_9447;
   wire n_257_76_9448;
   wire n_257_76_9449;
   wire n_257_76_9450;
   wire n_257_76_9451;
   wire n_257_76_9452;
   wire n_257_76_9453;
   wire n_257_76_9454;
   wire n_257_76_9455;
   wire n_257_76_9456;
   wire n_257_76_9457;
   wire n_257_76_9458;
   wire n_257_76_9459;
   wire n_257_76_9460;
   wire n_257_76_9461;
   wire n_257_76_9462;
   wire n_257_76_9463;
   wire n_257_76_9464;
   wire n_257_76_9465;
   wire n_257_76_9466;
   wire n_257_76_9467;
   wire n_257_76_9468;
   wire n_257_76_9469;
   wire n_257_76_9470;
   wire n_257_76_9471;
   wire n_257_76_9472;
   wire n_257_76_9473;
   wire n_257_76_9474;
   wire n_257_76_9475;
   wire n_257_76_9476;
   wire n_257_76_9477;
   wire n_257_76_9478;
   wire n_257_76_9479;
   wire n_257_76_9480;
   wire n_257_76_9481;
   wire n_257_76_9482;
   wire n_257_76_9483;
   wire n_257_76_9484;
   wire n_257_76_9485;
   wire n_257_76_9486;
   wire n_257_76_9487;
   wire n_257_76_9488;
   wire n_257_76_9489;
   wire n_257_76_9490;
   wire n_257_76_9491;
   wire n_257_76_9492;
   wire n_257_76_9493;
   wire n_257_76_9494;
   wire n_257_76_9495;
   wire n_257_76_9496;
   wire n_257_76_9497;
   wire n_257_76_9498;
   wire n_257_76_9499;
   wire n_257_76_9500;
   wire n_257_76_9501;
   wire n_257_76_9502;
   wire n_257_76_9503;
   wire n_257_76_9504;
   wire n_257_76_9505;
   wire n_257_76_9506;
   wire n_257_76_9507;
   wire n_257_76_9508;
   wire n_257_76_9509;
   wire n_257_76_9510;
   wire n_257_76_9511;
   wire n_257_76_9512;
   wire n_257_76_9513;
   wire n_257_76_9514;
   wire n_257_76_9515;
   wire n_257_76_9516;
   wire n_257_76_9517;
   wire n_257_76_9518;
   wire n_257_76_9519;
   wire n_257_76_9520;
   wire n_257_76_9521;
   wire n_257_76_9522;
   wire n_257_76_9523;
   wire n_257_76_9524;
   wire n_257_76_9525;
   wire n_257_76_9526;
   wire n_257_76_9527;
   wire n_257_76_9528;
   wire n_257_76_9529;
   wire n_257_76_9530;
   wire n_257_76_9531;
   wire n_257_76_9532;
   wire n_257_76_9533;
   wire n_257_76_9534;
   wire n_257_76_9535;
   wire n_257_76_9536;
   wire n_257_76_9537;
   wire n_257_76_9538;
   wire n_257_76_9539;
   wire n_257_76_9540;
   wire n_257_76_9541;
   wire n_257_76_9542;
   wire n_257_76_9543;
   wire n_257_76_9544;
   wire n_257_76_9545;
   wire n_257_76_9546;
   wire n_257_76_9547;
   wire n_257_76_9548;
   wire n_257_76_9549;
   wire n_257_76_9550;
   wire n_257_76_9551;
   wire n_257_76_9552;
   wire n_257_76_9553;
   wire n_257_76_9554;
   wire n_257_76_9555;
   wire n_257_76_9556;
   wire n_257_76_9557;
   wire n_257_76_9558;
   wire n_257_76_9559;
   wire n_257_76_9560;
   wire n_257_76_9561;
   wire n_257_76_9562;
   wire n_257_76_9563;
   wire n_257_76_9564;
   wire n_257_76_9565;
   wire n_257_76_9566;
   wire n_257_76_9567;
   wire n_257_76_9568;
   wire n_257_76_9569;
   wire n_257_76_9570;
   wire n_257_76_9571;
   wire n_257_76_9572;
   wire n_257_76_9573;
   wire n_257_76_9574;
   wire n_257_76_9575;
   wire n_257_76_9576;
   wire n_257_76_9577;
   wire n_257_76_9578;
   wire n_257_76_9579;
   wire n_257_76_9580;
   wire n_257_76_9581;
   wire n_257_76_9582;
   wire n_257_76_9583;
   wire n_257_76_9584;
   wire n_257_76_9585;
   wire n_257_76_9586;
   wire n_257_76_9587;
   wire n_257_76_9588;
   wire n_257_76_9589;
   wire n_257_76_9590;
   wire n_257_76_9591;
   wire n_257_76_9592;
   wire n_257_76_9593;
   wire n_257_76_9594;
   wire n_257_76_9595;
   wire n_257_76_9596;
   wire n_257_76_9597;
   wire n_257_76_9598;
   wire n_257_76_9599;
   wire n_257_76_9600;
   wire n_257_76_9601;
   wire n_257_76_9602;
   wire n_257_76_9603;
   wire n_257_76_9604;
   wire n_257_76_9605;
   wire n_257_76_9606;
   wire n_257_76_9607;
   wire n_257_76_9608;
   wire n_257_76_9609;
   wire n_257_76_9610;
   wire n_257_76_9611;
   wire n_257_76_9612;
   wire n_257_76_9613;
   wire n_257_76_9614;
   wire n_257_76_9615;
   wire n_257_76_9616;
   wire n_257_76_9617;
   wire n_257_76_9618;
   wire n_257_76_9619;
   wire n_257_76_9620;
   wire n_257_76_9621;
   wire n_257_76_9622;
   wire n_257_76_9623;
   wire n_257_76_9624;
   wire n_257_76_9625;
   wire n_257_76_9626;
   wire n_257_76_9627;
   wire n_257_76_9628;
   wire n_257_76_9629;
   wire n_257_76_9630;
   wire n_257_76_9631;
   wire n_257_76_9632;
   wire n_257_76_9633;
   wire n_257_76_9634;
   wire n_257_76_9635;
   wire n_257_76_9636;
   wire n_257_76_9637;
   wire n_257_76_9638;
   wire n_257_76_9639;
   wire n_257_76_9640;
   wire n_257_76_9641;
   wire n_257_76_9642;
   wire n_257_76_9643;
   wire n_257_76_9644;
   wire n_257_76_9645;
   wire n_257_76_9646;
   wire n_257_76_9647;
   wire n_257_76_9648;
   wire n_257_76_9649;
   wire n_257_76_9650;
   wire n_257_76_9651;
   wire n_257_76_9652;
   wire n_257_76_9653;
   wire n_257_76_9654;
   wire n_257_76_9655;
   wire n_257_76_9656;
   wire n_257_76_9657;
   wire n_257_76_9658;
   wire n_257_76_9659;
   wire n_257_76_9660;
   wire n_257_76_9661;
   wire n_257_76_9662;
   wire n_257_76_9663;
   wire n_257_76_9664;
   wire n_257_76_9665;
   wire n_257_76_9666;
   wire n_257_76_9667;
   wire n_257_76_9668;
   wire n_257_76_9669;
   wire n_257_76_9670;
   wire n_257_76_9671;
   wire n_257_76_9672;
   wire n_257_76_9673;
   wire n_257_76_9674;
   wire n_257_76_9675;
   wire n_257_76_9676;
   wire n_257_76_9677;
   wire n_257_76_9678;
   wire n_257_76_9679;
   wire n_257_76_9680;
   wire n_257_76_9681;
   wire n_257_76_9682;
   wire n_257_76_9683;
   wire n_257_76_9684;
   wire n_257_76_9685;
   wire n_257_76_9686;
   wire n_257_76_9687;
   wire n_257_76_9688;
   wire n_257_76_9689;
   wire n_257_76_9690;
   wire n_257_76_9691;
   wire n_257_76_9692;
   wire n_257_76_9693;
   wire n_257_76_9694;
   wire n_257_76_9695;
   wire n_257_76_9696;
   wire n_257_76_9697;
   wire n_257_76_9698;
   wire n_257_76_9699;
   wire n_257_76_9700;
   wire n_257_76_9701;
   wire n_257_76_9702;
   wire n_257_76_9703;
   wire n_257_76_9704;
   wire n_257_76_9705;
   wire n_257_76_9706;
   wire n_257_76_9707;
   wire n_257_76_9708;
   wire n_257_76_9709;
   wire n_257_76_9710;
   wire n_257_76_9711;
   wire n_257_76_9712;
   wire n_257_76_9713;
   wire n_257_76_9714;
   wire n_257_76_9715;
   wire n_257_76_9716;
   wire n_257_76_9717;
   wire n_257_76_9718;
   wire n_257_76_9719;
   wire n_257_76_9720;
   wire n_257_76_9721;
   wire n_257_76_9722;
   wire n_257_76_9723;
   wire n_257_76_9724;
   wire n_257_76_9725;
   wire n_257_76_9726;
   wire n_257_76_9727;
   wire n_257_76_9728;
   wire n_257_76_9729;
   wire n_257_76_9730;
   wire n_257_76_9731;
   wire n_257_76_9732;
   wire n_257_76_9733;
   wire n_257_76_9734;
   wire n_257_76_9735;
   wire n_257_76_9736;
   wire n_257_76_9737;
   wire n_257_76_9738;
   wire n_257_76_9739;
   wire n_257_76_9740;
   wire n_257_76_9741;
   wire n_257_76_9742;
   wire n_257_76_9743;
   wire n_257_76_9744;
   wire n_257_76_9745;
   wire n_257_76_9746;
   wire n_257_76_9747;
   wire n_257_76_9748;
   wire n_257_76_9749;
   wire n_257_76_9750;
   wire n_257_76_9751;
   wire n_257_76_9752;
   wire n_257_76_9753;
   wire n_257_76_9754;
   wire n_257_76_9755;
   wire n_257_76_9756;
   wire n_257_76_9757;
   wire n_257_76_9758;
   wire n_257_76_9759;
   wire n_257_76_9760;
   wire n_257_76_9761;
   wire n_257_76_9762;
   wire n_257_76_9763;
   wire n_257_76_9764;
   wire n_257_76_9765;
   wire n_257_76_9766;
   wire n_257_76_9767;
   wire n_257_76_9768;
   wire n_257_76_9769;
   wire n_257_76_9770;
   wire n_257_76_9771;
   wire n_257_76_9772;
   wire n_257_76_9773;
   wire n_257_76_9774;
   wire n_257_76_9775;
   wire n_257_76_9776;
   wire n_257_76_9777;
   wire n_257_76_9778;
   wire n_257_76_9779;
   wire n_257_76_9780;
   wire n_257_76_9781;
   wire n_257_76_9782;
   wire n_257_76_9783;
   wire n_257_76_9784;
   wire n_257_76_9785;
   wire n_257_76_9786;
   wire n_257_76_9787;
   wire n_257_76_9788;
   wire n_257_76_9789;
   wire n_257_76_9790;
   wire n_257_76_9791;
   wire n_257_76_9792;
   wire n_257_76_9793;
   wire n_257_76_9794;
   wire n_257_76_9795;
   wire n_257_76_9796;
   wire n_257_76_9797;
   wire n_257_76_9798;
   wire n_257_76_9799;
   wire n_257_76_9800;
   wire n_257_76_9801;
   wire n_257_76_9802;
   wire n_257_76_9803;
   wire n_257_76_9804;
   wire n_257_76_9805;
   wire n_257_76_9806;
   wire n_257_76_9807;
   wire n_257_76_9808;
   wire n_257_76_9809;
   wire n_257_76_9810;
   wire n_257_76_9811;
   wire n_257_76_9812;
   wire n_257_76_9813;
   wire n_257_76_9814;
   wire n_257_76_9815;
   wire n_257_76_9816;
   wire n_257_76_9817;
   wire n_257_76_9818;
   wire n_257_76_9819;
   wire n_257_76_9820;
   wire n_257_76_9821;
   wire n_257_76_9822;
   wire n_257_76_9823;
   wire n_257_76_9824;
   wire n_257_76_9825;
   wire n_257_76_9826;
   wire n_257_76_9827;
   wire n_257_76_9828;
   wire n_257_76_9829;
   wire n_257_76_9830;
   wire n_257_76_9831;
   wire n_257_76_9832;
   wire n_257_76_9833;
   wire n_257_76_9834;
   wire n_257_76_9835;
   wire n_257_76_9836;
   wire n_257_76_9837;
   wire n_257_76_9838;
   wire n_257_76_9839;
   wire n_257_76_9840;
   wire n_257_76_9841;
   wire n_257_76_9842;
   wire n_257_76_9843;
   wire n_257_76_9844;
   wire n_257_76_9845;
   wire n_257_76_9846;
   wire n_257_76_9847;
   wire n_257_76_9848;
   wire n_257_76_9849;
   wire n_257_76_9850;
   wire n_257_76_9851;
   wire n_257_76_9852;
   wire n_257_76_9853;
   wire n_257_76_9854;
   wire n_257_76_9855;
   wire n_257_76_9856;
   wire n_257_76_9857;
   wire n_257_76_9858;
   wire n_257_76_9859;
   wire n_257_76_9860;
   wire n_257_76_9861;
   wire n_257_76_9862;
   wire n_257_76_9863;
   wire n_257_76_9864;
   wire n_257_76_9865;
   wire n_257_76_9866;
   wire n_257_76_9867;
   wire n_257_76_9868;
   wire n_257_76_9869;
   wire n_257_76_9870;
   wire n_257_76_9871;
   wire n_257_76_9872;
   wire n_257_76_9873;
   wire n_257_76_9874;
   wire n_257_76_9875;
   wire n_257_76_9876;
   wire n_257_76_9877;
   wire n_257_76_9878;
   wire n_257_76_9879;
   wire n_257_76_9880;
   wire n_257_76_9881;
   wire n_257_76_9882;
   wire n_257_76_9883;
   wire n_257_76_9884;
   wire n_257_76_9885;
   wire n_257_76_9886;
   wire n_257_76_9887;
   wire n_257_76_9888;
   wire n_257_76_9889;
   wire n_257_76_9890;
   wire n_257_76_9891;
   wire n_257_76_9892;
   wire n_257_76_9893;
   wire n_257_76_9894;
   wire n_257_76_9895;
   wire n_257_76_9896;
   wire n_257_76_9897;
   wire n_257_76_9898;
   wire n_257_76_9899;
   wire n_257_76_9900;
   wire n_257_76_9901;
   wire n_257_76_9902;
   wire n_257_76_9903;
   wire n_257_76_9904;
   wire n_257_76_9905;
   wire n_257_76_9906;
   wire n_257_76_9907;
   wire n_257_76_9908;
   wire n_257_76_9909;
   wire n_257_76_9910;
   wire n_257_76_9911;
   wire n_257_76_9912;
   wire n_257_76_9913;
   wire n_257_76_9914;
   wire n_257_76_9915;
   wire n_257_76_9916;
   wire n_257_76_9917;
   wire n_257_76_9918;
   wire n_257_76_9919;
   wire n_257_76_9920;
   wire n_257_76_9921;
   wire n_257_76_9922;
   wire n_257_76_9923;
   wire n_257_76_9924;
   wire n_257_76_9925;
   wire n_257_76_9926;
   wire n_257_76_9927;
   wire n_257_76_9928;
   wire n_257_76_9929;
   wire n_257_76_9930;
   wire n_257_76_9931;
   wire n_257_76_9932;
   wire n_257_76_9933;
   wire n_257_76_9934;
   wire n_257_76_9935;
   wire n_257_76_9936;
   wire n_257_76_9937;
   wire n_257_76_9938;
   wire n_257_76_9939;
   wire n_257_76_9940;
   wire n_257_76_9941;
   wire n_257_76_9942;
   wire n_257_76_9943;
   wire n_257_76_9944;
   wire n_257_76_9945;
   wire n_257_76_9946;
   wire n_257_76_9947;
   wire n_257_76_9948;
   wire n_257_76_9949;
   wire n_257_76_9950;
   wire n_257_76_9951;
   wire n_257_76_9952;
   wire n_257_76_9953;
   wire n_257_76_9954;
   wire n_257_76_9955;
   wire n_257_76_9956;
   wire n_257_76_9957;
   wire n_257_76_9958;
   wire n_257_76_9959;
   wire n_257_76_9960;
   wire n_257_76_9961;
   wire n_257_76_9962;
   wire n_257_76_9963;
   wire n_257_76_9964;
   wire n_257_76_9965;
   wire n_257_76_9966;
   wire n_257_76_9967;
   wire n_257_76_9968;
   wire n_257_76_9969;
   wire n_257_76_9970;
   wire n_257_76_9971;
   wire n_257_76_9972;
   wire n_257_76_9973;
   wire n_257_76_9974;
   wire n_257_76_9975;
   wire n_257_76_9976;
   wire n_257_76_9977;
   wire n_257_76_9978;
   wire n_257_76_9979;
   wire n_257_76_9980;
   wire n_257_76_9981;
   wire n_257_76_9982;
   wire n_257_76_9983;
   wire n_257_76_9984;
   wire n_257_76_9985;
   wire n_257_76_9986;
   wire n_257_76_9987;
   wire n_257_76_9988;
   wire n_257_76_9989;
   wire n_257_76_9990;
   wire n_257_76_9991;
   wire n_257_76_9992;
   wire n_257_76_9993;
   wire n_257_76_9994;
   wire n_257_76_9995;
   wire n_257_76_9996;
   wire n_257_76_9997;
   wire n_257_76_9998;
   wire n_257_76_9999;
   wire n_257_76_10000;
   wire n_257_76_10001;
   wire n_257_76_10002;
   wire n_257_76_10003;
   wire n_257_76_10004;
   wire n_257_76_10005;
   wire n_257_76_10006;
   wire n_257_76_10007;
   wire n_257_76_10008;
   wire n_257_76_10009;
   wire n_257_76_10010;
   wire n_257_76_10011;
   wire n_257_76_10012;
   wire n_257_76_10013;
   wire n_257_76_10014;
   wire n_257_76_10015;
   wire n_257_76_10016;
   wire n_257_76_10017;
   wire n_257_76_10018;
   wire n_257_76_10019;
   wire n_257_76_10020;
   wire n_257_76_10021;
   wire n_257_76_10022;
   wire n_257_76_10023;
   wire n_257_76_10024;
   wire n_257_76_10025;
   wire n_257_76_10026;
   wire n_257_76_10027;
   wire n_257_76_10028;
   wire n_257_76_10029;
   wire n_257_76_10030;
   wire n_257_76_10031;
   wire n_257_76_10032;
   wire n_257_76_10033;
   wire n_257_76_10034;
   wire n_257_76_10035;
   wire n_257_76_10036;
   wire n_257_76_10037;
   wire n_257_76_10038;
   wire n_257_76_10039;
   wire n_257_76_10040;
   wire n_257_76_10041;
   wire n_257_76_10042;
   wire n_257_76_10043;
   wire n_257_76_10044;
   wire n_257_76_10045;
   wire n_257_76_10046;
   wire n_257_76_10047;
   wire n_257_76_10048;
   wire n_257_76_10049;
   wire n_257_76_10050;
   wire n_257_76_10051;
   wire n_257_76_10052;
   wire n_257_76_10053;
   wire n_257_76_10054;
   wire n_257_76_10055;
   wire n_257_76_10056;
   wire n_257_76_10057;
   wire n_257_76_10058;
   wire n_257_76_10059;
   wire n_257_76_10060;
   wire n_257_76_10061;
   wire n_257_76_10062;
   wire n_257_76_10063;
   wire n_257_76_10064;
   wire n_257_76_10065;
   wire n_257_76_10066;
   wire n_257_76_10067;
   wire n_257_76_10068;
   wire n_257_76_10069;
   wire n_257_76_10070;
   wire n_257_76_10071;
   wire n_257_76_10072;
   wire n_257_76_10073;
   wire n_257_76_10074;
   wire n_257_76_10075;
   wire n_257_76_10076;
   wire n_257_76_10077;
   wire n_257_76_10078;
   wire n_257_76_10079;
   wire n_257_76_10080;
   wire n_257_76_10081;
   wire n_257_76_10082;
   wire n_257_76_10083;
   wire n_257_76_10084;
   wire n_257_76_10085;
   wire n_257_76_10086;
   wire n_257_76_10087;
   wire n_257_76_10088;
   wire n_257_76_10089;
   wire n_257_76_10090;
   wire n_257_76_10091;
   wire n_257_76_10092;
   wire n_257_76_10093;
   wire n_257_76_10094;
   wire n_257_76_10095;
   wire n_257_76_10096;
   wire n_257_76_10097;
   wire n_257_76_10098;
   wire n_257_76_10099;
   wire n_257_76_10100;
   wire n_257_76_10101;
   wire n_257_76_10102;
   wire n_257_76_10103;
   wire n_257_76_10104;
   wire n_257_76_10105;
   wire n_257_76_10106;
   wire n_257_76_10107;
   wire n_257_76_10108;
   wire n_257_76_10109;
   wire n_257_76_10110;
   wire n_257_76_10111;
   wire n_257_76_10112;
   wire n_257_76_10113;
   wire n_257_76_10114;
   wire n_257_76_10115;
   wire n_257_76_10116;
   wire n_257_76_10117;
   wire n_257_76_10118;
   wire n_257_76_10119;
   wire n_257_76_10120;
   wire n_257_76_10121;
   wire n_257_76_10122;
   wire n_257_76_10123;
   wire n_257_76_10124;
   wire n_257_76_10125;
   wire n_257_76_10126;
   wire n_257_76_10127;
   wire n_257_76_10128;
   wire n_257_76_10129;
   wire n_257_76_10130;
   wire n_257_76_10131;
   wire n_257_76_10132;
   wire n_257_76_10133;
   wire n_257_76_10134;
   wire n_257_76_10135;
   wire n_257_76_10136;
   wire n_257_76_10137;
   wire n_257_76_10138;
   wire n_257_76_10139;
   wire n_257_76_10140;
   wire n_257_76_10141;
   wire n_257_76_10142;
   wire n_257_76_10143;
   wire n_257_76_10144;
   wire n_257_76_10145;
   wire n_257_76_10146;
   wire n_257_76_10147;
   wire n_257_76_10148;
   wire n_257_76_10149;
   wire n_257_76_10150;
   wire n_257_76_10151;
   wire n_257_76_10152;
   wire n_257_76_10153;
   wire n_257_76_10154;
   wire n_257_76_10155;
   wire n_257_76_10156;
   wire n_257_76_10157;
   wire n_257_76_10158;
   wire n_257_76_10159;
   wire n_257_76_10160;
   wire n_257_76_10161;
   wire n_257_76_10162;
   wire n_257_76_10163;
   wire n_257_76_10164;
   wire n_257_76_10165;
   wire n_257_76_10166;
   wire n_257_76_10167;
   wire n_257_76_10168;
   wire n_257_76_10169;
   wire n_257_76_10170;
   wire n_257_76_10171;
   wire n_257_76_10172;
   wire n_257_76_10173;
   wire n_257_76_10174;
   wire n_257_76_10175;
   wire n_257_76_10176;
   wire n_257_76_10177;
   wire n_257_76_10178;
   wire n_257_76_10179;
   wire n_257_76_10180;
   wire n_257_76_10181;
   wire n_257_76_10182;
   wire n_257_76_10183;
   wire n_257_76_10184;
   wire n_257_76_10185;
   wire n_257_76_10186;
   wire n_257_76_10187;
   wire n_257_76_10188;
   wire n_257_76_10189;
   wire n_257_76_10190;
   wire n_257_76_10191;
   wire n_257_76_10192;
   wire n_257_76_10193;
   wire n_257_76_10194;
   wire n_257_76_10195;
   wire n_257_76_10196;
   wire n_257_76_10197;
   wire n_257_76_10198;
   wire n_257_76_10199;
   wire n_257_76_10200;
   wire n_257_76_10201;
   wire n_257_76_10202;
   wire n_257_76_10203;
   wire n_257_76_10204;
   wire n_257_76_10205;
   wire n_257_76_10206;
   wire n_257_76_10207;
   wire n_257_76_10208;
   wire n_257_76_10209;
   wire n_257_76_10210;
   wire n_257_76_10211;
   wire n_257_76_10212;
   wire n_257_76_10213;
   wire n_257_76_10214;
   wire n_257_76_10215;
   wire n_257_76_10216;
   wire n_257_76_10217;
   wire n_257_76_10218;
   wire n_257_76_10219;
   wire n_257_76_10220;
   wire n_257_76_10221;
   wire n_257_76_10222;
   wire n_257_76_10223;
   wire n_257_76_10224;
   wire n_257_76_10225;
   wire n_257_76_10226;
   wire n_257_76_10227;
   wire n_257_76_10228;
   wire n_257_76_10229;
   wire n_257_76_10230;
   wire n_257_76_10231;
   wire n_257_76_10232;
   wire n_257_76_10233;
   wire n_257_76_10234;
   wire n_257_76_10235;
   wire n_257_76_10236;
   wire n_257_76_10237;
   wire n_257_76_10238;
   wire n_257_76_10239;
   wire n_257_76_10240;
   wire n_257_76_10241;
   wire n_257_76_10242;
   wire n_257_76_10243;
   wire n_257_76_10244;
   wire n_257_76_10245;
   wire n_257_76_10246;
   wire n_257_76_10247;
   wire n_257_76_10248;
   wire n_257_76_10249;
   wire n_257_76_10250;
   wire n_257_76_10251;
   wire n_257_76_10252;
   wire n_257_76_10253;
   wire n_257_76_10254;
   wire n_257_76_10255;
   wire n_257_76_10256;
   wire n_257_76_10257;
   wire n_257_76_10258;
   wire n_257_76_10259;
   wire n_257_76_10260;
   wire n_257_76_10261;
   wire n_257_76_10262;
   wire n_257_76_10263;
   wire n_257_76_10264;
   wire n_257_76_10265;
   wire n_257_76_10266;
   wire n_257_76_10267;
   wire n_257_76_10268;
   wire n_257_76_10269;
   wire n_257_76_10270;
   wire n_257_76_10271;
   wire n_257_76_10272;
   wire n_257_76_10273;
   wire n_257_76_10274;
   wire n_257_76_10275;
   wire n_257_76_10276;
   wire n_257_76_10277;
   wire n_257_76_10278;
   wire n_257_76_10279;
   wire n_257_76_10280;
   wire n_257_76_10281;
   wire n_257_76_10282;
   wire n_257_76_10283;
   wire n_257_76_10284;
   wire n_257_76_10285;
   wire n_257_76_10286;
   wire n_257_76_10287;
   wire n_257_76_10288;
   wire n_257_76_10289;
   wire n_257_76_10290;
   wire n_257_76_10291;
   wire n_257_76_10292;
   wire n_257_76_10293;
   wire n_257_76_10294;
   wire n_257_76_10295;
   wire n_257_76_10296;
   wire n_257_76_10297;
   wire n_257_76_10298;
   wire n_257_76_10299;
   wire n_257_76_10300;
   wire n_257_76_10301;
   wire n_257_76_10302;
   wire n_257_76_10303;
   wire n_257_76_10304;
   wire n_257_76_10305;
   wire n_257_76_10306;
   wire n_257_76_10307;
   wire n_257_76_10308;
   wire n_257_76_10309;
   wire n_257_76_10310;
   wire n_257_76_10311;
   wire n_257_76_10312;
   wire n_257_76_10313;
   wire n_257_76_10314;
   wire n_257_76_10315;
   wire n_257_76_10316;
   wire n_257_76_10317;
   wire n_257_76_10318;
   wire n_257_76_10319;
   wire n_257_76_10320;
   wire n_257_76_10321;
   wire n_257_76_10322;
   wire n_257_76_10323;
   wire n_257_76_10324;
   wire n_257_76_10325;
   wire n_257_76_10326;
   wire n_257_76_10327;
   wire n_257_76_10328;
   wire n_257_76_10329;
   wire n_257_76_10330;
   wire n_257_76_10331;
   wire n_257_76_10332;
   wire n_257_76_10333;
   wire n_257_76_10334;
   wire n_257_76_10335;
   wire n_257_76_10336;
   wire n_257_76_10337;
   wire n_257_76_10338;
   wire n_257_76_10339;
   wire n_257_76_10340;
   wire n_257_76_10341;
   wire n_257_76_10342;
   wire n_257_76_10343;
   wire n_257_76_10344;
   wire n_257_76_10345;
   wire n_257_76_10346;
   wire n_257_76_10347;
   wire n_257_76_10348;
   wire n_257_76_10349;
   wire n_257_76_10350;
   wire n_257_76_10351;
   wire n_257_76_10352;
   wire n_257_76_10353;
   wire n_257_76_10354;
   wire n_257_76_10355;
   wire n_257_76_10356;
   wire n_257_76_10357;
   wire n_257_76_10358;
   wire n_257_76_10359;
   wire n_257_76_10360;
   wire n_257_76_10361;
   wire n_257_76_10362;
   wire n_257_76_10363;
   wire n_257_76_10364;
   wire n_257_76_10365;
   wire n_257_76_10366;
   wire n_257_76_10367;
   wire n_257_76_10368;
   wire n_257_76_10369;
   wire n_257_76_10370;
   wire n_257_76_10371;
   wire n_257_76_10372;
   wire n_257_76_10373;
   wire n_257_76_10374;
   wire n_257_76_10375;
   wire n_257_76_10376;
   wire n_257_76_10377;
   wire n_257_76_10378;
   wire n_257_76_10379;
   wire n_257_76_10380;
   wire n_257_76_10381;
   wire n_257_76_10382;
   wire n_257_76_10383;
   wire n_257_76_10384;
   wire n_257_76_10385;
   wire n_257_76_10386;
   wire n_257_76_10387;
   wire n_257_76_10388;
   wire n_257_76_10389;
   wire n_257_76_10390;
   wire n_257_76_10391;
   wire n_257_76_10392;
   wire n_257_76_10393;
   wire n_257_76_10394;
   wire n_257_76_10395;
   wire n_257_76_10396;
   wire n_257_76_10397;
   wire n_257_76_10398;
   wire n_257_76_10399;
   wire n_257_76_10400;
   wire n_257_76_10401;
   wire n_257_76_10402;
   wire n_257_76_10403;
   wire n_257_76_10404;
   wire n_257_76_10405;
   wire n_257_76_10406;
   wire n_257_76_10407;
   wire n_257_76_10408;
   wire n_257_76_10409;
   wire n_257_76_10410;
   wire n_257_76_10411;
   wire n_257_76_10412;
   wire n_257_76_10413;
   wire n_257_76_10414;
   wire n_257_76_10415;
   wire n_257_76_10416;
   wire n_257_76_10417;
   wire n_257_76_10418;
   wire n_257_76_10419;
   wire n_257_76_10420;
   wire n_257_76_10421;
   wire n_257_76_10422;
   wire n_257_76_10423;
   wire n_257_76_10424;
   wire n_257_76_10425;
   wire n_257_76_10426;
   wire n_257_76_10427;
   wire n_257_76_10428;
   wire n_257_76_10429;
   wire n_257_76_10430;
   wire n_257_76_10431;
   wire n_257_76_10432;
   wire n_257_76_10433;
   wire n_257_76_10434;
   wire n_257_76_10435;
   wire n_257_76_10436;
   wire n_257_76_10437;
   wire n_257_76_10438;
   wire n_257_76_10439;
   wire n_257_76_10440;
   wire n_257_76_10441;
   wire n_257_76_10442;
   wire n_257_76_10443;
   wire n_257_76_10444;
   wire n_257_76_10445;
   wire n_257_76_10446;
   wire n_257_76_10447;
   wire n_257_76_10448;
   wire n_257_76_10449;
   wire n_257_76_10450;
   wire n_257_76_10451;
   wire n_257_76_10452;
   wire n_257_76_10453;
   wire n_257_76_10454;
   wire n_257_76_10455;
   wire n_257_76_10456;
   wire n_257_76_10457;
   wire n_257_76_10458;
   wire n_257_76_10459;
   wire n_257_76_10460;
   wire n_257_76_10461;
   wire n_257_76_10462;
   wire n_257_76_10463;
   wire n_257_76_10464;
   wire n_257_76_10465;
   wire n_257_76_10466;
   wire n_257_76_10467;
   wire n_257_76_10468;
   wire n_257_76_10469;
   wire n_257_76_10470;
   wire n_257_76_10471;
   wire n_257_76_10472;
   wire n_257_76_10473;
   wire n_257_76_10474;
   wire n_257_76_10475;
   wire n_257_76_10476;
   wire n_257_76_10477;
   wire n_257_76_10478;
   wire n_257_76_10479;
   wire n_257_76_10480;
   wire n_257_76_10481;
   wire n_257_76_10482;
   wire n_257_76_10483;
   wire n_257_76_10484;
   wire n_257_76_10485;
   wire n_257_76_10486;
   wire n_257_76_10487;
   wire n_257_76_10488;
   wire n_257_76_10489;
   wire n_257_76_10490;
   wire n_257_76_10491;
   wire n_257_76_10492;
   wire n_257_76_10493;
   wire n_257_76_10494;
   wire n_257_76_10495;
   wire n_257_76_10496;
   wire n_257_76_10497;
   wire n_257_76_10498;
   wire n_257_76_10499;
   wire n_257_76_10500;
   wire n_257_76_10501;
   wire n_257_76_10502;
   wire n_257_76_10503;
   wire n_257_76_10504;
   wire n_257_76_10505;
   wire n_257_76_10506;
   wire n_257_76_10507;
   wire n_257_76_10508;
   wire n_257_76_10509;
   wire n_257_76_10510;
   wire n_257_76_10511;
   wire n_257_76_10512;
   wire n_257_76_10513;
   wire n_257_76_10514;
   wire n_257_76_10515;
   wire n_257_76_10516;
   wire n_257_76_10517;
   wire n_257_76_10518;
   wire n_257_76_10519;
   wire n_257_76_10520;
   wire n_257_76_10521;
   wire n_257_76_10522;
   wire n_257_76_10523;
   wire n_257_76_10524;
   wire n_257_76_10525;
   wire n_257_76_10526;
   wire n_257_76_10527;
   wire n_257_76_10528;
   wire n_257_76_10529;
   wire n_257_76_10530;
   wire n_257_76_10531;
   wire n_257_76_10532;
   wire n_257_76_10533;
   wire n_257_76_10534;
   wire n_257_76_10535;
   wire n_257_76_10536;
   wire n_257_76_10537;
   wire n_257_76_10538;
   wire n_257_76_10539;
   wire n_257_76_10540;
   wire n_257_76_10541;
   wire n_257_76_10542;
   wire n_257_76_10543;
   wire n_257_76_10544;
   wire n_257_76_10545;
   wire n_257_76_10546;
   wire n_257_76_10547;
   wire n_257_76_10548;
   wire n_257_76_10549;
   wire n_257_76_10550;
   wire n_257_76_10551;
   wire n_257_76_10552;
   wire n_257_76_10553;
   wire n_257_76_10554;
   wire n_257_76_10555;
   wire n_257_76_10556;
   wire n_257_76_10557;
   wire n_257_76_10558;
   wire n_257_76_10559;
   wire n_257_76_10560;
   wire n_257_76_10561;
   wire n_257_76_10562;
   wire n_257_76_10563;
   wire n_257_76_10564;
   wire n_257_76_10565;
   wire n_257_76_10566;
   wire n_257_76_10567;
   wire n_257_76_10568;
   wire n_257_76_10569;
   wire n_257_76_10570;
   wire n_257_76_10571;
   wire n_257_76_10572;
   wire n_257_76_10573;
   wire n_257_76_10574;
   wire n_257_76_10575;
   wire n_257_76_10576;
   wire n_257_76_10577;
   wire n_257_76_10578;
   wire n_257_76_10579;
   wire n_257_76_10580;
   wire n_257_76_10581;
   wire n_257_76_10582;
   wire n_257_76_10583;
   wire n_257_76_10584;
   wire n_257_76_10585;
   wire n_257_76_10586;
   wire n_257_76_10587;
   wire n_257_76_10588;
   wire n_257_76_10589;
   wire n_257_76_10590;
   wire n_257_76_10591;
   wire n_257_76_10592;
   wire n_257_76_10593;
   wire n_257_76_10594;
   wire n_257_76_10595;
   wire n_257_76_10596;
   wire n_257_76_10597;
   wire n_257_76_10598;
   wire n_257_76_10599;
   wire n_257_76_10600;
   wire n_257_76_10601;
   wire n_257_76_10602;
   wire n_257_76_10603;
   wire n_257_76_10604;
   wire n_257_76_10605;
   wire n_257_76_10606;
   wire n_257_76_10607;
   wire n_257_76_10608;
   wire n_257_76_10609;
   wire n_257_76_10610;
   wire n_257_76_10611;
   wire n_257_76_10612;
   wire n_257_76_10613;
   wire n_257_76_10614;
   wire n_257_76_10615;
   wire n_257_76_10616;
   wire n_257_76_10617;
   wire n_257_76_10618;
   wire n_257_76_10619;
   wire n_257_76_10620;
   wire n_257_76_10621;
   wire n_257_76_10622;
   wire n_257_76_10623;
   wire n_257_76_10624;
   wire n_257_76_10625;
   wire n_257_76_10626;
   wire n_257_76_10627;
   wire n_257_76_10628;
   wire n_257_76_10629;
   wire n_257_76_10630;
   wire n_257_76_10631;
   wire n_257_76_10632;
   wire n_257_76_10633;
   wire n_257_76_10634;
   wire n_257_76_10635;
   wire n_257_76_10636;
   wire n_257_76_10637;
   wire n_257_76_10638;
   wire n_257_76_10639;
   wire n_257_76_10640;
   wire n_257_76_10641;
   wire n_257_76_10642;
   wire n_257_76_10643;
   wire n_257_76_10644;
   wire n_257_76_10645;
   wire n_257_76_10646;
   wire n_257_76_10647;
   wire n_257_76_10648;
   wire n_257_76_10649;
   wire n_257_76_10650;
   wire n_257_76_10651;
   wire n_257_76_10652;
   wire n_257_76_10653;
   wire n_257_76_10654;
   wire n_257_76_10655;
   wire n_257_76_10656;
   wire n_257_76_10657;
   wire n_257_76_10658;
   wire n_257_76_10659;
   wire n_257_76_10660;
   wire n_257_76_10661;
   wire n_257_76_10662;
   wire n_257_76_10663;
   wire n_257_76_10664;
   wire n_257_76_10665;
   wire n_257_76_10666;
   wire n_257_76_10667;
   wire n_257_76_10668;
   wire n_257_76_10669;
   wire n_257_76_10670;
   wire n_257_76_10671;
   wire n_257_76_10672;
   wire n_257_76_10673;
   wire n_257_76_10674;
   wire n_257_76_10675;
   wire n_257_76_10676;
   wire n_257_76_10677;
   wire n_257_76_10678;
   wire n_257_76_10679;
   wire n_257_76_10680;
   wire n_257_76_10681;
   wire n_257_76_10682;
   wire n_257_76_10683;
   wire n_257_76_10684;
   wire n_257_76_10685;
   wire n_257_76_10686;
   wire n_257_76_10687;
   wire n_257_76_10688;
   wire n_257_76_10689;
   wire n_257_76_10690;
   wire n_257_76_10691;
   wire n_257_76_10692;
   wire n_257_76_10693;
   wire n_257_76_10694;
   wire n_257_76_10695;
   wire n_257_76_10696;
   wire n_257_76_10697;
   wire n_257_76_10698;
   wire n_257_76_10699;
   wire n_257_76_10700;
   wire n_257_76_10701;
   wire n_257_76_10702;
   wire n_257_76_10703;
   wire n_257_76_10704;
   wire n_257_76_10705;
   wire n_257_76_10706;
   wire n_257_76_10707;
   wire n_257_76_10708;
   wire n_257_76_10709;
   wire n_257_76_10710;
   wire n_257_76_10711;
   wire n_257_76_10712;
   wire n_257_76_10713;
   wire n_257_76_10714;
   wire n_257_76_10715;
   wire n_257_76_10716;
   wire n_257_76_10717;
   wire n_257_76_10718;
   wire n_257_76_10719;
   wire n_257_76_10720;
   wire n_257_76_10721;
   wire n_257_76_10722;
   wire n_257_76_10723;
   wire n_257_76_10724;
   wire n_257_76_10725;
   wire n_257_76_10726;
   wire n_257_76_10727;
   wire n_257_76_10728;
   wire n_257_76_10729;
   wire n_257_76_10730;
   wire n_257_76_10731;
   wire n_257_76_10732;
   wire n_257_76_10733;
   wire n_257_76_10734;
   wire n_257_76_10735;
   wire n_257_76_10736;
   wire n_257_76_10737;
   wire n_257_76_10738;
   wire n_257_76_10739;
   wire n_257_76_10740;
   wire n_257_76_10741;
   wire n_257_76_10742;
   wire n_257_76_10743;
   wire n_257_76_10744;
   wire n_257_76_10745;
   wire n_257_76_10746;
   wire n_257_76_10747;
   wire n_257_76_10748;
   wire n_257_76_10749;
   wire n_257_76_10750;
   wire n_257_76_10751;
   wire n_257_76_10752;
   wire n_257_76_10753;
   wire n_257_76_10754;
   wire n_257_76_10755;
   wire n_257_76_10756;
   wire n_257_76_10757;
   wire n_257_76_10758;
   wire n_257_76_10759;
   wire n_257_76_10760;
   wire n_257_76_10761;
   wire n_257_76_10762;
   wire n_257_76_10763;
   wire n_257_76_10764;
   wire n_257_76_10765;
   wire n_257_76_10766;
   wire n_257_76_10767;
   wire n_257_76_10768;
   wire n_257_76_10769;
   wire n_257_76_10770;
   wire n_257_76_10771;
   wire n_257_76_10772;
   wire n_257_76_10773;
   wire n_257_76_10774;
   wire n_257_76_10775;
   wire n_257_76_10776;
   wire n_257_76_10777;
   wire n_257_76_10778;
   wire n_257_76_10779;
   wire n_257_76_10780;
   wire n_257_76_10781;
   wire n_257_76_10782;
   wire n_257_76_10783;
   wire n_257_76_10784;
   wire n_257_76_10785;
   wire n_257_76_10786;
   wire n_257_76_10787;
   wire n_257_76_10788;
   wire n_257_76_10789;
   wire n_257_76_10790;
   wire n_257_76_10791;
   wire n_257_76_10792;
   wire n_257_76_10793;
   wire n_257_76_10794;
   wire n_257_76_10795;
   wire n_257_76_10796;
   wire n_257_76_10797;
   wire n_257_76_10798;
   wire n_257_76_10799;
   wire n_257_76_10800;
   wire n_257_76_10801;
   wire n_257_76_10802;
   wire n_257_76_10803;
   wire n_257_76_10804;
   wire n_257_76_10805;
   wire n_257_76_10806;
   wire n_257_76_10807;
   wire n_257_76_10808;
   wire n_257_76_10809;
   wire n_257_76_10810;
   wire n_257_76_10811;
   wire n_257_76_10812;
   wire n_257_76_10813;
   wire n_257_76_10814;
   wire n_257_76_10815;
   wire n_257_76_10816;
   wire n_257_76_10817;
   wire n_257_76_10818;
   wire n_257_76_10819;
   wire n_257_76_10820;
   wire n_257_76_10821;
   wire n_257_76_10822;
   wire n_257_76_10823;
   wire n_257_76_10824;
   wire n_257_76_10825;
   wire n_257_76_10826;
   wire n_257_76_10827;
   wire n_257_76_10828;
   wire n_257_76_10829;
   wire n_257_76_10830;
   wire n_257_76_10831;
   wire n_257_76_10832;
   wire n_257_76_10833;
   wire n_257_76_10834;
   wire n_257_76_10835;
   wire n_257_76_10836;
   wire n_257_76_10837;
   wire n_257_76_10838;
   wire n_257_76_10839;
   wire n_257_76_10840;
   wire n_257_76_10841;
   wire n_257_76_10842;
   wire n_257_76_10843;
   wire n_257_76_10844;
   wire n_257_76_10845;
   wire n_257_76_10846;
   wire n_257_76_10847;
   wire n_257_76_10848;
   wire n_257_76_10849;
   wire n_257_76_10850;
   wire n_257_76_10851;
   wire n_257_76_10852;
   wire n_257_76_10853;
   wire n_257_76_10854;
   wire n_257_76_10855;
   wire n_257_76_10856;
   wire n_257_76_10857;
   wire n_257_76_10858;
   wire n_257_76_10859;
   wire n_257_76_10860;
   wire n_257_76_10861;
   wire n_257_76_10862;
   wire n_257_76_10863;
   wire n_257_76_10864;
   wire n_257_76_10865;
   wire n_257_76_10866;
   wire n_257_76_10867;
   wire n_257_76_10868;
   wire n_257_76_10869;
   wire n_257_76_10870;
   wire n_257_76_10871;
   wire n_257_76_10872;
   wire n_257_76_10873;
   wire n_257_76_10874;
   wire n_257_76_10875;
   wire n_257_76_10876;
   wire n_257_76_10877;
   wire n_257_76_10878;
   wire n_257_76_10879;
   wire n_257_76_10880;
   wire n_257_76_10881;
   wire n_257_76_10882;
   wire n_257_76_10883;
   wire n_257_76_10884;
   wire n_257_76_10885;
   wire n_257_76_10886;
   wire n_257_76_10887;
   wire n_257_76_10888;
   wire n_257_76_10889;
   wire n_257_76_10890;
   wire n_257_76_10891;
   wire n_257_76_10892;
   wire n_257_76_10893;
   wire n_257_76_10894;
   wire n_257_76_10895;
   wire n_257_76_10896;
   wire n_257_76_10897;
   wire n_257_76_10898;
   wire n_257_76_10899;
   wire n_257_76_10900;
   wire n_257_76_10901;
   wire n_257_76_10902;
   wire n_257_76_10903;
   wire n_257_76_10904;
   wire n_257_76_10905;
   wire n_257_76_10906;
   wire n_257_76_10907;
   wire n_257_76_10908;
   wire n_257_76_10909;
   wire n_257_76_10910;
   wire n_257_76_10911;
   wire n_257_76_10912;
   wire n_257_76_10913;
   wire n_257_76_10914;
   wire n_257_76_10915;
   wire n_257_76_10916;
   wire n_257_76_10917;
   wire n_257_76_10918;
   wire n_257_76_10919;
   wire n_257_76_10920;
   wire n_257_76_10921;
   wire n_257_76_10922;
   wire n_257_76_10923;
   wire n_257_76_10924;
   wire n_257_76_10925;
   wire n_257_76_10926;
   wire n_257_76_10927;
   wire n_257_76_10928;
   wire n_257_76_10929;
   wire n_257_76_10930;
   wire n_257_76_10931;
   wire n_257_76_10932;
   wire n_257_76_10933;
   wire n_257_76_10934;
   wire n_257_76_10935;
   wire n_257_76_10936;
   wire n_257_76_10937;
   wire n_257_76_10938;
   wire n_257_76_10939;
   wire n_257_76_10940;
   wire n_257_76_10941;
   wire n_257_76_10942;
   wire n_257_76_10943;
   wire n_257_76_10944;
   wire n_257_76_10945;
   wire n_257_76_10946;
   wire n_257_76_10947;
   wire n_257_76_10948;
   wire n_257_76_10949;
   wire n_257_76_10950;
   wire n_257_76_10951;
   wire n_257_76_10952;
   wire n_257_76_10953;
   wire n_257_76_10954;
   wire n_257_76_10955;
   wire n_257_76_10956;
   wire n_257_76_10957;
   wire n_257_76_10958;
   wire n_257_76_10959;
   wire n_257_76_10960;
   wire n_257_76_10961;
   wire n_257_76_10962;
   wire n_257_76_10963;
   wire n_257_76_10964;
   wire n_257_76_10965;
   wire n_257_76_10966;
   wire n_257_76_10967;
   wire n_257_76_10968;
   wire n_257_76_10969;
   wire n_257_76_10970;
   wire n_257_76_10971;
   wire n_257_76_10972;
   wire n_257_76_10973;
   wire n_257_76_10974;
   wire n_257_76_10975;
   wire n_257_76_10976;
   wire n_257_76_10977;
   wire n_257_76_10978;
   wire n_257_76_10979;
   wire n_257_76_10980;
   wire n_257_76_10981;
   wire n_257_76_10982;
   wire n_257_76_10983;
   wire n_257_76_10984;
   wire n_257_76_10985;
   wire n_257_76_10986;
   wire n_257_76_10987;
   wire n_257_76_10988;
   wire n_257_76_10989;
   wire n_257_76_10990;
   wire n_257_76_10991;
   wire n_257_76_10992;
   wire n_257_76_10993;
   wire n_257_76_10994;
   wire n_257_76_10995;
   wire n_257_76_10996;
   wire n_257_76_10997;
   wire n_257_76_10998;
   wire n_257_76_10999;
   wire n_257_76_11000;
   wire n_257_76_11001;
   wire n_257_76_11002;
   wire n_257_76_11003;
   wire n_257_76_11004;
   wire n_257_76_11005;
   wire n_257_76_11006;
   wire n_257_76_11007;
   wire n_257_76_11008;
   wire n_257_76_11009;
   wire n_257_76_11010;
   wire n_257_76_11011;
   wire n_257_76_11012;
   wire n_257_76_11013;
   wire n_257_76_11014;
   wire n_257_76_11015;
   wire n_257_76_11016;
   wire n_257_76_11017;
   wire n_257_76_11018;
   wire n_257_76_11019;
   wire n_257_76_11020;
   wire n_257_76_11021;
   wire n_257_76_11022;
   wire n_257_76_11023;
   wire n_257_76_11024;
   wire n_257_76_11025;
   wire n_257_76_11026;
   wire n_257_76_11027;
   wire n_257_76_11028;
   wire n_257_76_11029;
   wire n_257_76_11030;
   wire n_257_76_11031;
   wire n_257_76_11032;
   wire n_257_76_11033;
   wire n_257_76_11034;
   wire n_257_76_11035;
   wire n_257_76_11036;
   wire n_257_76_11037;
   wire n_257_76_11038;
   wire n_257_76_11039;
   wire n_257_76_11040;
   wire n_257_76_11041;
   wire n_257_76_11042;
   wire n_257_76_11043;
   wire n_257_76_11044;
   wire n_257_76_11045;
   wire n_257_76_11046;
   wire n_257_76_11047;
   wire n_257_76_11048;
   wire n_257_76_11049;
   wire n_257_76_11050;
   wire n_257_76_11051;
   wire n_257_76_11052;
   wire n_257_76_11053;
   wire n_257_76_11054;
   wire n_257_76_11055;
   wire n_257_76_11056;
   wire n_257_76_11057;
   wire n_257_76_11058;
   wire n_257_76_11059;
   wire n_257_76_11060;
   wire n_257_76_11061;
   wire n_257_76_11062;
   wire n_257_76_11063;
   wire n_257_76_11064;
   wire n_257_76_11065;
   wire n_257_76_11066;
   wire n_257_76_11067;
   wire n_257_76_11068;
   wire n_257_76_11069;
   wire n_257_76_11070;
   wire n_257_76_11071;
   wire n_257_76_11072;
   wire n_257_76_11073;
   wire n_257_76_11074;
   wire n_257_76_11075;
   wire n_257_76_11076;
   wire n_257_76_11077;
   wire n_257_76_11078;
   wire n_257_76_11079;
   wire n_257_76_11080;
   wire n_257_76_11081;
   wire n_257_76_11082;
   wire n_257_76_11083;
   wire n_257_76_11084;
   wire n_257_76_11085;
   wire n_257_76_11086;
   wire n_257_76_11087;
   wire n_257_76_11088;
   wire n_257_76_11089;
   wire n_257_76_11090;
   wire n_257_76_11091;
   wire n_257_76_11092;
   wire n_257_76_11093;
   wire n_257_76_11094;
   wire n_257_76_11095;
   wire n_257_76_11096;
   wire n_257_76_11097;
   wire n_257_76_11098;
   wire n_257_76_11099;
   wire n_257_76_11100;
   wire n_257_76_11101;
   wire n_257_76_11102;
   wire n_257_76_11103;
   wire n_257_76_11104;
   wire n_257_76_11105;
   wire n_257_76_11106;
   wire n_257_76_11107;
   wire n_257_76_11108;
   wire n_257_76_11109;
   wire n_257_76_11110;
   wire n_257_76_11111;
   wire n_257_76_11112;
   wire n_257_76_11113;
   wire n_257_76_11114;
   wire n_257_76_11115;
   wire n_257_76_11116;
   wire n_257_76_11117;
   wire n_257_76_11118;
   wire n_257_76_11119;
   wire n_257_76_11120;
   wire n_257_76_11121;
   wire n_257_76_11122;
   wire n_257_76_11123;
   wire n_257_76_11124;
   wire n_257_76_11125;
   wire n_257_76_11126;
   wire n_257_76_11127;
   wire n_257_76_11128;
   wire n_257_76_11129;
   wire n_257_76_11130;
   wire n_257_76_11131;
   wire n_257_76_11132;
   wire n_257_76_11133;
   wire n_257_76_11134;
   wire n_257_76_11135;
   wire n_257_76_11136;
   wire n_257_76_11137;
   wire n_257_76_11138;
   wire n_257_76_11139;
   wire n_257_76_11140;
   wire n_257_76_11141;
   wire n_257_76_11142;
   wire n_257_76_11143;
   wire n_257_76_11144;
   wire n_257_76_11145;
   wire n_257_76_11146;
   wire n_257_76_11147;
   wire n_257_76_11148;
   wire n_257_76_11149;
   wire n_257_76_11150;
   wire n_257_76_11151;
   wire n_257_76_11152;
   wire n_257_76_11153;
   wire n_257_76_11154;
   wire n_257_76_11155;
   wire n_257_76_11156;
   wire n_257_76_11157;
   wire n_257_76_11158;
   wire n_257_76_11159;
   wire n_257_76_11160;
   wire n_257_76_11161;
   wire n_257_76_11162;
   wire n_257_76_11163;
   wire n_257_76_11164;
   wire n_257_76_11165;
   wire n_257_76_11166;
   wire n_257_76_11167;
   wire n_257_76_11168;
   wire n_257_76_11169;
   wire n_257_76_11170;
   wire n_257_76_11171;
   wire n_257_76_11172;
   wire n_257_76_11173;
   wire n_257_76_11174;
   wire n_257_76_11175;
   wire n_257_76_11176;
   wire n_257_76_11177;
   wire n_257_76_11178;
   wire n_257_76_11179;
   wire n_257_76_11180;
   wire n_257_76_11181;
   wire n_257_76_11182;
   wire n_257_76_11183;
   wire n_257_76_11184;
   wire n_257_76_11185;
   wire n_257_76_11186;
   wire n_257_76_11187;
   wire n_257_76_11188;
   wire n_257_76_11189;
   wire n_257_76_11190;
   wire n_257_76_11191;
   wire n_257_76_11192;
   wire n_257_76_11193;
   wire n_257_76_11194;
   wire n_257_76_11195;
   wire n_257_76_11196;
   wire n_257_76_11197;
   wire n_257_76_11198;
   wire n_257_76_11199;
   wire n_257_76_11200;
   wire n_257_76_11201;
   wire n_257_76_11202;
   wire n_257_76_11203;
   wire n_257_76_11204;
   wire n_257_76_11205;
   wire n_257_76_11206;
   wire n_257_76_11207;
   wire n_257_76_11208;
   wire n_257_76_11209;
   wire n_257_76_11210;
   wire n_257_76_11211;
   wire n_257_76_11212;
   wire n_257_76_11213;
   wire n_257_76_11214;
   wire n_257_76_11215;
   wire n_257_76_11216;
   wire n_257_76_11217;
   wire n_257_76_11218;
   wire n_257_76_11219;
   wire n_257_76_11220;
   wire n_257_76_11221;
   wire n_257_76_11222;
   wire n_257_76_11223;
   wire n_257_76_11224;
   wire n_257_76_11225;
   wire n_257_76_11226;
   wire n_257_76_11227;
   wire n_257_76_11228;
   wire n_257_76_11229;
   wire n_257_76_11230;
   wire n_257_76_11231;
   wire n_257_76_11232;
   wire n_257_76_11233;
   wire n_257_76_11234;
   wire n_257_76_11235;
   wire n_257_76_11236;
   wire n_257_76_11237;
   wire n_257_76_11238;
   wire n_257_76_11239;
   wire n_257_76_11240;
   wire n_257_76_11241;
   wire n_257_76_11242;
   wire n_257_76_11243;
   wire n_257_76_11244;
   wire n_257_76_11245;
   wire n_257_76_11246;
   wire n_257_76_11247;
   wire n_257_76_11248;
   wire n_257_76_11249;
   wire n_257_76_11250;
   wire n_257_76_11251;
   wire n_257_76_11252;
   wire n_257_76_11253;
   wire n_257_76_11254;
   wire n_257_76_11255;
   wire n_257_76_11256;
   wire n_257_76_11257;
   wire n_257_76_11258;
   wire n_257_76_11259;
   wire n_257_76_11260;
   wire n_257_76_11261;
   wire n_257_76_11262;
   wire n_257_76_11263;
   wire n_257_76_11264;
   wire n_257_76_11265;
   wire n_257_76_11266;
   wire n_257_76_11267;
   wire n_257_76_11268;
   wire n_257_76_11269;
   wire n_257_76_11270;
   wire n_257_76_11271;
   wire n_257_76_11272;
   wire n_257_76_11273;
   wire n_257_76_11274;
   wire n_257_76_11275;
   wire n_257_76_11276;
   wire n_257_76_11277;
   wire n_257_76_11278;
   wire n_257_76_11279;
   wire n_257_76_11280;
   wire n_257_76_11281;
   wire n_257_76_11282;
   wire n_257_76_11283;
   wire n_257_76_11284;
   wire n_257_76_11285;
   wire n_257_76_11286;
   wire n_257_76_11287;
   wire n_257_76_11288;
   wire n_257_76_11289;
   wire n_257_76_11290;
   wire n_257_76_11291;
   wire n_257_76_11292;
   wire n_257_76_11293;
   wire n_257_76_11294;
   wire n_257_76_11295;
   wire n_257_76_11296;
   wire n_257_76_11297;
   wire n_257_76_11298;
   wire n_257_76_11299;
   wire n_257_76_11300;
   wire n_257_76_11301;
   wire n_257_76_11302;
   wire n_257_76_11303;
   wire n_257_76_11304;
   wire n_257_76_11305;
   wire n_257_76_11306;
   wire n_257_76_11307;
   wire n_257_76_11308;
   wire n_257_76_11309;
   wire n_257_76_11310;
   wire n_257_76_11311;
   wire n_257_76_11312;
   wire n_257_76_11313;
   wire n_257_76_11314;
   wire n_257_76_11315;
   wire n_257_76_11316;
   wire n_257_76_11317;
   wire n_257_76_11318;
   wire n_257_76_11319;
   wire n_257_76_11320;
   wire n_257_76_11321;
   wire n_257_76_11322;
   wire n_257_76_11323;
   wire n_257_76_11324;
   wire n_257_76_11325;
   wire n_257_76_11326;
   wire n_257_76_11327;
   wire n_257_76_11328;
   wire n_257_76_11329;
   wire n_257_76_11330;
   wire n_257_76_11331;
   wire n_257_76_11332;
   wire n_257_76_11333;
   wire n_257_76_11334;
   wire n_257_76_11335;
   wire n_257_76_11336;
   wire n_257_76_11337;
   wire n_257_76_11338;
   wire n_257_76_11339;
   wire n_257_76_11340;
   wire n_257_76_11341;
   wire n_257_76_11342;
   wire n_257_76_11343;
   wire n_257_76_11344;
   wire n_257_76_11345;
   wire n_257_76_11346;
   wire n_257_76_11347;
   wire n_257_76_11348;
   wire n_257_76_11349;
   wire n_257_76_11350;
   wire n_257_76_11351;
   wire n_257_76_11352;
   wire n_257_76_11353;
   wire n_257_76_11354;
   wire n_257_76_11355;
   wire n_257_76_11356;
   wire n_257_76_11357;
   wire n_257_76_11358;
   wire n_257_76_11359;
   wire n_257_76_11360;
   wire n_257_76_11361;
   wire n_257_76_11362;
   wire n_257_76_11363;
   wire n_257_76_11364;
   wire n_257_76_11365;
   wire n_257_76_11366;
   wire n_257_76_11367;
   wire n_257_76_11368;
   wire n_257_76_11369;
   wire n_257_76_11370;
   wire n_257_76_11371;
   wire n_257_76_11372;
   wire n_257_76_11373;
   wire n_257_76_11374;
   wire n_257_76_11375;
   wire n_257_76_11376;
   wire n_257_76_11377;
   wire n_257_76_11378;
   wire n_257_76_11379;
   wire n_257_76_11380;
   wire n_257_76_11381;
   wire n_257_76_11382;
   wire n_257_76_11383;
   wire n_257_76_11384;
   wire n_257_76_11385;
   wire n_257_76_11386;
   wire n_257_76_11387;
   wire n_257_76_11388;
   wire n_257_76_11389;
   wire n_257_76_11390;
   wire n_257_76_11391;
   wire n_257_76_11392;
   wire n_257_76_11393;
   wire n_257_76_11394;
   wire n_257_76_11395;
   wire n_257_76_11396;
   wire n_257_76_11397;
   wire n_257_76_11398;
   wire n_257_76_11399;
   wire n_257_76_11400;
   wire n_257_76_11401;
   wire n_257_76_11402;
   wire n_257_76_11403;
   wire n_257_76_11404;
   wire n_257_76_11405;
   wire n_257_76_11406;
   wire n_257_76_11407;
   wire n_257_76_11408;
   wire n_257_76_11409;
   wire n_257_76_11410;
   wire n_257_76_11411;
   wire n_257_76_11412;
   wire n_257_76_11413;
   wire n_257_76_11414;
   wire n_257_76_11415;
   wire n_257_76_11416;
   wire n_257_76_11417;
   wire n_257_76_11418;
   wire n_257_76_11419;
   wire n_257_76_11420;
   wire n_257_76_11421;
   wire n_257_76_11422;
   wire n_257_76_11423;
   wire n_257_76_11424;
   wire n_257_76_11425;
   wire n_257_76_11426;
   wire n_257_76_11427;
   wire n_257_76_11428;
   wire n_257_76_11429;
   wire n_257_76_11430;
   wire n_257_76_11431;
   wire n_257_76_11432;
   wire n_257_76_11433;
   wire n_257_76_11434;
   wire n_257_76_11435;
   wire n_257_76_11436;
   wire n_257_76_11437;
   wire n_257_76_11438;
   wire n_257_76_11439;
   wire n_257_76_11440;
   wire n_257_76_11441;
   wire n_257_76_11442;
   wire n_257_76_11443;
   wire n_257_76_11444;
   wire n_257_76_11445;
   wire n_257_76_11446;
   wire n_257_76_11447;
   wire n_257_76_11448;
   wire n_257_76_11449;
   wire n_257_76_11450;
   wire n_257_76_11451;
   wire n_257_76_11452;
   wire n_257_76_11453;
   wire n_257_76_11454;
   wire n_257_76_11455;
   wire n_257_76_11456;
   wire n_257_76_11457;
   wire n_257_76_11458;
   wire n_257_76_11459;
   wire n_257_76_11460;
   wire n_257_76_11461;
   wire n_257_76_11462;
   wire n_257_76_11463;
   wire n_257_76_11464;
   wire n_257_76_11465;
   wire n_257_76_11466;
   wire n_257_76_11467;
   wire n_257_76_11468;
   wire n_257_76_11469;
   wire n_257_76_11470;
   wire n_257_76_11471;
   wire n_257_76_11472;
   wire n_257_76_11473;
   wire n_257_76_11474;
   wire n_257_76_11475;
   wire n_257_76_11476;
   wire n_257_76_11477;
   wire n_257_76_11478;
   wire n_257_76_11479;
   wire n_257_76_11480;
   wire n_257_76_11481;
   wire n_257_76_11482;
   wire n_257_76_11483;
   wire n_257_76_11484;
   wire n_257_76_11485;
   wire n_257_76_11486;
   wire n_257_76_11487;
   wire n_257_76_11488;
   wire n_257_76_11489;
   wire n_257_76_11490;
   wire n_257_76_11491;
   wire n_257_76_11492;
   wire n_257_76_11493;
   wire n_257_76_11494;
   wire n_257_76_11495;
   wire n_257_76_11496;
   wire n_257_76_11497;
   wire n_257_76_11498;
   wire n_257_76_11499;
   wire n_257_76_11500;
   wire n_257_76_11501;
   wire n_257_76_11502;
   wire n_257_76_11503;
   wire n_257_76_11504;
   wire n_257_76_11505;
   wire n_257_76_11506;
   wire n_257_76_11507;
   wire n_257_76_11508;
   wire n_257_76_11509;
   wire n_257_76_11510;
   wire n_257_76_11511;
   wire n_257_76_11512;
   wire n_257_76_11513;
   wire n_257_76_11514;
   wire n_257_76_11515;
   wire n_257_76_11516;
   wire n_257_76_11517;
   wire n_257_76_11518;
   wire n_257_76_11519;
   wire n_257_76_11520;
   wire n_257_76_11521;
   wire n_257_76_11522;
   wire n_257_76_11523;
   wire n_257_76_11524;
   wire n_257_76_11525;
   wire n_257_76_11526;
   wire n_257_76_11527;
   wire n_257_76_11528;
   wire n_257_76_11529;
   wire n_257_76_11530;
   wire n_257_76_11531;
   wire n_257_76_11532;
   wire n_257_76_11533;
   wire n_257_76_11534;
   wire n_257_76_11535;
   wire n_257_76_11536;
   wire n_257_76_11537;
   wire n_257_76_11538;
   wire n_257_76_11539;
   wire n_257_76_11540;
   wire n_257_76_11541;
   wire n_257_76_11542;
   wire n_257_76_11543;
   wire n_257_76_11544;
   wire n_257_76_11545;
   wire n_257_76_11546;
   wire n_257_76_11547;
   wire n_257_76_11548;
   wire n_257_76_11549;
   wire n_257_76_11550;
   wire n_257_76_11551;
   wire n_257_76_11552;
   wire n_257_76_11553;
   wire n_257_76_11554;
   wire n_257_76_11555;
   wire n_257_76_11556;
   wire n_257_76_11557;
   wire n_257_76_11558;
   wire n_257_76_11559;
   wire n_257_76_11560;
   wire n_257_76_11561;
   wire n_257_76_11562;
   wire n_257_76_11563;
   wire n_257_76_11564;
   wire n_257_76_11565;
   wire n_257_76_11566;
   wire n_257_76_11567;
   wire n_257_76_11568;
   wire n_257_76_11569;
   wire n_257_76_11570;
   wire n_257_76_11571;
   wire n_257_76_11572;
   wire n_257_76_11573;
   wire n_257_76_11574;
   wire n_257_76_11575;
   wire n_257_76_11576;
   wire n_257_76_11577;
   wire n_257_76_11578;
   wire n_257_76_11579;
   wire n_257_76_11580;
   wire n_257_76_11581;
   wire n_257_76_11582;
   wire n_257_76_11583;
   wire n_257_76_11584;
   wire n_257_76_11585;
   wire n_257_76_11586;
   wire n_257_76_11587;
   wire n_257_76_11588;
   wire n_257_76_11589;
   wire n_257_76_11590;
   wire n_257_76_11591;
   wire n_257_76_11592;
   wire n_257_76_11593;
   wire n_257_76_11594;
   wire n_257_76_11595;
   wire n_257_76_11596;
   wire n_257_76_11597;
   wire n_257_76_11598;
   wire n_257_76_11599;
   wire n_257_76_11600;
   wire n_257_76_11601;
   wire n_257_76_11602;
   wire n_257_76_11603;
   wire n_257_76_11604;
   wire n_257_76_11605;
   wire n_257_76_11606;
   wire n_257_76_11607;
   wire n_257_76_11608;
   wire n_257_76_11609;
   wire n_257_76_11610;
   wire n_257_76_11611;
   wire n_257_76_11612;
   wire n_257_76_11613;
   wire n_257_76_11614;
   wire n_257_76_11615;
   wire n_257_76_11616;
   wire n_257_76_11617;
   wire n_257_76_11618;
   wire n_257_76_11619;
   wire n_257_76_11620;
   wire n_257_76_11621;
   wire n_257_76_11622;
   wire n_257_76_11623;
   wire n_257_76_11624;
   wire n_257_76_11625;
   wire n_257_76_11626;
   wire n_257_76_11627;
   wire n_257_76_11628;
   wire n_257_76_11629;
   wire n_257_76_11630;
   wire n_257_76_11631;
   wire n_257_76_11632;
   wire n_257_76_11633;
   wire n_257_76_11634;
   wire n_257_76_11635;
   wire n_257_76_11636;
   wire n_257_76_11637;
   wire n_257_76_11638;
   wire n_257_76_11639;
   wire n_257_76_11640;
   wire n_257_76_11641;
   wire n_257_76_11642;
   wire n_257_76_11643;
   wire n_257_76_11644;
   wire n_257_76_11645;
   wire n_257_76_11646;
   wire n_257_76_11647;
   wire n_257_76_11648;
   wire n_257_76_11649;
   wire n_257_76_11650;
   wire n_257_76_11651;
   wire n_257_76_11652;
   wire n_257_76_11653;
   wire n_257_76_11654;
   wire n_257_76_11655;
   wire n_257_76_11656;
   wire n_257_76_11657;
   wire n_257_76_11658;
   wire n_257_76_11659;
   wire n_257_76_11660;
   wire n_257_76_11661;
   wire n_257_76_11662;
   wire n_257_76_11663;
   wire n_257_76_11664;
   wire n_257_76_11665;
   wire n_257_76_11666;
   wire n_257_76_11667;
   wire n_257_76_11668;
   wire n_257_76_11669;
   wire n_257_76_11670;
   wire n_257_76_11671;
   wire n_257_76_11672;
   wire n_257_76_11673;
   wire n_257_76_11674;
   wire n_257_76_11675;
   wire n_257_76_11676;
   wire n_257_76_11677;
   wire n_257_76_11678;
   wire n_257_76_11679;
   wire n_257_76_11680;
   wire n_257_76_11681;
   wire n_257_76_11682;
   wire n_257_76_11683;
   wire n_257_76_11684;
   wire n_257_76_11685;
   wire n_257_76_11686;
   wire n_257_76_11687;
   wire n_257_76_11688;
   wire n_257_76_11689;
   wire n_257_76_11690;
   wire n_257_76_11691;
   wire n_257_76_11692;
   wire n_257_76_11693;
   wire n_257_76_11694;
   wire n_257_76_11695;
   wire n_257_76_11696;
   wire n_257_76_11697;
   wire n_257_76_11698;
   wire n_257_76_11699;
   wire n_257_76_11700;
   wire n_257_76_11701;
   wire n_257_76_11702;
   wire n_257_76_11703;
   wire n_257_76_11704;
   wire n_257_76_11705;
   wire n_257_76_11706;
   wire n_257_76_11707;
   wire n_257_76_11708;
   wire n_257_76_11709;
   wire n_257_76_11710;
   wire n_257_76_11711;
   wire n_257_76_11712;
   wire n_257_76_11713;
   wire n_257_76_11714;
   wire n_257_76_11715;
   wire n_257_76_11716;
   wire n_257_76_11717;
   wire n_257_76_11718;
   wire n_257_76_11719;
   wire n_257_76_11720;
   wire n_257_76_11721;
   wire n_257_76_11722;
   wire n_257_76_11723;
   wire n_257_76_11724;
   wire n_257_76_11725;
   wire n_257_76_11726;
   wire n_257_76_11727;
   wire n_257_76_11728;
   wire n_257_76_11729;
   wire n_257_76_11730;
   wire n_257_76_11731;
   wire n_257_76_11732;
   wire n_257_76_11733;
   wire n_257_76_11734;
   wire n_257_76_11735;
   wire n_257_76_11736;
   wire n_257_76_11737;
   wire n_257_76_11738;
   wire n_257_76_11739;
   wire n_257_76_11740;
   wire n_257_76_11741;
   wire n_257_76_11742;
   wire n_257_76_11743;
   wire n_257_76_11744;
   wire n_257_76_11745;
   wire n_257_76_11746;
   wire n_257_76_11747;
   wire n_257_76_11748;
   wire n_257_76_11749;
   wire n_257_76_11750;
   wire n_257_76_11751;
   wire n_257_76_11752;
   wire n_257_76_11753;
   wire n_257_76_11754;
   wire n_257_76_11755;
   wire n_257_76_11756;
   wire n_257_76_11757;
   wire n_257_76_11758;
   wire n_257_76_11759;
   wire n_257_76_11760;
   wire n_257_76_11761;
   wire n_257_76_11762;
   wire n_257_76_11763;
   wire n_257_76_11764;
   wire n_257_76_11765;
   wire n_257_76_11766;
   wire n_257_76_11767;
   wire n_257_76_11768;
   wire n_257_76_11769;
   wire n_257_76_11770;
   wire n_257_76_11771;
   wire n_257_76_11772;
   wire n_257_76_11773;
   wire n_257_76_11774;
   wire n_257_76_11775;
   wire n_257_76_11776;
   wire n_257_76_11777;
   wire n_257_76_11778;
   wire n_257_76_11779;
   wire n_257_76_11780;
   wire n_257_76_11781;
   wire n_257_76_11782;
   wire n_257_76_11783;
   wire n_257_76_11784;
   wire n_257_76_11785;
   wire n_257_76_11786;
   wire n_257_76_11787;
   wire n_257_76_11788;
   wire n_257_76_11789;
   wire n_257_76_11790;
   wire n_257_76_11791;
   wire n_257_76_11792;
   wire n_257_76_11793;
   wire n_257_76_11794;
   wire n_257_76_11795;
   wire n_257_76_11796;
   wire n_257_76_11797;
   wire n_257_76_11798;
   wire n_257_76_11799;
   wire n_257_76_11800;
   wire n_257_76_11801;
   wire n_257_76_11802;
   wire n_257_76_11803;
   wire n_257_76_11804;
   wire n_257_76_11805;
   wire n_257_76_11806;
   wire n_257_76_11807;
   wire n_257_76_11808;
   wire n_257_76_11809;
   wire n_257_76_11810;
   wire n_257_76_11811;
   wire n_257_76_11812;
   wire n_257_76_11813;
   wire n_257_76_11814;
   wire n_257_76_11815;
   wire n_257_76_11816;
   wire n_257_76_11817;
   wire n_257_76_11818;
   wire n_257_76_11819;
   wire n_257_76_11820;
   wire n_257_76_11821;
   wire n_257_76_11822;
   wire n_257_76_11823;
   wire n_257_76_11824;
   wire n_257_76_11825;
   wire n_257_76_11826;
   wire n_257_76_11827;
   wire n_257_76_11828;
   wire n_257_76_11829;
   wire n_257_76_11830;
   wire n_257_76_11831;
   wire n_257_76_11832;
   wire n_257_76_11833;
   wire n_257_76_11834;
   wire n_257_76_11835;
   wire n_257_76_11836;
   wire n_257_76_11837;
   wire n_257_76_11838;
   wire n_257_76_11839;
   wire n_257_76_11840;
   wire n_257_76_11841;
   wire n_257_76_11842;
   wire n_257_76_11843;
   wire n_257_76_11844;
   wire n_257_76_11845;
   wire n_257_76_11846;
   wire n_257_76_11847;
   wire n_257_76_11848;
   wire n_257_76_11849;
   wire n_257_76_11850;
   wire n_257_76_11851;
   wire n_257_76_11852;
   wire n_257_76_11853;
   wire n_257_76_11854;
   wire n_257_76_11855;
   wire n_257_76_11856;
   wire n_257_76_11857;
   wire n_257_76_11858;
   wire n_257_76_11859;
   wire n_257_76_11860;
   wire n_257_76_11861;
   wire n_257_76_11862;
   wire n_257_76_11863;
   wire n_257_76_11864;
   wire n_257_76_11865;
   wire n_257_76_11866;
   wire n_257_76_11867;
   wire n_257_76_11868;
   wire n_257_76_11869;
   wire n_257_76_11870;
   wire n_257_76_11871;
   wire n_257_76_11872;
   wire n_257_76_11873;
   wire n_257_76_11874;
   wire n_257_76_11875;
   wire n_257_76_11876;
   wire n_257_76_11877;
   wire n_257_76_11878;
   wire n_257_76_11879;
   wire n_257_76_11880;
   wire n_257_76_11881;
   wire n_257_76_11882;
   wire n_257_76_11883;
   wire n_257_76_11884;
   wire n_257_76_11885;
   wire n_257_76_11886;
   wire n_257_76_11887;
   wire n_257_76_11888;
   wire n_257_76_11889;
   wire n_257_76_11890;
   wire n_257_76_11891;
   wire n_257_76_11892;
   wire n_257_76_11893;
   wire n_257_76_11894;
   wire n_257_76_11895;
   wire n_257_76_11896;
   wire n_257_76_11897;
   wire n_257_76_11898;
   wire n_257_76_11899;
   wire n_257_76_11900;
   wire n_257_76_11901;
   wire n_257_76_11902;
   wire n_257_76_11903;
   wire n_257_76_11904;
   wire n_257_76_11905;
   wire n_257_76_11906;
   wire n_257_76_11907;
   wire n_257_76_11908;
   wire n_257_76_11909;
   wire n_257_76_11910;
   wire n_257_76_11911;
   wire n_257_76_11912;
   wire n_257_76_11913;
   wire n_257_76_11914;
   wire n_257_76_11915;
   wire n_257_76_11916;
   wire n_257_76_11917;
   wire n_257_76_11918;
   wire n_257_76_11919;
   wire n_257_76_11920;
   wire n_257_76_11921;
   wire n_257_76_11922;
   wire n_257_76_11923;
   wire n_257_76_11924;
   wire n_257_76_11925;
   wire n_257_76_11926;
   wire n_257_76_11927;
   wire n_257_76_11928;
   wire n_257_76_11929;
   wire n_257_76_11930;
   wire n_257_76_11931;
   wire n_257_76_11932;
   wire n_257_76_11933;
   wire n_257_76_11934;
   wire n_257_76_11935;
   wire n_257_76_11936;
   wire n_257_76_11937;
   wire n_257_76_11938;
   wire n_257_76_11939;
   wire n_257_76_11940;
   wire n_257_76_11941;
   wire n_257_76_11942;
   wire n_257_76_11943;
   wire n_257_76_11944;
   wire n_257_76_11945;
   wire n_257_76_11946;
   wire n_257_76_11947;
   wire n_257_76_11948;
   wire n_257_76_11949;
   wire n_257_76_11950;
   wire n_257_76_11951;
   wire n_257_76_11952;
   wire n_257_76_11953;
   wire n_257_76_11954;
   wire n_257_76_11955;
   wire n_257_76_11956;
   wire n_257_76_11957;
   wire n_257_76_11958;
   wire n_257_76_11959;
   wire n_257_76_11960;
   wire n_257_76_11961;
   wire n_257_76_11962;
   wire n_257_76_11963;
   wire n_257_76_11964;
   wire n_257_76_11965;
   wire n_257_76_11966;
   wire n_257_76_11967;
   wire n_257_76_11968;
   wire n_257_76_11969;
   wire n_257_76_11970;
   wire n_257_76_11971;
   wire n_257_76_11972;
   wire n_257_76_11973;
   wire n_257_76_11974;
   wire n_257_76_11975;
   wire n_257_76_11976;
   wire n_257_76_11977;
   wire n_257_76_11978;
   wire n_257_76_11979;
   wire n_257_76_11980;
   wire n_257_76_11981;
   wire n_257_76_11982;
   wire n_257_76_11983;
   wire n_257_76_11984;
   wire n_257_76_11985;
   wire n_257_76_11986;
   wire n_257_76_11987;
   wire n_257_76_11988;
   wire n_257_76_11989;
   wire n_257_76_11990;
   wire n_257_76_11991;
   wire n_257_76_11992;
   wire n_257_76_11993;
   wire n_257_76_11994;
   wire n_257_76_11995;
   wire n_257_76_11996;
   wire n_257_76_11997;
   wire n_257_76_11998;
   wire n_257_76_11999;
   wire n_257_76_12000;
   wire n_257_76_12001;
   wire n_257_76_12002;
   wire n_257_76_12003;
   wire n_257_76_12004;
   wire n_257_76_12005;
   wire n_257_76_12006;
   wire n_257_76_12007;
   wire n_257_76_12008;
   wire n_257_76_12009;
   wire n_257_76_12010;
   wire n_257_76_12011;
   wire n_257_76_12012;
   wire n_257_76_12013;
   wire n_257_76_12014;
   wire n_257_76_12015;
   wire n_257_76_12016;
   wire n_257_76_12017;
   wire n_257_76_12018;
   wire n_257_76_12019;
   wire n_257_76_12020;
   wire n_257_76_12021;
   wire n_257_76_12022;
   wire n_257_76_12023;
   wire n_257_76_12024;
   wire n_257_76_12025;
   wire n_257_76_12026;
   wire n_257_76_12027;
   wire n_257_76_12028;
   wire n_257_76_12029;
   wire n_257_76_12030;
   wire n_257_76_12031;
   wire n_257_76_12032;
   wire n_257_76_12033;
   wire n_257_76_12034;
   wire n_257_76_12035;
   wire n_257_76_12036;
   wire n_257_76_12037;
   wire n_257_76_12038;
   wire n_257_76_12039;
   wire n_257_76_12040;
   wire n_257_76_12041;
   wire n_257_76_12042;
   wire n_257_76_12043;
   wire n_257_76_12044;
   wire n_257_76_12045;
   wire n_257_76_12046;
   wire n_257_76_12047;
   wire n_257_76_12048;
   wire n_257_76_12049;
   wire n_257_76_12050;
   wire n_257_76_12051;
   wire n_257_76_12052;
   wire n_257_76_12053;
   wire n_257_76_12054;
   wire n_257_76_12055;
   wire n_257_76_12056;
   wire n_257_76_12057;
   wire n_257_76_12058;
   wire n_257_76_12059;
   wire n_257_76_12060;
   wire n_257_76_12061;
   wire n_257_76_12062;
   wire n_257_76_12063;
   wire n_257_76_12064;
   wire n_257_76_12065;
   wire n_257_76_12066;
   wire n_257_76_12067;
   wire n_257_76_12068;
   wire n_257_76_12069;
   wire n_257_76_12070;
   wire n_257_76_12071;
   wire n_257_76_12072;
   wire n_257_76_12073;
   wire n_257_76_12074;
   wire n_257_76_12075;
   wire n_257_76_12076;
   wire n_257_76_12077;
   wire n_257_76_12078;
   wire n_257_76_12079;
   wire n_257_76_12080;
   wire n_257_76_12081;
   wire n_257_76_12082;
   wire n_257_76_12083;
   wire n_257_76_12084;
   wire n_257_76_12085;
   wire n_257_76_12086;
   wire n_257_76_12087;
   wire n_257_76_12088;
   wire n_257_76_12089;
   wire n_257_76_12090;
   wire n_257_76_12091;
   wire n_257_76_12092;
   wire n_257_76_12093;
   wire n_257_76_12094;
   wire n_257_76_12095;
   wire n_257_76_12096;
   wire n_257_76_12097;
   wire n_257_76_12098;
   wire n_257_76_12099;
   wire n_257_76_12100;
   wire n_257_76_12101;
   wire n_257_76_12102;
   wire n_257_76_12103;
   wire n_257_76_12104;
   wire n_257_76_12105;
   wire n_257_76_12106;
   wire n_257_76_12107;
   wire n_257_76_12108;
   wire n_257_76_12109;
   wire n_257_76_12110;
   wire n_257_76_12111;
   wire n_257_76_12112;
   wire n_257_76_12113;
   wire n_257_76_12114;
   wire n_257_76_12115;
   wire n_257_76_12116;
   wire n_257_76_12117;
   wire n_257_76_12118;
   wire n_257_76_12119;
   wire n_257_76_12120;
   wire n_257_76_12121;
   wire n_257_76_12122;
   wire n_257_76_12123;
   wire n_257_76_12124;
   wire n_257_76_12125;
   wire n_257_76_12126;
   wire n_257_76_12127;
   wire n_257_76_12128;
   wire n_257_76_12129;
   wire n_257_76_12130;
   wire n_257_76_12131;
   wire n_257_76_12132;
   wire n_257_76_12133;
   wire n_257_76_12134;
   wire n_257_76_12135;
   wire n_257_76_12136;
   wire n_257_76_12137;
   wire n_257_76_12138;
   wire n_257_76_12139;
   wire n_257_76_12140;
   wire n_257_76_12141;
   wire n_257_76_12142;
   wire n_257_76_12143;
   wire n_257_76_12144;
   wire n_257_76_12145;
   wire n_257_76_12146;
   wire n_257_76_12147;
   wire n_257_76_12148;
   wire n_257_76_12149;
   wire n_257_76_12150;
   wire n_257_76_12151;
   wire n_257_76_12152;
   wire n_257_76_12153;
   wire n_257_76_12154;
   wire n_257_76_12155;
   wire n_257_76_12156;
   wire n_257_76_12157;
   wire n_257_76_12158;
   wire n_257_76_12159;
   wire n_257_76_12160;
   wire n_257_76_12161;
   wire n_257_76_12162;
   wire n_257_76_12163;
   wire n_257_76_12164;
   wire n_257_76_12165;
   wire n_257_76_12166;
   wire n_257_76_12167;
   wire n_257_76_12168;
   wire n_257_76_12169;
   wire n_257_76_12170;
   wire n_257_76_12171;
   wire n_257_76_12172;
   wire n_257_76_12173;
   wire n_257_76_12174;
   wire n_257_76_12175;
   wire n_257_76_12176;
   wire n_257_76_12177;
   wire n_257_76_12178;
   wire n_257_76_12179;
   wire n_257_76_12180;
   wire n_257_76_12181;
   wire n_257_76_12182;
   wire n_257_76_12183;
   wire n_257_76_12184;
   wire n_257_76_12185;
   wire n_257_76_12186;
   wire n_257_76_12187;
   wire n_257_76_12188;
   wire n_257_76_12189;
   wire n_257_76_12190;
   wire n_257_76_12191;
   wire n_257_76_12192;
   wire n_257_76_12193;
   wire n_257_76_12194;
   wire n_257_76_12195;
   wire n_257_76_12196;
   wire n_257_76_12197;
   wire n_257_76_12198;
   wire n_257_76_12199;
   wire n_257_76_12200;
   wire n_257_76_12201;
   wire n_257_76_12202;
   wire n_257_76_12203;
   wire n_257_76_12204;
   wire n_257_76_12205;
   wire n_257_76_12206;
   wire n_257_76_12207;
   wire n_257_76_12208;
   wire n_257_76_12209;
   wire n_257_76_12210;
   wire n_257_76_12211;
   wire n_257_76_12212;
   wire n_257_76_12213;
   wire n_257_76_12214;
   wire n_257_76_12215;
   wire n_257_76_12216;
   wire n_257_76_12217;
   wire n_257_76_12218;
   wire n_257_76_12219;
   wire n_257_76_12220;
   wire n_257_76_12221;
   wire n_257_76_12222;
   wire n_257_76_12223;
   wire n_257_76_12224;
   wire n_257_76_12225;
   wire n_257_76_12226;
   wire n_257_76_12227;
   wire n_257_76_12228;
   wire n_257_76_12229;
   wire n_257_76_12230;
   wire n_257_76_12231;
   wire n_257_76_12232;
   wire n_257_76_12233;
   wire n_257_76_12234;
   wire n_257_76_12235;
   wire n_257_76_12236;
   wire n_257_76_12237;
   wire n_257_76_12238;
   wire n_257_76_12239;
   wire n_257_76_12240;
   wire n_257_76_12241;
   wire n_257_76_12242;
   wire n_257_76_12243;
   wire n_257_76_12244;
   wire n_257_76_12245;
   wire n_257_76_12246;
   wire n_257_76_12247;
   wire n_257_76_12248;
   wire n_257_76_12249;
   wire n_257_76_12250;
   wire n_257_76_12251;
   wire n_257_76_12252;
   wire n_257_76_12253;
   wire n_257_76_12254;
   wire n_257_76_12255;
   wire n_257_76_12256;
   wire n_257_76_12257;
   wire n_257_76_12258;
   wire n_257_76_12259;
   wire n_257_76_12260;
   wire n_257_76_12261;
   wire n_257_76_12262;
   wire n_257_76_12263;
   wire n_257_76_12264;
   wire n_257_76_12265;
   wire n_257_76_12266;
   wire n_257_76_12267;
   wire n_257_76_12268;
   wire n_257_76_12269;
   wire n_257_76_12270;
   wire n_257_76_12271;
   wire n_257_76_12272;
   wire n_257_76_12273;
   wire n_257_76_12274;
   wire n_257_76_12275;
   wire n_257_76_12276;
   wire n_257_76_12277;
   wire n_257_76_12278;
   wire n_257_76_12279;
   wire n_257_76_12280;
   wire n_257_76_12281;
   wire n_257_76_12282;
   wire n_257_76_12283;
   wire n_257_76_12284;
   wire n_257_76_12285;
   wire n_257_76_12286;
   wire n_257_76_12287;
   wire n_257_76_12288;
   wire n_257_76_12289;
   wire n_257_76_12290;
   wire n_257_76_12291;
   wire n_257_76_12292;
   wire n_257_76_12293;
   wire n_257_76_12294;
   wire n_257_76_12295;
   wire n_257_76_12296;
   wire n_257_76_12297;
   wire n_257_76_12298;
   wire n_257_76_12299;
   wire n_257_76_12300;
   wire n_257_76_12301;
   wire n_257_76_12302;
   wire n_257_76_12303;
   wire n_257_76_12304;
   wire n_257_76_12305;
   wire n_257_76_12306;
   wire n_257_76_12307;
   wire n_257_76_12308;
   wire n_257_76_12309;
   wire n_257_76_12310;
   wire n_257_76_12311;
   wire n_257_76_12312;
   wire n_257_76_12313;
   wire n_257_76_12314;
   wire n_257_76_12315;
   wire n_257_76_12316;
   wire n_257_76_12317;
   wire n_257_76_12318;
   wire n_257_76_12319;
   wire n_257_76_12320;
   wire n_257_76_12321;
   wire n_257_76_12322;
   wire n_257_76_12323;
   wire n_257_76_12324;
   wire n_257_76_12325;
   wire n_257_76_12326;
   wire n_257_76_12327;
   wire n_257_76_12328;
   wire n_257_76_12329;
   wire n_257_76_12330;
   wire n_257_76_12331;
   wire n_257_76_12332;
   wire n_257_76_12333;
   wire n_257_76_12334;
   wire n_257_76_12335;
   wire n_257_76_12336;
   wire n_257_76_12337;
   wire n_257_76_12338;
   wire n_257_76_12339;
   wire n_257_76_12340;
   wire n_257_76_12341;
   wire n_257_76_12342;
   wire n_257_76_12343;
   wire n_257_76_12344;
   wire n_257_76_12345;
   wire n_257_76_12346;
   wire n_257_76_12347;
   wire n_257_76_12348;
   wire n_257_76_12349;
   wire n_257_76_12350;
   wire n_257_76_12351;
   wire n_257_76_12352;
   wire n_257_76_12353;
   wire n_257_76_12354;
   wire n_257_76_12355;
   wire n_257_76_12356;
   wire n_257_76_12357;
   wire n_257_76_12358;
   wire n_257_76_12359;
   wire n_257_76_12360;
   wire n_257_76_12361;
   wire n_257_76_12362;
   wire n_257_76_12363;
   wire n_257_76_12364;
   wire n_257_76_12365;
   wire n_257_76_12366;
   wire n_257_76_12367;
   wire n_257_76_12368;
   wire n_257_76_12369;
   wire n_257_76_12370;
   wire n_257_76_12371;
   wire n_257_76_12372;
   wire n_257_76_12373;
   wire n_257_76_12374;
   wire n_257_76_12375;
   wire n_257_76_12376;
   wire n_257_76_12377;
   wire n_257_76_12378;
   wire n_257_76_12379;
   wire n_257_76_12380;
   wire n_257_76_12381;
   wire n_257_76_12382;
   wire n_257_76_12383;
   wire n_257_76_12384;
   wire n_257_76_12385;
   wire n_257_76_12386;
   wire n_257_76_12387;
   wire n_257_76_12388;
   wire n_257_76_12389;
   wire n_257_76_12390;
   wire n_257_76_12391;
   wire n_257_76_12392;
   wire n_257_76_12393;
   wire n_257_76_12394;
   wire n_257_76_12395;
   wire n_257_76_12396;
   wire n_257_76_12397;
   wire n_257_76_12398;
   wire n_257_76_12399;
   wire n_257_76_12400;
   wire n_257_76_12401;
   wire n_257_76_12402;
   wire n_257_76_12403;
   wire n_257_76_12404;
   wire n_257_76_12405;
   wire n_257_76_12406;
   wire n_257_76_12407;
   wire n_257_76_12408;
   wire n_257_76_12409;
   wire n_257_76_12410;
   wire n_257_76_12411;
   wire n_257_76_12412;
   wire n_257_76_12413;
   wire n_257_76_12414;
   wire n_257_76_12415;
   wire n_257_76_12416;
   wire n_257_76_12417;
   wire n_257_76_12418;
   wire n_257_76_12419;
   wire n_257_76_12420;
   wire n_257_76_12421;
   wire n_257_76_12422;
   wire n_257_76_12423;
   wire n_257_76_12424;
   wire n_257_76_12425;
   wire n_257_76_12426;
   wire n_257_76_12427;
   wire n_257_76_12428;
   wire n_257_76_12429;
   wire n_257_76_12430;
   wire n_257_76_12431;
   wire n_257_76_12432;
   wire n_257_76_12433;
   wire n_257_76_12434;
   wire n_257_76_12435;
   wire n_257_76_12436;
   wire n_257_76_12437;
   wire n_257_76_12438;
   wire n_257_76_12439;
   wire n_257_76_12440;
   wire n_257_76_12441;
   wire n_257_76_12442;
   wire n_257_76_12443;
   wire n_257_76_12444;
   wire n_257_76_12445;
   wire n_257_76_12446;
   wire n_257_76_12447;
   wire n_257_76_12448;
   wire n_257_76_12449;
   wire n_257_76_12450;
   wire n_257_76_12451;
   wire n_257_76_12452;
   wire n_257_76_12453;
   wire n_257_76_12454;
   wire n_257_76_12455;
   wire n_257_76_12456;
   wire n_257_76_12457;
   wire n_257_76_12458;
   wire n_257_76_12459;
   wire n_257_76_12460;
   wire n_257_76_12461;
   wire n_257_76_12462;
   wire n_257_76_12463;
   wire n_257_76_12464;
   wire n_257_76_12465;
   wire n_257_76_12466;
   wire n_257_76_12467;
   wire n_257_76_12468;
   wire n_257_76_12469;
   wire n_257_76_12470;
   wire n_257_76_12471;
   wire n_257_76_12472;
   wire n_257_76_12473;
   wire n_257_76_12474;
   wire n_257_76_12475;
   wire n_257_76_12476;
   wire n_257_76_12477;
   wire n_257_76_12478;
   wire n_257_76_12479;
   wire n_257_76_12480;
   wire n_257_76_12481;
   wire n_257_76_12482;
   wire n_257_76_12483;
   wire n_257_76_12484;
   wire n_257_76_12485;
   wire n_257_76_12486;
   wire n_257_76_12487;
   wire n_257_76_12488;
   wire n_257_76_12489;
   wire n_257_76_12490;
   wire n_257_76_12491;
   wire n_257_76_12492;
   wire n_257_76_12493;
   wire n_257_76_12494;
   wire n_257_76_12495;
   wire n_257_76_12496;
   wire n_257_76_12497;
   wire n_257_76_12498;
   wire n_257_76_12499;
   wire n_257_76_12500;
   wire n_257_76_12501;
   wire n_257_76_12502;
   wire n_257_76_12503;
   wire n_257_76_12504;
   wire n_257_76_12505;
   wire n_257_76_12506;
   wire n_257_76_12507;
   wire n_257_76_12508;
   wire n_257_76_12509;
   wire n_257_76_12510;
   wire n_257_76_12511;
   wire n_257_76_12512;
   wire n_257_76_12513;
   wire n_257_76_12514;
   wire n_257_76_12515;
   wire n_257_76_12516;
   wire n_257_76_12517;
   wire n_257_76_12518;
   wire n_257_76_12519;
   wire n_257_76_12520;
   wire n_257_76_12521;
   wire n_257_76_12522;
   wire n_257_76_12523;
   wire n_257_76_12524;
   wire n_257_76_12525;
   wire n_257_76_12526;
   wire n_257_76_12527;
   wire n_257_76_12528;
   wire n_257_76_12529;
   wire n_257_76_12530;
   wire n_257_76_12531;
   wire n_257_76_12532;
   wire n_257_76_12533;
   wire n_257_76_12534;
   wire n_257_76_12535;
   wire n_257_76_12536;
   wire n_257_76_12537;
   wire n_257_76_12538;
   wire n_257_76_12539;
   wire n_257_76_12540;
   wire n_257_76_12541;
   wire n_257_76_12542;
   wire n_257_76_12543;
   wire n_257_76_12544;
   wire n_257_76_12545;
   wire n_257_76_12546;
   wire n_257_76_12547;
   wire n_257_76_12548;
   wire n_257_76_12549;
   wire n_257_76_12550;
   wire n_257_76_12551;
   wire n_257_76_12552;
   wire n_257_76_12553;
   wire n_257_76_12554;
   wire n_257_76_12555;
   wire n_257_76_12556;
   wire n_257_76_12557;
   wire n_257_76_12558;
   wire n_257_76_12559;
   wire n_257_76_12560;
   wire n_257_76_12561;
   wire n_257_76_12562;
   wire n_257_76_12563;
   wire n_257_76_12564;
   wire n_257_76_12565;
   wire n_257_76_12566;
   wire n_257_76_12567;
   wire n_257_76_12568;
   wire n_257_76_12569;
   wire n_257_76_12570;
   wire n_257_76_12571;
   wire n_257_76_12572;
   wire n_257_76_12573;
   wire n_257_76_12574;
   wire n_257_76_12575;
   wire n_257_76_12576;
   wire n_257_76_12577;
   wire n_257_76_12578;
   wire n_257_76_12579;
   wire n_257_76_12580;
   wire n_257_76_12581;
   wire n_257_76_12582;
   wire n_257_76_12583;
   wire n_257_76_12584;
   wire n_257_76_12585;
   wire n_257_76_12586;
   wire n_257_76_12587;
   wire n_257_76_12588;
   wire n_257_76_12589;
   wire n_257_76_12590;
   wire n_257_76_12591;
   wire n_257_76_12592;
   wire n_257_76_12593;
   wire n_257_76_12594;
   wire n_257_76_12595;
   wire n_257_76_12596;
   wire n_257_76_12597;
   wire n_257_76_12598;
   wire n_257_76_12599;
   wire n_257_76_12600;
   wire n_257_76_12601;
   wire n_257_76_12602;
   wire n_257_76_12603;
   wire n_257_76_12604;
   wire n_257_76_12605;
   wire n_257_76_12606;
   wire n_257_76_12607;
   wire n_257_76_12608;
   wire n_257_76_12609;
   wire n_257_76_12610;
   wire n_257_76_12611;
   wire n_257_76_12612;
   wire n_257_76_12613;
   wire n_257_76_12614;
   wire n_257_76_12615;
   wire n_257_76_12616;
   wire n_257_76_12617;
   wire n_257_76_12618;
   wire n_257_76_12619;
   wire n_257_76_12620;
   wire n_257_76_12621;
   wire n_257_76_12622;
   wire n_257_76_12623;
   wire n_257_76_12624;
   wire n_257_76_12625;
   wire n_257_76_12626;
   wire n_257_76_12627;
   wire n_257_76_12628;
   wire n_257_76_12629;
   wire n_257_76_12630;
   wire n_257_76_12631;
   wire n_257_76_12632;
   wire n_257_76_12633;
   wire n_257_76_12634;
   wire n_257_76_12635;
   wire n_257_76_12636;
   wire n_257_76_12637;
   wire n_257_76_12638;
   wire n_257_76_12639;
   wire n_257_76_12640;
   wire n_257_76_12641;
   wire n_257_76_12642;
   wire n_257_76_12643;
   wire n_257_76_12644;
   wire n_257_76_12645;
   wire n_257_76_12646;
   wire n_257_76_12647;
   wire n_257_76_12648;
   wire n_257_76_12649;
   wire n_257_76_12650;
   wire n_257_76_12651;
   wire n_257_76_12652;
   wire n_257_76_12653;
   wire n_257_76_12654;
   wire n_257_76_12655;
   wire n_257_76_12656;
   wire n_257_76_12657;
   wire n_257_76_12658;
   wire n_257_76_12659;
   wire n_257_76_12660;
   wire n_257_76_12661;
   wire n_257_76_12662;
   wire n_257_76_12663;
   wire n_257_76_12664;
   wire n_257_76_12665;
   wire n_257_76_12666;
   wire n_257_76_12667;
   wire n_257_76_12668;
   wire n_257_76_12669;
   wire n_257_76_12670;
   wire n_257_76_12671;
   wire n_257_76_12672;
   wire n_257_76_12673;
   wire n_257_76_12674;
   wire n_257_76_12675;
   wire n_257_76_12676;
   wire n_257_76_12677;
   wire n_257_76_12678;
   wire n_257_76_12679;
   wire n_257_76_12680;
   wire n_257_76_12681;
   wire n_257_76_12682;
   wire n_257_76_12683;
   wire n_257_76_12684;
   wire n_257_76_12685;
   wire n_257_76_12686;
   wire n_257_76_12687;
   wire n_257_76_12688;
   wire n_257_76_12689;
   wire n_257_76_12690;
   wire n_257_76_12691;
   wire n_257_76_12692;
   wire n_257_76_12693;
   wire n_257_76_12694;
   wire n_257_76_12695;
   wire n_257_76_12696;
   wire n_257_76_12697;
   wire n_257_76_12698;
   wire n_257_76_12699;
   wire n_257_76_12700;
   wire n_257_76_12701;
   wire n_257_76_12702;
   wire n_257_76_12703;
   wire n_257_76_12704;
   wire n_257_76_12705;
   wire n_257_76_12706;
   wire n_257_76_12707;
   wire n_257_76_12708;
   wire n_257_76_12709;
   wire n_257_76_12710;
   wire n_257_76_12711;
   wire n_257_76_12712;
   wire n_257_76_12713;
   wire n_257_76_12714;
   wire n_257_76_12715;
   wire n_257_76_12716;
   wire n_257_76_12717;
   wire n_257_76_12718;
   wire n_257_76_12719;
   wire n_257_76_12720;
   wire n_257_76_12721;
   wire n_257_76_12722;
   wire n_257_76_12723;
   wire n_257_76_12724;
   wire n_257_76_12725;
   wire n_257_76_12726;
   wire n_257_76_12727;
   wire n_257_76_12728;
   wire n_257_76_12729;
   wire n_257_76_12730;
   wire n_257_76_12731;
   wire n_257_76_12732;
   wire n_257_76_12733;
   wire n_257_76_12734;
   wire n_257_76_12735;
   wire n_257_76_12736;
   wire n_257_76_12737;
   wire n_257_76_12738;
   wire n_257_76_12739;
   wire n_257_76_12740;
   wire n_257_76_12741;
   wire n_257_76_12742;
   wire n_257_76_12743;
   wire n_257_76_12744;
   wire n_257_76_12745;
   wire n_257_76_12746;
   wire n_257_76_12747;
   wire n_257_76_12748;
   wire n_257_76_12749;
   wire n_257_76_12750;
   wire n_257_76_12751;
   wire n_257_76_12752;
   wire n_257_76_12753;
   wire n_257_76_12754;
   wire n_257_76_12755;
   wire n_257_76_12756;
   wire n_257_76_12757;
   wire n_257_76_12758;
   wire n_257_76_12759;
   wire n_257_76_12760;
   wire n_257_76_12761;
   wire n_257_76_12762;
   wire n_257_76_12763;
   wire n_257_76_12764;
   wire n_257_76_12765;
   wire n_257_76_12766;
   wire n_257_76_12767;
   wire n_257_76_12768;
   wire n_257_76_12769;
   wire n_257_76_12770;
   wire n_257_76_12771;
   wire n_257_76_12772;
   wire n_257_76_12773;
   wire n_257_76_12774;
   wire n_257_76_12775;
   wire n_257_76_12776;
   wire n_257_76_12777;
   wire n_257_76_12778;
   wire n_257_76_12779;
   wire n_257_76_12780;
   wire n_257_76_12781;
   wire n_257_76_12782;
   wire n_257_76_12783;
   wire n_257_76_12784;
   wire n_257_76_12785;
   wire n_257_76_12786;
   wire n_257_76_12787;
   wire n_257_76_12788;
   wire n_257_76_12789;
   wire n_257_76_12790;
   wire n_257_76_12791;
   wire n_257_76_12792;
   wire n_257_76_12793;
   wire n_257_76_12794;
   wire n_257_76_12795;
   wire n_257_76_12796;
   wire n_257_76_12797;
   wire n_257_76_12798;
   wire n_257_76_12799;
   wire n_257_76_12800;
   wire n_257_76_12801;
   wire n_257_76_12802;
   wire n_257_76_12803;
   wire n_257_76_12804;
   wire n_257_76_12805;
   wire n_257_76_12806;
   wire n_257_76_12807;
   wire n_257_76_12808;
   wire n_257_76_12809;
   wire n_257_76_12810;
   wire n_257_76_12811;
   wire n_257_76_12812;
   wire n_257_76_12813;
   wire n_257_76_12814;
   wire n_257_76_12815;
   wire n_257_76_12816;
   wire n_257_76_12817;
   wire n_257_76_12818;
   wire n_257_76_12819;
   wire n_257_76_12820;
   wire n_257_76_12821;
   wire n_257_76_12822;
   wire n_257_76_12823;
   wire n_257_76_12824;
   wire n_257_76_12825;
   wire n_257_76_12826;
   wire n_257_76_12827;
   wire n_257_76_12828;
   wire n_257_76_12829;
   wire n_257_76_12830;
   wire n_257_76_12831;
   wire n_257_76_12832;
   wire n_257_76_12833;
   wire n_257_76_12834;
   wire n_257_76_12835;
   wire n_257_76_12836;
   wire n_257_76_12837;
   wire n_257_76_12838;
   wire n_257_76_12839;
   wire n_257_76_12840;
   wire n_257_76_12841;
   wire n_257_76_12842;
   wire n_257_76_12843;
   wire n_257_76_12844;
   wire n_257_76_12845;
   wire n_257_76_12846;
   wire n_257_76_12847;
   wire n_257_76_12848;
   wire n_257_76_12849;
   wire n_257_76_12850;
   wire n_257_76_12851;
   wire n_257_76_12852;
   wire n_257_76_12853;
   wire n_257_76_12854;
   wire n_257_76_12855;
   wire n_257_76_12856;
   wire n_257_76_12857;
   wire n_257_76_12858;
   wire n_257_76_12859;
   wire n_257_76_12860;
   wire n_257_76_12861;
   wire n_257_76_12862;
   wire n_257_76_12863;
   wire n_257_76_12864;
   wire n_257_76_12865;
   wire n_257_76_12866;
   wire n_257_76_12867;
   wire n_257_76_12868;
   wire n_257_76_12869;
   wire n_257_76_12870;
   wire n_257_76_12871;
   wire n_257_76_12872;
   wire n_257_76_12873;
   wire n_257_76_12874;
   wire n_257_76_12875;
   wire n_257_76_12876;
   wire n_257_76_12877;
   wire n_257_76_12878;
   wire n_257_76_12879;
   wire n_257_76_12880;
   wire n_257_76_12881;
   wire n_257_76_12882;
   wire n_257_76_12883;
   wire n_257_76_12884;
   wire n_257_76_12885;
   wire n_257_76_12886;
   wire n_257_76_12887;
   wire n_257_76_12888;
   wire n_257_76_12889;
   wire n_257_76_12890;
   wire n_257_76_12891;
   wire n_257_76_12892;
   wire n_257_76_12893;
   wire n_257_76_12894;
   wire n_257_76_12895;
   wire n_257_76_12896;
   wire n_257_76_12897;
   wire n_257_76_12898;
   wire n_257_76_12899;
   wire n_257_76_12900;
   wire n_257_76_12901;
   wire n_257_76_12902;
   wire n_257_76_12903;
   wire n_257_76_12904;
   wire n_257_76_12905;
   wire n_257_76_12906;
   wire n_257_76_12907;
   wire n_257_76_12908;
   wire n_257_76_12909;
   wire n_257_76_12910;
   wire n_257_76_12911;
   wire n_257_76_12912;
   wire n_257_76_12913;
   wire n_257_76_12914;
   wire n_257_76_12915;
   wire n_257_76_12916;
   wire n_257_76_12917;
   wire n_257_76_12918;
   wire n_257_76_12919;
   wire n_257_76_12920;
   wire n_257_76_12921;
   wire n_257_76_12922;
   wire n_257_76_12923;
   wire n_257_76_12924;
   wire n_257_76_12925;
   wire n_257_76_12926;
   wire n_257_76_12927;
   wire n_257_76_12928;
   wire n_257_76_12929;
   wire n_257_76_12930;
   wire n_257_76_12931;
   wire n_257_76_12932;
   wire n_257_76_12933;
   wire n_257_76_12934;
   wire n_257_76_12935;
   wire n_257_76_12936;
   wire n_257_76_12937;
   wire n_257_76_12938;
   wire n_257_76_12939;
   wire n_257_76_12940;
   wire n_257_76_12941;
   wire n_257_76_12942;
   wire n_257_76_12943;
   wire n_257_76_12944;
   wire n_257_76_12945;
   wire n_257_76_12946;
   wire n_257_76_12947;
   wire n_257_76_12948;
   wire n_257_76_12949;
   wire n_257_76_12950;
   wire n_257_76_12951;
   wire n_257_76_12952;
   wire n_257_76_12953;
   wire n_257_76_12954;
   wire n_257_76_12955;
   wire n_257_76_12956;
   wire n_257_76_12957;
   wire n_257_76_12958;
   wire n_257_76_12959;
   wire n_257_76_12960;
   wire n_257_76_12961;
   wire n_257_76_12962;
   wire n_257_76_12963;
   wire n_257_76_12964;
   wire n_257_76_12965;
   wire n_257_76_12966;
   wire n_257_76_12967;
   wire n_257_76_12968;
   wire n_257_76_12969;
   wire n_257_76_12970;
   wire n_257_76_12971;
   wire n_257_76_12972;
   wire n_257_76_12973;
   wire n_257_76_12974;
   wire n_257_76_12975;
   wire n_257_76_12976;
   wire n_257_76_12977;
   wire n_257_76_12978;
   wire n_257_76_12979;
   wire n_257_76_12980;
   wire n_257_76_12981;
   wire n_257_76_12982;
   wire n_257_76_12983;
   wire n_257_76_12984;
   wire n_257_76_12985;
   wire n_257_76_12986;
   wire n_257_76_12987;
   wire n_257_76_12988;
   wire n_257_76_12989;
   wire n_257_76_12990;
   wire n_257_76_12991;
   wire n_257_76_12992;
   wire n_257_76_12993;
   wire n_257_76_12994;
   wire n_257_76_12995;
   wire n_257_76_12996;
   wire n_257_76_12997;
   wire n_257_76_12998;
   wire n_257_76_12999;
   wire n_257_76_13000;
   wire n_257_76_13001;
   wire n_257_76_13002;
   wire n_257_76_13003;
   wire n_257_76_13004;
   wire n_257_76_13005;
   wire n_257_76_13006;
   wire n_257_76_13007;
   wire n_257_76_13008;
   wire n_257_76_13009;
   wire n_257_76_13010;
   wire n_257_76_13011;
   wire n_257_76_13012;
   wire n_257_76_13013;
   wire n_257_76_13014;
   wire n_257_76_13015;
   wire n_257_76_13016;
   wire n_257_76_13017;
   wire n_257_76_13018;
   wire n_257_76_13019;
   wire n_257_76_13020;
   wire n_257_76_13021;
   wire n_257_76_13022;
   wire n_257_76_13023;
   wire n_257_76_13024;
   wire n_257_76_13025;
   wire n_257_76_13026;
   wire n_257_76_13027;
   wire n_257_76_13028;
   wire n_257_76_13029;
   wire n_257_76_13030;
   wire n_257_76_13031;
   wire n_257_76_13032;
   wire n_257_76_13033;
   wire n_257_76_13034;
   wire n_257_76_13035;
   wire n_257_76_13036;
   wire n_257_76_13037;
   wire n_257_76_13038;
   wire n_257_76_13039;
   wire n_257_76_13040;
   wire n_257_76_13041;
   wire n_257_76_13042;
   wire n_257_76_13043;
   wire n_257_76_13044;
   wire n_257_76_13045;
   wire n_257_76_13046;
   wire n_257_76_13047;
   wire n_257_76_13048;
   wire n_257_76_13049;
   wire n_257_76_13050;
   wire n_257_76_13051;
   wire n_257_76_13052;
   wire n_257_76_13053;
   wire n_257_76_13054;
   wire n_257_76_13055;
   wire n_257_76_13056;
   wire n_257_76_13057;
   wire n_257_76_13058;
   wire n_257_76_13059;
   wire n_257_76_13060;
   wire n_257_76_13061;
   wire n_257_76_13062;
   wire n_257_76_13063;
   wire n_257_76_13064;
   wire n_257_76_13065;
   wire n_257_76_13066;
   wire n_257_76_13067;
   wire n_257_76_13068;
   wire n_257_76_13069;
   wire n_257_76_13070;
   wire n_257_76_13071;
   wire n_257_76_13072;
   wire n_257_76_13073;
   wire n_257_76_13074;
   wire n_257_76_13075;
   wire n_257_76_13076;
   wire n_257_76_13077;
   wire n_257_76_13078;
   wire n_257_76_13079;
   wire n_257_76_13080;
   wire n_257_76_13081;
   wire n_257_76_13082;
   wire n_257_76_13083;
   wire n_257_76_13084;
   wire n_257_76_13085;
   wire n_257_76_13086;
   wire n_257_76_13087;
   wire n_257_76_13088;
   wire n_257_76_13089;
   wire n_257_76_13090;
   wire n_257_76_13091;
   wire n_257_76_13092;
   wire n_257_76_13093;
   wire n_257_76_13094;
   wire n_257_76_13095;
   wire n_257_76_13096;
   wire n_257_76_13097;
   wire n_257_76_13098;
   wire n_257_76_13099;
   wire n_257_76_13100;
   wire n_257_76_13101;
   wire n_257_76_13102;
   wire n_257_76_13103;
   wire n_257_76_13104;
   wire n_257_76_13105;
   wire n_257_76_13106;
   wire n_257_76_13107;
   wire n_257_76_13108;
   wire n_257_76_13109;
   wire n_257_76_13110;
   wire n_257_76_13111;
   wire n_257_76_13112;
   wire n_257_76_13113;
   wire n_257_76_13114;
   wire n_257_76_13115;
   wire n_257_76_13116;
   wire n_257_76_13117;
   wire n_257_76_13118;
   wire n_257_76_13119;
   wire n_257_76_13120;
   wire n_257_76_13121;
   wire n_257_76_13122;
   wire n_257_76_13123;
   wire n_257_76_13124;
   wire n_257_76_13125;
   wire n_257_76_13126;
   wire n_257_76_13127;
   wire n_257_76_13128;
   wire n_257_76_13129;
   wire n_257_76_13130;
   wire n_257_76_13131;
   wire n_257_76_13132;
   wire n_257_76_13133;
   wire n_257_76_13134;
   wire n_257_76_13135;
   wire n_257_76_13136;
   wire n_257_76_13137;
   wire n_257_76_13138;
   wire n_257_76_13139;
   wire n_257_76_13140;
   wire n_257_76_13141;
   wire n_257_76_13142;
   wire n_257_76_13143;
   wire n_257_76_13144;
   wire n_257_76_13145;
   wire n_257_76_13146;
   wire n_257_76_13147;
   wire n_257_76_13148;
   wire n_257_76_13149;
   wire n_257_76_13150;
   wire n_257_76_13151;
   wire n_257_76_13152;
   wire n_257_76_13153;
   wire n_257_76_13154;
   wire n_257_76_13155;
   wire n_257_76_13156;
   wire n_257_76_13157;
   wire n_257_76_13158;
   wire n_257_76_13159;
   wire n_257_76_13160;
   wire n_257_76_13161;
   wire n_257_76_13162;
   wire n_257_76_13163;
   wire n_257_76_13164;
   wire n_257_76_13165;
   wire n_257_76_13166;
   wire n_257_76_13167;
   wire n_257_76_13168;
   wire n_257_76_13169;
   wire n_257_76_13170;
   wire n_257_76_13171;
   wire n_257_76_13172;
   wire n_257_76_13173;
   wire n_257_76_13174;
   wire n_257_76_13175;
   wire n_257_76_13176;
   wire n_257_76_13177;
   wire n_257_76_13178;
   wire n_257_76_13179;
   wire n_257_76_13180;
   wire n_257_76_13181;
   wire n_257_76_13182;
   wire n_257_76_13183;
   wire n_257_76_13184;
   wire n_257_76_13185;
   wire n_257_76_13186;
   wire n_257_76_13187;
   wire n_257_76_13188;
   wire n_257_76_13189;
   wire n_257_76_13190;
   wire n_257_76_13191;
   wire n_257_76_13192;
   wire n_257_76_13193;
   wire n_257_76_13194;
   wire n_257_76_13195;
   wire n_257_76_13196;
   wire n_257_76_13197;
   wire n_257_76_13198;
   wire n_257_76_13199;
   wire n_257_76_13200;
   wire n_257_76_13201;
   wire n_257_76_13202;
   wire n_257_76_13203;
   wire n_257_76_13204;
   wire n_257_76_13205;
   wire n_257_76_13206;
   wire n_257_76_13207;
   wire n_257_76_13208;
   wire n_257_76_13209;
   wire n_257_76_13210;
   wire n_257_76_13211;
   wire n_257_76_13212;
   wire n_257_76_13213;
   wire n_257_76_13214;
   wire n_257_76_13215;
   wire n_257_76_13216;
   wire n_257_76_13217;
   wire n_257_76_13218;
   wire n_257_76_13219;
   wire n_257_76_13220;
   wire n_257_76_13221;
   wire n_257_76_13222;
   wire n_257_76_13223;
   wire n_257_76_13224;
   wire n_257_76_13225;
   wire n_257_76_13226;
   wire n_257_76_13227;
   wire n_257_76_13228;
   wire n_257_76_13229;
   wire n_257_76_13230;
   wire n_257_76_13231;
   wire n_257_76_13232;
   wire n_257_76_13233;
   wire n_257_76_13234;
   wire n_257_76_13235;
   wire n_257_76_13236;
   wire n_257_76_13237;
   wire n_257_76_13238;
   wire n_257_76_13239;
   wire n_257_76_13240;
   wire n_257_76_13241;
   wire n_257_76_13242;
   wire n_257_76_13243;
   wire n_257_76_13244;
   wire n_257_76_13245;
   wire n_257_76_13246;
   wire n_257_76_13247;
   wire n_257_76_13248;
   wire n_257_76_13249;
   wire n_257_76_13250;
   wire n_257_76_13251;
   wire n_257_76_13252;
   wire n_257_76_13253;
   wire n_257_76_13254;
   wire n_257_76_13255;
   wire n_257_76_13256;
   wire n_257_76_13257;
   wire n_257_76_13258;
   wire n_257_76_13259;
   wire n_257_76_13260;
   wire n_257_76_13261;
   wire n_257_76_13262;
   wire n_257_76_13263;
   wire n_257_76_13264;
   wire n_257_76_13265;
   wire n_257_76_13266;
   wire n_257_76_13267;
   wire n_257_76_13268;
   wire n_257_76_13269;
   wire n_257_76_13270;
   wire n_257_76_13271;
   wire n_257_76_13272;
   wire n_257_76_13273;
   wire n_257_76_13274;
   wire n_257_76_13275;
   wire n_257_76_13276;
   wire n_257_76_13277;
   wire n_257_76_13278;
   wire n_257_76_13279;
   wire n_257_76_13280;
   wire n_257_76_13281;
   wire n_257_76_13282;
   wire n_257_76_13283;
   wire n_257_76_13284;
   wire n_257_76_13285;
   wire n_257_76_13286;
   wire n_257_76_13287;
   wire n_257_76_13288;
   wire n_257_76_13289;
   wire n_257_76_13290;
   wire n_257_76_13291;
   wire n_257_76_13292;
   wire n_257_76_13293;
   wire n_257_76_13294;
   wire n_257_76_13295;
   wire n_257_76_13296;
   wire n_257_76_13297;
   wire n_257_76_13298;
   wire n_257_76_13299;
   wire n_257_76_13300;
   wire n_257_76_13301;
   wire n_257_76_13302;
   wire n_257_76_13303;
   wire n_257_76_13304;
   wire n_257_76_13305;
   wire n_257_76_13306;
   wire n_257_76_13307;
   wire n_257_76_13308;
   wire n_257_76_13309;
   wire n_257_76_13310;
   wire n_257_76_13311;
   wire n_257_76_13312;
   wire n_257_76_13313;
   wire n_257_76_13314;
   wire n_257_76_13315;
   wire n_257_76_13316;
   wire n_257_76_13317;
   wire n_257_76_13318;
   wire n_257_76_13319;
   wire n_257_76_13320;
   wire n_257_76_13321;
   wire n_257_76_13322;
   wire n_257_76_13323;
   wire n_257_76_13324;
   wire n_257_76_13325;
   wire n_257_76_13326;
   wire n_257_76_13327;
   wire n_257_76_13328;
   wire n_257_76_13329;
   wire n_257_76_13330;
   wire n_257_76_13331;
   wire n_257_76_13332;
   wire n_257_76_13333;
   wire n_257_76_13334;
   wire n_257_76_13335;
   wire n_257_76_13336;
   wire n_257_76_13337;
   wire n_257_76_13338;
   wire n_257_76_13339;
   wire n_257_76_13340;
   wire n_257_76_13341;
   wire n_257_76_13342;
   wire n_257_76_13343;
   wire n_257_76_13344;
   wire n_257_76_13345;
   wire n_257_76_13346;
   wire n_257_76_13347;
   wire n_257_76_13348;
   wire n_257_76_13349;
   wire n_257_76_13350;
   wire n_257_76_13351;
   wire n_257_76_13352;
   wire n_257_76_13353;
   wire n_257_76_13354;
   wire n_257_76_13355;
   wire n_257_76_13356;
   wire n_257_76_13357;
   wire n_257_76_13358;
   wire n_257_76_13359;
   wire n_257_76_13360;
   wire n_257_76_13361;
   wire n_257_76_13362;
   wire n_257_76_13363;
   wire n_257_76_13364;
   wire n_257_76_13365;
   wire n_257_76_13366;
   wire n_257_76_13367;
   wire n_257_76_13368;
   wire n_257_76_13369;
   wire n_257_76_13370;
   wire n_257_76_13371;
   wire n_257_76_13372;
   wire n_257_76_13373;
   wire n_257_76_13374;
   wire n_257_76_13375;
   wire n_257_76_13376;
   wire n_257_76_13377;
   wire n_257_76_13378;
   wire n_257_76_13379;
   wire n_257_76_13380;
   wire n_257_76_13381;
   wire n_257_76_13382;
   wire n_257_76_13383;
   wire n_257_76_13384;
   wire n_257_76_13385;
   wire n_257_76_13386;
   wire n_257_76_13387;
   wire n_257_76_13388;
   wire n_257_76_13389;
   wire n_257_76_13390;
   wire n_257_76_13391;
   wire n_257_76_13392;
   wire n_257_76_13393;
   wire n_257_76_13394;
   wire n_257_76_13395;
   wire n_257_76_13396;
   wire n_257_76_13397;
   wire n_257_76_13398;
   wire n_257_76_13399;
   wire n_257_76_13400;
   wire n_257_76_13401;
   wire n_257_76_13402;
   wire n_257_76_13403;
   wire n_257_76_13404;
   wire n_257_76_13405;
   wire n_257_76_13406;
   wire n_257_76_13407;
   wire n_257_76_13408;
   wire n_257_76_13409;
   wire n_257_76_13410;
   wire n_257_76_13411;
   wire n_257_76_13412;
   wire n_257_76_13413;
   wire n_257_76_13414;
   wire n_257_76_13415;
   wire n_257_76_13416;
   wire n_257_76_13417;
   wire n_257_76_13418;
   wire n_257_76_13419;
   wire n_257_76_13420;
   wire n_257_76_13421;
   wire n_257_76_13422;
   wire n_257_76_13423;
   wire n_257_76_13424;
   wire n_257_76_13425;
   wire n_257_76_13426;
   wire n_257_76_13427;
   wire n_257_76_13428;
   wire n_257_76_13429;
   wire n_257_76_13430;
   wire n_257_76_13431;
   wire n_257_76_13432;
   wire n_257_76_13433;
   wire n_257_76_13434;
   wire n_257_76_13435;
   wire n_257_76_13436;
   wire n_257_76_13437;
   wire n_257_76_13438;
   wire n_257_76_13439;
   wire n_257_76_13440;
   wire n_257_76_13441;
   wire n_257_76_13442;
   wire n_257_76_13443;
   wire n_257_76_13444;
   wire n_257_76_13445;
   wire n_257_76_13446;
   wire n_257_76_13447;
   wire n_257_76_13448;
   wire n_257_76_13449;
   wire n_257_76_13450;
   wire n_257_76_13451;
   wire n_257_76_13452;
   wire n_257_76_13453;
   wire n_257_76_13454;
   wire n_257_76_13455;
   wire n_257_76_13456;
   wire n_257_76_13457;
   wire n_257_76_13458;
   wire n_257_76_13459;
   wire n_257_76_13460;
   wire n_257_76_13461;
   wire n_257_76_13462;
   wire n_257_76_13463;
   wire n_257_76_13464;
   wire n_257_76_13465;
   wire n_257_76_13466;
   wire n_257_76_13467;
   wire n_257_76_13468;
   wire n_257_76_13469;
   wire n_257_76_13470;
   wire n_257_76_13471;
   wire n_257_76_13472;
   wire n_257_76_13473;
   wire n_257_76_13474;
   wire n_257_76_13475;
   wire n_257_76_13476;
   wire n_257_76_13477;
   wire n_257_76_13478;
   wire n_257_76_13479;
   wire n_257_76_13480;
   wire n_257_76_13481;
   wire n_257_76_13482;
   wire n_257_76_13483;
   wire n_257_76_13484;
   wire n_257_76_13485;
   wire n_257_76_13486;
   wire n_257_76_13487;
   wire n_257_76_13488;
   wire n_257_76_13489;
   wire n_257_76_13490;
   wire n_257_76_13491;
   wire n_257_76_13492;
   wire n_257_76_13493;
   wire n_257_76_13494;
   wire n_257_76_13495;
   wire n_257_76_13496;
   wire n_257_76_13497;
   wire n_257_76_13498;
   wire n_257_76_13499;
   wire n_257_76_13500;
   wire n_257_76_13501;
   wire n_257_76_13502;
   wire n_257_76_13503;
   wire n_257_76_13504;
   wire n_257_76_13505;
   wire n_257_76_13506;
   wire n_257_76_13507;
   wire n_257_76_13508;
   wire n_257_76_13509;
   wire n_257_76_13510;
   wire n_257_76_13511;
   wire n_257_76_13512;
   wire n_257_76_13513;
   wire n_257_76_13514;
   wire n_257_76_13515;
   wire n_257_76_13516;
   wire n_257_76_13517;
   wire n_257_76_13518;
   wire n_257_76_13519;
   wire n_257_76_13520;
   wire n_257_76_13521;
   wire n_257_76_13522;
   wire n_257_76_13523;
   wire n_257_76_13524;
   wire n_257_76_13525;
   wire n_257_76_13526;
   wire n_257_76_13527;
   wire n_257_76_13528;
   wire n_257_76_13529;
   wire n_257_76_13530;
   wire n_257_76_13531;
   wire n_257_76_13532;
   wire n_257_76_13533;
   wire n_257_76_13534;
   wire n_257_76_13535;
   wire n_257_76_13536;
   wire n_257_76_13537;
   wire n_257_76_13538;
   wire n_257_76_13539;
   wire n_257_76_13540;
   wire n_257_76_13541;
   wire n_257_76_13542;
   wire n_257_76_13543;
   wire n_257_76_13544;
   wire n_257_76_13545;
   wire n_257_76_13546;
   wire n_257_76_13547;
   wire n_257_76_13548;
   wire n_257_76_13549;
   wire n_257_76_13550;
   wire n_257_76_13551;
   wire n_257_76_13552;
   wire n_257_76_13553;
   wire n_257_76_13554;
   wire n_257_76_13555;
   wire n_257_76_13556;
   wire n_257_76_13557;
   wire n_257_76_13558;
   wire n_257_76_13559;
   wire n_257_76_13560;
   wire n_257_76_13561;
   wire n_257_76_13562;
   wire n_257_76_13563;
   wire n_257_76_13564;
   wire n_257_76_13565;
   wire n_257_76_13566;
   wire n_257_76_13567;
   wire n_257_76_13568;
   wire n_257_76_13569;
   wire n_257_76_13570;
   wire n_257_76_13571;
   wire n_257_76_13572;
   wire n_257_76_13573;
   wire n_257_76_13574;
   wire n_257_76_13575;
   wire n_257_76_13576;
   wire n_257_76_13577;
   wire n_257_76_13578;
   wire n_257_76_13579;
   wire n_257_76_13580;
   wire n_257_76_13581;
   wire n_257_76_13582;
   wire n_257_76_13583;
   wire n_257_76_13584;
   wire n_257_76_13585;
   wire n_257_76_13586;
   wire n_257_76_13587;
   wire n_257_76_13588;
   wire n_257_76_13589;
   wire n_257_76_13590;
   wire n_257_76_13591;
   wire n_257_76_13592;
   wire n_257_76_13593;
   wire n_257_76_13594;
   wire n_257_76_13595;
   wire n_257_76_13596;
   wire n_257_76_13597;
   wire n_257_76_13598;
   wire n_257_76_13599;
   wire n_257_76_13600;
   wire n_257_76_13601;
   wire n_257_76_13602;
   wire n_257_76_13603;
   wire n_257_76_13604;
   wire n_257_76_13605;
   wire n_257_76_13606;
   wire n_257_76_13607;
   wire n_257_76_13608;
   wire n_257_76_13609;
   wire n_257_76_13610;
   wire n_257_76_13611;
   wire n_257_76_13612;
   wire n_257_76_13613;
   wire n_257_76_13614;
   wire n_257_76_13615;
   wire n_257_76_13616;
   wire n_257_76_13617;
   wire n_257_76_13618;
   wire n_257_76_13619;
   wire n_257_76_13620;
   wire n_257_76_13621;
   wire n_257_76_13622;
   wire n_257_76_13623;
   wire n_257_76_13624;
   wire n_257_76_13625;
   wire n_257_76_13626;
   wire n_257_76_13627;
   wire n_257_76_13628;
   wire n_257_76_13629;
   wire n_257_76_13630;
   wire n_257_76_13631;
   wire n_257_76_13632;
   wire n_257_76_13633;
   wire n_257_76_13634;
   wire n_257_76_13635;
   wire n_257_76_13636;
   wire n_257_76_13637;
   wire n_257_76_13638;
   wire n_257_76_13639;
   wire n_257_76_13640;
   wire n_257_76_13641;
   wire n_257_76_13642;
   wire n_257_76_13643;
   wire n_257_76_13644;
   wire n_257_76_13645;
   wire n_257_76_13646;
   wire n_257_76_13647;
   wire n_257_76_13648;
   wire n_257_76_13649;
   wire n_257_76_13650;
   wire n_257_76_13651;
   wire n_257_76_13652;
   wire n_257_76_13653;
   wire n_257_76_13654;
   wire n_257_76_13655;
   wire n_257_76_13656;
   wire n_257_76_13657;
   wire n_257_76_13658;
   wire n_257_76_13659;
   wire n_257_76_13660;
   wire n_257_76_13661;
   wire n_257_76_13662;
   wire n_257_76_13663;
   wire n_257_76_13664;
   wire n_257_76_13665;
   wire n_257_76_13666;
   wire n_257_76_13667;
   wire n_257_76_13668;
   wire n_257_76_13669;
   wire n_257_76_13670;
   wire n_257_76_13671;
   wire n_257_76_13672;
   wire n_257_76_13673;
   wire n_257_76_13674;
   wire n_257_76_13675;
   wire n_257_76_13676;
   wire n_257_76_13677;
   wire n_257_76_13678;
   wire n_257_76_13679;
   wire n_257_76_13680;
   wire n_257_76_13681;
   wire n_257_76_13682;
   wire n_257_76_13683;
   wire n_257_76_13684;
   wire n_257_76_13685;
   wire n_257_76_13686;
   wire n_257_76_13687;
   wire n_257_76_13688;
   wire n_257_76_13689;
   wire n_257_76_13690;
   wire n_257_76_13691;
   wire n_257_76_13692;
   wire n_257_76_13693;
   wire n_257_76_13694;
   wire n_257_76_13695;
   wire n_257_76_13696;
   wire n_257_76_13697;
   wire n_257_76_13698;
   wire n_257_76_13699;
   wire n_257_76_13700;
   wire n_257_76_13701;
   wire n_257_76_13702;
   wire n_257_76_13703;
   wire n_257_76_13704;
   wire n_257_76_13705;
   wire n_257_76_13706;
   wire n_257_76_13707;
   wire n_257_76_13708;
   wire n_257_76_13709;
   wire n_257_76_13710;
   wire n_257_76_13711;
   wire n_257_76_13712;
   wire n_257_76_13713;
   wire n_257_76_13714;
   wire n_257_76_13715;
   wire n_257_76_13716;
   wire n_257_76_13717;
   wire n_257_76_13718;
   wire n_257_76_13719;
   wire n_257_76_13720;
   wire n_257_76_13721;
   wire n_257_76_13722;
   wire n_257_76_13723;
   wire n_257_76_13724;
   wire n_257_76_13725;
   wire n_257_76_13726;
   wire n_257_76_13727;
   wire n_257_76_13728;
   wire n_257_76_13729;
   wire n_257_76_13730;
   wire n_257_76_13731;
   wire n_257_76_13732;
   wire n_257_76_13733;
   wire n_257_76_13734;
   wire n_257_76_13735;
   wire n_257_76_13736;
   wire n_257_76_13737;
   wire n_257_76_13738;
   wire n_257_76_13739;
   wire n_257_76_13740;
   wire n_257_76_13741;
   wire n_257_76_13742;
   wire n_257_76_13743;
   wire n_257_76_13744;
   wire n_257_76_13745;
   wire n_257_76_13746;
   wire n_257_76_13747;
   wire n_257_76_13748;
   wire n_257_76_13749;
   wire n_257_76_13750;
   wire n_257_76_13751;
   wire n_257_76_13752;
   wire n_257_76_13753;
   wire n_257_76_13754;
   wire n_257_76_13755;
   wire n_257_76_13756;
   wire n_257_76_13757;
   wire n_257_76_13758;
   wire n_257_76_13759;
   wire n_257_76_13760;
   wire n_257_76_13761;
   wire n_257_76_13762;
   wire n_257_76_13763;
   wire n_257_76_13764;
   wire n_257_76_13765;
   wire n_257_76_13766;
   wire n_257_76_13767;
   wire n_257_76_13768;
   wire n_257_76_13769;
   wire n_257_76_13770;
   wire n_257_76_13771;
   wire n_257_76_13772;
   wire n_257_76_13773;
   wire n_257_76_13774;
   wire n_257_76_13775;
   wire n_257_76_13776;
   wire n_257_76_13777;
   wire n_257_76_13778;
   wire n_257_76_13779;
   wire n_257_76_13780;
   wire n_257_76_13781;
   wire n_257_76_13782;
   wire n_257_76_13783;
   wire n_257_76_13784;
   wire n_257_76_13785;
   wire n_257_76_13786;
   wire n_257_76_13787;
   wire n_257_76_13788;
   wire n_257_76_13789;
   wire n_257_76_13790;
   wire n_257_76_13791;
   wire n_257_76_13792;
   wire n_257_76_13793;
   wire n_257_76_13794;
   wire n_257_76_13795;
   wire n_257_76_13796;
   wire n_257_76_13797;
   wire n_257_76_13798;
   wire n_257_76_13799;
   wire n_257_76_13800;
   wire n_257_76_13801;
   wire n_257_76_13802;
   wire n_257_76_13803;
   wire n_257_76_13804;
   wire n_257_76_13805;
   wire n_257_76_13806;
   wire n_257_76_13807;
   wire n_257_76_13808;
   wire n_257_76_13809;
   wire n_257_76_13810;
   wire n_257_76_13811;
   wire n_257_76_13812;
   wire n_257_76_13813;
   wire n_257_76_13814;
   wire n_257_76_13815;
   wire n_257_76_13816;
   wire n_257_76_13817;
   wire n_257_76_13818;
   wire n_257_76_13819;
   wire n_257_76_13820;
   wire n_257_76_13821;
   wire n_257_76_13822;
   wire n_257_76_13823;
   wire n_257_76_13824;
   wire n_257_76_13825;
   wire n_257_76_13826;
   wire n_257_76_13827;
   wire n_257_76_13828;
   wire n_257_76_13829;
   wire n_257_76_13830;
   wire n_257_76_13831;
   wire n_257_76_13832;
   wire n_257_76_13833;
   wire n_257_76_13834;
   wire n_257_76_13835;
   wire n_257_76_13836;
   wire n_257_76_13837;
   wire n_257_76_13838;
   wire n_257_76_13839;
   wire n_257_76_13840;
   wire n_257_76_13841;
   wire n_257_76_13842;
   wire n_257_76_13843;
   wire n_257_76_13844;
   wire n_257_76_13845;
   wire n_257_76_13846;
   wire n_257_76_13847;
   wire n_257_76_13848;
   wire n_257_76_13849;
   wire n_257_76_13850;
   wire n_257_76_13851;
   wire n_257_76_13852;
   wire n_257_76_13853;
   wire n_257_76_13854;
   wire n_257_76_13855;
   wire n_257_76_13856;
   wire n_257_76_13857;
   wire n_257_76_13858;
   wire n_257_76_13859;
   wire n_257_76_13860;
   wire n_257_76_13861;
   wire n_257_76_13862;
   wire n_257_76_13863;
   wire n_257_76_13864;
   wire n_257_76_13865;
   wire n_257_76_13866;
   wire n_257_76_13867;
   wire n_257_76_13868;
   wire n_257_76_13869;
   wire n_257_76_13870;
   wire n_257_76_13871;
   wire n_257_76_13872;
   wire n_257_76_13873;
   wire n_257_76_13874;
   wire n_257_76_13875;
   wire n_257_76_13876;
   wire n_257_76_13877;
   wire n_257_76_13878;
   wire n_257_76_13879;
   wire n_257_76_13880;
   wire n_257_76_13881;
   wire n_257_76_13882;
   wire n_257_76_13883;
   wire n_257_76_13884;
   wire n_257_76_13885;
   wire n_257_76_13886;
   wire n_257_76_13887;
   wire n_257_76_13888;
   wire n_257_76_13889;
   wire n_257_76_13890;
   wire n_257_76_13891;
   wire n_257_76_13892;
   wire n_257_76_13893;
   wire n_257_76_13894;
   wire n_257_76_13895;
   wire n_257_76_13896;
   wire n_257_76_13897;
   wire n_257_76_13898;
   wire n_257_76_13899;
   wire n_257_76_13900;
   wire n_257_76_13901;
   wire n_257_76_13902;
   wire n_257_76_13903;
   wire n_257_76_13904;
   wire n_257_76_13905;
   wire n_257_76_13906;
   wire n_257_76_13907;
   wire n_257_76_13908;
   wire n_257_76_13909;
   wire n_257_76_13910;
   wire n_257_76_13911;
   wire n_257_76_13912;
   wire n_257_76_13913;
   wire n_257_76_13914;
   wire n_257_76_13915;
   wire n_257_76_13916;
   wire n_257_76_13917;
   wire n_257_76_13918;
   wire n_257_76_13919;
   wire n_257_76_13920;
   wire n_257_76_13921;
   wire n_257_76_13922;
   wire n_257_76_13923;
   wire n_257_76_13924;
   wire n_257_76_13925;
   wire n_257_76_13926;
   wire n_257_76_13927;
   wire n_257_76_13928;
   wire n_257_76_13929;
   wire n_257_76_13930;
   wire n_257_76_13931;
   wire n_257_76_13932;
   wire n_257_76_13933;
   wire n_257_76_13934;
   wire n_257_76_13935;
   wire n_257_76_13936;
   wire n_257_76_13937;
   wire n_257_76_13938;
   wire n_257_76_13939;
   wire n_257_76_13940;
   wire n_257_76_13941;
   wire n_257_76_13942;
   wire n_257_76_13943;
   wire n_257_76_13944;
   wire n_257_76_13945;
   wire n_257_76_13946;
   wire n_257_76_13947;
   wire n_257_76_13948;
   wire n_257_76_13949;
   wire n_257_76_13950;
   wire n_257_76_13951;
   wire n_257_76_13952;
   wire n_257_76_13953;
   wire n_257_76_13954;
   wire n_257_76_13955;
   wire n_257_76_13956;
   wire n_257_76_13957;
   wire n_257_76_13958;
   wire n_257_76_13959;
   wire n_257_76_13960;
   wire n_257_76_13961;
   wire n_257_76_13962;
   wire n_257_76_13963;
   wire n_257_76_13964;
   wire n_257_76_13965;
   wire n_257_76_13966;
   wire n_257_76_13967;
   wire n_257_76_13968;
   wire n_257_76_13969;
   wire n_257_76_13970;
   wire n_257_76_13971;
   wire n_257_76_13972;
   wire n_257_76_13973;
   wire n_257_76_13974;
   wire n_257_76_13975;
   wire n_257_76_13976;
   wire n_257_76_13977;
   wire n_257_76_13978;
   wire n_257_76_13979;
   wire n_257_76_13980;
   wire n_257_76_13981;
   wire n_257_76_13982;
   wire n_257_76_13983;
   wire n_257_76_13984;
   wire n_257_76_13985;
   wire n_257_76_13986;
   wire n_257_76_13987;
   wire n_257_76_13988;
   wire n_257_76_13989;
   wire n_257_76_13990;
   wire n_257_76_13991;
   wire n_257_76_13992;
   wire n_257_76_13993;
   wire n_257_76_13994;
   wire n_257_76_13995;
   wire n_257_76_13996;
   wire n_257_76_13997;
   wire n_257_76_13998;
   wire n_257_76_13999;
   wire n_257_76_14000;
   wire n_257_76_14001;
   wire n_257_76_14002;
   wire n_257_76_14003;
   wire n_257_76_14004;
   wire n_257_76_14005;
   wire n_257_76_14006;
   wire n_257_76_14007;
   wire n_257_76_14008;
   wire n_257_76_14009;
   wire n_257_76_14010;
   wire n_257_76_14011;
   wire n_257_76_14012;
   wire n_257_76_14013;
   wire n_257_76_14014;
   wire n_257_76_14015;
   wire n_257_76_14016;
   wire n_257_76_14017;
   wire n_257_76_14018;
   wire n_257_76_14019;
   wire n_257_76_14020;
   wire n_257_76_14021;
   wire n_257_76_14022;
   wire n_257_76_14023;
   wire n_257_76_14024;
   wire n_257_76_14025;
   wire n_257_76_14026;
   wire n_257_76_14027;
   wire n_257_76_14028;
   wire n_257_76_14029;
   wire n_257_76_14030;
   wire n_257_76_14031;
   wire n_257_76_14032;
   wire n_257_76_14033;
   wire n_257_76_14034;
   wire n_257_76_14035;
   wire n_257_76_14036;
   wire n_257_76_14037;
   wire n_257_76_14038;
   wire n_257_76_14039;
   wire n_257_76_14040;
   wire n_257_76_14041;
   wire n_257_76_14042;
   wire n_257_76_14043;
   wire n_257_76_14044;
   wire n_257_76_14045;
   wire n_257_76_14046;
   wire n_257_76_14047;
   wire n_257_76_14048;
   wire n_257_76_14049;
   wire n_257_76_14050;
   wire n_257_76_14051;
   wire n_257_76_14052;
   wire n_257_76_14053;
   wire n_257_76_14054;
   wire n_257_76_14055;
   wire n_257_76_14056;
   wire n_257_76_14057;
   wire n_257_76_14058;
   wire n_257_76_14059;
   wire n_257_76_14060;
   wire n_257_76_14061;
   wire n_257_76_14062;
   wire n_257_76_14063;
   wire n_257_76_14064;
   wire n_257_76_14065;
   wire n_257_76_14066;
   wire n_257_76_14067;
   wire n_257_76_14068;
   wire n_257_76_14069;
   wire n_257_76_14070;
   wire n_257_76_14071;
   wire n_257_76_14072;
   wire n_257_76_14073;
   wire n_257_76_14074;
   wire n_257_76_14075;
   wire n_257_76_14076;
   wire n_257_76_14077;
   wire n_257_76_14078;
   wire n_257_76_14079;
   wire n_257_76_14080;
   wire n_257_76_14081;
   wire n_257_76_14082;
   wire n_257_76_14083;
   wire n_257_76_14084;
   wire n_257_76_14085;
   wire n_257_76_14086;
   wire n_257_76_14087;
   wire n_257_76_14088;
   wire n_257_76_14089;
   wire n_257_76_14090;
   wire n_257_76_14091;
   wire n_257_76_14092;
   wire n_257_76_14093;
   wire n_257_76_14094;
   wire n_257_76_14095;
   wire n_257_76_14096;
   wire n_257_76_14097;
   wire n_257_76_14098;
   wire n_257_76_14099;
   wire n_257_76_14100;
   wire n_257_76_14101;
   wire n_257_76_14102;
   wire n_257_76_14103;
   wire n_257_76_14104;
   wire n_257_76_14105;
   wire n_257_76_14106;
   wire n_257_76_14107;
   wire n_257_76_14108;
   wire n_257_76_14109;
   wire n_257_76_14110;
   wire n_257_76_14111;
   wire n_257_76_14112;
   wire n_257_76_14113;
   wire n_257_76_14114;
   wire n_257_76_14115;
   wire n_257_76_14116;
   wire n_257_76_14117;
   wire n_257_76_14118;
   wire n_257_76_14119;
   wire n_257_76_14120;
   wire n_257_76_14121;
   wire n_257_76_14122;
   wire n_257_76_14123;
   wire n_257_76_14124;
   wire n_257_76_14125;
   wire n_257_76_14126;
   wire n_257_76_14127;
   wire n_257_76_14128;
   wire n_257_76_14129;
   wire n_257_76_14130;
   wire n_257_76_14131;
   wire n_257_76_14132;
   wire n_257_76_14133;
   wire n_257_76_14134;
   wire n_257_76_14135;
   wire n_257_76_14136;
   wire n_257_76_14137;
   wire n_257_76_14138;
   wire n_257_76_14139;
   wire n_257_76_14140;
   wire n_257_76_14141;
   wire n_257_76_14142;
   wire n_257_76_14143;
   wire n_257_76_14144;
   wire n_257_76_14145;
   wire n_257_76_14146;
   wire n_257_76_14147;
   wire n_257_76_14148;
   wire n_257_76_14149;
   wire n_257_76_14150;
   wire n_257_76_14151;
   wire n_257_76_14152;
   wire n_257_76_14153;
   wire n_257_76_14154;
   wire n_257_76_14155;
   wire n_257_76_14156;
   wire n_257_76_14157;
   wire n_257_76_14158;
   wire n_257_76_14159;
   wire n_257_76_14160;
   wire n_257_76_14161;
   wire n_257_76_14162;
   wire n_257_76_14163;
   wire n_257_76_14164;
   wire n_257_76_14165;
   wire n_257_76_14166;
   wire n_257_76_14167;
   wire n_257_76_14168;
   wire n_257_76_14169;
   wire n_257_76_14170;
   wire n_257_76_14171;
   wire n_257_76_14172;
   wire n_257_76_14173;
   wire n_257_76_14174;
   wire n_257_76_14175;
   wire n_257_76_14176;
   wire n_257_76_14177;
   wire n_257_76_14178;
   wire n_257_76_14179;
   wire n_257_76_14180;
   wire n_257_76_14181;
   wire n_257_76_14182;
   wire n_257_76_14183;
   wire n_257_76_14184;
   wire n_257_76_14185;
   wire n_257_76_14186;
   wire n_257_76_14187;
   wire n_257_76_14188;
   wire n_257_76_14189;
   wire n_257_76_14190;
   wire n_257_76_14191;
   wire n_257_76_14192;
   wire n_257_76_14193;
   wire n_257_76_14194;
   wire n_257_76_14195;
   wire n_257_76_14196;
   wire n_257_76_14197;
   wire n_257_76_14198;
   wire n_257_76_14199;
   wire n_257_76_14200;
   wire n_257_76_14201;
   wire n_257_76_14202;
   wire n_257_76_14203;
   wire n_257_76_14204;
   wire n_257_76_14205;
   wire n_257_76_14206;
   wire n_257_76_14207;
   wire n_257_76_14208;
   wire n_257_76_14209;
   wire n_257_76_14210;
   wire n_257_76_14211;
   wire n_257_76_14212;
   wire n_257_76_14213;
   wire n_257_76_14214;
   wire n_257_76_14215;
   wire n_257_76_14216;
   wire n_257_76_14217;
   wire n_257_76_14218;
   wire n_257_76_14219;
   wire n_257_76_14220;
   wire n_257_76_14221;
   wire n_257_76_14222;
   wire n_257_76_14223;
   wire n_257_76_14224;
   wire n_257_76_14225;
   wire n_257_76_14226;
   wire n_257_76_14227;
   wire n_257_76_14228;
   wire n_257_76_14229;
   wire n_257_76_14230;
   wire n_257_76_14231;
   wire n_257_76_14232;
   wire n_257_76_14233;
   wire n_257_76_14234;
   wire n_257_76_14235;
   wire n_257_76_14236;
   wire n_257_76_14237;
   wire n_257_76_14238;
   wire n_257_76_14239;
   wire n_257_76_14240;
   wire n_257_76_14241;
   wire n_257_76_14242;
   wire n_257_76_14243;
   wire n_257_76_14244;
   wire n_257_76_14245;
   wire n_257_76_14246;
   wire n_257_76_14247;
   wire n_257_76_14248;
   wire n_257_76_14249;
   wire n_257_76_14250;
   wire n_257_76_14251;
   wire n_257_76_14252;
   wire n_257_76_14253;
   wire n_257_76_14254;
   wire n_257_76_14255;
   wire n_257_76_14256;
   wire n_257_76_14257;
   wire n_257_76_14258;
   wire n_257_76_14259;
   wire n_257_76_14260;
   wire n_257_76_14261;
   wire n_257_76_14262;
   wire n_257_76_14263;
   wire n_257_76_14264;
   wire n_257_76_14265;
   wire n_257_76_14266;
   wire n_257_76_14267;
   wire n_257_76_14268;
   wire n_257_76_14269;
   wire n_257_76_14270;
   wire n_257_76_14271;
   wire n_257_76_14272;
   wire n_257_76_14273;
   wire n_257_76_14274;
   wire n_257_76_14275;
   wire n_257_76_14276;
   wire n_257_76_14277;
   wire n_257_76_14278;
   wire n_257_76_14279;
   wire n_257_76_14280;
   wire n_257_76_14281;
   wire n_257_76_14282;
   wire n_257_76_14283;
   wire n_257_76_14284;
   wire n_257_76_14285;
   wire n_257_76_14286;
   wire n_257_76_14287;
   wire n_257_76_14288;
   wire n_257_76_14289;
   wire n_257_76_14290;
   wire n_257_76_14291;
   wire n_257_76_14292;
   wire n_257_76_14293;
   wire n_257_76_14294;
   wire n_257_76_14295;
   wire n_257_76_14296;
   wire n_257_76_14297;
   wire n_257_76_14298;
   wire n_257_76_14299;
   wire n_257_76_14300;
   wire n_257_76_14301;
   wire n_257_76_14302;
   wire n_257_76_14303;
   wire n_257_76_14304;
   wire n_257_76_14305;
   wire n_257_76_14306;
   wire n_257_76_14307;
   wire n_257_76_14308;
   wire n_257_76_14309;
   wire n_257_76_14310;
   wire n_257_76_14311;
   wire n_257_76_14312;
   wire n_257_76_14313;
   wire n_257_76_14314;
   wire n_257_76_14315;
   wire n_257_76_14316;
   wire n_257_76_14317;
   wire n_257_76_14318;
   wire n_257_76_14319;
   wire n_257_76_14320;
   wire n_257_76_14321;
   wire n_257_76_14322;
   wire n_257_76_14323;
   wire n_257_76_14324;
   wire n_257_76_14325;
   wire n_257_76_14326;
   wire n_257_76_14327;
   wire n_257_76_14328;
   wire n_257_76_14329;
   wire n_257_76_14330;
   wire n_257_76_14331;
   wire n_257_76_14332;
   wire n_257_76_14333;
   wire n_257_76_14334;
   wire n_257_76_14335;
   wire n_257_76_14336;
   wire n_257_76_14337;
   wire n_257_76_14338;
   wire n_257_76_14339;
   wire n_257_76_14340;
   wire n_257_76_14341;
   wire n_257_76_14342;
   wire n_257_76_14343;
   wire n_257_76_14344;
   wire n_257_76_14345;
   wire n_257_76_14346;
   wire n_257_76_14347;
   wire n_257_76_14348;
   wire n_257_76_14349;
   wire n_257_76_14350;
   wire n_257_76_14351;
   wire n_257_76_14352;
   wire n_257_76_14353;
   wire n_257_76_14354;
   wire n_257_76_14355;
   wire n_257_76_14356;
   wire n_257_76_14357;
   wire n_257_76_14358;
   wire n_257_76_14359;
   wire n_257_76_14360;
   wire n_257_76_14361;
   wire n_257_76_14362;
   wire n_257_76_14363;
   wire n_257_76_14364;
   wire n_257_76_14365;
   wire n_257_76_14366;
   wire n_257_76_14367;
   wire n_257_76_14368;
   wire n_257_76_14369;
   wire n_257_76_14370;
   wire n_257_76_14371;
   wire n_257_76_14372;
   wire n_257_76_14373;
   wire n_257_76_14374;
   wire n_257_76_14375;
   wire n_257_76_14376;
   wire n_257_76_14377;
   wire n_257_76_14378;
   wire n_257_76_14379;
   wire n_257_76_14380;
   wire n_257_76_14381;
   wire n_257_76_14382;
   wire n_257_76_14383;
   wire n_257_76_14384;
   wire n_257_76_14385;
   wire n_257_76_14386;
   wire n_257_76_14387;
   wire n_257_76_14388;
   wire n_257_76_14389;
   wire n_257_76_14390;
   wire n_257_76_14391;
   wire n_257_76_14392;
   wire n_257_76_14393;
   wire n_257_76_14394;
   wire n_257_76_14395;
   wire n_257_76_14396;
   wire n_257_76_14397;
   wire n_257_76_14398;
   wire n_257_76_14399;
   wire n_257_76_14400;
   wire n_257_76_14401;
   wire n_257_76_14402;
   wire n_257_76_14403;
   wire n_257_76_14404;
   wire n_257_76_14405;
   wire n_257_76_14406;
   wire n_257_76_14407;
   wire n_257_76_14408;
   wire n_257_76_14409;
   wire n_257_76_14410;
   wire n_257_76_14411;
   wire n_257_76_14412;
   wire n_257_76_14413;
   wire n_257_76_14414;
   wire n_257_76_14415;
   wire n_257_76_14416;
   wire n_257_76_14417;
   wire n_257_76_14418;
   wire n_257_76_14419;
   wire n_257_76_14420;
   wire n_257_76_14421;
   wire n_257_76_14422;
   wire n_257_76_14423;
   wire n_257_76_14424;
   wire n_257_76_14425;
   wire n_257_76_14426;
   wire n_257_76_14427;
   wire n_257_76_14428;
   wire n_257_76_14429;
   wire n_257_76_14430;
   wire n_257_76_14431;
   wire n_257_76_14432;
   wire n_257_76_14433;
   wire n_257_76_14434;
   wire n_257_76_14435;
   wire n_257_76_14436;
   wire n_257_76_14437;
   wire n_257_76_14438;
   wire n_257_76_14439;
   wire n_257_76_14440;
   wire n_257_76_14441;
   wire n_257_76_14442;
   wire n_257_76_14443;
   wire n_257_76_14444;
   wire n_257_76_14445;
   wire n_257_76_14446;
   wire n_257_76_14447;
   wire n_257_76_14448;
   wire n_257_76_14449;
   wire n_257_76_14450;
   wire n_257_76_14451;
   wire n_257_76_14452;
   wire n_257_76_14453;
   wire n_257_76_14454;
   wire n_257_76_14455;
   wire n_257_76_14456;
   wire n_257_76_14457;
   wire n_257_76_14458;
   wire n_257_76_14459;
   wire n_257_76_14460;
   wire n_257_76_14461;
   wire n_257_76_14462;
   wire n_257_76_14463;
   wire n_257_76_14464;
   wire n_257_76_14465;
   wire n_257_76_14466;
   wire n_257_76_14467;
   wire n_257_76_14468;
   wire n_257_76_14469;
   wire n_257_76_14470;
   wire n_257_76_14471;
   wire n_257_76_14472;
   wire n_257_76_14473;
   wire n_257_76_14474;
   wire n_257_76_14475;
   wire n_257_76_14476;
   wire n_257_76_14477;
   wire n_257_76_14478;
   wire n_257_76_14479;
   wire n_257_76_14480;
   wire n_257_76_14481;
   wire n_257_76_14482;
   wire n_257_76_14483;
   wire n_257_76_14484;
   wire n_257_76_14485;
   wire n_257_76_14486;
   wire n_257_76_14487;
   wire n_257_76_14488;
   wire n_257_76_14489;
   wire n_257_76_14490;
   wire n_257_76_14491;
   wire n_257_76_14492;
   wire n_257_76_14493;
   wire n_257_76_14494;
   wire n_257_76_14495;
   wire n_257_76_14496;
   wire n_257_76_14497;
   wire n_257_76_14498;
   wire n_257_76_14499;
   wire n_257_76_14500;
   wire n_257_76_14501;
   wire n_257_76_14502;
   wire n_257_76_14503;
   wire n_257_76_14504;
   wire n_257_76_14505;
   wire n_257_76_14506;
   wire n_257_76_14507;
   wire n_257_76_14508;
   wire n_257_76_14509;
   wire n_257_76_14510;
   wire n_257_76_14511;
   wire n_257_76_14512;
   wire n_257_76_14513;
   wire n_257_76_14514;
   wire n_257_76_14515;
   wire n_257_76_14516;
   wire n_257_76_14517;
   wire n_257_76_14518;
   wire n_257_76_14519;
   wire n_257_76_14520;
   wire n_257_76_14521;
   wire n_257_76_14522;
   wire n_257_76_14523;
   wire n_257_76_14524;
   wire n_257_76_14525;
   wire n_257_76_14526;
   wire n_257_76_14527;
   wire n_257_76_14528;
   wire n_257_76_14529;
   wire n_257_76_14530;
   wire n_257_76_14531;
   wire n_257_76_14532;
   wire n_257_76_14533;
   wire n_257_76_14534;
   wire n_257_76_14535;
   wire n_257_76_14536;
   wire n_257_76_14537;
   wire n_257_76_14538;
   wire n_257_76_14539;
   wire n_257_76_14540;
   wire n_257_76_14541;
   wire n_257_76_14542;
   wire n_257_76_14543;
   wire n_257_76_14544;
   wire n_257_76_14545;
   wire n_257_76_14546;
   wire n_257_76_14547;
   wire n_257_76_14548;
   wire n_257_76_14549;
   wire n_257_76_14550;
   wire n_257_76_14551;
   wire n_257_76_14552;
   wire n_257_76_14553;
   wire n_257_76_14554;
   wire n_257_76_14555;
   wire n_257_76_14556;
   wire n_257_76_14557;
   wire n_257_76_14558;
   wire n_257_76_14559;
   wire n_257_76_14560;
   wire n_257_76_14561;
   wire n_257_76_14562;
   wire n_257_76_14563;
   wire n_257_76_14564;
   wire n_257_76_14565;
   wire n_257_76_14566;
   wire n_257_76_14567;
   wire n_257_76_14568;
   wire n_257_76_14569;
   wire n_257_76_14570;
   wire n_257_76_14571;
   wire n_257_76_14572;
   wire n_257_76_14573;
   wire n_257_76_14574;
   wire n_257_76_14575;
   wire n_257_76_14576;
   wire n_257_76_14577;
   wire n_257_76_14578;
   wire n_257_76_14579;
   wire n_257_76_14580;
   wire n_257_76_14581;
   wire n_257_76_14582;
   wire n_257_76_14583;
   wire n_257_76_14584;
   wire n_257_76_14585;
   wire n_257_76_14586;
   wire n_257_76_14587;
   wire n_257_76_14588;
   wire n_257_76_14589;
   wire n_257_76_14590;
   wire n_257_76_14591;
   wire n_257_76_14592;
   wire n_257_76_14593;
   wire n_257_76_14594;
   wire n_257_76_14595;
   wire n_257_76_14596;
   wire n_257_76_14597;
   wire n_257_76_14598;
   wire n_257_76_14599;
   wire n_257_76_14600;
   wire n_257_76_14601;
   wire n_257_76_14602;
   wire n_257_76_14603;
   wire n_257_76_14604;
   wire n_257_76_14605;
   wire n_257_76_14606;
   wire n_257_76_14607;
   wire n_257_76_14608;
   wire n_257_76_14609;
   wire n_257_76_14610;
   wire n_257_76_14611;
   wire n_257_76_14612;
   wire n_257_76_14613;
   wire n_257_76_14614;
   wire n_257_76_14615;
   wire n_257_76_14616;
   wire n_257_76_14617;
   wire n_257_76_14618;
   wire n_257_76_14619;
   wire n_257_76_14620;
   wire n_257_76_14621;
   wire n_257_76_14622;
   wire n_257_76_14623;
   wire n_257_76_14624;
   wire n_257_76_14625;
   wire n_257_76_14626;
   wire n_257_76_14627;
   wire n_257_76_14628;
   wire n_257_76_14629;
   wire n_257_76_14630;
   wire n_257_76_14631;
   wire n_257_76_14632;
   wire n_257_76_14633;
   wire n_257_76_14634;
   wire n_257_76_14635;
   wire n_257_76_14636;
   wire n_257_76_14637;
   wire n_257_76_14638;
   wire n_257_76_14639;
   wire n_257_76_14640;
   wire n_257_76_14641;
   wire n_257_76_14642;
   wire n_257_76_14643;
   wire n_257_76_14644;
   wire n_257_76_14645;
   wire n_257_76_14646;
   wire n_257_76_14647;
   wire n_257_76_14648;
   wire n_257_76_14649;
   wire n_257_76_14650;
   wire n_257_76_14651;
   wire n_257_76_14652;
   wire n_257_76_14653;
   wire n_257_76_14654;
   wire n_257_76_14655;
   wire n_257_76_14656;
   wire n_257_76_14657;
   wire n_257_76_14658;
   wire n_257_76_14659;
   wire n_257_76_14660;
   wire n_257_76_14661;
   wire n_257_76_14662;
   wire n_257_76_14663;
   wire n_257_76_14664;
   wire n_257_76_14665;
   wire n_257_76_14666;
   wire n_257_76_14667;
   wire n_257_76_14668;
   wire n_257_76_14669;
   wire n_257_76_14670;
   wire n_257_76_14671;
   wire n_257_76_14672;
   wire n_257_76_14673;
   wire n_257_76_14674;
   wire n_257_76_14675;
   wire n_257_76_14676;
   wire n_257_76_14677;
   wire n_257_76_14678;
   wire n_257_76_14679;
   wire n_257_76_14680;
   wire n_257_76_14681;
   wire n_257_76_14682;
   wire n_257_76_14683;
   wire n_257_76_14684;
   wire n_257_76_14685;
   wire n_257_76_14686;
   wire n_257_76_14687;
   wire n_257_76_14688;
   wire n_257_76_14689;
   wire n_257_76_14690;
   wire n_257_76_14691;
   wire n_257_76_14692;
   wire n_257_76_14693;
   wire n_257_76_14694;
   wire n_257_76_14695;
   wire n_257_76_14696;
   wire n_257_76_14697;
   wire n_257_76_14698;
   wire n_257_76_14699;
   wire n_257_76_14700;
   wire n_257_76_14701;
   wire n_257_76_14702;
   wire n_257_76_14703;
   wire n_257_76_14704;
   wire n_257_76_14705;
   wire n_257_76_14706;
   wire n_257_76_14707;
   wire n_257_76_14708;
   wire n_257_76_14709;
   wire n_257_76_14710;
   wire n_257_76_14711;
   wire n_257_76_14712;
   wire n_257_76_14713;
   wire n_257_76_14714;
   wire n_257_76_14715;
   wire n_257_76_14716;
   wire n_257_76_14717;
   wire n_257_76_14718;
   wire n_257_76_14719;
   wire n_257_76_14720;
   wire n_257_76_14721;
   wire n_257_76_14722;
   wire n_257_76_14723;
   wire n_257_76_14724;
   wire n_257_76_14725;
   wire n_257_76_14726;
   wire n_257_76_14727;
   wire n_257_76_14728;
   wire n_257_76_14729;
   wire n_257_76_14730;
   wire n_257_76_14731;
   wire n_257_76_14732;
   wire n_257_76_14733;
   wire n_257_76_14734;
   wire n_257_76_14735;
   wire n_257_76_14736;
   wire n_257_76_14737;
   wire n_257_76_14738;
   wire n_257_76_14739;
   wire n_257_76_14740;
   wire n_257_76_14741;
   wire n_257_76_14742;
   wire n_257_76_14743;
   wire n_257_76_14744;
   wire n_257_76_14745;
   wire n_257_76_14746;
   wire n_257_76_14747;
   wire n_257_76_14748;
   wire n_257_76_14749;
   wire n_257_76_14750;
   wire n_257_76_14751;
   wire n_257_76_14752;
   wire n_257_76_14753;
   wire n_257_76_14754;
   wire n_257_76_14755;
   wire n_257_76_14756;
   wire n_257_76_14757;
   wire n_257_76_14758;
   wire n_257_76_14759;
   wire n_257_76_14760;
   wire n_257_76_14761;
   wire n_257_76_14762;
   wire n_257_76_14763;
   wire n_257_76_14764;
   wire n_257_76_14765;
   wire n_257_76_14766;
   wire n_257_76_14767;
   wire n_257_76_14768;
   wire n_257_76_14769;
   wire n_257_76_14770;
   wire n_257_76_14771;
   wire n_257_76_14772;
   wire n_257_76_14773;
   wire n_257_76_14774;
   wire n_257_76_14775;
   wire n_257_76_14776;
   wire n_257_76_14777;
   wire n_257_76_14778;
   wire n_257_76_14779;
   wire n_257_76_14780;
   wire n_257_76_14781;
   wire n_257_76_14782;
   wire n_257_76_14783;
   wire n_257_76_14784;
   wire n_257_76_14785;
   wire n_257_76_14786;
   wire n_257_76_14787;
   wire n_257_76_14788;
   wire n_257_76_14789;
   wire n_257_76_14790;
   wire n_257_76_14791;
   wire n_257_76_14792;
   wire n_257_76_14793;
   wire n_257_76_14794;
   wire n_257_76_14795;
   wire n_257_76_14796;
   wire n_257_76_14797;
   wire n_257_76_14798;
   wire n_257_76_14799;
   wire n_257_76_14800;
   wire n_257_76_14801;
   wire n_257_76_14802;
   wire n_257_76_14803;
   wire n_257_76_14804;
   wire n_257_76_14805;
   wire n_257_76_14806;
   wire n_257_76_14807;
   wire n_257_76_14808;
   wire n_257_76_14809;
   wire n_257_76_14810;
   wire n_257_76_14811;
   wire n_257_76_14812;
   wire n_257_76_14813;
   wire n_257_76_14814;
   wire n_257_76_14815;
   wire n_257_76_14816;
   wire n_257_76_14817;
   wire n_257_76_14818;
   wire n_257_76_14819;
   wire n_257_76_14820;
   wire n_257_76_14821;
   wire n_257_76_14822;
   wire n_257_76_14823;
   wire n_257_76_14824;
   wire n_257_76_14825;
   wire n_257_76_14826;
   wire n_257_76_14827;
   wire n_257_76_14828;
   wire n_257_76_14829;
   wire n_257_76_14830;
   wire n_257_76_14831;
   wire n_257_76_14832;
   wire n_257_76_14833;
   wire n_257_76_14834;
   wire n_257_76_14835;
   wire n_257_76_14836;
   wire n_257_76_14837;
   wire n_257_76_14838;
   wire n_257_76_14839;
   wire n_257_76_14840;
   wire n_257_76_14841;
   wire n_257_76_14842;
   wire n_257_76_14843;
   wire n_257_76_14844;
   wire n_257_76_14845;
   wire n_257_76_14846;
   wire n_257_76_14847;
   wire n_257_76_14848;
   wire n_257_76_14849;
   wire n_257_76_14850;
   wire n_257_76_14851;
   wire n_257_76_14852;
   wire n_257_76_14853;
   wire n_257_76_14854;
   wire n_257_76_14855;
   wire n_257_76_14856;
   wire n_257_76_14857;
   wire n_257_76_14858;
   wire n_257_76_14859;
   wire n_257_76_14860;
   wire n_257_76_14861;
   wire n_257_76_14862;
   wire n_257_76_14863;
   wire n_257_76_14864;
   wire n_257_76_14865;
   wire n_257_76_14866;
   wire n_257_76_14867;
   wire n_257_76_14868;
   wire n_257_76_14869;
   wire n_257_76_14870;
   wire n_257_76_14871;
   wire n_257_76_14872;
   wire n_257_76_14873;
   wire n_257_76_14874;
   wire n_257_76_14875;
   wire n_257_76_14876;
   wire n_257_76_14877;
   wire n_257_76_14878;
   wire n_257_76_14879;
   wire n_257_76_14880;
   wire n_257_76_14881;
   wire n_257_76_14882;
   wire n_257_76_14883;
   wire n_257_76_14884;
   wire n_257_76_14885;
   wire n_257_76_14886;
   wire n_257_76_14887;
   wire n_257_76_14888;
   wire n_257_76_14889;
   wire n_257_76_14890;
   wire n_257_76_14891;
   wire n_257_76_14892;
   wire n_257_76_14893;
   wire n_257_76_14894;
   wire n_257_76_14895;
   wire n_257_76_14896;
   wire n_257_76_14897;
   wire n_257_76_14898;
   wire n_257_76_14899;
   wire n_257_76_14900;
   wire n_257_76_14901;
   wire n_257_76_14902;
   wire n_257_76_14903;
   wire n_257_76_14904;
   wire n_257_76_14905;
   wire n_257_76_14906;
   wire n_257_76_14907;
   wire n_257_76_14908;
   wire n_257_76_14909;
   wire n_257_76_14910;
   wire n_257_76_14911;
   wire n_257_76_14912;
   wire n_257_76_14913;
   wire n_257_76_14914;
   wire n_257_76_14915;
   wire n_257_76_14916;
   wire n_257_76_14917;
   wire n_257_76_14918;
   wire n_257_76_14919;
   wire n_257_76_14920;
   wire n_257_76_14921;
   wire n_257_76_14922;
   wire n_257_76_14923;
   wire n_257_76_14924;
   wire n_257_76_14925;
   wire n_257_76_14926;
   wire n_257_76_14927;
   wire n_257_76_14928;
   wire n_257_76_14929;
   wire n_257_76_14930;
   wire n_257_76_14931;
   wire n_257_76_14932;
   wire n_257_76_14933;
   wire n_257_76_14934;
   wire n_257_76_14935;
   wire n_257_76_14936;
   wire n_257_76_14937;
   wire n_257_76_14938;
   wire n_257_76_14939;
   wire n_257_76_14940;
   wire n_257_76_14941;
   wire n_257_76_14942;
   wire n_257_76_14943;
   wire n_257_76_14944;
   wire n_257_76_14945;
   wire n_257_76_14946;
   wire n_257_76_14947;
   wire n_257_76_14948;
   wire n_257_76_14949;
   wire n_257_76_14950;
   wire n_257_76_14951;
   wire n_257_76_14952;
   wire n_257_76_14953;
   wire n_257_76_14954;
   wire n_257_76_14955;
   wire n_257_76_14956;
   wire n_257_76_14957;
   wire n_257_76_14958;
   wire n_257_76_14959;
   wire n_257_76_14960;
   wire n_257_76_14961;
   wire n_257_76_14962;
   wire n_257_76_14963;
   wire n_257_76_14964;
   wire n_257_76_14965;
   wire n_257_76_14966;
   wire n_257_76_14967;
   wire n_257_76_14968;
   wire n_257_76_14969;
   wire n_257_76_14970;
   wire n_257_76_14971;
   wire n_257_76_14972;
   wire n_257_76_14973;
   wire n_257_76_14974;
   wire n_257_76_14975;
   wire n_257_76_14976;
   wire n_257_76_14977;
   wire n_257_76_14978;
   wire n_257_76_14979;
   wire n_257_76_14980;
   wire n_257_76_14981;
   wire n_257_76_14982;
   wire n_257_76_14983;
   wire n_257_76_14984;
   wire n_257_76_14985;
   wire n_257_76_14986;
   wire n_257_76_14987;
   wire n_257_76_14988;
   wire n_257_76_14989;
   wire n_257_76_14990;
   wire n_257_76_14991;
   wire n_257_76_14992;
   wire n_257_76_14993;
   wire n_257_76_14994;
   wire n_257_76_14995;
   wire n_257_76_14996;
   wire n_257_76_14997;
   wire n_257_76_14998;
   wire n_257_76_14999;
   wire n_257_76_15000;
   wire n_257_76_15001;
   wire n_257_76_15002;
   wire n_257_76_15003;
   wire n_257_76_15004;
   wire n_257_76_15005;
   wire n_257_76_15006;
   wire n_257_76_15007;
   wire n_257_76_15008;
   wire n_257_76_15009;
   wire n_257_76_15010;
   wire n_257_76_15011;
   wire n_257_76_15012;
   wire n_257_76_15013;
   wire n_257_76_15014;
   wire n_257_76_15015;
   wire n_257_76_15016;
   wire n_257_76_15017;
   wire n_257_76_15018;
   wire n_257_76_15019;
   wire n_257_76_15020;
   wire n_257_76_15021;
   wire n_257_76_15022;
   wire n_257_76_15023;
   wire n_257_76_15024;
   wire n_257_76_15025;
   wire n_257_76_15026;
   wire n_257_76_15027;
   wire n_257_76_15028;
   wire n_257_76_15029;
   wire n_257_76_15030;
   wire n_257_76_15031;
   wire n_257_76_15032;
   wire n_257_76_15033;
   wire n_257_76_15034;
   wire n_257_76_15035;
   wire n_257_76_15036;
   wire n_257_76_15037;
   wire n_257_76_15038;
   wire n_257_76_15039;
   wire n_257_76_15040;
   wire n_257_76_15041;
   wire n_257_76_15042;
   wire n_257_76_15043;
   wire n_257_76_15044;
   wire n_257_76_15045;
   wire n_257_76_15046;
   wire n_257_76_15047;
   wire n_257_76_15048;
   wire n_257_76_15049;
   wire n_257_76_15050;
   wire n_257_76_15051;
   wire n_257_76_15052;
   wire n_257_76_15053;
   wire n_257_76_15054;
   wire n_257_76_15055;
   wire n_257_76_15056;
   wire n_257_76_15057;
   wire n_257_76_15058;
   wire n_257_76_15059;
   wire n_257_76_15060;
   wire n_257_76_15061;
   wire n_257_76_15062;
   wire n_257_76_15063;
   wire n_257_76_15064;
   wire n_257_76_15065;
   wire n_257_76_15066;
   wire n_257_76_15067;
   wire n_257_76_15068;
   wire n_257_76_15069;
   wire n_257_76_15070;
   wire n_257_76_15071;
   wire n_257_76_15072;
   wire n_257_76_15073;
   wire n_257_76_15074;
   wire n_257_76_15075;
   wire n_257_76_15076;
   wire n_257_76_15077;
   wire n_257_76_15078;
   wire n_257_76_15079;
   wire n_257_76_15080;
   wire n_257_76_15081;
   wire n_257_76_15082;
   wire n_257_76_15083;
   wire n_257_76_15084;
   wire n_257_76_15085;
   wire n_257_76_15086;
   wire n_257_76_15087;
   wire n_257_76_15088;
   wire n_257_76_15089;
   wire n_257_76_15090;
   wire n_257_76_15091;
   wire n_257_76_15092;
   wire n_257_76_15093;
   wire n_257_76_15094;
   wire n_257_76_15095;
   wire n_257_76_15096;
   wire n_257_76_15097;
   wire n_257_76_15098;
   wire n_257_76_15099;
   wire n_257_76_15100;
   wire n_257_76_15101;
   wire n_257_76_15102;
   wire n_257_76_15103;
   wire n_257_76_15104;
   wire n_257_76_15105;
   wire n_257_76_15106;
   wire n_257_76_15107;
   wire n_257_76_15108;
   wire n_257_76_15109;
   wire n_257_76_15110;
   wire n_257_76_15111;
   wire n_257_76_15112;
   wire n_257_76_15113;
   wire n_257_76_15114;
   wire n_257_76_15115;
   wire n_257_76_15116;
   wire n_257_76_15117;
   wire n_257_76_15118;
   wire n_257_76_15119;
   wire n_257_76_15120;
   wire n_257_76_15121;
   wire n_257_76_15122;
   wire n_257_76_15123;
   wire n_257_76_15124;
   wire n_257_76_15125;
   wire n_257_76_15126;
   wire n_257_76_15127;
   wire n_257_76_15128;
   wire n_257_76_15129;
   wire n_257_76_15130;
   wire n_257_76_15131;
   wire n_257_76_15132;
   wire n_257_76_15133;
   wire n_257_76_15134;
   wire n_257_76_15135;
   wire n_257_76_15136;
   wire n_257_76_15137;
   wire n_257_76_15138;
   wire n_257_76_15139;
   wire n_257_76_15140;
   wire n_257_76_15141;
   wire n_257_76_15142;
   wire n_257_76_15143;
   wire n_257_76_15144;
   wire n_257_76_15145;
   wire n_257_76_15146;
   wire n_257_76_15147;
   wire n_257_76_15148;
   wire n_257_76_15149;
   wire n_257_76_15150;
   wire n_257_76_15151;
   wire n_257_76_15152;
   wire n_257_76_15153;
   wire n_257_76_15154;
   wire n_257_76_15155;
   wire n_257_76_15156;
   wire n_257_76_15157;
   wire n_257_76_15158;
   wire n_257_76_15159;
   wire n_257_76_15160;
   wire n_257_76_15161;
   wire n_257_76_15162;
   wire n_257_76_15163;
   wire n_257_76_15164;
   wire n_257_76_15165;
   wire n_257_76_15166;
   wire n_257_76_15167;
   wire n_257_76_15168;
   wire n_257_76_15169;
   wire n_257_76_15170;
   wire n_257_76_15171;
   wire n_257_76_15172;
   wire n_257_76_15173;
   wire n_257_76_15174;
   wire n_257_76_15175;
   wire n_257_76_15176;
   wire n_257_76_15177;
   wire n_257_76_15178;
   wire n_257_76_15179;
   wire n_257_76_15180;
   wire n_257_76_15181;
   wire n_257_76_15182;
   wire n_257_76_15183;
   wire n_257_76_15184;
   wire n_257_76_15185;
   wire n_257_76_15186;
   wire n_257_76_15187;
   wire n_257_76_15188;
   wire n_257_76_15189;
   wire n_257_76_15190;
   wire n_257_76_15191;
   wire n_257_76_15192;
   wire n_257_76_15193;
   wire n_257_76_15194;
   wire n_257_76_15195;
   wire n_257_76_15196;
   wire n_257_76_15197;
   wire n_257_76_15198;
   wire n_257_76_15199;
   wire n_257_76_15200;
   wire n_257_76_15201;
   wire n_257_76_15202;
   wire n_257_76_15203;
   wire n_257_76_15204;
   wire n_257_76_15205;
   wire n_257_76_15206;
   wire n_257_76_15207;
   wire n_257_76_15208;
   wire n_257_76_15209;
   wire n_257_76_15210;
   wire n_257_76_15211;
   wire n_257_76_15212;
   wire n_257_76_15213;
   wire n_257_76_15214;
   wire n_257_76_15215;
   wire n_257_76_15216;
   wire n_257_76_15217;
   wire n_257_76_15218;
   wire n_257_76_15219;
   wire n_257_76_15220;
   wire n_257_76_15221;
   wire n_257_76_15222;
   wire n_257_76_15223;
   wire n_257_76_15224;
   wire n_257_76_15225;
   wire n_257_76_15226;
   wire n_257_76_15227;
   wire n_257_76_15228;
   wire n_257_76_15229;
   wire n_257_76_15230;
   wire n_257_76_15231;
   wire n_257_76_15232;
   wire n_257_76_15233;
   wire n_257_76_15234;
   wire n_257_76_15235;
   wire n_257_76_15236;
   wire n_257_76_15237;
   wire n_257_76_15238;
   wire n_257_76_15239;
   wire n_257_76_15240;
   wire n_257_76_15241;
   wire n_257_76_15242;
   wire n_257_76_15243;
   wire n_257_76_15244;
   wire n_257_76_15245;
   wire n_257_76_15246;
   wire n_257_76_15247;
   wire n_257_76_15248;
   wire n_257_76_15249;
   wire n_257_76_15250;
   wire n_257_76_15251;
   wire n_257_76_15252;
   wire n_257_76_15253;
   wire n_257_76_15254;
   wire n_257_76_15255;
   wire n_257_76_15256;
   wire n_257_76_15257;
   wire n_257_76_15258;
   wire n_257_76_15259;
   wire n_257_76_15260;
   wire n_257_76_15261;
   wire n_257_76_15262;
   wire n_257_76_15263;
   wire n_257_76_15264;
   wire n_257_76_15265;
   wire n_257_76_15266;
   wire n_257_76_15267;
   wire n_257_76_15268;
   wire n_257_76_15269;
   wire n_257_76_15270;
   wire n_257_76_15271;
   wire n_257_76_15272;
   wire n_257_76_15273;
   wire n_257_76_15274;
   wire n_257_76_15275;
   wire n_257_76_15276;
   wire n_257_76_15277;
   wire n_257_76_15278;
   wire n_257_76_15279;
   wire n_257_76_15280;
   wire n_257_76_15281;
   wire n_257_76_15282;
   wire n_257_76_15283;
   wire n_257_76_15284;
   wire n_257_76_15285;
   wire n_257_76_15286;
   wire n_257_76_15287;
   wire n_257_76_15288;
   wire n_257_76_15289;
   wire n_257_76_15290;
   wire n_257_76_15291;
   wire n_257_76_15292;
   wire n_257_76_15293;
   wire n_257_76_15294;
   wire n_257_76_15295;
   wire n_257_76_15296;
   wire n_257_76_15297;
   wire n_257_76_15298;
   wire n_257_76_15299;
   wire n_257_76_15300;
   wire n_257_76_15301;
   wire n_257_76_15302;
   wire n_257_76_15303;
   wire n_257_76_15304;
   wire n_257_76_15305;
   wire n_257_76_15306;
   wire n_257_76_15307;
   wire n_257_76_15308;
   wire n_257_76_15309;
   wire n_257_76_15310;
   wire n_257_76_15311;
   wire n_257_76_15312;
   wire n_257_76_15313;
   wire n_257_76_15314;
   wire n_257_76_15315;
   wire n_257_76_15316;
   wire n_257_76_15317;
   wire n_257_76_15318;
   wire n_257_76_15319;
   wire n_257_76_15320;
   wire n_257_76_15321;
   wire n_257_76_15322;
   wire n_257_76_15323;
   wire n_257_76_15324;
   wire n_257_76_15325;
   wire n_257_76_15326;
   wire n_257_76_15327;
   wire n_257_76_15328;
   wire n_257_76_15329;
   wire n_257_76_15330;
   wire n_257_76_15331;
   wire n_257_76_15332;
   wire n_257_76_15333;
   wire n_257_76_15334;
   wire n_257_76_15335;
   wire n_257_76_15336;
   wire n_257_76_15337;
   wire n_257_76_15338;
   wire n_257_76_15339;
   wire n_257_76_15340;
   wire n_257_76_15341;
   wire n_257_76_15342;
   wire n_257_76_15343;
   wire n_257_76_15344;
   wire n_257_76_15345;
   wire n_257_76_15346;
   wire n_257_76_15347;
   wire n_257_76_15348;
   wire n_257_76_15349;
   wire n_257_76_15350;
   wire n_257_76_15351;
   wire n_257_76_15352;
   wire n_257_76_15353;
   wire n_257_76_15354;
   wire n_257_76_15355;
   wire n_257_76_15356;
   wire n_257_76_15357;
   wire n_257_76_15358;
   wire n_257_76_15359;
   wire n_257_76_15360;
   wire n_257_76_15361;
   wire n_257_76_15362;
   wire n_257_76_15363;
   wire n_257_76_15364;
   wire n_257_76_15365;
   wire n_257_76_15366;
   wire n_257_76_15367;
   wire n_257_76_15368;
   wire n_257_76_15369;
   wire n_257_76_15370;
   wire n_257_76_15371;
   wire n_257_76_15372;
   wire n_257_76_15373;
   wire n_257_76_15374;
   wire n_257_76_15375;
   wire n_257_76_15376;
   wire n_257_76_15377;
   wire n_257_76_15378;
   wire n_257_76_15379;
   wire n_257_76_15380;
   wire n_257_76_15381;
   wire n_257_76_15382;
   wire n_257_76_15383;
   wire n_257_76_15384;
   wire n_257_76_15385;
   wire n_257_76_15386;
   wire n_257_76_15387;
   wire n_257_76_15388;
   wire n_257_76_15389;
   wire n_257_76_15390;
   wire n_257_76_15391;
   wire n_257_76_15392;
   wire n_257_76_15393;
   wire n_257_76_15394;
   wire n_257_76_15395;
   wire n_257_76_15396;
   wire n_257_76_15397;
   wire n_257_76_15398;
   wire n_257_76_15399;
   wire n_257_76_15400;
   wire n_257_76_15401;
   wire n_257_76_15402;
   wire n_257_76_15403;
   wire n_257_76_15404;
   wire n_257_76_15405;
   wire n_257_76_15406;
   wire n_257_76_15407;
   wire n_257_76_15408;
   wire n_257_76_15409;
   wire n_257_76_15410;
   wire n_257_76_15411;
   wire n_257_76_15412;
   wire n_257_76_15413;
   wire n_257_76_15414;
   wire n_257_76_15415;
   wire n_257_76_15416;
   wire n_257_76_15417;
   wire n_257_76_15418;
   wire n_257_76_15419;
   wire n_257_76_15420;
   wire n_257_76_15421;
   wire n_257_76_15422;
   wire n_257_76_15423;
   wire n_257_76_15424;
   wire n_257_76_15425;
   wire n_257_76_15426;
   wire n_257_76_15427;
   wire n_257_76_15428;
   wire n_257_76_15429;
   wire n_257_76_15430;
   wire n_257_76_15431;
   wire n_257_76_15432;
   wire n_257_76_15433;
   wire n_257_76_15434;
   wire n_257_76_15435;
   wire n_257_76_15436;
   wire n_257_76_15437;
   wire n_257_76_15438;
   wire n_257_76_15439;
   wire n_257_76_15440;
   wire n_257_76_15441;
   wire n_257_76_15442;
   wire n_257_76_15443;
   wire n_257_76_15444;
   wire n_257_76_15445;
   wire n_257_76_15446;
   wire n_257_76_15447;
   wire n_257_76_15448;
   wire n_257_76_15449;
   wire n_257_76_15450;
   wire n_257_76_15451;
   wire n_257_76_15452;
   wire n_257_76_15453;
   wire n_257_76_15454;
   wire n_257_76_15455;
   wire n_257_76_15456;
   wire n_257_76_15457;
   wire n_257_76_15458;
   wire n_257_76_15459;
   wire n_257_76_15460;
   wire n_257_76_15461;
   wire n_257_76_15462;
   wire n_257_76_15463;
   wire n_257_76_15464;
   wire n_257_76_15465;
   wire n_257_76_15466;
   wire n_257_76_15467;
   wire n_257_76_15468;
   wire n_257_76_15469;
   wire n_257_76_15470;
   wire n_257_76_15471;
   wire n_257_76_15472;
   wire n_257_76_15473;
   wire n_257_76_15474;
   wire n_257_76_15475;
   wire n_257_76_15476;
   wire n_257_76_15477;
   wire n_257_76_15478;
   wire n_257_76_15479;
   wire n_257_76_15480;
   wire n_257_76_15481;
   wire n_257_76_15482;
   wire n_257_76_15483;
   wire n_257_76_15484;
   wire n_257_76_15485;
   wire n_257_76_15486;
   wire n_257_76_15487;
   wire n_257_76_15488;
   wire n_257_76_15489;
   wire n_257_76_15490;
   wire n_257_76_15491;
   wire n_257_76_15492;
   wire n_257_76_15493;
   wire n_257_76_15494;
   wire n_257_76_15495;
   wire n_257_76_15496;
   wire n_257_76_15497;
   wire n_257_76_15498;
   wire n_257_76_15499;
   wire n_257_76_15500;
   wire n_257_76_15501;
   wire n_257_76_15502;
   wire n_257_76_15503;
   wire n_257_76_15504;
   wire n_257_76_15505;
   wire n_257_76_15506;
   wire n_257_76_15507;
   wire n_257_76_15508;
   wire n_257_76_15509;
   wire n_257_76_15510;
   wire n_257_76_15511;
   wire n_257_76_15512;
   wire n_257_76_15513;
   wire n_257_76_15514;
   wire n_257_76_15515;
   wire n_257_76_15516;
   wire n_257_76_15517;
   wire n_257_76_15518;
   wire n_257_76_15519;
   wire n_257_76_15520;
   wire n_257_76_15521;
   wire n_257_76_15522;
   wire n_257_76_15523;
   wire n_257_76_15524;
   wire n_257_76_15525;
   wire n_257_76_15526;
   wire n_257_76_15527;
   wire n_257_76_15528;
   wire n_257_76_15529;
   wire n_257_76_15530;
   wire n_257_76_15531;
   wire n_257_76_15532;
   wire n_257_76_15533;
   wire n_257_76_15534;
   wire n_257_76_15535;
   wire n_257_76_15536;
   wire n_257_76_15537;
   wire n_257_76_15538;
   wire n_257_76_15539;
   wire n_257_76_15540;
   wire n_257_76_15541;
   wire n_257_76_15542;
   wire n_257_76_15543;
   wire n_257_76_15544;
   wire n_257_76_15545;
   wire n_257_76_15546;
   wire n_257_76_15547;
   wire n_257_76_15548;
   wire n_257_76_15549;
   wire n_257_76_15550;
   wire n_257_76_15551;
   wire n_257_76_15552;
   wire n_257_76_15553;
   wire n_257_76_15554;
   wire n_257_76_15555;
   wire n_257_76_15556;
   wire n_257_76_15557;
   wire n_257_76_15558;
   wire n_257_76_15559;
   wire n_257_76_15560;
   wire n_257_76_15561;
   wire n_257_76_15562;
   wire n_257_76_15563;
   wire n_257_76_15564;
   wire n_257_76_15565;
   wire n_257_76_15566;
   wire n_257_76_15567;
   wire n_257_76_15568;
   wire n_257_76_15569;
   wire n_257_76_15570;
   wire n_257_76_15571;
   wire n_257_76_15572;
   wire n_257_76_15573;
   wire n_257_76_15574;
   wire n_257_76_15575;
   wire n_257_76_15576;
   wire n_257_76_15577;
   wire n_257_76_15578;
   wire n_257_76_15579;
   wire n_257_76_15580;
   wire n_257_76_15581;
   wire n_257_76_15582;
   wire n_257_76_15583;
   wire n_257_76_15584;
   wire n_257_76_15585;
   wire n_257_76_15586;
   wire n_257_76_15587;
   wire n_257_76_15588;
   wire n_257_76_15589;
   wire n_257_76_15590;
   wire n_257_76_15591;
   wire n_257_76_15592;
   wire n_257_76_15593;
   wire n_257_76_15594;
   wire n_257_76_15595;
   wire n_257_76_15596;
   wire n_257_76_15597;
   wire n_257_76_15598;
   wire n_257_76_15599;
   wire n_257_76_15600;
   wire n_257_76_15601;
   wire n_257_76_15602;
   wire n_257_76_15603;
   wire n_257_76_15604;
   wire n_257_76_15605;
   wire n_257_76_15606;
   wire n_257_76_15607;
   wire n_257_76_15608;
   wire n_257_76_15609;
   wire n_257_76_15610;
   wire n_257_76_15611;
   wire n_257_76_15612;
   wire n_257_76_15613;
   wire n_257_76_15614;
   wire n_257_76_15615;
   wire n_257_76_15616;
   wire n_257_76_15617;
   wire n_257_76_15618;
   wire n_257_76_15619;
   wire n_257_76_15620;
   wire n_257_76_15621;
   wire n_257_76_15622;
   wire n_257_76_15623;
   wire n_257_76_15624;
   wire n_257_76_15625;
   wire n_257_76_15626;
   wire n_257_76_15627;
   wire n_257_76_15628;
   wire n_257_76_15629;
   wire n_257_76_15630;
   wire n_257_76_15631;
   wire n_257_76_15632;
   wire n_257_76_15633;
   wire n_257_76_15634;
   wire n_257_76_15635;
   wire n_257_76_15636;
   wire n_257_76_15637;
   wire n_257_76_15638;
   wire n_257_76_15639;
   wire n_257_76_15640;
   wire n_257_76_15641;
   wire n_257_76_15642;
   wire n_257_76_15643;
   wire n_257_76_15644;
   wire n_257_76_15645;
   wire n_257_76_15646;
   wire n_257_76_15647;
   wire n_257_76_15648;
   wire n_257_76_15649;
   wire n_257_76_15650;
   wire n_257_76_15651;
   wire n_257_76_15652;
   wire n_257_76_15653;
   wire n_257_76_15654;
   wire n_257_76_15655;
   wire n_257_76_15656;
   wire n_257_76_15657;
   wire n_257_76_15658;
   wire n_257_76_15659;
   wire n_257_76_15660;
   wire n_257_76_15661;
   wire n_257_76_15662;
   wire n_257_76_15663;
   wire n_257_76_15664;
   wire n_257_76_15665;
   wire n_257_76_15666;
   wire n_257_76_15667;
   wire n_257_76_15668;
   wire n_257_76_15669;
   wire n_257_76_15670;
   wire n_257_76_15671;
   wire n_257_76_15672;
   wire n_257_76_15673;
   wire n_257_76_15674;
   wire n_257_76_15675;
   wire n_257_76_15676;
   wire n_257_76_15677;
   wire n_257_76_15678;
   wire n_257_76_15679;
   wire n_257_76_15680;
   wire n_257_76_15681;
   wire n_257_76_15682;
   wire n_257_76_15683;
   wire n_257_76_15684;
   wire n_257_76_15685;
   wire n_257_76_15686;
   wire n_257_76_15687;
   wire n_257_76_15688;
   wire n_257_76_15689;
   wire n_257_76_15690;
   wire n_257_76_15691;
   wire n_257_76_15692;
   wire n_257_76_15693;
   wire n_257_76_15694;
   wire n_257_76_15695;
   wire n_257_76_15696;
   wire n_257_76_15697;
   wire n_257_76_15698;
   wire n_257_76_15699;
   wire n_257_76_15700;
   wire n_257_76_15701;
   wire n_257_76_15702;
   wire n_257_76_15703;
   wire n_257_76_15704;
   wire n_257_76_15705;
   wire n_257_76_15706;
   wire n_257_76_15707;
   wire n_257_76_15708;
   wire n_257_76_15709;
   wire n_257_76_15710;
   wire n_257_76_15711;
   wire n_257_76_15712;
   wire n_257_76_15713;
   wire n_257_76_15714;
   wire n_257_76_15715;
   wire n_257_76_15716;
   wire n_257_76_15717;
   wire n_257_76_15718;
   wire n_257_76_15719;
   wire n_257_76_15720;
   wire n_257_76_15721;
   wire n_257_76_15722;
   wire n_257_76_15723;
   wire n_257_76_15724;
   wire n_257_76_15725;
   wire n_257_76_15726;
   wire n_257_76_15727;
   wire n_257_76_15728;
   wire n_257_76_15729;
   wire n_257_76_15730;
   wire n_257_76_15731;
   wire n_257_76_15732;
   wire n_257_76_15733;
   wire n_257_76_15734;
   wire n_257_76_15735;
   wire n_257_76_15736;
   wire n_257_76_15737;
   wire n_257_76_15738;
   wire n_257_76_15739;
   wire n_257_76_15740;
   wire n_257_76_15741;
   wire n_257_76_15742;
   wire n_257_76_15743;
   wire n_257_76_15744;
   wire n_257_76_15745;
   wire n_257_76_15746;
   wire n_257_76_15747;
   wire n_257_76_15748;
   wire n_257_76_15749;
   wire n_257_76_15750;
   wire n_257_76_15751;
   wire n_257_76_15752;
   wire n_257_76_15753;
   wire n_257_76_15754;
   wire n_257_76_15755;
   wire n_257_76_15756;
   wire n_257_76_15757;
   wire n_257_76_15758;
   wire n_257_76_15759;
   wire n_257_76_15760;
   wire n_257_76_15761;
   wire n_257_76_15762;
   wire n_257_76_15763;
   wire n_257_76_15764;
   wire n_257_76_15765;
   wire n_257_76_15766;
   wire n_257_76_15767;
   wire n_257_76_15768;
   wire n_257_76_15769;
   wire n_257_76_15770;
   wire n_257_76_15771;
   wire n_257_76_15772;
   wire n_257_76_15773;
   wire n_257_76_15774;
   wire n_257_76_15775;
   wire n_257_76_15776;
   wire n_257_76_15777;
   wire n_257_76_15778;
   wire n_257_76_15779;
   wire n_257_76_15780;
   wire n_257_76_15781;
   wire n_257_76_15782;
   wire n_257_76_15783;
   wire n_257_76_15784;
   wire n_257_76_15785;
   wire n_257_76_15786;
   wire n_257_76_15787;
   wire n_257_76_15788;
   wire n_257_76_15789;
   wire n_257_76_15790;
   wire n_257_76_15791;
   wire n_257_76_15792;
   wire n_257_76_15793;
   wire n_257_76_15794;
   wire n_257_76_15795;
   wire n_257_76_15796;
   wire n_257_76_15797;
   wire n_257_76_15798;
   wire n_257_76_15799;
   wire n_257_76_15800;
   wire n_257_76_15801;
   wire n_257_76_15802;
   wire n_257_76_15803;
   wire n_257_76_15804;
   wire n_257_76_15805;
   wire n_257_76_15806;
   wire n_257_76_15807;
   wire n_257_76_15808;
   wire n_257_76_15809;
   wire n_257_76_15810;
   wire n_257_76_15811;
   wire n_257_76_15812;
   wire n_257_76_15813;
   wire n_257_76_15814;
   wire n_257_76_15815;
   wire n_257_76_15816;
   wire n_257_76_15817;
   wire n_257_76_15818;
   wire n_257_76_15819;
   wire n_257_76_15820;
   wire n_257_76_15821;
   wire n_257_76_15822;
   wire n_257_76_15823;
   wire n_257_76_15824;
   wire n_257_76_15825;
   wire n_257_76_15826;
   wire n_257_76_15827;
   wire n_257_76_15828;
   wire n_257_76_15829;
   wire n_257_76_15830;
   wire n_257_76_15831;
   wire n_257_76_15832;
   wire n_257_76_15833;
   wire n_257_76_15834;
   wire n_257_76_15835;
   wire n_257_76_15836;
   wire n_257_76_15837;
   wire n_257_76_15838;
   wire n_257_76_15839;
   wire n_257_76_15840;
   wire n_257_76_15841;
   wire n_257_76_15842;
   wire n_257_76_15843;
   wire n_257_76_15844;
   wire n_257_76_15845;
   wire n_257_76_15846;
   wire n_257_76_15847;
   wire n_257_76_15848;
   wire n_257_76_15849;
   wire n_257_76_15850;
   wire n_257_76_15851;
   wire n_257_76_15852;
   wire n_257_76_15853;
   wire n_257_76_15854;
   wire n_257_76_15855;
   wire n_257_76_15856;
   wire n_257_76_15857;
   wire n_257_76_15858;
   wire n_257_76_15859;
   wire n_257_76_15860;
   wire n_257_76_15861;
   wire n_257_76_15862;
   wire n_257_76_15863;
   wire n_257_76_15864;
   wire n_257_76_15865;
   wire n_257_76_15866;
   wire n_257_76_15867;
   wire n_257_76_15868;
   wire n_257_76_15869;
   wire n_257_76_15870;
   wire n_257_76_15871;
   wire n_257_76_15872;
   wire n_257_76_15873;
   wire n_257_76_15874;
   wire n_257_76_15875;
   wire n_257_76_15876;
   wire n_257_76_15877;
   wire n_257_76_15878;
   wire n_257_76_15879;
   wire n_257_76_15880;
   wire n_257_76_15881;
   wire n_257_76_15882;
   wire n_257_76_15883;
   wire n_257_76_15884;
   wire n_257_76_15885;
   wire n_257_76_15886;
   wire n_257_76_15887;
   wire n_257_76_15888;
   wire n_257_76_15889;
   wire n_257_76_15890;
   wire n_257_76_15891;
   wire n_257_76_15892;
   wire n_257_76_15893;
   wire n_257_76_15894;
   wire n_257_76_15895;
   wire n_257_76_15896;
   wire n_257_76_15897;
   wire n_257_76_15898;
   wire n_257_76_15899;
   wire n_257_76_15900;
   wire n_257_76_15901;
   wire n_257_76_15902;
   wire n_257_76_15903;
   wire n_257_76_15904;
   wire n_257_76_15905;
   wire n_257_76_15906;
   wire n_257_76_15907;
   wire n_257_76_15908;
   wire n_257_76_15909;
   wire n_257_76_15910;
   wire n_257_76_15911;
   wire n_257_76_15912;
   wire n_257_76_15913;
   wire n_257_76_15914;
   wire n_257_76_15915;
   wire n_257_76_15916;
   wire n_257_76_15917;
   wire n_257_76_15918;
   wire n_257_76_15919;
   wire n_257_76_15920;
   wire n_257_76_15921;
   wire n_257_76_15922;
   wire n_257_76_15923;
   wire n_257_76_15924;
   wire n_257_76_15925;
   wire n_257_76_15926;
   wire n_257_76_15927;
   wire n_257_76_15928;
   wire n_257_76_15929;
   wire n_257_76_15930;
   wire n_257_76_15931;
   wire n_257_76_15932;
   wire n_257_76_15933;
   wire n_257_76_15934;
   wire n_257_76_15935;
   wire n_257_76_15936;
   wire n_257_76_15937;
   wire n_257_76_15938;
   wire n_257_76_15939;
   wire n_257_76_15940;
   wire n_257_76_15941;
   wire n_257_76_15942;
   wire n_257_76_15943;
   wire n_257_76_15944;
   wire n_257_76_15945;
   wire n_257_76_15946;
   wire n_257_76_15947;
   wire n_257_76_15948;
   wire n_257_76_15949;
   wire n_257_76_15950;
   wire n_257_76_15951;
   wire n_257_76_15952;
   wire n_257_76_15953;
   wire n_257_76_15954;
   wire n_257_76_15955;
   wire n_257_76_15956;
   wire n_257_76_15957;
   wire n_257_76_15958;
   wire n_257_76_15959;
   wire n_257_76_15960;
   wire n_257_76_15961;
   wire n_257_76_15962;
   wire n_257_76_15963;
   wire n_257_76_15964;
   wire n_257_76_15965;
   wire n_257_76_15966;
   wire n_257_76_15967;
   wire n_257_76_15968;
   wire n_257_76_15969;
   wire n_257_76_15970;
   wire n_257_76_15971;
   wire n_257_76_15972;
   wire n_257_76_15973;
   wire n_257_76_15974;
   wire n_257_76_15975;
   wire n_257_76_15976;
   wire n_257_76_15977;
   wire n_257_76_15978;
   wire n_257_76_15979;
   wire n_257_76_15980;
   wire n_257_76_15981;
   wire n_257_76_15982;
   wire n_257_76_15983;
   wire n_257_76_15984;
   wire n_257_76_15985;
   wire n_257_76_15986;
   wire n_257_76_15987;
   wire n_257_76_15988;
   wire n_257_76_15989;
   wire n_257_76_15990;
   wire n_257_76_15991;
   wire n_257_76_15992;
   wire n_257_76_15993;
   wire n_257_76_15994;
   wire n_257_76_15995;
   wire n_257_76_15996;
   wire n_257_76_15997;
   wire n_257_76_15998;
   wire n_257_76_15999;
   wire n_257_76_16000;
   wire n_257_76_16001;
   wire n_257_76_16002;
   wire n_257_76_16003;
   wire n_257_76_16004;
   wire n_257_76_16005;
   wire n_257_76_16006;
   wire n_257_76_16007;
   wire n_257_76_16008;
   wire n_257_76_16009;
   wire n_257_76_16010;
   wire n_257_76_16011;
   wire n_257_76_16012;
   wire n_257_76_16013;
   wire n_257_76_16014;
   wire n_257_76_16015;
   wire n_257_76_16016;
   wire n_257_76_16017;
   wire n_257_76_16018;
   wire n_257_76_16019;
   wire n_257_76_16020;
   wire n_257_76_16021;
   wire n_257_76_16022;
   wire n_257_76_16023;
   wire n_257_76_16024;
   wire n_257_76_16025;
   wire n_257_76_16026;
   wire n_257_76_16027;
   wire n_257_76_16028;
   wire n_257_76_16029;
   wire n_257_76_16030;
   wire n_257_76_16031;
   wire n_257_76_16032;
   wire n_257_76_16033;
   wire n_257_76_16034;
   wire n_257_76_16035;
   wire n_257_76_16036;
   wire n_257_76_16037;
   wire n_257_76_16038;
   wire n_257_76_16039;
   wire n_257_76_16040;
   wire n_257_76_16041;
   wire n_257_76_16042;
   wire n_257_76_16043;
   wire n_257_76_16044;
   wire n_257_76_16045;
   wire n_257_76_16046;
   wire n_257_76_16047;
   wire n_257_76_16048;
   wire n_257_76_16049;
   wire n_257_76_16050;
   wire n_257_76_16051;
   wire n_257_76_16052;
   wire n_257_76_16053;
   wire n_257_76_16054;
   wire n_257_76_16055;
   wire n_257_76_16056;
   wire n_257_76_16057;
   wire n_257_76_16058;
   wire n_257_76_16059;
   wire n_257_76_16060;
   wire n_257_76_16061;
   wire n_257_76_16062;
   wire n_257_76_16063;
   wire n_257_76_16064;
   wire n_257_76_16065;
   wire n_257_76_16066;
   wire n_257_76_16067;
   wire n_257_76_16068;
   wire n_257_76_16069;
   wire n_257_76_16070;
   wire n_257_76_16071;
   wire n_257_76_16072;
   wire n_257_76_16073;
   wire n_257_76_16074;
   wire n_257_76_16075;
   wire n_257_76_16076;
   wire n_257_76_16077;
   wire n_257_76_16078;
   wire n_257_76_16079;
   wire n_257_76_16080;
   wire n_257_76_16081;
   wire n_257_76_16082;
   wire n_257_76_16083;
   wire n_257_76_16084;
   wire n_257_76_16085;
   wire n_257_76_16086;
   wire n_257_76_16087;
   wire n_257_76_16088;
   wire n_257_76_16089;
   wire n_257_76_16090;
   wire n_257_76_16091;
   wire n_257_76_16092;
   wire n_257_76_16093;
   wire n_257_76_16094;
   wire n_257_76_16095;
   wire n_257_76_16096;
   wire n_257_76_16097;
   wire n_257_76_16098;
   wire n_257_76_16099;
   wire n_257_76_16100;
   wire n_257_76_16101;
   wire n_257_76_16102;
   wire n_257_76_16103;
   wire n_257_76_16104;
   wire n_257_76_16105;
   wire n_257_76_16106;
   wire n_257_76_16107;
   wire n_257_76_16108;
   wire n_257_76_16109;
   wire n_257_76_16110;
   wire n_257_76_16111;
   wire n_257_76_16112;
   wire n_257_76_16113;
   wire n_257_76_16114;
   wire n_257_76_16115;
   wire n_257_76_16116;
   wire n_257_76_16117;
   wire n_257_76_16118;
   wire n_257_76_16119;
   wire n_257_76_16120;
   wire n_257_76_16121;
   wire n_257_76_16122;
   wire n_257_76_16123;
   wire n_257_76_16124;
   wire n_257_76_16125;
   wire n_257_76_16126;
   wire n_257_76_16127;
   wire n_257_76_16128;
   wire n_257_76_16129;
   wire n_257_76_16130;
   wire n_257_76_16131;
   wire n_257_76_16132;
   wire n_257_76_16133;
   wire n_257_76_16134;
   wire n_257_76_16135;
   wire n_257_76_16136;
   wire n_257_76_16137;
   wire n_257_76_16138;
   wire n_257_76_16139;
   wire n_257_76_16140;
   wire n_257_76_16141;
   wire n_257_76_16142;
   wire n_257_76_16143;
   wire n_257_76_16144;
   wire n_257_76_16145;
   wire n_257_76_16146;
   wire n_257_76_16147;
   wire n_257_76_16148;
   wire n_257_76_16149;
   wire n_257_76_16150;
   wire n_257_76_16151;
   wire n_257_76_16152;
   wire n_257_76_16153;
   wire n_257_76_16154;
   wire n_257_76_16155;
   wire n_257_76_16156;
   wire n_257_76_16157;
   wire n_257_76_16158;
   wire n_257_76_16159;
   wire n_257_76_16160;
   wire n_257_76_16161;
   wire n_257_76_16162;
   wire n_257_76_16163;
   wire n_257_76_16164;
   wire n_257_76_16165;
   wire n_257_76_16166;
   wire n_257_76_16167;
   wire n_257_76_16168;
   wire n_257_76_16169;
   wire n_257_76_16170;
   wire n_257_76_16171;
   wire n_257_76_16172;
   wire n_257_76_16173;
   wire n_257_76_16174;
   wire n_257_76_16175;
   wire n_257_76_16176;
   wire n_257_76_16177;
   wire n_257_76_16178;
   wire n_257_76_16179;
   wire n_257_76_16180;
   wire n_257_76_16181;
   wire n_257_76_16182;
   wire n_257_76_16183;
   wire n_257_76_16184;
   wire n_257_76_16185;
   wire n_257_76_16186;
   wire n_257_76_16187;
   wire n_257_76_16188;
   wire n_257_76_16189;
   wire n_257_76_16190;
   wire n_257_76_16191;
   wire n_257_76_16192;
   wire n_257_76_16193;
   wire n_257_76_16194;
   wire n_257_76_16195;
   wire n_257_76_16196;
   wire n_257_76_16197;
   wire n_257_76_16198;
   wire n_257_76_16199;
   wire n_257_76_16200;
   wire n_257_76_16201;
   wire n_257_76_16202;
   wire n_257_76_16203;
   wire n_257_76_16204;
   wire n_257_76_16205;
   wire n_257_76_16206;
   wire n_257_76_16207;
   wire n_257_76_16208;
   wire n_257_76_16209;
   wire n_257_76_16210;
   wire n_257_76_16211;
   wire n_257_76_16212;
   wire n_257_76_16213;
   wire n_257_76_16214;
   wire n_257_76_16215;
   wire n_257_76_16216;
   wire n_257_76_16217;
   wire n_257_76_16218;
   wire n_257_76_16219;
   wire n_257_76_16220;
   wire n_257_76_16221;
   wire n_257_76_16222;
   wire n_257_76_16223;
   wire n_257_76_16224;
   wire n_257_76_16225;
   wire n_257_76_16226;
   wire n_257_76_16227;
   wire n_257_76_16228;
   wire n_257_76_16229;
   wire n_257_76_16230;
   wire n_257_76_16231;
   wire n_257_76_16232;
   wire n_257_76_16233;
   wire n_257_76_16234;
   wire n_257_76_16235;
   wire n_257_76_16236;
   wire n_257_76_16237;
   wire n_257_76_16238;
   wire n_257_76_16239;
   wire n_257_76_16240;
   wire n_257_76_16241;
   wire n_257_76_16242;
   wire n_257_76_16243;
   wire n_257_76_16244;
   wire n_257_76_16245;
   wire n_257_76_16246;
   wire n_257_76_16247;
   wire n_257_76_16248;
   wire n_257_76_16249;
   wire n_257_76_16250;
   wire n_257_76_16251;
   wire n_257_76_16252;
   wire n_257_76_16253;
   wire n_257_76_16254;
   wire n_257_76_16255;
   wire n_257_76_16256;
   wire n_257_76_16257;
   wire n_257_76_16258;
   wire n_257_76_16259;
   wire n_257_76_16260;
   wire n_257_76_16261;
   wire n_257_76_16262;
   wire n_257_76_16263;
   wire n_257_76_16264;
   wire n_257_76_16265;
   wire n_257_76_16266;
   wire n_257_76_16267;
   wire n_257_76_16268;
   wire n_257_76_16269;
   wire n_257_76_16270;
   wire n_257_76_16271;
   wire n_257_76_16272;
   wire n_257_76_16273;
   wire n_257_76_16274;
   wire n_257_76_16275;
   wire n_257_76_16276;
   wire n_257_76_16277;
   wire n_257_76_16278;
   wire n_257_76_16279;
   wire n_257_76_16280;
   wire n_257_76_16281;
   wire n_257_76_16282;
   wire n_257_76_16283;
   wire n_257_76_16284;
   wire n_257_76_16285;
   wire n_257_76_16286;
   wire n_257_76_16287;
   wire n_257_76_16288;
   wire n_257_76_16289;
   wire n_257_76_16290;
   wire n_257_76_16291;
   wire n_257_76_16292;
   wire n_257_76_16293;
   wire n_257_76_16294;
   wire n_257_76_16295;
   wire n_257_76_16296;
   wire n_257_76_16297;
   wire n_257_76_16298;
   wire n_257_76_16299;
   wire n_257_76_16300;
   wire n_257_76_16301;
   wire n_257_76_16302;
   wire n_257_76_16303;
   wire n_257_76_16304;
   wire n_257_76_16305;
   wire n_257_76_16306;
   wire n_257_76_16307;
   wire n_257_76_16308;
   wire n_257_76_16309;
   wire n_257_76_16310;
   wire n_257_76_16311;
   wire n_257_76_16312;
   wire n_257_76_16313;
   wire n_257_76_16314;
   wire n_257_76_16315;
   wire n_257_76_16316;
   wire n_257_76_16317;
   wire n_257_76_16318;
   wire n_257_76_16319;
   wire n_257_76_16320;
   wire n_257_76_16321;
   wire n_257_76_16322;
   wire n_257_76_16323;
   wire n_257_76_16324;
   wire n_257_76_16325;
   wire n_257_76_16326;
   wire n_257_76_16327;
   wire n_257_76_16328;
   wire n_257_76_16329;
   wire n_257_76_16330;
   wire n_257_76_16331;
   wire n_257_76_16332;
   wire n_257_76_16333;
   wire n_257_76_16334;
   wire n_257_76_16335;
   wire n_257_76_16336;
   wire n_257_76_16337;
   wire n_257_76_16338;
   wire n_257_76_16339;
   wire n_257_76_16340;
   wire n_257_76_16341;
   wire n_257_76_16342;
   wire n_257_76_16343;
   wire n_257_76_16344;
   wire n_257_76_16345;
   wire n_257_76_16346;
   wire n_257_76_16347;
   wire n_257_76_16348;
   wire n_257_76_16349;
   wire n_257_76_16350;
   wire n_257_76_16351;
   wire n_257_76_16352;
   wire n_257_76_16353;
   wire n_257_76_16354;
   wire n_257_76_16355;
   wire n_257_76_16356;
   wire n_257_76_16357;
   wire n_257_76_16358;
   wire n_257_76_16359;
   wire n_257_76_16360;
   wire n_257_76_16361;
   wire n_257_76_16362;
   wire n_257_76_16363;
   wire n_257_76_16364;
   wire n_257_76_16365;
   wire n_257_76_16366;
   wire n_257_76_16367;
   wire n_257_76_16368;
   wire n_257_76_16369;
   wire n_257_76_16370;
   wire n_257_76_16371;
   wire n_257_76_16372;
   wire n_257_76_16373;
   wire n_257_76_16374;
   wire n_257_76_16375;
   wire n_257_76_16376;
   wire n_257_76_16377;
   wire n_257_76_16378;
   wire n_257_76_16379;
   wire n_257_76_16380;
   wire n_257_76_16381;
   wire n_257_76_16382;
   wire n_257_76_16383;
   wire n_257_76_16384;
   wire n_257_76_16385;
   wire n_257_76_16386;
   wire n_257_76_16387;
   wire n_257_76_16388;
   wire n_257_76_16389;
   wire n_257_76_16390;
   wire n_257_76_16391;
   wire n_257_76_16392;
   wire n_257_76_16393;
   wire n_257_76_16394;
   wire n_257_76_16395;
   wire n_257_76_16396;
   wire n_257_76_16397;
   wire n_257_76_16398;
   wire n_257_76_16399;
   wire n_257_76_16400;
   wire n_257_76_16401;
   wire n_257_76_16402;
   wire n_257_76_16403;
   wire n_257_76_16404;
   wire n_257_76_16405;
   wire n_257_76_16406;
   wire n_257_76_16407;
   wire n_257_76_16408;
   wire n_257_76_16409;
   wire n_257_76_16410;
   wire n_257_76_16411;
   wire n_257_76_16412;
   wire n_257_76_16413;
   wire n_257_76_16414;
   wire n_257_76_16415;
   wire n_257_76_16416;
   wire n_257_76_16417;
   wire n_257_76_16418;
   wire n_257_76_16419;
   wire n_257_76_16420;
   wire n_257_76_16421;
   wire n_257_76_16422;
   wire n_257_76_16423;
   wire n_257_76_16424;
   wire n_257_76_16425;
   wire n_257_76_16426;
   wire n_257_76_16427;
   wire n_257_76_16428;
   wire n_257_76_16429;
   wire n_257_76_16430;
   wire n_257_76_16431;
   wire n_257_76_16432;
   wire n_257_76_16433;
   wire n_257_76_16434;
   wire n_257_76_16435;
   wire n_257_76_16436;
   wire n_257_76_16437;
   wire n_257_76_16438;
   wire n_257_76_16439;
   wire n_257_76_16440;
   wire n_257_76_16441;
   wire n_257_76_16442;
   wire n_257_76_16443;
   wire n_257_76_16444;
   wire n_257_76_16445;
   wire n_257_76_16446;
   wire n_257_76_16447;
   wire n_257_76_16448;
   wire n_257_76_16449;
   wire n_257_76_16450;
   wire n_257_76_16451;
   wire n_257_76_16452;
   wire n_257_76_16453;
   wire n_257_76_16454;
   wire n_257_76_16455;
   wire n_257_76_16456;
   wire n_257_76_16457;
   wire n_257_76_16458;
   wire n_257_76_16459;
   wire n_257_76_16460;
   wire n_257_76_16461;
   wire n_257_76_16462;
   wire n_257_76_16463;
   wire n_257_76_16464;
   wire n_257_76_16465;
   wire n_257_76_16466;
   wire n_257_76_16467;
   wire n_257_76_16468;
   wire n_257_76_16469;
   wire n_257_76_16470;
   wire n_257_76_16471;
   wire n_257_76_16472;
   wire n_257_76_16473;
   wire n_257_76_16474;
   wire n_257_76_16475;
   wire n_257_76_16476;
   wire n_257_76_16477;
   wire n_257_76_16478;
   wire n_257_76_16479;
   wire n_257_76_16480;
   wire n_257_76_16481;
   wire n_257_76_16482;
   wire n_257_76_16483;
   wire n_257_76_16484;
   wire n_257_76_16485;
   wire n_257_76_16486;
   wire n_257_76_16487;
   wire n_257_76_16488;
   wire n_257_76_16489;
   wire n_257_76_16490;
   wire n_257_76_16491;
   wire n_257_76_16492;
   wire n_257_76_16493;
   wire n_257_76_16494;
   wire n_257_76_16495;
   wire n_257_76_16496;
   wire n_257_76_16497;
   wire n_257_76_16498;
   wire n_257_76_16499;
   wire n_257_76_16500;
   wire n_257_76_16501;
   wire n_257_76_16502;
   wire n_257_76_16503;
   wire n_257_76_16504;
   wire n_257_76_16505;
   wire n_257_76_16506;
   wire n_257_76_16507;
   wire n_257_76_16508;
   wire n_257_76_16509;
   wire n_257_76_16510;
   wire n_257_76_16511;
   wire n_257_76_16512;
   wire n_257_76_16513;
   wire n_257_76_16514;
   wire n_257_76_16515;
   wire n_257_76_16516;
   wire n_257_76_16517;
   wire n_257_76_16518;
   wire n_257_76_16519;
   wire n_257_76_16520;
   wire n_257_76_16521;
   wire n_257_76_16522;
   wire n_257_76_16523;
   wire n_257_76_16524;
   wire n_257_76_16525;
   wire n_257_76_16526;
   wire n_257_76_16527;
   wire n_257_76_16528;
   wire n_257_76_16529;
   wire n_257_76_16530;
   wire n_257_76_16531;
   wire n_257_76_16532;
   wire n_257_76_16533;
   wire n_257_76_16534;
   wire n_257_76_16535;
   wire n_257_76_16536;
   wire n_257_76_16537;
   wire n_257_76_16538;
   wire n_257_76_16539;
   wire n_257_76_16540;
   wire n_257_76_16541;
   wire n_257_76_16542;
   wire n_257_76_16543;
   wire n_257_76_16544;
   wire n_257_76_16545;
   wire n_257_76_16546;
   wire n_257_76_16547;
   wire n_257_76_16548;
   wire n_257_76_16549;
   wire n_257_76_16550;
   wire n_257_76_16551;
   wire n_257_76_16552;
   wire n_257_76_16553;
   wire n_257_76_16554;
   wire n_257_76_16555;
   wire n_257_76_16556;
   wire n_257_76_16557;
   wire n_257_76_16558;
   wire n_257_76_16559;
   wire n_257_76_16560;
   wire n_257_76_16561;
   wire n_257_76_16562;
   wire n_257_76_16563;
   wire n_257_76_16564;
   wire n_257_76_16565;
   wire n_257_76_16566;
   wire n_257_76_16567;
   wire n_257_76_16568;
   wire n_257_76_16569;
   wire n_257_76_16570;
   wire n_257_76_16571;
   wire n_257_76_16572;
   wire n_257_76_16573;
   wire n_257_76_16574;
   wire n_257_76_16575;
   wire n_257_76_16576;
   wire n_257_76_16577;
   wire n_257_76_16578;
   wire n_257_76_16579;
   wire n_257_76_16580;
   wire n_257_76_16581;
   wire n_257_76_16582;
   wire n_257_76_16583;
   wire n_257_76_16584;
   wire n_257_76_16585;
   wire n_257_76_16586;
   wire n_257_76_16587;
   wire n_257_76_16588;
   wire n_257_76_16589;
   wire n_257_76_16590;
   wire n_257_76_16591;
   wire n_257_76_16592;
   wire n_257_76_16593;
   wire n_257_76_16594;
   wire n_257_76_16595;
   wire n_257_76_16596;
   wire n_257_76_16597;
   wire n_257_76_16598;
   wire n_257_76_16599;
   wire n_257_76_16600;
   wire n_257_76_16601;
   wire n_257_76_16602;
   wire n_257_76_16603;
   wire n_257_76_16604;
   wire n_257_76_16605;
   wire n_257_76_16606;
   wire n_257_76_16607;
   wire n_257_76_16608;
   wire n_257_76_16609;
   wire n_257_76_16610;
   wire n_257_76_16611;
   wire n_257_76_16612;
   wire n_257_76_16613;
   wire n_257_76_16614;
   wire n_257_76_16615;
   wire n_257_76_16616;
   wire n_257_76_16617;
   wire n_257_76_16618;
   wire n_257_76_16619;
   wire n_257_76_16620;
   wire n_257_76_16621;
   wire n_257_76_16622;
   wire n_257_76_16623;
   wire n_257_76_16624;
   wire n_257_76_16625;
   wire n_257_76_16626;
   wire n_257_76_16627;
   wire n_257_76_16628;
   wire n_257_76_16629;
   wire n_257_76_16630;
   wire n_257_76_16631;
   wire n_257_76_16632;
   wire n_257_76_16633;
   wire n_257_76_16634;
   wire n_257_76_16635;
   wire n_257_76_16636;
   wire n_257_76_16637;
   wire n_257_76_16638;
   wire n_257_76_16639;
   wire n_257_76_16640;
   wire n_257_76_16641;
   wire n_257_76_16642;
   wire n_257_76_16643;
   wire n_257_76_16644;
   wire n_257_76_16645;
   wire n_257_76_16646;
   wire n_257_76_16647;
   wire n_257_76_16648;
   wire n_257_76_16649;
   wire n_257_76_16650;
   wire n_257_76_16651;
   wire n_257_76_16652;
   wire n_257_76_16653;
   wire n_257_76_16654;
   wire n_257_76_16655;
   wire n_257_76_16656;
   wire n_257_76_16657;
   wire n_257_76_16658;
   wire n_257_76_16659;
   wire n_257_76_16660;
   wire n_257_76_16661;
   wire n_257_76_16662;
   wire n_257_76_16663;
   wire n_257_76_16664;
   wire n_257_76_16665;
   wire n_257_76_16666;
   wire n_257_76_16667;
   wire n_257_76_16668;
   wire n_257_76_16669;
   wire n_257_76_16670;
   wire n_257_76_16671;
   wire n_257_76_16672;
   wire n_257_76_16673;
   wire n_257_76_16674;
   wire n_257_76_16675;
   wire n_257_76_16676;
   wire n_257_76_16677;
   wire n_257_76_16678;
   wire n_257_76_16679;
   wire n_257_76_16680;
   wire n_257_76_16681;
   wire n_257_76_16682;
   wire n_257_76_16683;
   wire n_257_76_16684;
   wire n_257_76_16685;
   wire n_257_76_16686;
   wire n_257_76_16687;
   wire n_257_76_16688;
   wire n_257_76_16689;
   wire n_257_76_16690;
   wire n_257_76_16691;
   wire n_257_76_16692;
   wire n_257_76_16693;
   wire n_257_76_16694;
   wire n_257_76_16695;
   wire n_257_76_16696;
   wire n_257_76_16697;
   wire n_257_76_16698;
   wire n_257_76_16699;
   wire n_257_76_16700;
   wire n_257_76_16701;
   wire n_257_76_16702;
   wire n_257_76_16703;
   wire n_257_76_16704;
   wire n_257_76_16705;
   wire n_257_76_16706;
   wire n_257_76_16707;
   wire n_257_76_16708;
   wire n_257_76_16709;
   wire n_257_76_16710;
   wire n_257_76_16711;
   wire n_257_76_16712;
   wire n_257_76_16713;
   wire n_257_76_16714;
   wire n_257_76_16715;
   wire n_257_76_16716;
   wire n_257_76_16717;
   wire n_257_76_16718;
   wire n_257_76_16719;
   wire n_257_76_16720;
   wire n_257_76_16721;
   wire n_257_76_16722;
   wire n_257_76_16723;
   wire n_257_76_16724;
   wire n_257_76_16725;
   wire n_257_76_16726;
   wire n_257_76_16727;
   wire n_257_76_16728;
   wire n_257_76_16729;
   wire n_257_76_16730;
   wire n_257_76_16731;
   wire n_257_76_16732;
   wire n_257_76_16733;
   wire n_257_76_16734;
   wire n_257_76_16735;
   wire n_257_76_16736;
   wire n_257_76_16737;
   wire n_257_76_16738;
   wire n_257_76_16739;
   wire n_257_76_16740;
   wire n_257_76_16741;
   wire n_257_76_16742;
   wire n_257_76_16743;
   wire n_257_76_16744;
   wire n_257_76_16745;
   wire n_257_76_16746;
   wire n_257_76_16747;
   wire n_257_76_16748;
   wire n_257_76_16749;
   wire n_257_76_16750;
   wire n_257_76_16751;
   wire n_257_76_16752;
   wire n_257_76_16753;
   wire n_257_76_16754;
   wire n_257_76_16755;
   wire n_257_76_16756;
   wire n_257_76_16757;
   wire n_257_76_16758;
   wire n_257_76_16759;
   wire n_257_76_16760;
   wire n_257_76_16761;
   wire n_257_76_16762;
   wire n_257_76_16763;
   wire n_257_76_16764;
   wire n_257_76_16765;
   wire n_257_76_16766;
   wire n_257_76_16767;
   wire n_257_76_16768;
   wire n_257_76_16769;
   wire n_257_76_16770;
   wire n_257_76_16771;
   wire n_257_76_16772;
   wire n_257_76_16773;
   wire n_257_76_16774;
   wire n_257_76_16775;
   wire n_257_76_16776;
   wire n_257_76_16777;
   wire n_257_76_16778;
   wire n_257_76_16779;
   wire n_257_76_16780;
   wire n_257_76_16781;
   wire n_257_76_16782;
   wire n_257_76_16783;
   wire n_257_76_16784;
   wire n_257_76_16785;
   wire n_257_76_16786;
   wire n_257_76_16787;
   wire n_257_76_16788;
   wire n_257_76_16789;
   wire n_257_76_16790;
   wire n_257_76_16791;
   wire n_257_76_16792;
   wire n_257_76_16793;
   wire n_257_76_16794;
   wire n_257_76_16795;
   wire n_257_76_16796;
   wire n_257_76_16797;
   wire n_257_76_16798;
   wire n_257_76_16799;
   wire n_257_76_16800;
   wire n_257_76_16801;
   wire n_257_76_16802;
   wire n_257_76_16803;
   wire n_257_76_16804;
   wire n_257_76_16805;
   wire n_257_76_16806;
   wire n_257_76_16807;
   wire n_257_76_16808;
   wire n_257_76_16809;
   wire n_257_76_16810;
   wire n_257_76_16811;
   wire n_257_76_16812;
   wire n_257_76_16813;
   wire n_257_76_16814;
   wire n_257_76_16815;
   wire n_257_76_16816;
   wire n_257_76_16817;
   wire n_257_76_16818;
   wire n_257_76_16819;
   wire n_257_76_16820;
   wire n_257_76_16821;
   wire n_257_76_16822;
   wire n_257_76_16823;
   wire n_257_76_16824;
   wire n_257_76_16825;
   wire n_257_76_16826;
   wire n_257_76_16827;
   wire n_257_76_16828;
   wire n_257_76_16829;
   wire n_257_76_16830;
   wire n_257_76_16831;
   wire n_257_76_16832;
   wire n_257_76_16833;
   wire n_257_76_16834;
   wire n_257_76_16835;
   wire n_257_76_16836;
   wire n_257_76_16837;
   wire n_257_76_16838;
   wire n_257_76_16839;
   wire n_257_76_16840;
   wire n_257_76_16841;
   wire n_257_76_16842;
   wire n_257_76_16843;
   wire n_257_76_16844;
   wire n_257_76_16845;
   wire n_257_76_16846;
   wire n_257_76_16847;
   wire n_257_76_16848;
   wire n_257_76_16849;
   wire n_257_76_16850;
   wire n_257_76_16851;
   wire n_257_76_16852;
   wire n_257_76_16853;
   wire n_257_76_16854;
   wire n_257_76_16855;
   wire n_257_76_16856;
   wire n_257_76_16857;
   wire n_257_76_16858;
   wire n_257_76_16859;
   wire n_257_76_16860;
   wire n_257_76_16861;
   wire n_257_76_16862;
   wire n_257_76_16863;
   wire n_257_76_16864;
   wire n_257_76_16865;
   wire n_257_76_16866;
   wire n_257_76_16867;
   wire n_257_76_16868;
   wire n_257_76_16869;
   wire n_257_76_16870;
   wire n_257_76_16871;
   wire n_257_76_16872;
   wire n_257_76_16873;
   wire n_257_76_16874;
   wire n_257_76_16875;
   wire n_257_76_16876;
   wire n_257_76_16877;
   wire n_257_76_16878;
   wire n_257_76_16879;
   wire n_257_76_16880;
   wire n_257_76_16881;
   wire n_257_76_16882;
   wire n_257_76_16883;
   wire n_257_76_16884;
   wire n_257_76_16885;
   wire n_257_76_16886;
   wire n_257_76_16887;
   wire n_257_76_16888;
   wire n_257_76_16889;
   wire n_257_76_16890;
   wire n_257_76_16891;
   wire n_257_76_16892;
   wire n_257_76_16893;
   wire n_257_76_16894;
   wire n_257_76_16895;
   wire n_257_76_16896;
   wire n_257_76_16897;
   wire n_257_76_16898;
   wire n_257_76_16899;
   wire n_257_76_16900;
   wire n_257_76_16901;
   wire n_257_76_16902;
   wire n_257_76_16903;
   wire n_257_76_16904;
   wire n_257_76_16905;
   wire n_257_76_16906;
   wire n_257_76_16907;
   wire n_257_76_16908;
   wire n_257_76_16909;
   wire n_257_76_16910;
   wire n_257_76_16911;
   wire n_257_76_16912;
   wire n_257_76_16913;
   wire n_257_76_16914;
   wire n_257_76_16915;
   wire n_257_76_16916;
   wire n_257_76_16917;
   wire n_257_76_16918;
   wire n_257_76_16919;
   wire n_257_76_16920;
   wire n_257_76_16921;
   wire n_257_76_16922;
   wire n_257_76_16923;
   wire n_257_76_16924;
   wire n_257_76_16925;
   wire n_257_76_16926;
   wire n_257_76_16927;
   wire n_257_76_16928;
   wire n_257_76_16929;
   wire n_257_76_16930;
   wire n_257_76_16931;
   wire n_257_76_16932;
   wire n_257_76_16933;
   wire n_257_76_16934;
   wire n_257_76_16935;
   wire n_257_76_16936;
   wire n_257_76_16937;
   wire n_257_76_16938;
   wire n_257_76_16939;
   wire n_257_76_16940;
   wire n_257_76_16941;
   wire n_257_76_16942;
   wire n_257_76_16943;
   wire n_257_76_16944;
   wire n_257_76_16945;
   wire n_257_76_16946;
   wire n_257_76_16947;
   wire n_257_76_16948;
   wire n_257_76_16949;
   wire n_257_76_16950;
   wire n_257_76_16951;
   wire n_257_76_16952;
   wire n_257_76_16953;
   wire n_257_76_16954;
   wire n_257_76_16955;
   wire n_257_76_16956;
   wire n_257_76_16957;
   wire n_257_76_16958;
   wire n_257_76_16959;
   wire n_257_76_16960;
   wire n_257_76_16961;
   wire n_257_76_16962;
   wire n_257_76_16963;
   wire n_257_76_16964;
   wire n_257_76_16965;
   wire n_257_76_16966;
   wire n_257_76_16967;
   wire n_257_76_16968;
   wire n_257_76_16969;
   wire n_257_76_16970;
   wire n_257_76_16971;
   wire n_257_76_16972;
   wire n_257_76_16973;
   wire n_257_76_16974;
   wire n_257_76_16975;
   wire n_257_76_16976;
   wire n_257_76_16977;
   wire n_257_76_16978;
   wire n_257_76_16979;
   wire n_257_76_16980;
   wire n_257_76_16981;
   wire n_257_76_16982;
   wire n_257_76_16983;
   wire n_257_76_16984;
   wire n_257_76_16985;
   wire n_257_76_16986;
   wire n_257_76_16987;
   wire n_257_76_16988;
   wire n_257_76_16989;
   wire n_257_76_16990;
   wire n_257_76_16991;
   wire n_257_76_16992;
   wire n_257_76_16993;
   wire n_257_76_16994;
   wire n_257_76_16995;
   wire n_257_76_16996;
   wire n_257_76_16997;
   wire n_257_76_16998;
   wire n_257_76_16999;
   wire n_257_76_17000;
   wire n_257_76_17001;
   wire n_257_76_17002;
   wire n_257_76_17003;
   wire n_257_76_17004;
   wire n_257_76_17005;
   wire n_257_76_17006;
   wire n_257_76_17007;
   wire n_257_76_17008;
   wire n_257_76_17009;
   wire n_257_76_17010;
   wire n_257_76_17011;
   wire n_257_76_17012;
   wire n_257_76_17013;
   wire n_257_76_17014;
   wire n_257_76_17015;
   wire n_257_76_17016;
   wire n_257_76_17017;
   wire n_257_76_17018;
   wire n_257_76_17019;
   wire n_257_76_17020;
   wire n_257_76_17021;
   wire n_257_76_17022;
   wire n_257_76_17023;
   wire n_257_76_17024;
   wire n_257_76_17025;
   wire n_257_76_17026;
   wire n_257_76_17027;
   wire n_257_76_17028;
   wire n_257_76_17029;
   wire n_257_76_17030;
   wire n_257_76_17031;
   wire n_257_76_17032;
   wire n_257_76_17033;
   wire n_257_76_17034;
   wire n_257_76_17035;
   wire n_257_76_17036;
   wire n_257_76_17037;
   wire n_257_76_17038;
   wire n_257_76_17039;
   wire n_257_76_17040;
   wire n_257_76_17041;
   wire n_257_76_17042;
   wire n_257_76_17043;
   wire n_257_76_17044;
   wire n_257_76_17045;
   wire n_257_76_17046;
   wire n_257_76_17047;
   wire n_257_76_17048;
   wire n_257_76_17049;
   wire n_257_76_17050;
   wire n_257_76_17051;
   wire n_257_76_17052;
   wire n_257_76_17053;
   wire n_257_76_17054;
   wire n_257_76_17055;
   wire n_257_76_17056;
   wire n_257_76_17057;
   wire n_257_76_17058;
   wire n_257_76_17059;
   wire n_257_76_17060;
   wire n_257_76_17061;
   wire n_257_76_17062;
   wire n_257_76_17063;
   wire n_257_76_17064;
   wire n_257_76_17065;
   wire n_257_76_17066;
   wire n_257_76_17067;
   wire n_257_76_17068;
   wire n_257_76_17069;
   wire n_257_76_17070;
   wire n_257_76_17071;
   wire n_257_76_17072;
   wire n_257_76_17073;
   wire n_257_76_17074;
   wire n_257_76_17075;
   wire n_257_76_17076;
   wire n_257_76_17077;
   wire n_257_76_17078;
   wire n_257_76_17079;
   wire n_257_76_17080;
   wire n_257_76_17081;
   wire n_257_76_17082;
   wire n_257_76_17083;
   wire n_257_76_17084;
   wire n_257_76_17085;
   wire n_257_76_17086;
   wire n_257_76_17087;
   wire n_257_76_17088;
   wire n_257_76_17089;
   wire n_257_76_17090;
   wire n_257_76_17091;
   wire n_257_76_17092;
   wire n_257_76_17093;
   wire n_257_76_17094;
   wire n_257_76_17095;
   wire n_257_76_17096;
   wire n_257_76_17097;
   wire n_257_76_17098;
   wire n_257_76_17099;
   wire n_257_76_17100;
   wire n_257_76_17101;
   wire n_257_76_17102;
   wire n_257_76_17103;
   wire n_257_76_17104;
   wire n_257_76_17105;
   wire n_257_76_17106;
   wire n_257_76_17107;
   wire n_257_76_17108;
   wire n_257_76_17109;
   wire n_257_76_17110;
   wire n_257_76_17111;
   wire n_257_76_17112;
   wire n_257_76_17113;
   wire n_257_76_17114;
   wire n_257_76_17115;
   wire n_257_76_17116;
   wire n_257_76_17117;
   wire n_257_76_17118;
   wire n_257_76_17119;
   wire n_257_76_17120;
   wire n_257_76_17121;
   wire n_257_76_17122;
   wire n_257_76_17123;
   wire n_257_76_17124;
   wire n_257_76_17125;
   wire n_257_76_17126;
   wire n_257_76_17127;
   wire n_257_76_17128;
   wire n_257_76_17129;
   wire n_257_76_17130;
   wire n_257_76_17131;
   wire n_257_76_17132;
   wire n_257_76_17133;
   wire n_257_76_17134;
   wire n_257_76_17135;
   wire n_257_76_17136;
   wire n_257_76_17137;
   wire n_257_76_17138;
   wire n_257_76_17139;
   wire n_257_76_17140;
   wire n_257_76_17141;
   wire n_257_76_17142;
   wire n_257_76_17143;
   wire n_257_76_17144;
   wire n_257_76_17145;
   wire n_257_76_17146;
   wire n_257_76_17147;
   wire n_257_76_17148;
   wire n_257_76_17149;
   wire n_257_76_17150;
   wire n_257_76_17151;
   wire n_257_76_17152;
   wire n_257_76_17153;
   wire n_257_76_17154;
   wire n_257_76_17155;
   wire n_257_76_17156;
   wire n_257_76_17157;
   wire n_257_76_17158;
   wire n_257_76_17159;
   wire n_257_76_17160;
   wire n_257_76_17161;
   wire n_257_76_17162;
   wire n_257_76_17163;
   wire n_257_76_17164;
   wire n_257_76_17165;
   wire n_257_76_17166;
   wire n_257_76_17167;
   wire n_257_76_17168;
   wire n_257_76_17169;
   wire n_257_76_17170;
   wire n_257_76_17171;
   wire n_257_76_17172;
   wire n_257_76_17173;
   wire n_257_76_17174;
   wire n_257_76_17175;
   wire n_257_76_17176;
   wire n_257_76_17177;
   wire n_257_76_17178;
   wire n_257_76_17179;
   wire n_257_76_17180;
   wire n_257_76_17181;
   wire n_257_76_17182;
   wire n_257_76_17183;
   wire n_257_76_17184;
   wire n_257_76_17185;
   wire n_257_76_17186;
   wire n_257_76_17187;
   wire n_257_76_17188;
   wire n_257_76_17189;
   wire n_257_76_17190;
   wire n_257_76_17191;
   wire n_257_76_17192;
   wire n_257_76_17193;
   wire n_257_76_17194;
   wire n_257_76_17195;
   wire n_257_76_17196;
   wire n_257_76_17197;
   wire n_257_76_17198;
   wire n_257_76_17199;
   wire n_257_76_17200;
   wire n_257_76_17201;
   wire n_257_76_17202;
   wire n_257_76_17203;
   wire n_257_76_17204;
   wire n_257_76_17205;
   wire n_257_76_17206;
   wire n_257_76_17207;
   wire n_257_76_17208;
   wire n_257_76_17209;
   wire n_257_76_17210;
   wire n_257_76_17211;
   wire n_257_76_17212;
   wire n_257_76_17213;
   wire n_257_76_17214;
   wire n_257_76_17215;
   wire n_257_76_17216;
   wire n_257_76_17217;
   wire n_257_76_17218;
   wire n_257_76_17219;
   wire n_257_76_17220;
   wire n_257_76_17221;
   wire n_257_76_17222;
   wire n_257_76_17223;
   wire n_257_76_17224;
   wire n_257_76_17225;
   wire n_257_76_17226;
   wire n_257_76_17227;
   wire n_257_76_17228;
   wire n_257_76_17229;
   wire n_257_76_17230;
   wire n_257_76_17231;
   wire n_257_76_17232;
   wire n_257_76_17233;
   wire n_257_76_17234;
   wire n_257_76_17235;
   wire n_257_76_17236;
   wire n_257_76_17237;
   wire n_257_76_17238;
   wire n_257_76_17239;
   wire n_257_76_17240;
   wire n_257_76_17241;
   wire n_257_76_17242;
   wire n_257_76_17243;
   wire n_257_76_17244;
   wire n_257_76_17245;
   wire n_257_76_17246;
   wire n_257_76_17247;
   wire n_257_76_17248;
   wire n_257_76_17249;
   wire n_257_76_17250;
   wire n_257_76_17251;
   wire n_257_76_17252;
   wire n_257_76_17253;
   wire n_257_76_17254;
   wire n_257_76_17255;
   wire n_257_76_17256;
   wire n_257_76_17257;
   wire n_257_76_17258;
   wire n_257_76_17259;
   wire n_257_76_17260;
   wire n_257_76_17261;
   wire n_257_76_17262;
   wire n_257_76_17263;
   wire n_257_76_17264;
   wire n_257_76_17265;
   wire n_257_76_17266;
   wire n_257_76_17267;
   wire n_257_76_17268;
   wire n_257_76_17269;
   wire n_257_76_17270;
   wire n_257_76_17271;
   wire n_257_76_17272;
   wire n_257_76_17273;
   wire n_257_76_17274;
   wire n_257_76_17275;
   wire n_257_76_17276;
   wire n_257_76_17277;
   wire n_257_76_17278;
   wire n_257_76_17279;
   wire n_257_76_17280;
   wire n_257_76_17281;
   wire n_257_76_17282;
   wire n_257_76_17283;
   wire n_257_76_17284;
   wire n_257_76_17285;
   wire n_257_76_17286;
   wire n_257_76_17287;
   wire n_257_76_17288;
   wire n_257_76_17289;
   wire n_257_76_17290;
   wire n_257_76_17291;
   wire n_257_76_17292;
   wire n_257_76_17293;
   wire n_257_76_17294;
   wire n_257_76_17295;
   wire n_257_76_17296;
   wire n_257_76_17297;
   wire n_257_76_17298;
   wire n_257_76_17299;
   wire n_257_76_17300;
   wire n_257_76_17301;
   wire n_257_76_17302;
   wire n_257_76_17303;
   wire n_257_76_17304;
   wire n_257_76_17305;
   wire n_257_76_17306;
   wire n_257_76_17307;
   wire n_257_76_17308;
   wire n_257_76_17309;
   wire n_257_76_17310;
   wire n_257_76_17311;
   wire n_257_76_17312;
   wire n_257_76_17313;
   wire n_257_76_17314;
   wire n_257_76_17315;
   wire n_257_76_17316;
   wire n_257_76_17317;
   wire n_257_76_17318;
   wire n_257_76_17319;
   wire n_257_76_17320;
   wire n_257_76_17321;
   wire n_257_76_17322;
   wire n_257_76_17323;
   wire n_257_76_17324;
   wire n_257_76_17325;
   wire n_257_76_17326;
   wire n_257_76_17327;
   wire n_257_76_17328;
   wire n_257_76_17329;
   wire n_257_76_17330;
   wire n_257_76_17331;
   wire n_257_76_17332;
   wire n_257_76_17333;
   wire n_257_76_17334;
   wire n_257_76_17335;
   wire n_257_76_17336;
   wire n_257_76_17337;
   wire n_257_76_17338;
   wire n_257_76_17339;
   wire n_257_76_17340;
   wire n_257_76_17341;
   wire n_257_76_17342;
   wire n_257_76_17343;
   wire n_257_76_17344;
   wire n_257_76_17345;
   wire n_257_76_17346;
   wire n_257_76_17347;
   wire n_257_76_17348;
   wire n_257_76_17349;
   wire n_257_76_17350;
   wire n_257_76_17351;
   wire n_257_76_17352;
   wire n_257_76_17353;
   wire n_257_76_17354;
   wire n_257_76_17355;
   wire n_257_76_17356;
   wire n_257_76_17357;
   wire n_257_76_17358;
   wire n_257_76_17359;
   wire n_257_76_17360;
   wire n_257_76_17361;
   wire n_257_76_17362;
   wire n_257_76_17363;
   wire n_257_76_17364;
   wire n_257_76_17365;
   wire n_257_76_17366;
   wire n_257_76_17367;
   wire n_257_76_17368;
   wire n_257_76_17369;
   wire n_257_76_17370;
   wire n_257_76_17371;
   wire n_257_76_17372;
   wire n_257_76_17373;
   wire n_257_76_17374;
   wire n_257_76_17375;
   wire n_257_76_17376;
   wire n_257_76_17377;
   wire n_257_76_17378;
   wire n_257_76_17379;
   wire n_257_76_17380;
   wire n_257_76_17381;
   wire n_257_76_17382;
   wire n_257_76_17383;
   wire n_257_76_17384;
   wire n_257_76_17385;
   wire n_257_76_17386;
   wire n_257_76_17387;
   wire n_257_76_17388;
   wire n_257_76_17389;
   wire n_257_76_17390;
   wire n_257_76_17391;
   wire n_257_76_17392;
   wire n_257_76_17393;
   wire n_257_76_17394;
   wire n_257_76_17395;
   wire n_257_76_17396;
   wire n_257_76_17397;
   wire n_257_76_17398;
   wire n_257_76_17399;
   wire n_257_76_17400;
   wire n_257_76_17401;
   wire n_257_76_17402;
   wire n_257_76_17403;
   wire n_257_76_17404;
   wire n_257_76_17405;
   wire n_257_76_17406;
   wire n_257_76_17407;
   wire n_257_76_17408;
   wire n_257_76_17409;
   wire n_257_76_17410;
   wire n_257_76_17411;
   wire n_257_76_17412;
   wire n_257_76_17413;
   wire n_257_76_17414;
   wire n_257_76_17415;
   wire n_257_76_17416;
   wire n_257_76_17417;
   wire n_257_76_17418;
   wire n_257_76_17419;
   wire n_257_76_17420;
   wire n_257_76_17421;
   wire n_257_76_17422;
   wire n_257_76_17423;
   wire n_257_76_17424;
   wire n_257_76_17425;
   wire n_257_76_17426;
   wire n_257_76_17427;
   wire n_257_76_17428;
   wire n_257_76_17429;
   wire n_257_76_17430;
   wire n_257_76_17431;
   wire n_257_76_17432;
   wire n_257_76_17433;
   wire n_257_76_17434;
   wire n_257_76_17435;
   wire n_257_76_17436;
   wire n_257_76_17437;
   wire n_257_76_17438;
   wire n_257_76_17439;
   wire n_257_76_17440;
   wire n_257_76_17441;
   wire n_257_76_17442;
   wire n_257_76_17443;
   wire n_257_76_17444;
   wire n_257_76_17445;
   wire n_257_76_17446;
   wire n_257_76_17447;
   wire n_257_76_17448;
   wire n_257_76_17449;
   wire n_257_76_17450;
   wire n_257_76_17451;
   wire n_257_76_17452;
   wire n_257_76_17453;
   wire n_257_76_17454;
   wire n_257_76_17455;
   wire n_257_76_17456;
   wire n_257_76_17457;
   wire n_257_76_17458;
   wire n_257_76_17459;
   wire n_257_76_17460;
   wire n_257_76_17461;
   wire n_257_76_17462;
   wire n_257_76_17463;
   wire n_257_76_17464;
   wire n_257_76_17465;
   wire n_257_76_17466;
   wire n_257_76_17467;
   wire n_257_76_17468;
   wire n_257_76_17469;
   wire n_257_76_17470;
   wire n_257_76_17471;
   wire n_257_76_17472;
   wire n_257_76_17473;
   wire n_257_76_17474;
   wire n_257_76_17475;
   wire n_257_76_17476;
   wire n_257_76_17477;
   wire n_257_76_17478;
   wire n_257_76_17479;
   wire n_257_76_17480;
   wire n_257_76_17481;
   wire n_257_76_17482;
   wire n_257_76_17483;
   wire n_257_76_17484;
   wire n_257_76_17485;
   wire n_257_76_17486;
   wire n_257_76_17487;
   wire n_257_76_17488;
   wire n_257_76_17489;
   wire n_257_76_17490;
   wire n_257_76_17491;
   wire n_257_76_17492;
   wire n_257_76_17493;
   wire n_257_76_17494;
   wire n_257_76_17495;
   wire n_257_76_17496;
   wire n_257_76_17497;
   wire n_257_76_17498;
   wire n_257_76_17499;
   wire n_257_76_17500;
   wire n_257_76_17501;
   wire n_257_76_17502;
   wire n_257_76_17503;
   wire n_257_76_17504;
   wire n_257_76_17505;
   wire n_257_76_17506;
   wire n_257_76_17507;
   wire n_257_76_17508;
   wire n_257_76_17509;
   wire n_257_76_17510;
   wire n_257_76_17511;
   wire n_257_76_17512;
   wire n_257_76_17513;
   wire n_257_76_17514;
   wire n_257_76_17515;
   wire n_257_76_17516;
   wire n_257_76_17517;
   wire n_257_76_17518;
   wire n_257_76_17519;
   wire n_257_76_17520;
   wire n_257_76_17521;
   wire n_257_76_17522;
   wire n_257_76_17523;
   wire n_257_76_17524;
   wire n_257_76_17525;
   wire n_257_76_17526;
   wire n_257_76_17527;
   wire n_257_76_17528;
   wire n_257_76_17529;
   wire n_257_76_17530;
   wire n_257_76_17531;
   wire n_257_76_17532;
   wire n_257_76_17533;
   wire n_257_76_17534;
   wire n_257_76_17535;
   wire n_257_76_17536;
   wire n_257_76_17537;
   wire n_257_76_17538;
   wire n_257_76_17539;
   wire n_257_76_17540;
   wire n_257_76_17541;
   wire n_257_76_17542;
   wire n_257_76_17543;
   wire n_257_76_17544;
   wire n_257_76_17545;
   wire n_257_76_17546;
   wire n_257_76_17547;
   wire n_257_76_17548;
   wire n_257_76_17549;
   wire n_257_76_17550;
   wire n_257_76_17551;
   wire n_257_76_17552;
   wire n_257_76_17553;
   wire n_257_76_17554;
   wire n_257_76_17555;
   wire n_257_76_17556;
   wire n_257_76_17557;
   wire n_257_76_17558;
   wire n_257_76_17559;
   wire n_257_76_17560;
   wire n_257_76_17561;
   wire n_257_76_17562;
   wire n_257_76_17563;
   wire n_257_76_17564;
   wire n_257_76_17565;
   wire n_257_76_17566;
   wire n_257_76_17567;
   wire n_257_76_17568;
   wire n_257_76_17569;
   wire n_257_76_17570;
   wire n_257_76_17571;
   wire n_257_76_17572;
   wire n_257_76_17573;
   wire n_257_76_17574;
   wire n_257_76_17575;
   wire n_257_76_17576;
   wire n_257_76_17577;
   wire n_257_76_17578;
   wire n_257_76_17579;
   wire n_257_76_17580;
   wire n_257_76_17581;
   wire n_257_76_17582;
   wire n_257_76_17583;
   wire n_257_76_17584;
   wire n_257_76_17585;
   wire n_257_76_17586;
   wire n_257_76_17587;
   wire n_257_76_17588;
   wire n_257_76_17589;
   wire n_257_76_17590;
   wire n_257_76_17591;
   wire n_257_76_17592;
   wire n_257_76_17593;
   wire n_257_76_17594;
   wire n_257_76_17595;
   wire n_257_76_17596;
   wire n_257_76_17597;
   wire n_257_76_17598;
   wire n_257_76_17599;
   wire n_257_76_17600;
   wire n_257_76_17601;
   wire n_257_76_17602;
   wire n_257_76_17603;
   wire n_257_76_17604;
   wire n_257_76_17605;
   wire n_257_76_17606;
   wire n_257_76_17607;
   wire n_257_76_17608;
   wire n_257_76_17609;
   wire n_257_76_17610;
   wire n_257_76_17611;
   wire n_257_76_17612;
   wire n_257_76_17613;
   wire n_257_76_17614;
   wire n_257_76_17615;
   wire n_257_76_17616;
   wire n_257_76_17617;
   wire n_257_76_17618;
   wire n_257_76_17619;
   wire n_257_76_17620;
   wire n_257_76_17621;
   wire n_257_76_17622;
   wire n_257_76_17623;
   wire n_257_76_17624;
   wire n_257_76_17625;
   wire n_257_76_17626;
   wire n_257_76_17627;
   wire n_257_76_17628;
   wire n_257_76_17629;
   wire n_257_76_17630;
   wire n_257_76_17631;
   wire n_257_76_17632;
   wire n_257_76_17633;
   wire n_257_76_17634;
   wire n_257_76_17635;
   wire n_257_76_17636;
   wire n_257_76_17637;
   wire n_257_76_17638;
   wire n_257_76_17639;
   wire n_257_76_17640;
   wire n_257_76_17641;
   wire n_257_76_17642;
   wire n_257_76_17643;
   wire n_257_76_17644;
   wire n_257_76_17645;
   wire n_257_76_17646;
   wire n_257_76_17647;
   wire n_257_76_17648;
   wire n_257_76_17649;
   wire n_257_76_17650;
   wire n_257_76_17651;
   wire n_257_76_17652;
   wire n_257_76_17653;
   wire n_257_76_17654;
   wire n_257_76_17655;
   wire n_257_76_17656;
   wire n_257_76_17657;
   wire n_257_76_17658;
   wire n_257_76_17659;
   wire n_257_76_17660;
   wire n_257_76_17661;
   wire n_257_76_17662;
   wire n_257_76_17663;
   wire n_257_76_17664;
   wire n_257_76_17665;
   wire n_257_76_17666;
   wire n_257_76_17667;
   wire n_257_76_17668;
   wire n_257_76_17669;
   wire n_257_76_17670;
   wire n_257_76_17671;
   wire n_257_76_17672;
   wire n_257_76_17673;
   wire n_257_76_17674;
   wire n_257_76_17675;
   wire n_257_76_17676;
   wire n_257_76_17677;
   wire n_257_76_17678;
   wire n_257_76_17679;
   wire n_257_76_17680;
   wire n_257_76_17681;
   wire n_257_76_17682;
   wire n_257_76_17683;
   wire n_257_76_17684;
   wire n_257_76_17685;
   wire n_257_76_17686;
   wire n_257_76_17687;
   wire n_257_76_17688;
   wire n_257_76_17689;
   wire n_257_76_17690;
   wire n_257_76_17691;
   wire n_257_76_17692;
   wire n_257_76_17693;
   wire n_257_76_17694;
   wire n_257_76_17695;
   wire n_257_76_17696;
   wire n_257_76_17697;
   wire n_257_76_17698;
   wire n_257_76_17699;
   wire n_257_76_17700;
   wire n_257_76_17701;
   wire n_257_76_17702;
   wire n_257_76_17703;
   wire n_257_76_17704;
   wire n_257_76_17705;
   wire n_257_76_17706;
   wire n_257_76_17707;
   wire n_257_76_17708;
   wire n_257_76_17709;
   wire n_257_76_17710;
   wire n_257_76_17711;
   wire n_257_76_17712;
   wire n_257_76_17713;
   wire n_257_76_17714;
   wire n_257_76_17715;
   wire n_257_76_17716;
   wire n_257_76_17717;
   wire n_257_76_17718;
   wire n_257_76_17719;
   wire n_257_76_17720;
   wire n_257_76_17721;
   wire n_257_76_17722;
   wire n_257_76_17723;
   wire n_257_76_17724;
   wire n_257_76_17725;
   wire n_257_76_17726;
   wire n_257_76_17727;
   wire n_257_76_17728;
   wire n_257_76_17729;
   wire n_257_76_17730;
   wire n_257_76_17731;
   wire n_257_76_17732;
   wire n_257_76_17733;
   wire n_257_76_17734;
   wire n_257_76_17735;
   wire n_257_76_17736;
   wire n_257_76_17737;
   wire n_257_76_17738;
   wire n_257_76_17739;
   wire n_257_76_17740;
   wire n_257_76_17741;
   wire n_257_76_17742;
   wire n_257_76_17743;
   wire n_257_76_17744;
   wire n_257_76_17745;
   wire n_257_76_17746;
   wire n_257_76_17747;
   wire n_257_76_17748;
   wire n_257_76_17749;
   wire n_257_76_17750;
   wire n_257_76_17751;
   wire n_257_76_17752;
   wire n_257_76_17753;
   wire n_257_76_17754;
   wire n_257_76_17755;
   wire n_257_76_17756;
   wire n_257_76_17757;
   wire n_257_76_17758;
   wire n_257_76_17759;
   wire n_257_76_17760;
   wire n_257_76_17761;
   wire n_257_76_17762;
   wire n_257_76_17763;
   wire n_257_76_17764;
   wire n_257_76_17765;
   wire n_257_76_17766;
   wire n_257_76_17767;
   wire n_257_76_17768;
   wire n_257_76_17769;
   wire n_257_76_17770;
   wire n_257_76_17771;
   wire n_257_76_17772;
   wire n_257_76_17773;
   wire n_257_76_17774;
   wire n_257_76_17775;
   wire n_257_76_17776;
   wire n_257_76_17777;
   wire n_257_76_17778;
   wire n_257_76_17779;
   wire n_257_76_17780;
   wire n_257_76_17781;
   wire n_257_76_17782;
   wire n_257_76_17783;
   wire n_257_76_17784;
   wire n_257_76_17785;
   wire n_257_76_17786;
   wire n_257_76_17787;
   wire n_257_76_17788;
   wire n_257_76_17789;
   wire n_257_76_17790;
   wire n_257_76_17791;
   wire n_257_76_17792;
   wire n_257_76_17793;
   wire n_257_76_17794;
   wire n_257_76_17795;
   wire n_257_76_17796;
   wire n_257_76_17797;
   wire n_257_76_17798;
   wire n_257_76_17799;
   wire n_257_76_17800;
   wire n_257_76_17801;
   wire n_257_76_17802;
   wire n_257_76_17803;
   wire n_257_76_17804;
   wire n_257_76_17805;
   wire n_257_76_17806;
   wire n_257_76_17807;
   wire n_257_76_17808;
   wire n_257_76_17809;
   wire n_257_76_17810;
   wire n_257_76_17811;
   wire n_257_76_17812;
   wire n_257_76_17813;
   wire n_257_76_17814;
   wire n_257_76_17815;
   wire n_257_76_17816;
   wire n_257_76_17817;
   wire n_257_76_17818;
   wire n_257_76_17819;
   wire n_257_76_17820;
   wire n_257_76_17821;
   wire n_257_76_17822;
   wire n_257_76_17823;
   wire n_257_76_17824;
   wire n_257_76_17825;
   wire n_257_76_17826;
   wire n_257_76_17827;
   wire n_257_76_17828;
   wire n_257_76_17829;
   wire n_257_76_17830;
   wire n_257_76_17831;
   wire n_257_76_17832;
   wire n_257_76_17833;
   wire n_257_76_17834;
   wire n_257_76_17835;
   wire n_257_76_17836;
   wire n_257_76_17837;
   wire n_257_76_17838;
   wire n_257_76_17839;
   wire n_257_76_17840;
   wire n_257_76_17841;
   wire n_257_76_17842;
   wire n_257_76_17843;
   wire n_257_76_17844;
   wire n_257_76_17845;
   wire n_257_76_17846;
   wire n_257_76_17847;
   wire n_257_76_17848;
   wire n_257_76_17849;
   wire n_257_76_17850;
   wire n_257_76_17851;
   wire n_257_76_17852;
   wire n_257_76_17853;
   wire n_257_76_17854;
   wire n_257_76_17855;
   wire n_257_76_17856;
   wire n_257_76_17857;
   wire n_257_76_17858;
   wire n_257_76_17859;
   wire n_257_76_17860;
   wire n_257_76_17861;
   wire n_257_76_17862;
   wire n_257_76_17863;
   wire n_257_76_17864;
   wire n_257_76_17865;
   wire n_257_76_17866;
   wire n_257_76_17867;
   wire n_257_76_17868;
   wire n_257_76_17869;
   wire n_257_76_17870;
   wire n_257_76_17871;
   wire n_257_76_17872;
   wire n_257_76_17873;
   wire n_257_76_17874;
   wire n_257_76_17875;
   wire n_257_76_17876;
   wire n_257_76_17877;
   wire n_257_76_17878;
   wire n_257_76_17879;
   wire n_257_76_17880;
   wire n_257_76_17881;
   wire n_257_76_17882;
   wire n_257_76_17883;
   wire n_257_76_17884;
   wire n_257_76_17885;
   wire n_257_76_17886;
   wire n_257_76_17887;
   wire n_257_76_17888;
   wire n_257_76_17889;
   wire n_257_76_17890;
   wire n_257_76_17891;
   wire n_257_76_17892;
   wire n_257_76_17893;
   wire n_257_76_17894;
   wire n_257_76_17895;
   wire n_257_76_17896;
   wire n_257_76_17897;
   wire n_257_76_17898;
   wire n_257_76_17899;
   wire n_257_76_17900;
   wire n_257_76_17901;
   wire n_257_76_17902;
   wire n_257_76_17903;
   wire n_257_76_17904;
   wire n_257_76_17905;
   wire n_257_76_17906;
   wire n_257_76_17907;
   wire n_257_76_17908;
   wire n_257_76_17909;
   wire n_257_76_17910;
   wire n_257_76_17911;
   wire n_257_76_17912;
   wire n_257_76_17913;
   wire n_257_76_17914;
   wire n_257_76_17915;
   wire n_257_76_17916;
   wire n_257_76_17917;
   wire n_257_76_17918;
   wire n_257_76_17919;
   wire n_257_76_17920;
   wire n_257_76_17921;
   wire n_257_76_17922;
   wire n_257_76_17923;
   wire n_257_76_17924;
   wire n_257_76_17925;
   wire n_257_76_17926;
   wire n_257_76_17927;
   wire n_257_76_17928;
   wire n_257_76_17929;
   wire n_257_76_17930;
   wire n_257_76_17931;
   wire n_257_76_17932;
   wire n_257_76_17933;
   wire n_257_76_17934;
   wire n_257_76_17935;
   wire n_257_76_17936;
   wire n_257_76_17937;
   wire n_257_76_17938;
   wire n_257_76_17939;
   wire n_257_76_17940;
   wire n_257_76_17941;
   wire n_257_76_17942;
   wire n_257_76_17943;
   wire n_257_76_17944;
   wire n_257_76_17945;
   wire n_257_76_17946;
   wire n_257_76_17947;
   wire n_257_76_17948;
   wire n_257_76_17949;
   wire n_257_76_17950;
   wire n_257_76_17951;
   wire n_257_76_17952;
   wire n_257_76_17953;
   wire n_257_76_17954;
   wire n_257_76_17955;
   wire n_257_76_17956;
   wire n_257_76_17957;
   wire n_257_76_17958;
   wire n_257_76_17959;
   wire n_257_76_17960;
   wire n_257_76_17961;
   wire n_257_76_17962;
   wire n_257_76_17963;
   wire n_257_76_17964;
   wire n_257_76_17965;
   wire n_257_76_17966;
   wire n_257_76_17967;
   wire n_257_76_17968;
   wire n_257_76_17969;
   wire n_257_76_17970;
   wire n_257_76_17971;
   wire n_257_76_17972;
   wire n_257_76_17973;
   wire n_257_76_17974;
   wire n_257_76_17975;
   wire n_257_76_17976;
   wire n_257_76_17977;
   wire n_257_76_17978;
   wire n_257_76_17979;
   wire n_257_76_17980;
   wire n_257_76_17981;
   wire n_257_76_17982;
   wire n_257_76_17983;
   wire n_257_76_17984;
   wire n_257_76_17985;
   wire n_257_76_17986;
   wire n_257_76_17987;
   wire n_257_76_17988;
   wire n_257_76_17989;
   wire n_257_76_17990;
   wire n_257_76_17991;
   wire n_257_76_17992;
   wire n_257_76_17993;
   wire n_257_76_17994;
   wire n_257_76_17995;
   wire n_257_76_17996;
   wire n_257_76_17997;
   wire n_257_76_17998;
   wire n_257_76_17999;
   wire n_257_76_18000;
   wire n_257_76_18001;
   wire n_257_76_18002;
   wire n_257_76_18003;
   wire n_257_76_18004;
   wire n_257_76_18005;
   wire n_257_76_18006;
   wire n_257_76_18007;
   wire n_257_76_18008;
   wire n_257_76_18009;
   wire n_257_76_18010;
   wire n_257_76_18011;
   wire n_257_76_18012;
   wire n_257_76_18013;
   wire n_257_76_18014;
   wire n_257_76_18015;
   wire n_257_76_18016;
   wire n_257_76_18017;
   wire n_257_76_18018;
   wire n_257_76_18019;
   wire n_257_76_18020;
   wire n_257_76_18021;
   wire n_257_76_18022;
   wire n_257_76_18023;
   wire n_257_76_18024;
   wire n_257_76_18025;
   wire n_257_76_18026;
   wire n_257_76_18027;
   wire n_257_76_18028;
   wire n_257_76_18029;
   wire n_257_76_18030;
   wire n_257_76_18031;
   wire n_257_76_18032;
   wire n_257_76_18033;
   wire n_257_76_18034;
   wire n_257_76_18035;
   wire n_257_76_18036;
   wire n_257_76_18037;
   wire n_257_76_18038;
   wire n_257_76_18039;
   wire n_257_76_18040;
   wire n_257_76_18041;
   wire n_257_76_18042;
   wire n_257_76_18043;
   wire n_257_76_18044;
   wire n_257_76_18045;
   wire n_257_76_18046;
   wire n_257_76_18047;
   wire n_257_76_18048;
   wire n_257_76_18049;
   wire n_257_76_18050;
   wire n_257_76_18051;
   wire n_257_76_18052;
   wire n_257_76_18053;
   wire n_257_76_18054;
   wire n_257_76_18055;
   wire n_257_76_18056;
   wire n_257_76_18057;
   wire n_257_76_18058;
   wire n_257_76_18059;
   wire n_257_76_18060;
   wire n_257_76_18061;
   wire n_257_76_18062;
   wire n_257_76_18063;
   wire n_257_76_18064;
   wire n_257_76_18065;
   wire n_257_76_18066;
   wire n_257_76_18067;
   wire n_257_76_18068;
   wire n_257_76_18069;
   wire n_257_76_18070;
   wire n_257_76_18071;
   wire n_257_76_18072;
   wire n_257_76_18073;
   wire n_257_76_18074;
   wire n_257_76_18075;
   wire n_257_76_18076;
   wire n_257_76_18077;
   wire n_257_76_18078;
   wire n_257_76_18079;
   wire n_257_76_18080;
   wire n_257_76_18081;
   wire n_257_76_18082;
   wire n_257_76_18083;
   wire n_257_76_18084;
   wire n_257_76_18085;
   wire n_2_0;
   wire n_2_1;
   wire n_2_2;
   wire n_2_3;
   wire n_2_4;
   wire n_2_5;
   wire n_2_6;
   wire n_2_7;
   wire n_2_8;
   wire n_2_9;
   wire n_2_10;
   wire n_2_11;
   wire n_2_12;
   wire n_2_13;
   wire n_2_14;
   wire n_2_15;
   wire n_2_16;
   wire n_2_17;
   wire n_2_18;
   wire n_2_19;
   wire n_2_20;
   wire n_2_21;
   wire n_2_22;
   wire n_2_23;
   wire n_2_24;
   wire n_2_25;
   wire n_2_26;
   wire n_2_27;
   wire n_2_28;
   wire n_2_29;
   wire n_2_30;
   wire n_2_31;
   wire n_2_32;
   wire n_2_33;
   wire n_2_34;
   wire n_2_35;
   wire n_2_36;
   wire n_2_37;
   wire n_2_38;
   wire n_2_39;
   wire n_2_40;
   wire n_2_41;
   wire n_2_42;
   wire n_2_43;
   wire n_2_44;
   wire n_2_45;
   wire n_2_46;
   wire n_2_47;
   wire n_2_48;
   wire n_2_49;
   wire n_2_50;
   wire n_2_51;
   wire n_2_52;
   wire n_2_53;
   wire n_2_54;
   wire n_2_55;
   wire n_2_56;
   wire n_2_57;
   wire n_2_58;
   wire n_2_59;
   wire n_2_60;
   wire n_2_61;
   wire n_2_62;
   wire n_2_63;
   wire n_2_64;
   wire n_2_65;
   wire n_2_66;
   wire n_2_67;
   wire n_2_68;
   wire n_2_69;
   wire n_2_70;
   wire n_2_2_0;
   wire n_2_71;
   wire n_2_2_1;
   wire n_2_72;
   wire n_2_2_2;
   wire n_2_73;
   wire n_2_2_3;
   wire n_2_74;
   wire n_2_2_4;
   wire n_2_75;
   wire n_2_2_5;
   wire n_2_76;
   wire n_2_2_6;
   wire n_2_77;
   wire n_2_2_7;
   wire n_2_78;
   wire n_2_2_8;
   wire n_2_79;
   wire n_2_2_9;
   wire n_2_80;
   wire n_2_2_10;
   wire n_2_81;
   wire n_2_2_11;
   wire n_2_82;
   wire n_2_2_12;
   wire n_2_83;
   wire n_2_2_13;
   wire n_2_84;
   wire n_2_2_14;
   wire n_2_85;
   wire n_2_2_15;
   wire n_2_86;
   wire n_2_2_16;
   wire n_2_87;
   wire n_2_2_17;
   wire n_2_88;
   wire n_2_2_18;
   wire n_2_91;
   wire n_2_2_19;
   wire n_2_95;
   wire n_2_2_20;
   wire n_2_98;
   wire n_2_89;
   wire n_2_90;
   wire n_2_92;
   wire n_2_2_21;
   wire n_2_2_22;
   wire n_2_93;
   wire n_2_2_23;
   wire n_2_2_24;
   wire n_2_94;
   wire n_2_96;
   wire n_2_2_25;
   wire n_2_2_26;
   wire n_2_97;
   wire n_2_99;
   wire n_2_2_27;
   wire n_2_2_28;
   wire n_2_100;
   wire n_2_2_29;
   wire n_2_2_30;
   wire n_2_101;
   wire n_2_2_31;
   wire n_2_2_32;
   wire n_2_2_33;
   wire n_2_102;
   wire n_2_4_0;
   wire n_2_4_1;
   wire n_2_4_2;
   wire n_2_4_3;
   wire n_2_4_4;
   wire n_2_4_5;
   wire n_2_4_6;
   wire n_2_4_7;
   wire n_2_4_8;
   wire n_2_4_9;
   wire n_2_4_10;
   wire n_2_4_11;
   wire n_2_4_12;
   wire n_2_4_13;
   wire n_2_4_14;
   wire n_2_4_15;
   wire n_2_4_16;
   wire n_2_4_17;
   wire n_2_4_18;
   wire n_2_4_19;
   wire n_2_4_20;
   wire n_2_4_21;
   wire n_2_4_22;
   wire n_2_4_23;
   wire n_2_4_24;
   wire n_2_4_25;
   wire n_2_4_26;
   wire n_2_4_27;
   wire n_2_4_28;
   wire n_2_4_29;
   wire n_2_4_30;
   wire n_2_4_31;
   wire n_2_4_32;
   wire n_2_4_33;
   wire n_2_4_34;
   wire n_2_103;
   wire n_2_104;
   wire n_2_105;
   wire n_2_6_0;
   wire n_2_106;
   wire n_2_6_1;
   wire n_2_107;
   wire n_2_6_2;
   wire n_2_108;
   wire n_2_6_3;
   wire n_2_109;
   wire n_2_6_4;
   wire n_2_110;
   wire n_2_7_0;
   wire n_2_7_1;
   wire n_2_7_2;
   wire n_2_7_3;
   wire n_2_7_4;
   wire n_2_7_5;
   wire n_2_111;
   wire n_2_8_0;
   wire n_2_8_1;
   wire n_2_8_2;
   wire n_2_9_0;
   wire n_2_117;
   wire n_2_9_1;
   wire n_2_118;
   wire n_2_9_2;
   wire n_2_119;
   wire n_2_9_3;
   wire n_2_120;
   wire n_2_9_4;
   wire n_2_121;
   wire n_2_9_5;
   wire n_2_122;
   wire n_2_9_6;
   wire n_2_123;
   wire n_2_9_7;
   wire n_2_9_8;
   wire n_2_112;
   wire n_2_9_9;
   wire n_2_113;
   wire n_2_9_10;
   wire n_2_114;
   wire n_2_9_11;
   wire n_2_115;
   wire n_2_9_12;
   wire n_2_116;
   wire n_2_9_13;
   wire n_2_10_0;
   wire n_2_124;
   wire n_2_10_1;
   wire n_2_127;
   wire n_2_10_2;
   wire n_2_128;
   wire n_2_10_3;
   wire n_2_132;
   wire n_2_10_4;
   wire n_2_135;
   wire n_2_10_5;
   wire n_2_137;
   wire n_2_10_6;
   wire n_2_138;
   wire n_2_10_7;
   wire n_2_140;
   wire n_2_10_8;
   wire n_2_141;
   wire n_2_10_9;
   wire n_2_142;
   wire n_2_10_10;
   wire n_2_143;
   wire n_2_10_11;
   wire n_2_144;
   wire n_2_10_12;
   wire n_2_145;
   wire n_2_10_13;
   wire n_2_146;
   wire n_2_10_14;
   wire n_2_147;
   wire n_2_10_15;
   wire n_2_148;
   wire n_2_10_16;
   wire n_2_150;
   wire n_2_10_17;
   wire n_2_152;
   wire n_2_10_18;
   wire n_2_153;
   wire n_2_10_19;
   wire n_2_154;
   wire n_2_10_20;
   wire n_2_155;
   wire n_2_125;
   wire n_2_10_21;
   wire n_2_10_22;
   wire n_2_126;
   wire n_2_10_23;
   wire n_2_10_24;
   wire n_2_129;
   wire n_2_10_25;
   wire n_2_10_26;
   wire n_2_130;
   wire n_2_10_27;
   wire n_2_10_28;
   wire n_2_131;
   wire n_2_10_29;
   wire n_2_10_30;
   wire n_2_133;
   wire n_2_10_31;
   wire n_2_10_32;
   wire n_2_134;
   wire n_2_10_33;
   wire n_2_10_34;
   wire n_2_136;
   wire n_2_10_35;
   wire n_2_10_36;
   wire n_2_139;
   wire n_2_10_37;
   wire n_2_10_38;
   wire n_2_149;
   wire n_2_10_39;
   wire n_2_10_40;
   wire n_2_151;
   wire n_2_10_41;
   wire n_2_10_42;
   wire n_2_10_43;
   wire n_2_156;
   wire n_2_157;
   wire n_2_158;
   wire n_2_159;
   wire n_2_160;
   wire n_2_161;
   wire n_2_162;
   wire n_2_163;
   wire n_2_164;
   wire n_2_165;
   wire n_2_166;
   wire n_2_167;
   wire n_2_168;
   wire n_2_169;
   wire n_2_15_0;
   wire n_2_15_1;
   wire n_2_15_2;
   wire n_2_15_3;
   wire n_2_15_4;
   wire n_2_16_0;
   wire n_2_16_1;
   wire n_2_16_2;
   wire n_2_16_3;
   wire n_2_16_4;
   wire n_2_16_5;
   wire n_2_16_6;
   wire n_2_16_7;
   wire n_2_17_0;
   wire n_2_17_1;
   wire n_2_17_2;
   wire n_2_17_3;
   wire n_2_17_4;
   wire n_2_17_5;
   wire n_2_17_6;
   wire n_2_17_7;
   wire n_2_17_8;
   wire n_2_17_9;
   wire n_2_17_10;
   wire n_2_17_11;
   wire n_2_17_12;
   wire n_2_17_13;
   wire n_2_17_14;
   wire n_2_17_15;
   wire n_2_17_16;
   wire n_2_17_17;
   wire n_2_17_18;
   wire n_2_17_19;
   wire n_2_17_20;
   wire n_2_17_21;
   wire n_2_17_22;
   wire n_2_17_23;
   wire n_2_17_24;
   wire n_2_17_25;
   wire n_2_17_26;
   wire n_2_17_27;
   wire n_2_17_28;
   wire n_2_17_29;
   wire n_2_17_30;
   wire n_2_17_31;
   wire n_2_17_32;
   wire n_2_17_33;
   wire n_2_17_34;
   wire n_2_17_35;
   wire n_2_17_36;
   wire n_2_17_37;
   wire n_2_17_38;
   wire n_2_17_39;
   wire n_2_17_40;
   wire n_2_17_41;
   wire n_2_17_42;
   wire n_2_17_43;
   wire n_2_17_44;
   wire n_2_17_45;
   wire n_2_17_46;
   wire n_2_17_47;
   wire n_2_17_48;
   wire n_2_17_49;
   wire n_2_17_50;
   wire n_2_17_51;
   wire n_2_17_52;
   wire n_2_17_53;
   wire n_2_17_54;
   wire n_2_17_55;
   wire n_2_17_56;
   wire n_2_17_57;
   wire n_2_17_58;
   wire n_2_17_59;
   wire n_2_17_60;
   wire n_2_17_61;
   wire n_2_17_62;
   wire n_2_17_63;
   wire n_2_17_64;
   wire n_2_17_65;
   wire n_2_17_66;
   wire n_2_17_67;
   wire n_2_17_68;
   wire n_2_17_69;
   wire n_2_17_70;
   wire n_2_17_71;
   wire n_2_17_72;
   wire n_2_17_73;
   wire n_2_17_74;
   wire n_2_17_75;
   wire n_2_17_76;
   wire n_2_17_77;
   wire n_2_17_78;
   wire n_2_17_79;
   wire n_2_17_80;
   wire n_2_17_81;
   wire n_2_17_82;
   wire n_2_17_83;
   wire n_2_17_84;
   wire n_2_17_85;
   wire n_2_17_86;
   wire n_2_17_87;
   wire n_2_17_88;
   wire n_2_17_89;
   wire n_2_17_90;
   wire n_2_17_91;
   wire n_2_17_92;
   wire n_2_17_93;
   wire n_2_17_94;
   wire n_2_17_95;
   wire n_2_17_96;
   wire n_2_17_97;
   wire n_2_17_98;
   wire n_2_17_99;
   wire n_2_17_100;
   wire n_2_17_101;
   wire n_2_17_102;
   wire n_2_17_103;
   wire n_2_17_104;
   wire n_2_17_105;
   wire n_2_17_106;
   wire n_2_17_107;
   wire n_2_17_108;
   wire n_2_17_109;
   wire n_2_17_110;
   wire n_2_17_111;
   wire n_2_17_112;
   wire n_2_17_113;
   wire n_2_17_114;
   wire n_2_17_115;
   wire n_2_17_116;
   wire n_2_17_117;
   wire n_2_17_118;
   wire n_2_17_119;
   wire n_2_17_120;
   wire n_2_17_121;
   wire n_2_209;
   wire n_2_18_0;
   wire n_2_210;
   wire n_2_18_1;
   wire n_2_211;
   wire n_2_18_2;
   wire n_2_212;
   wire n_2_18_3;
   wire n_2_185;
   wire n_2_18_4;
   wire n_2_186;
   wire n_2_18_5;
   wire n_2_189;
   wire n_2_18_6;
   wire n_2_190;
   wire n_2_18_7;
   wire n_2_191;
   wire n_2_18_8;
   wire n_2_192;
   wire n_2_18_9;
   wire n_2_193;
   wire n_2_18_10;
   wire n_2_194;
   wire n_2_18_11;
   wire n_2_195;
   wire n_2_18_12;
   wire n_2_18_13;
   wire n_2_18_14;
   wire n_2_18_15;
   wire n_2_18_16;
   wire n_2_172;
   wire n_2_18_17;
   wire n_2_173;
   wire n_2_18_18;
   wire n_2_174;
   wire n_2_18_19;
   wire n_2_175;
   wire n_2_18_20;
   wire n_2_176;
   wire n_2_18_21;
   wire n_2_177;
   wire n_2_18_22;
   wire n_2_178;
   wire n_2_18_23;
   wire n_2_179;
   wire n_2_18_24;
   wire n_2_180;
   wire n_2_18_25;
   wire n_2_181;
   wire n_2_18_26;
   wire n_2_182;
   wire n_2_18_27;
   wire n_2_18_28;
   wire n_2_199;
   wire n_2_18_29;
   wire n_2_18_30;
   wire n_2_198;
   wire n_2_18_31;
   wire n_2_18_32;
   wire n_2_18_33;
   wire n_2_18_34;
   wire n_2_18_35;
   wire n_2_18_36;
   wire n_2_18_37;
   wire n_2_18_38;
   wire n_2_18_39;
   wire n_2_18_40;
   wire n_2_18_41;
   wire n_2_18_42;
   wire n_2_18_43;
   wire n_2_18_44;
   wire n_2_18_45;
   wire n_2_18_46;
   wire n_2_18_47;
   wire n_2_18_48;
   wire n_2_18_49;
   wire n_2_18_50;
   wire n_2_18_51;
   wire n_2_18_52;
   wire n_2_18_53;
   wire n_2_18_54;
   wire n_2_18_55;
   wire n_2_18_56;
   wire n_2_18_57;
   wire n_2_18_58;
   wire n_2_18_59;
   wire n_2_18_60;
   wire n_2_18_61;
   wire n_2_18_62;
   wire n_2_18_63;
   wire n_2_18_64;
   wire n_2_18_65;
   wire n_2_18_66;
   wire n_2_18_67;
   wire n_2_18_68;
   wire n_2_18_69;
   wire n_2_18_70;
   wire n_2_18_71;
   wire n_2_18_72;
   wire n_2_18_73;
   wire n_2_18_74;
   wire n_2_18_75;
   wire n_2_18_76;
   wire n_2_18_77;
   wire n_2_18_78;
   wire n_2_18_79;
   wire n_2_18_80;
   wire n_2_18_81;
   wire n_2_18_82;
   wire n_2_18_83;
   wire n_2_18_84;
   wire n_2_18_85;
   wire n_2_18_86;
   wire n_2_18_87;
   wire n_2_18_88;
   wire n_2_18_89;
   wire n_2_18_90;
   wire n_2_18_91;
   wire n_2_18_92;
   wire n_2_18_93;
   wire n_2_18_94;
   wire n_2_18_95;
   wire n_2_18_96;
   wire n_2_18_97;
   wire n_2_18_98;
   wire n_2_18_99;
   wire n_2_18_100;
   wire n_2_18_101;
   wire n_2_18_102;
   wire n_2_18_103;
   wire n_2_18_104;
   wire n_2_18_105;
   wire n_2_18_106;
   wire n_2_18_107;
   wire n_2_18_108;
   wire n_2_18_109;
   wire n_2_18_110;
   wire n_2_18_111;
   wire n_2_18_112;
   wire n_2_18_113;
   wire n_2_18_114;
   wire n_2_18_115;
   wire n_2_18_116;
   wire n_2_18_117;
   wire n_2_18_118;
   wire n_2_18_119;
   wire n_2_18_120;
   wire n_2_18_121;
   wire n_2_18_122;
   wire n_2_18_123;
   wire n_2_18_124;
   wire n_2_18_125;
   wire n_2_18_126;
   wire n_2_18_127;
   wire n_2_18_128;
   wire n_2_18_129;
   wire n_2_18_130;
   wire n_2_18_131;
   wire n_2_18_132;
   wire n_2_18_133;
   wire n_2_18_134;
   wire n_2_18_135;
   wire n_2_18_136;
   wire n_2_18_137;
   wire n_2_183;
   wire n_2_18_138;
   wire n_2_18_139;
   wire n_2_18_140;
   wire n_2_18_141;
   wire n_2_18_142;
   wire n_2_18_143;
   wire n_2_18_144;
   wire n_2_18_145;
   wire n_2_18_146;
   wire n_2_18_147;
   wire n_2_18_148;
   wire n_2_18_149;
   wire n_2_18_150;
   wire n_2_18_151;
   wire n_2_18_152;
   wire n_2_18_153;
   wire n_2_18_154;
   wire n_2_18_155;
   wire n_2_188;
   wire n_2_18_156;
   wire n_2_18_157;
   wire n_2_187;
   wire n_2_18_158;
   wire n_2_18_159;
   wire n_2_18_160;
   wire n_2_18_161;
   wire n_2_18_162;
   wire n_2_18_163;
   wire n_2_18_164;
   wire n_2_18_165;
   wire n_2_18_166;
   wire n_2_18_167;
   wire n_2_18_168;
   wire n_2_18_169;
   wire n_2_18_170;
   wire n_2_18_171;
   wire n_2_18_172;
   wire n_2_18_173;
   wire n_2_18_174;
   wire n_2_18_175;
   wire n_2_18_176;
   wire n_2_18_177;
   wire n_2_196;
   wire n_2_197;
   wire n_2_18_178;
   wire n_2_18_179;
   wire n_2_18_180;
   wire n_2_18_181;
   wire n_2_18_182;
   wire n_2_18_183;
   wire n_2_18_184;
   wire n_2_18_185;
   wire n_2_18_186;
   wire n_2_18_187;
   wire n_2_18_188;
   wire n_2_18_189;
   wire n_2_18_190;
   wire n_2_217;
   wire n_2_18_191;
   wire n_2_18_192;
   wire n_2_18_193;
   wire n_2_18_194;
   wire n_2_218;
   wire n_2_18_195;
   wire n_2_18_196;
   wire n_2_18_197;
   wire n_2_18_198;
   wire n_2_18_199;
   wire n_2_18_200;
   wire n_2_18_201;
   wire n_2_18_202;
   wire n_2_18_203;
   wire n_2_18_204;
   wire n_2_219;
   wire n_2_18_205;
   wire n_2_18_206;
   wire n_2_18_207;
   wire n_2_18_208;
   wire n_2_18_209;
   wire n_2_220;
   wire n_2_18_210;
   wire n_2_18_211;
   wire n_2_18_212;
   wire n_2_18_213;
   wire n_2_18_214;
   wire n_2_18_215;
   wire n_2_221;
   wire n_2_18_216;
   wire n_2_18_217;
   wire n_2_18_218;
   wire n_2_18_219;
   wire n_2_18_220;
   wire n_2_222;
   wire n_2_18_221;
   wire n_2_18_222;
   wire n_2_18_223;
   wire n_2_18_224;
   wire n_2_18_225;
   wire n_2_18_226;
   wire n_2_18_227;
   wire n_2_18_228;
   wire n_2_223;
   wire n_2_18_229;
   wire n_2_18_230;
   wire n_2_18_231;
   wire n_2_18_232;
   wire n_2_18_233;
   wire n_2_18_234;
   wire n_2_18_235;
   wire n_2_224;
   wire n_2_18_236;
   wire n_2_18_237;
   wire n_2_18_238;
   wire n_2_18_239;
   wire n_2_18_240;
   wire n_2_18_241;
   wire n_2_18_242;
   wire n_2_18_243;
   wire n_2_18_244;
   wire n_2_225;
   wire n_2_18_245;
   wire n_2_18_246;
   wire n_2_18_247;
   wire n_2_18_248;
   wire n_2_18_249;
   wire n_2_18_250;
   wire n_2_18_251;
   wire n_2_18_252;
   wire n_2_18_253;
   wire n_2_18_254;
   wire n_2_18_255;
   wire n_2_18_256;
   wire n_2_18_257;
   wire n_2_18_258;
   wire n_2_18_259;
   wire n_2_18_260;
   wire n_2_18_261;
   wire n_2_18_262;
   wire n_2_18_263;
   wire n_2_18_264;
   wire n_2_18_265;
   wire n_2_18_266;
   wire n_2_18_267;
   wire n_2_18_268;
   wire n_2_18_269;
   wire n_2_18_270;
   wire n_2_18_271;
   wire n_2_18_272;
   wire n_2_18_273;
   wire n_2_18_274;
   wire n_2_18_275;
   wire n_2_18_276;
   wire n_2_18_277;
   wire n_2_18_278;
   wire n_2_18_279;
   wire n_2_18_280;
   wire n_2_18_281;
   wire n_2_18_282;
   wire n_2_18_283;
   wire n_2_18_284;
   wire n_2_18_285;
   wire n_2_18_286;
   wire n_2_18_287;
   wire n_2_18_288;
   wire n_2_18_289;
   wire n_2_18_290;
   wire n_2_18_291;
   wire n_2_18_292;
   wire n_2_18_293;
   wire n_2_18_294;
   wire n_2_18_295;
   wire n_2_18_296;
   wire n_2_18_297;
   wire n_2_18_298;
   wire n_2_18_299;
   wire n_2_18_300;
   wire n_2_18_301;
   wire n_2_18_302;
   wire n_2_18_303;
   wire n_2_18_304;
   wire n_2_18_305;
   wire n_2_18_306;
   wire n_2_18_307;
   wire n_2_18_308;
   wire n_2_18_309;
   wire n_2_18_310;
   wire n_2_18_311;
   wire n_2_18_312;
   wire n_2_18_313;
   wire n_2_18_314;
   wire n_2_18_315;
   wire n_2_18_316;
   wire n_2_18_317;
   wire n_2_18_318;
   wire n_2_18_319;
   wire n_2_18_320;
   wire n_2_18_321;
   wire n_2_18_322;
   wire n_2_18_323;
   wire n_2_18_324;
   wire n_2_18_325;
   wire n_2_18_326;
   wire n_2_18_327;
   wire n_2_18_328;
   wire n_2_18_329;
   wire n_2_18_330;
   wire n_2_18_331;
   wire n_2_18_332;
   wire n_2_18_333;
   wire n_2_18_334;
   wire n_2_18_335;
   wire n_2_18_336;
   wire n_2_18_337;
   wire n_2_18_338;
   wire n_2_18_339;
   wire n_2_18_340;
   wire n_2_18_341;
   wire n_2_18_342;
   wire n_2_18_343;
   wire n_2_18_344;
   wire n_2_18_345;
   wire n_2_18_346;
   wire n_2_18_347;
   wire n_2_18_348;
   wire n_2_18_349;
   wire n_2_18_350;
   wire n_2_18_351;
   wire n_2_18_352;
   wire n_2_18_353;
   wire n_2_18_354;
   wire n_2_18_355;
   wire n_2_18_356;
   wire n_2_18_357;
   wire n_2_18_358;
   wire n_2_18_359;
   wire n_2_18_360;
   wire n_2_18_361;
   wire n_2_18_362;
   wire n_2_18_363;
   wire n_2_18_364;
   wire n_2_18_365;
   wire n_2_18_366;
   wire n_2_18_367;
   wire n_2_18_368;
   wire n_2_18_369;
   wire n_2_18_370;
   wire n_2_18_371;
   wire n_2_18_372;
   wire n_2_18_373;
   wire n_2_18_374;
   wire n_2_18_375;
   wire n_2_18_376;
   wire n_2_18_377;
   wire n_2_18_378;
   wire n_2_18_379;
   wire n_2_18_380;
   wire n_2_18_381;
   wire n_2_18_382;
   wire n_2_18_383;
   wire n_2_18_384;
   wire n_2_18_385;
   wire n_2_18_386;
   wire n_2_18_387;
   wire n_2_18_388;
   wire n_2_18_389;
   wire n_2_18_390;
   wire n_2_18_391;
   wire n_2_18_392;
   wire n_2_18_393;
   wire n_2_18_394;
   wire n_2_18_395;
   wire n_2_18_396;
   wire n_2_18_397;
   wire n_2_18_398;
   wire n_2_18_399;
   wire n_2_18_400;
   wire n_2_18_401;
   wire n_2_18_402;
   wire n_2_18_403;
   wire n_2_18_404;
   wire n_2_18_405;
   wire n_2_18_406;
   wire n_2_18_407;
   wire n_2_18_408;
   wire n_2_18_409;
   wire n_2_18_410;
   wire n_2_18_411;
   wire n_2_18_412;
   wire n_2_18_413;
   wire n_2_18_414;
   wire n_2_18_415;
   wire n_2_200;
   wire n_2_201;
   wire n_2_202;
   wire n_2_203;
   wire n_2_204;
   wire n_2_205;
   wire n_2_206;
   wire n_2_207;
   wire n_2_213;
   wire n_2_18_416;
   wire n_2_18_417;
   wire n_2_18_418;
   wire n_2_18_419;
   wire n_2_18_420;
   wire n_2_18_421;
   wire n_2_18_422;
   wire n_2_18_423;
   wire n_2_214;
   wire n_2_171;
   wire n_2_184;
   wire n_2_170;
   wire n_2_18_424;
   wire n_2_18_425;
   wire n_2_18_426;
   wire n_2_18_427;
   wire n_2_18_428;
   wire n_2_208;
   wire n_2_18_429;
   wire n_2_18_430;
   wire n_2_18_431;
   wire n_2_18_432;
   wire n_2_216;
   wire n_2_18_433;
   wire n_2_18_434;
   wire n_2_215;
   wire n_2_18_435;
   wire n_2_18_436;
   wire n_2_18_437;
   wire n_2_18_438;
   wire n_2_18_439;
   wire n_2_18_440;
   wire n_2_18_441;
   wire n_2_18_442;
   wire n_2_18_443;
   wire n_2_18_444;
   wire n_2_18_445;
   wire n_2_18_446;
   wire n_2_226;
   wire n_2_227;
   wire n_2_228;
   wire n_2_19_0;
   wire n_2_19_1;
   wire n_2_19_2;
   wire n_2_19_3;
   wire n_2_19_4;
   wire n_2_19_5;
   wire n_2_19_6;
   wire n_2_19_7;
   wire n_2_229;
   wire n_2_19_8;
   wire n_3_0;
   wire [15:0]RowsNum;
   wire Start_Bit;
   wire Row_Done_Bit;
   wire n_3_1;
   wire [15:0]Relative_Address;
   wire Update_Address_Indication_Bit;
   wire Data_Bit;
   wire [5:0]Writing_Start_Index;
   wire [11:0]N;
   wire N_Indication_Bit;
   wire Row_Last_Bit;
   wire [5:0]Small_Packet_Indication_Bit_Location;
   wire [5:0]PacketSize;
   wire [31:0]Data_Size;
   wire [31:0]Small_Packet_Data_Size;
   wire n_3_2;
   wire n_3_3;
   wire [15:0]RowsCount;
   wire Done_Element_Delayed;
   wire [1:0]InitCount;
   wire Row_Done_Bit_Delayed;
   wire n_0_0;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_1;
   wire n_0_1_0;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_1_1;

   datapath__0_35 i_257_3 (.p_0({n_37, uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, 
      uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, 
      uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, n_36, n_35, n_34, n_33, 
      n_32, uc_25}), .p_1({uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, uc_32, 
      uc_33, uc_34, uc_35, uc_36, uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, 
      uc_43, uc_44, uc_45, n_257_5, uc_46, uc_47, uc_48, uc_49, n_257_4, n_257_3, 
      n_257_2, n_257_1, n_257_0, uc_50, uc_51}));
   datapath__0_39 i_257_6 (.p_0({n_257_1096, uc_52, uc_53, uc_54, uc_55, uc_56, 
      uc_57, uc_58, uc_59, uc_60, uc_61, uc_62, uc_63, uc_64, uc_65, uc_66, 
      uc_67, uc_68, uc_69, uc_70, uc_71, uc_72, uc_73, uc_74, uc_75, uc_76, 
      n_257_1095, n_257_1094, n_257_1093, n_257_1092, n_257_1091, uc_77}), 
      .p_1({uc_78, uc_79, uc_80, uc_81, uc_82, uc_83, uc_84, uc_85, uc_86, uc_87, 
      uc_88, uc_89, uc_90, uc_91, uc_92, uc_93, uc_94, uc_95, uc_96, uc_97, 
      n_257_11, uc_98, uc_99, uc_100, uc_101, n_257_10, n_257_9, n_257_8, 
      n_257_7, n_257_6, uc_102, uc_103}));
   NAND2_X1 i_257_0_0 (.A1(n_256), .A2(n_257), .ZN(n_257_0_0));
   INV_X1 i_257_0_1 (.A(n_258), .ZN(n_257_0_1));
   NOR2_X1 i_257_0_2 (.A1(n_257_0_0), .A2(n_257_0_1), .ZN(n_257_0_2));
   INV_X1 i_257_0_3 (.A(n_254), .ZN(n_257_0_3));
   NAND2_X1 i_257_0_4 (.A1(n_257_0_2), .A2(n_257_0_3), .ZN(n_257_0_4));
   INV_X1 i_257_0_5 (.A(n_255), .ZN(n_257_0_5));
   NOR2_X1 i_257_0_6 (.A1(n_257_0_4), .A2(n_257_0_5), .ZN(n_257_0_6));
   NAND2_X1 i_257_0_7 (.A1(CPU_Bus[30]), .A2(n_257_0_6), .ZN(n_257_0_7));
   NAND2_X1 i_257_0_8 (.A1(n_257_0_2), .A2(n_254), .ZN(n_257_0_8));
   NOR2_X1 i_257_0_9 (.A1(n_257_0_8), .A2(n_257_0_5), .ZN(n_257_0_9));
   NAND2_X1 i_257_0_10 (.A1(CPU_Bus[31]), .A2(n_257_0_9), .ZN(n_257_0_10));
   NAND2_X1 i_257_0_11 (.A1(n_257_0_7), .A2(n_257_0_10), .ZN(n_257_0_11));
   NOR2_X1 i_257_0_12 (.A1(n_257_0_8), .A2(n_255), .ZN(n_257_0_12));
   NAND2_X1 i_257_0_13 (.A1(CPU_Bus[29]), .A2(n_257_0_12), .ZN(n_257_0_13));
   NOR2_X1 i_257_0_14 (.A1(n_257_0_4), .A2(n_255), .ZN(n_257_0_14));
   NAND2_X1 i_257_0_15 (.A1(CPU_Bus[28]), .A2(n_257_0_14), .ZN(n_257_0_15));
   NAND2_X1 i_257_0_16 (.A1(n_257_0_13), .A2(n_257_0_15), .ZN(n_257_0_16));
   NOR2_X1 i_257_0_17 (.A1(n_257_0_11), .A2(n_257_0_16), .ZN(n_257_0_17));
   INV_X1 i_257_0_18 (.A(n_256), .ZN(n_257_0_18));
   NAND2_X1 i_257_0_19 (.A1(n_257_0_18), .A2(n_257), .ZN(n_257_0_19));
   NOR2_X1 i_257_0_20 (.A1(n_257_0_19), .A2(n_257_0_1), .ZN(n_257_0_20));
   NAND2_X1 i_257_0_21 (.A1(n_257_0_20), .A2(n_254), .ZN(n_257_0_21));
   NOR2_X1 i_257_0_22 (.A1(n_257_0_21), .A2(n_257_0_5), .ZN(n_257_0_22));
   NAND2_X1 i_257_0_23 (.A1(CPU_Bus[27]), .A2(n_257_0_22), .ZN(n_257_0_23));
   NAND2_X1 i_257_0_24 (.A1(n_257_0_20), .A2(n_257_0_3), .ZN(n_257_0_24));
   NOR2_X1 i_257_0_25 (.A1(n_257_0_24), .A2(n_257_0_5), .ZN(n_257_0_25));
   NAND2_X1 i_257_0_26 (.A1(CPU_Bus[26]), .A2(n_257_0_25), .ZN(n_257_0_26));
   NAND2_X1 i_257_0_27 (.A1(n_257_0_23), .A2(n_257_0_26), .ZN(n_257_0_27));
   NOR2_X1 i_257_0_28 (.A1(n_257_0_21), .A2(n_255), .ZN(n_257_0_28));
   NAND2_X1 i_257_0_29 (.A1(CPU_Bus[25]), .A2(n_257_0_28), .ZN(n_257_0_29));
   NOR2_X1 i_257_0_30 (.A1(n_257_0_24), .A2(n_255), .ZN(n_257_0_30));
   NAND2_X1 i_257_0_31 (.A1(CPU_Bus[24]), .A2(n_257_0_30), .ZN(n_257_0_31));
   NAND2_X1 i_257_0_32 (.A1(n_257_0_29), .A2(n_257_0_31), .ZN(n_257_0_32));
   NOR2_X1 i_257_0_33 (.A1(n_257_0_27), .A2(n_257_0_32), .ZN(n_257_0_33));
   NAND2_X1 i_257_0_34 (.A1(n_257_0_17), .A2(n_257_0_33), .ZN(n_257_0_34));
   INV_X1 i_257_0_35 (.A(n_257), .ZN(n_257_0_35));
   NAND2_X1 i_257_0_36 (.A1(n_257_0_35), .A2(n_256), .ZN(n_257_0_36));
   NOR2_X1 i_257_0_37 (.A1(n_257_0_36), .A2(n_257_0_1), .ZN(n_257_0_37));
   NAND2_X1 i_257_0_38 (.A1(n_257_0_37), .A2(n_254), .ZN(n_257_0_38));
   NOR2_X1 i_257_0_39 (.A1(n_257_0_38), .A2(n_257_0_5), .ZN(n_257_0_39));
   NAND2_X1 i_257_0_40 (.A1(CPU_Bus[23]), .A2(n_257_0_39), .ZN(n_257_0_40));
   NAND2_X1 i_257_0_41 (.A1(n_257_0_37), .A2(n_257_0_3), .ZN(n_257_0_41));
   NOR2_X1 i_257_0_42 (.A1(n_257_0_41), .A2(n_257_0_5), .ZN(n_257_0_42));
   NAND2_X1 i_257_0_43 (.A1(CPU_Bus[22]), .A2(n_257_0_42), .ZN(n_257_0_43));
   NAND2_X1 i_257_0_44 (.A1(n_257_0_40), .A2(n_257_0_43), .ZN(n_257_0_44));
   NOR2_X1 i_257_0_45 (.A1(n_257_0_38), .A2(n_255), .ZN(n_257_0_45));
   NAND2_X1 i_257_0_46 (.A1(CPU_Bus[21]), .A2(n_257_0_45), .ZN(n_257_0_46));
   NOR2_X1 i_257_0_47 (.A1(n_257_0_41), .A2(n_255), .ZN(n_257_0_47));
   NAND2_X1 i_257_0_48 (.A1(CPU_Bus[20]), .A2(n_257_0_47), .ZN(n_257_0_48));
   NAND2_X1 i_257_0_49 (.A1(n_257_0_46), .A2(n_257_0_48), .ZN(n_257_0_49));
   NOR2_X1 i_257_0_50 (.A1(n_257_0_44), .A2(n_257_0_49), .ZN(n_257_0_50));
   NAND2_X1 i_257_0_51 (.A1(n_257_0_18), .A2(n_257_0_35), .ZN(n_257_0_51));
   NOR2_X1 i_257_0_52 (.A1(n_257_0_51), .A2(n_257_0_1), .ZN(n_257_0_52));
   NAND2_X1 i_257_0_53 (.A1(n_257_0_52), .A2(n_254), .ZN(n_257_0_53));
   NOR2_X1 i_257_0_54 (.A1(n_257_0_53), .A2(n_257_0_5), .ZN(n_257_0_54));
   NAND2_X1 i_257_0_55 (.A1(CPU_Bus[19]), .A2(n_257_0_54), .ZN(n_257_0_55));
   NAND2_X1 i_257_0_56 (.A1(n_257_0_52), .A2(n_257_0_3), .ZN(n_257_0_56));
   NOR2_X1 i_257_0_57 (.A1(n_257_0_56), .A2(n_257_0_5), .ZN(n_257_0_57));
   NAND2_X1 i_257_0_58 (.A1(CPU_Bus[18]), .A2(n_257_0_57), .ZN(n_257_0_58));
   NAND2_X1 i_257_0_59 (.A1(n_257_0_55), .A2(n_257_0_58), .ZN(n_257_0_59));
   NOR2_X1 i_257_0_60 (.A1(n_257_0_53), .A2(n_255), .ZN(n_257_0_60));
   NAND2_X1 i_257_0_61 (.A1(CPU_Bus[17]), .A2(n_257_0_60), .ZN(n_257_0_61));
   NOR2_X1 i_257_0_62 (.A1(n_257_0_56), .A2(n_255), .ZN(n_257_0_62));
   NAND2_X1 i_257_0_63 (.A1(CPU_Bus[16]), .A2(n_257_0_62), .ZN(n_257_0_63));
   NAND2_X1 i_257_0_64 (.A1(n_257_0_61), .A2(n_257_0_63), .ZN(n_257_0_64));
   NOR2_X1 i_257_0_65 (.A1(n_257_0_59), .A2(n_257_0_64), .ZN(n_257_0_65));
   NAND2_X1 i_257_0_66 (.A1(n_257_0_50), .A2(n_257_0_65), .ZN(n_257_0_66));
   NOR2_X1 i_257_0_67 (.A1(n_257_0_34), .A2(n_257_0_66), .ZN(n_257_0_67));
   NOR2_X1 i_257_0_68 (.A1(n_257_0_0), .A2(n_258), .ZN(n_257_0_68));
   NAND2_X1 i_257_0_69 (.A1(n_257_0_68), .A2(n_254), .ZN(n_257_0_69));
   NOR2_X1 i_257_0_70 (.A1(n_257_0_69), .A2(n_257_0_5), .ZN(n_257_0_70));
   NAND2_X1 i_257_0_71 (.A1(CPU_Bus[15]), .A2(n_257_0_70), .ZN(n_257_0_71));
   NAND2_X1 i_257_0_72 (.A1(n_257_0_68), .A2(n_257_0_3), .ZN(n_257_0_72));
   NOR2_X1 i_257_0_73 (.A1(n_257_0_72), .A2(n_257_0_5), .ZN(n_257_0_73));
   NAND2_X1 i_257_0_74 (.A1(CPU_Bus[14]), .A2(n_257_0_73), .ZN(n_257_0_74));
   NAND2_X1 i_257_0_75 (.A1(n_257_0_71), .A2(n_257_0_74), .ZN(n_257_0_75));
   NOR2_X1 i_257_0_76 (.A1(n_257_0_69), .A2(n_255), .ZN(n_257_0_76));
   NAND2_X1 i_257_0_77 (.A1(CPU_Bus[13]), .A2(n_257_0_76), .ZN(n_257_0_77));
   NOR2_X1 i_257_0_78 (.A1(n_257_0_72), .A2(n_255), .ZN(n_257_0_78));
   NAND2_X1 i_257_0_79 (.A1(CPU_Bus[12]), .A2(n_257_0_78), .ZN(n_257_0_79));
   NAND2_X1 i_257_0_80 (.A1(n_257_0_77), .A2(n_257_0_79), .ZN(n_257_0_80));
   NOR2_X1 i_257_0_81 (.A1(n_257_0_75), .A2(n_257_0_80), .ZN(n_257_0_81));
   NOR2_X1 i_257_0_82 (.A1(n_257_0_19), .A2(n_258), .ZN(n_257_0_82));
   NAND2_X1 i_257_0_83 (.A1(n_257_0_82), .A2(n_254), .ZN(n_257_0_83));
   NOR2_X1 i_257_0_84 (.A1(n_257_0_83), .A2(n_257_0_5), .ZN(n_257_0_84));
   NAND2_X1 i_257_0_85 (.A1(CPU_Bus[11]), .A2(n_257_0_84), .ZN(n_257_0_85));
   NAND2_X1 i_257_0_86 (.A1(n_257_0_82), .A2(n_257_0_3), .ZN(n_257_0_86));
   NOR2_X1 i_257_0_87 (.A1(n_257_0_86), .A2(n_257_0_5), .ZN(n_257_0_87));
   NAND2_X1 i_257_0_88 (.A1(CPU_Bus[10]), .A2(n_257_0_87), .ZN(n_257_0_88));
   NAND2_X1 i_257_0_89 (.A1(n_257_0_85), .A2(n_257_0_88), .ZN(n_257_0_89));
   NOR2_X1 i_257_0_90 (.A1(n_257_0_83), .A2(n_255), .ZN(n_257_0_90));
   NAND2_X1 i_257_0_91 (.A1(CPU_Bus[9]), .A2(n_257_0_90), .ZN(n_257_0_91));
   NOR2_X1 i_257_0_92 (.A1(n_257_0_86), .A2(n_255), .ZN(n_257_0_92));
   NAND2_X1 i_257_0_93 (.A1(CPU_Bus[8]), .A2(n_257_0_92), .ZN(n_257_0_93));
   NAND2_X1 i_257_0_94 (.A1(n_257_0_91), .A2(n_257_0_93), .ZN(n_257_0_94));
   NOR2_X1 i_257_0_95 (.A1(n_257_0_89), .A2(n_257_0_94), .ZN(n_257_0_95));
   NAND2_X1 i_257_0_96 (.A1(n_257_0_81), .A2(n_257_0_95), .ZN(n_257_0_96));
   NOR2_X1 i_257_0_97 (.A1(n_257_0_36), .A2(n_258), .ZN(n_257_0_97));
   NAND2_X1 i_257_0_98 (.A1(n_257_0_97), .A2(n_254), .ZN(n_257_0_98));
   NOR2_X1 i_257_0_99 (.A1(n_257_0_98), .A2(n_257_0_5), .ZN(n_257_0_99));
   NAND2_X1 i_257_0_100 (.A1(CPU_Bus[7]), .A2(n_257_0_99), .ZN(n_257_0_100));
   NAND2_X1 i_257_0_101 (.A1(n_257_0_97), .A2(n_257_0_3), .ZN(n_257_0_101));
   NOR2_X1 i_257_0_102 (.A1(n_257_0_101), .A2(n_257_0_5), .ZN(n_257_0_102));
   NAND2_X1 i_257_0_103 (.A1(CPU_Bus[6]), .A2(n_257_0_102), .ZN(n_257_0_103));
   NAND2_X1 i_257_0_104 (.A1(n_257_0_100), .A2(n_257_0_103), .ZN(n_257_0_104));
   NOR2_X1 i_257_0_105 (.A1(n_257_0_98), .A2(n_255), .ZN(n_257_0_105));
   NAND2_X1 i_257_0_106 (.A1(CPU_Bus[5]), .A2(n_257_0_105), .ZN(n_257_0_106));
   NOR2_X1 i_257_0_107 (.A1(n_257_0_101), .A2(n_255), .ZN(n_257_0_107));
   NAND2_X1 i_257_0_108 (.A1(CPU_Bus[4]), .A2(n_257_0_107), .ZN(n_257_0_108));
   NAND2_X1 i_257_0_109 (.A1(n_257_0_106), .A2(n_257_0_108), .ZN(n_257_0_109));
   NOR2_X1 i_257_0_110 (.A1(n_257_0_104), .A2(n_257_0_109), .ZN(n_257_0_110));
   NOR2_X1 i_257_0_111 (.A1(n_257_0_51), .A2(n_258), .ZN(n_257_0_111));
   NAND2_X1 i_257_0_112 (.A1(n_257_0_111), .A2(n_254), .ZN(n_257_0_112));
   NOR2_X1 i_257_0_113 (.A1(n_257_0_112), .A2(n_257_0_5), .ZN(n_257_0_113));
   NAND2_X1 i_257_0_114 (.A1(CPU_Bus[3]), .A2(n_257_0_113), .ZN(n_257_0_114));
   NAND2_X1 i_257_0_115 (.A1(n_257_0_111), .A2(n_257_0_3), .ZN(n_257_0_115));
   NOR2_X1 i_257_0_116 (.A1(n_257_0_115), .A2(n_257_0_5), .ZN(n_257_0_116));
   NAND2_X1 i_257_0_117 (.A1(CPU_Bus[2]), .A2(n_257_0_116), .ZN(n_257_0_117));
   NAND2_X1 i_257_0_118 (.A1(n_257_0_114), .A2(n_257_0_117), .ZN(n_257_0_118));
   NOR2_X1 i_257_0_119 (.A1(n_257_0_112), .A2(n_255), .ZN(n_257_0_119));
   NAND2_X1 i_257_0_120 (.A1(CPU_Bus[1]), .A2(n_257_0_119), .ZN(n_257_0_120));
   NOR2_X1 i_257_0_121 (.A1(n_257_0_115), .A2(n_255), .ZN(n_257_0_121));
   NAND2_X1 i_257_0_122 (.A1(CPU_Bus[0]), .A2(n_257_0_121), .ZN(n_257_0_122));
   NAND2_X1 i_257_0_123 (.A1(n_257_0_120), .A2(n_257_0_122), .ZN(n_257_0_123));
   NOR2_X1 i_257_0_124 (.A1(n_257_0_118), .A2(n_257_0_123), .ZN(n_257_0_124));
   NAND2_X1 i_257_0_125 (.A1(n_257_0_110), .A2(n_257_0_124), .ZN(n_257_0_125));
   NOR2_X1 i_257_0_126 (.A1(n_257_0_96), .A2(n_257_0_125), .ZN(n_257_0_126));
   NAND2_X1 i_257_0_127 (.A1(n_257_0_67), .A2(n_257_0_126), .ZN(n_257_12));
   INV_X1 i_257_1_0 (.A(n_257_1_0), .ZN(n_257_13));
   NAND2_X1 i_257_1_1 (.A1(n_257_1_49), .A2(n_257_1_1), .ZN(n_257_1_0));
   NAND3_X1 i_257_1_2 (.A1(n_257_1_25), .A2(n_257_1_2), .A3(n_257_1_48), 
      .ZN(n_257_1_1));
   NAND3_X1 i_257_1_3 (.A1(n_257_1_14), .A2(n_257_1_3), .A3(n_257), .ZN(
      n_257_1_2));
   NAND3_X1 i_257_1_4 (.A1(n_257_1_9), .A2(n_257_1_4), .A3(n_257_1_85), .ZN(
      n_257_1_3));
   NAND3_X1 i_257_1_5 (.A1(n_257_1_7), .A2(n_257_1_5), .A3(n_257_1_96), .ZN(
      n_257_1_4));
   NAND2_X1 i_257_1_6 (.A1(n_257_1_6), .A2(n_257_1_95), .ZN(n_257_1_5));
   INV_X1 i_257_1_7 (.A(CPU_Bus[7]), .ZN(n_257_1_6));
   NAND2_X1 i_257_1_8 (.A1(n_257_1_8), .A2(n_254), .ZN(n_257_1_7));
   INV_X1 i_257_1_9 (.A(CPU_Bus[8]), .ZN(n_257_1_8));
   NAND3_X1 i_257_1_10 (.A1(n_257_1_12), .A2(n_257_1_10), .A3(n_255), .ZN(
      n_257_1_9));
   NAND2_X1 i_257_1_11 (.A1(n_257_1_11), .A2(n_257_1_95), .ZN(n_257_1_10));
   INV_X1 i_257_1_12 (.A(CPU_Bus[9]), .ZN(n_257_1_11));
   NAND2_X1 i_257_1_13 (.A1(n_257_1_13), .A2(n_254), .ZN(n_257_1_12));
   INV_X1 i_257_1_14 (.A(CPU_Bus[10]), .ZN(n_257_1_13));
   NAND3_X1 i_257_1_15 (.A1(n_257_1_20), .A2(n_257_1_15), .A3(n_256), .ZN(
      n_257_1_14));
   NAND3_X1 i_257_1_16 (.A1(n_257_1_18), .A2(n_257_1_16), .A3(n_257_1_96), 
      .ZN(n_257_1_15));
   NAND2_X1 i_257_1_17 (.A1(n_257_1_17), .A2(n_257_1_95), .ZN(n_257_1_16));
   INV_X1 i_257_1_18 (.A(CPU_Bus[11]), .ZN(n_257_1_17));
   NAND2_X1 i_257_1_19 (.A1(n_257_1_19), .A2(n_254), .ZN(n_257_1_18));
   INV_X1 i_257_1_20 (.A(CPU_Bus[12]), .ZN(n_257_1_19));
   NAND3_X1 i_257_1_21 (.A1(n_257_1_23), .A2(n_257_1_21), .A3(n_255), .ZN(
      n_257_1_20));
   NAND2_X1 i_257_1_22 (.A1(n_257_1_22), .A2(n_257_1_95), .ZN(n_257_1_21));
   INV_X1 i_257_1_23 (.A(CPU_Bus[13]), .ZN(n_257_1_22));
   NAND2_X1 i_257_1_24 (.A1(n_257_1_24), .A2(n_254), .ZN(n_257_1_23));
   INV_X1 i_257_1_25 (.A(CPU_Bus[14]), .ZN(n_257_1_24));
   NAND3_X1 i_257_1_26 (.A1(n_257_1_37), .A2(n_257_1_26), .A3(n_257_1_97), 
      .ZN(n_257_1_25));
   NAND3_X1 i_257_1_27 (.A1(n_257_1_32), .A2(n_257_1_27), .A3(n_256), .ZN(
      n_257_1_26));
   NAND3_X1 i_257_1_28 (.A1(n_257_1_30), .A2(n_257_1_28), .A3(n_255), .ZN(
      n_257_1_27));
   NAND2_X1 i_257_1_29 (.A1(n_257_1_29), .A2(n_254), .ZN(n_257_1_28));
   INV_X1 i_257_1_30 (.A(CPU_Bus[6]), .ZN(n_257_1_29));
   NAND2_X1 i_257_1_31 (.A1(n_257_1_31), .A2(n_257_1_95), .ZN(n_257_1_30));
   INV_X1 i_257_1_32 (.A(CPU_Bus[5]), .ZN(n_257_1_31));
   NAND3_X1 i_257_1_33 (.A1(n_257_1_35), .A2(n_257_1_33), .A3(n_257_1_96), 
      .ZN(n_257_1_32));
   NAND2_X1 i_257_1_34 (.A1(n_257_1_34), .A2(n_257_1_95), .ZN(n_257_1_33));
   INV_X1 i_257_1_35 (.A(CPU_Bus[3]), .ZN(n_257_1_34));
   NAND2_X1 i_257_1_36 (.A1(n_257_1_36), .A2(n_254), .ZN(n_257_1_35));
   INV_X1 i_257_1_37 (.A(CPU_Bus[4]), .ZN(n_257_1_36));
   NAND3_X1 i_257_1_38 (.A1(n_257_1_43), .A2(n_257_1_38), .A3(n_257_1_85), 
      .ZN(n_257_1_37));
   NAND3_X1 i_257_1_39 (.A1(n_257_1_41), .A2(n_257_1_39), .A3(n_255), .ZN(
      n_257_1_38));
   NAND2_X1 i_257_1_40 (.A1(n_257_1_40), .A2(n_254), .ZN(n_257_1_39));
   INV_X1 i_257_1_41 (.A(CPU_Bus[2]), .ZN(n_257_1_40));
   NAND2_X1 i_257_1_42 (.A1(n_257_1_42), .A2(n_257_1_95), .ZN(n_257_1_41));
   INV_X1 i_257_1_43 (.A(CPU_Bus[1]), .ZN(n_257_1_42));
   NAND3_X1 i_257_1_44 (.A1(n_257_1_46), .A2(n_257_1_44), .A3(n_257_1_96), 
      .ZN(n_257_1_43));
   NAND2_X1 i_257_1_45 (.A1(n_257_1_45), .A2(n_257_1_95), .ZN(n_257_1_44));
   INV_X1 i_257_1_46 (.A(CPU_Bus[31]), .ZN(n_257_1_45));
   NAND2_X1 i_257_1_47 (.A1(n_257_1_47), .A2(n_254), .ZN(n_257_1_46));
   INV_X1 i_257_1_48 (.A(CPU_Bus[0]), .ZN(n_257_1_47));
   INV_X1 i_257_1_49 (.A(n_258), .ZN(n_257_1_48));
   NAND3_X1 i_257_1_50 (.A1(n_257_1_73), .A2(n_257_1_50), .A3(n_258), .ZN(
      n_257_1_49));
   NAND3_X1 i_257_1_51 (.A1(n_257_1_62), .A2(n_257_1_51), .A3(n_257), .ZN(
      n_257_1_50));
   NAND3_X1 i_257_1_52 (.A1(n_257_1_57), .A2(n_257_1_52), .A3(n_257_1_85), 
      .ZN(n_257_1_51));
   NAND3_X1 i_257_1_53 (.A1(n_257_1_55), .A2(n_257_1_53), .A3(n_257_1_96), 
      .ZN(n_257_1_52));
   NAND2_X1 i_257_1_54 (.A1(n_257_1_54), .A2(n_257_1_95), .ZN(n_257_1_53));
   INV_X1 i_257_1_55 (.A(CPU_Bus[23]), .ZN(n_257_1_54));
   NAND2_X1 i_257_1_56 (.A1(n_257_1_56), .A2(n_254), .ZN(n_257_1_55));
   INV_X1 i_257_1_57 (.A(CPU_Bus[24]), .ZN(n_257_1_56));
   NAND3_X1 i_257_1_58 (.A1(n_257_1_60), .A2(n_257_1_58), .A3(n_255), .ZN(
      n_257_1_57));
   NAND2_X1 i_257_1_59 (.A1(n_257_1_59), .A2(n_254), .ZN(n_257_1_58));
   INV_X1 i_257_1_60 (.A(CPU_Bus[26]), .ZN(n_257_1_59));
   NAND2_X1 i_257_1_61 (.A1(n_257_1_61), .A2(n_257_1_95), .ZN(n_257_1_60));
   INV_X1 i_257_1_62 (.A(CPU_Bus[25]), .ZN(n_257_1_61));
   NAND3_X1 i_257_1_63 (.A1(n_257_1_68), .A2(n_257_1_63), .A3(n_256), .ZN(
      n_257_1_62));
   NAND3_X1 i_257_1_64 (.A1(n_257_1_66), .A2(n_257_1_64), .A3(n_257_1_96), 
      .ZN(n_257_1_63));
   NAND2_X1 i_257_1_65 (.A1(n_257_1_65), .A2(n_254), .ZN(n_257_1_64));
   INV_X1 i_257_1_66 (.A(CPU_Bus[28]), .ZN(n_257_1_65));
   NAND2_X1 i_257_1_67 (.A1(n_257_1_67), .A2(n_257_1_95), .ZN(n_257_1_66));
   INV_X1 i_257_1_68 (.A(CPU_Bus[27]), .ZN(n_257_1_67));
   NAND3_X1 i_257_1_69 (.A1(n_257_1_71), .A2(n_257_1_69), .A3(n_255), .ZN(
      n_257_1_68));
   NAND2_X1 i_257_1_70 (.A1(n_257_1_70), .A2(n_257_1_95), .ZN(n_257_1_69));
   INV_X1 i_257_1_71 (.A(CPU_Bus[29]), .ZN(n_257_1_70));
   NAND2_X1 i_257_1_72 (.A1(n_257_1_72), .A2(n_254), .ZN(n_257_1_71));
   INV_X1 i_257_1_73 (.A(CPU_Bus[30]), .ZN(n_257_1_72));
   NAND3_X1 i_257_1_74 (.A1(n_257_1_86), .A2(n_257_1_74), .A3(n_257_1_97), 
      .ZN(n_257_1_73));
   NAND3_X1 i_257_1_75 (.A1(n_257_1_80), .A2(n_257_1_75), .A3(n_257_1_85), 
      .ZN(n_257_1_74));
   NAND3_X1 i_257_1_76 (.A1(n_257_1_78), .A2(n_257_1_76), .A3(n_257_1_96), 
      .ZN(n_257_1_75));
   NAND2_X1 i_257_1_77 (.A1(n_257_1_77), .A2(n_254), .ZN(n_257_1_76));
   INV_X1 i_257_1_78 (.A(CPU_Bus[16]), .ZN(n_257_1_77));
   NAND2_X1 i_257_1_79 (.A1(n_257_1_79), .A2(n_257_1_95), .ZN(n_257_1_78));
   INV_X1 i_257_1_80 (.A(CPU_Bus[15]), .ZN(n_257_1_79));
   NAND3_X1 i_257_1_81 (.A1(n_257_1_83), .A2(n_257_1_81), .A3(n_255), .ZN(
      n_257_1_80));
   NAND2_X1 i_257_1_82 (.A1(n_257_1_82), .A2(n_254), .ZN(n_257_1_81));
   INV_X1 i_257_1_83 (.A(CPU_Bus[18]), .ZN(n_257_1_82));
   NAND2_X1 i_257_1_84 (.A1(n_257_1_84), .A2(n_257_1_95), .ZN(n_257_1_83));
   INV_X1 i_257_1_85 (.A(CPU_Bus[17]), .ZN(n_257_1_84));
   INV_X1 i_257_1_86 (.A(n_256), .ZN(n_257_1_85));
   NAND3_X1 i_257_1_87 (.A1(n_257_1_92), .A2(n_257_1_87), .A3(n_256), .ZN(
      n_257_1_86));
   NAND3_X1 i_257_1_88 (.A1(n_257_1_90), .A2(n_257_1_88), .A3(n_255), .ZN(
      n_257_1_87));
   NAND2_X1 i_257_1_89 (.A1(n_257_1_89), .A2(n_257_1_95), .ZN(n_257_1_88));
   INV_X1 i_257_1_90 (.A(CPU_Bus[21]), .ZN(n_257_1_89));
   NAND2_X1 i_257_1_91 (.A1(n_257_1_91), .A2(n_254), .ZN(n_257_1_90));
   INV_X1 i_257_1_92 (.A(CPU_Bus[22]), .ZN(n_257_1_91));
   OAI211_X1 i_257_1_93 (.A(n_257_1_93), .B(n_257_1_96), .C1(n_257_1_95), 
      .C2(CPU_Bus[20]), .ZN(n_257_1_92));
   NAND2_X1 i_257_1_94 (.A1(n_257_1_94), .A2(n_257_1_95), .ZN(n_257_1_93));
   INV_X1 i_257_1_95 (.A(CPU_Bus[19]), .ZN(n_257_1_94));
   INV_X1 i_257_1_96 (.A(n_254), .ZN(n_257_1_95));
   INV_X1 i_257_1_97 (.A(n_255), .ZN(n_257_1_96));
   INV_X1 i_257_1_98 (.A(n_257), .ZN(n_257_1_97));
   INV_X1 i_257_2_0 (.A(n_254), .ZN(n_257_2_0));
   NAND2_X1 i_257_2_1 (.A1(n_257_2_0), .A2(n_255), .ZN(n_257_2_1));
   INV_X1 i_257_2_2 (.A(n_256), .ZN(n_257_2_2));
   NOR2_X1 i_257_2_3 (.A1(n_257_2_1), .A2(n_257_2_2), .ZN(n_257_2_3));
   NAND2_X1 i_257_2_4 (.A1(n_257_2_3), .A2(n_257), .ZN(n_257_2_4));
   INV_X1 i_257_2_5 (.A(n_258), .ZN(n_257_2_5));
   NOR2_X1 i_257_2_6 (.A1(n_257_2_4), .A2(n_257_2_5), .ZN(n_257_2_6));
   NAND2_X1 i_257_2_7 (.A1(CPU_Bus[28]), .A2(n_257_2_6), .ZN(n_257_2_7));
   INV_X1 i_257_2_8 (.A(n_255), .ZN(n_257_2_8));
   NAND2_X1 i_257_2_9 (.A1(n_257_2_0), .A2(n_257_2_8), .ZN(n_257_2_9));
   NOR2_X1 i_257_2_10 (.A1(n_257_2_9), .A2(n_257_2_2), .ZN(n_257_2_10));
   NAND2_X1 i_257_2_11 (.A1(n_257_2_10), .A2(n_257), .ZN(n_257_2_11));
   NOR2_X1 i_257_2_12 (.A1(n_257_2_11), .A2(n_257_2_5), .ZN(n_257_2_12));
   NAND2_X1 i_257_2_13 (.A1(CPU_Bus[26]), .A2(n_257_2_12), .ZN(n_257_2_13));
   NAND2_X1 i_257_2_14 (.A1(n_257_2_7), .A2(n_257_2_13), .ZN(n_257_2_14));
   NOR2_X1 i_257_2_15 (.A1(n_257_2_1), .A2(n_256), .ZN(n_257_2_15));
   NAND2_X1 i_257_2_16 (.A1(n_257_2_15), .A2(n_257), .ZN(n_257_2_16));
   NOR2_X1 i_257_2_17 (.A1(n_257_2_16), .A2(n_257_2_5), .ZN(n_257_2_17));
   NAND2_X1 i_257_2_18 (.A1(CPU_Bus[24]), .A2(n_257_2_17), .ZN(n_257_2_18));
   NOR2_X1 i_257_2_19 (.A1(n_257_2_9), .A2(n_256), .ZN(n_257_2_19));
   NAND2_X1 i_257_2_20 (.A1(n_257_2_19), .A2(n_257), .ZN(n_257_2_20));
   NOR2_X1 i_257_2_21 (.A1(n_257_2_20), .A2(n_257_2_5), .ZN(n_257_2_21));
   NAND2_X1 i_257_2_22 (.A1(CPU_Bus[22]), .A2(n_257_2_21), .ZN(n_257_2_22));
   NAND2_X1 i_257_2_23 (.A1(n_257_2_18), .A2(n_257_2_22), .ZN(n_257_2_23));
   NOR2_X1 i_257_2_24 (.A1(n_257_2_14), .A2(n_257_2_23), .ZN(n_257_2_24));
   INV_X1 i_257_2_25 (.A(n_257), .ZN(n_257_2_25));
   NAND2_X1 i_257_2_26 (.A1(n_257_2_3), .A2(n_257_2_25), .ZN(n_257_2_26));
   NOR2_X1 i_257_2_27 (.A1(n_257_2_26), .A2(n_257_2_5), .ZN(n_257_2_27));
   NAND2_X1 i_257_2_28 (.A1(CPU_Bus[20]), .A2(n_257_2_27), .ZN(n_257_2_28));
   NAND2_X1 i_257_2_29 (.A1(n_257_2_10), .A2(n_257_2_25), .ZN(n_257_2_29));
   NOR2_X1 i_257_2_30 (.A1(n_257_2_29), .A2(n_257_2_5), .ZN(n_257_2_30));
   NAND2_X1 i_257_2_31 (.A1(CPU_Bus[18]), .A2(n_257_2_30), .ZN(n_257_2_31));
   NAND2_X1 i_257_2_32 (.A1(n_257_2_28), .A2(n_257_2_31), .ZN(n_257_2_32));
   NAND2_X1 i_257_2_33 (.A1(n_257_2_15), .A2(n_257_2_25), .ZN(n_257_2_33));
   NOR2_X1 i_257_2_34 (.A1(n_257_2_33), .A2(n_257_2_5), .ZN(n_257_2_34));
   NAND2_X1 i_257_2_35 (.A1(CPU_Bus[16]), .A2(n_257_2_34), .ZN(n_257_2_35));
   NAND2_X1 i_257_2_36 (.A1(n_257_2_19), .A2(n_257_2_25), .ZN(n_257_2_36));
   NOR2_X1 i_257_2_37 (.A1(n_257_2_36), .A2(n_257_2_5), .ZN(n_257_2_37));
   NAND2_X1 i_257_2_38 (.A1(CPU_Bus[14]), .A2(n_257_2_37), .ZN(n_257_2_38));
   NAND2_X1 i_257_2_39 (.A1(n_257_2_35), .A2(n_257_2_38), .ZN(n_257_2_39));
   NOR2_X1 i_257_2_40 (.A1(n_257_2_32), .A2(n_257_2_39), .ZN(n_257_2_40));
   NAND2_X1 i_257_2_41 (.A1(n_257_2_24), .A2(n_257_2_40), .ZN(n_257_2_41));
   NOR2_X1 i_257_2_42 (.A1(n_257_2_4), .A2(n_258), .ZN(n_257_2_42));
   NAND2_X1 i_257_2_43 (.A1(CPU_Bus[12]), .A2(n_257_2_42), .ZN(n_257_2_43));
   NOR2_X1 i_257_2_44 (.A1(n_257_2_11), .A2(n_258), .ZN(n_257_2_44));
   NAND2_X1 i_257_2_45 (.A1(CPU_Bus[10]), .A2(n_257_2_44), .ZN(n_257_2_45));
   NAND2_X1 i_257_2_46 (.A1(n_257_2_43), .A2(n_257_2_45), .ZN(n_257_2_46));
   NOR2_X1 i_257_2_47 (.A1(n_257_2_16), .A2(n_258), .ZN(n_257_2_47));
   NAND2_X1 i_257_2_48 (.A1(CPU_Bus[8]), .A2(n_257_2_47), .ZN(n_257_2_48));
   NOR2_X1 i_257_2_49 (.A1(n_257_2_20), .A2(n_258), .ZN(n_257_2_49));
   NAND2_X1 i_257_2_50 (.A1(CPU_Bus[6]), .A2(n_257_2_49), .ZN(n_257_2_50));
   NAND2_X1 i_257_2_51 (.A1(n_257_2_48), .A2(n_257_2_50), .ZN(n_257_2_51));
   NOR2_X1 i_257_2_52 (.A1(n_257_2_46), .A2(n_257_2_51), .ZN(n_257_2_52));
   NOR2_X1 i_257_2_53 (.A1(n_257_2_26), .A2(n_258), .ZN(n_257_2_53));
   NAND2_X1 i_257_2_54 (.A1(CPU_Bus[4]), .A2(n_257_2_53), .ZN(n_257_2_54));
   NOR2_X1 i_257_2_55 (.A1(n_257_2_29), .A2(n_258), .ZN(n_257_2_55));
   NAND2_X1 i_257_2_56 (.A1(CPU_Bus[2]), .A2(n_257_2_55), .ZN(n_257_2_56));
   NAND2_X1 i_257_2_57 (.A1(n_257_2_54), .A2(n_257_2_56), .ZN(n_257_2_57));
   NOR2_X1 i_257_2_58 (.A1(n_257_2_33), .A2(n_258), .ZN(n_257_2_58));
   NAND2_X1 i_257_2_59 (.A1(CPU_Bus[0]), .A2(n_257_2_58), .ZN(n_257_2_59));
   NOR2_X1 i_257_2_60 (.A1(n_257_2_36), .A2(n_258), .ZN(n_257_2_60));
   NAND2_X1 i_257_2_61 (.A1(CPU_Bus[30]), .A2(n_257_2_60), .ZN(n_257_2_61));
   NAND2_X1 i_257_2_62 (.A1(n_257_2_59), .A2(n_257_2_61), .ZN(n_257_2_62));
   NOR2_X1 i_257_2_63 (.A1(n_257_2_57), .A2(n_257_2_62), .ZN(n_257_2_63));
   NAND2_X1 i_257_2_64 (.A1(n_257_2_52), .A2(n_257_2_63), .ZN(n_257_2_64));
   NOR2_X1 i_257_2_65 (.A1(n_257_2_41), .A2(n_257_2_64), .ZN(n_257_2_65));
   NAND2_X1 i_257_2_66 (.A1(n_257_2_8), .A2(n_254), .ZN(n_257_2_66));
   NOR2_X1 i_257_2_67 (.A1(n_257_2_66), .A2(n_257_2_2), .ZN(n_257_2_67));
   NAND2_X1 i_257_2_68 (.A1(n_257_2_67), .A2(n_257), .ZN(n_257_2_68));
   NOR2_X1 i_257_2_69 (.A1(n_257_2_68), .A2(n_257_2_5), .ZN(n_257_2_69));
   NAND2_X1 i_257_2_70 (.A1(CPU_Bus[27]), .A2(n_257_2_69), .ZN(n_257_2_70));
   NOR2_X1 i_257_2_71 (.A1(n_257_2_66), .A2(n_256), .ZN(n_257_2_71));
   NAND2_X1 i_257_2_72 (.A1(n_257_2_71), .A2(n_257), .ZN(n_257_2_72));
   NOR2_X1 i_257_2_73 (.A1(n_257_2_72), .A2(n_257_2_5), .ZN(n_257_2_73));
   NAND2_X1 i_257_2_74 (.A1(CPU_Bus[23]), .A2(n_257_2_73), .ZN(n_257_2_74));
   NAND2_X1 i_257_2_75 (.A1(n_257_2_70), .A2(n_257_2_74), .ZN(n_257_2_75));
   NAND2_X1 i_257_2_76 (.A1(n_257_2_67), .A2(n_257_2_25), .ZN(n_257_2_76));
   NOR2_X1 i_257_2_77 (.A1(n_257_2_76), .A2(n_257_2_5), .ZN(n_257_2_77));
   NAND2_X1 i_257_2_78 (.A1(CPU_Bus[19]), .A2(n_257_2_77), .ZN(n_257_2_78));
   NAND2_X1 i_257_2_79 (.A1(n_257_2_71), .A2(n_257_2_25), .ZN(n_257_2_79));
   NOR2_X1 i_257_2_80 (.A1(n_257_2_79), .A2(n_257_2_5), .ZN(n_257_2_80));
   NAND2_X1 i_257_2_81 (.A1(CPU_Bus[15]), .A2(n_257_2_80), .ZN(n_257_2_81));
   NAND2_X1 i_257_2_82 (.A1(n_257_2_78), .A2(n_257_2_81), .ZN(n_257_2_82));
   NOR2_X1 i_257_2_83 (.A1(n_257_2_75), .A2(n_257_2_82), .ZN(n_257_2_83));
   NOR2_X1 i_257_2_84 (.A1(n_257_2_68), .A2(n_258), .ZN(n_257_2_84));
   NAND2_X1 i_257_2_85 (.A1(CPU_Bus[11]), .A2(n_257_2_84), .ZN(n_257_2_85));
   NOR2_X1 i_257_2_86 (.A1(n_257_2_72), .A2(n_258), .ZN(n_257_2_86));
   NAND2_X1 i_257_2_87 (.A1(CPU_Bus[7]), .A2(n_257_2_86), .ZN(n_257_2_87));
   NAND2_X1 i_257_2_88 (.A1(n_257_2_85), .A2(n_257_2_87), .ZN(n_257_2_88));
   NOR2_X1 i_257_2_89 (.A1(n_257_2_76), .A2(n_258), .ZN(n_257_2_89));
   NAND2_X1 i_257_2_90 (.A1(CPU_Bus[3]), .A2(n_257_2_89), .ZN(n_257_2_90));
   NOR2_X1 i_257_2_91 (.A1(n_257_2_79), .A2(n_258), .ZN(n_257_2_91));
   NAND2_X1 i_257_2_92 (.A1(CPU_Bus[31]), .A2(n_257_2_91), .ZN(n_257_2_92));
   NAND2_X1 i_257_2_93 (.A1(n_257_2_90), .A2(n_257_2_92), .ZN(n_257_2_93));
   NOR2_X1 i_257_2_94 (.A1(n_257_2_88), .A2(n_257_2_93), .ZN(n_257_2_94));
   NAND2_X1 i_257_2_95 (.A1(n_257_2_83), .A2(n_257_2_94), .ZN(n_257_2_95));
   NAND2_X1 i_257_2_96 (.A1(n_254), .A2(n_255), .ZN(n_257_2_96));
   NOR2_X1 i_257_2_97 (.A1(n_257_2_96), .A2(n_257_2_2), .ZN(n_257_2_97));
   NAND2_X1 i_257_2_98 (.A1(n_257_2_97), .A2(n_257), .ZN(n_257_2_98));
   NOR2_X1 i_257_2_99 (.A1(n_257_2_98), .A2(n_257_2_5), .ZN(n_257_2_99));
   NAND2_X1 i_257_2_100 (.A1(CPU_Bus[29]), .A2(n_257_2_99), .ZN(n_257_2_100));
   NOR2_X1 i_257_2_101 (.A1(n_257_2_96), .A2(n_256), .ZN(n_257_2_101));
   NAND2_X1 i_257_2_102 (.A1(n_257_2_101), .A2(n_257), .ZN(n_257_2_102));
   NOR2_X1 i_257_2_103 (.A1(n_257_2_102), .A2(n_257_2_5), .ZN(n_257_2_103));
   NAND2_X1 i_257_2_104 (.A1(CPU_Bus[25]), .A2(n_257_2_103), .ZN(n_257_2_104));
   NAND2_X1 i_257_2_105 (.A1(n_257_2_100), .A2(n_257_2_104), .ZN(n_257_2_105));
   NAND2_X1 i_257_2_106 (.A1(n_257_2_97), .A2(n_257_2_25), .ZN(n_257_2_106));
   NOR2_X1 i_257_2_107 (.A1(n_257_2_106), .A2(n_257_2_5), .ZN(n_257_2_107));
   NAND2_X1 i_257_2_108 (.A1(CPU_Bus[21]), .A2(n_257_2_107), .ZN(n_257_2_108));
   NAND2_X1 i_257_2_109 (.A1(n_257_2_101), .A2(n_257_2_25), .ZN(n_257_2_109));
   NOR2_X1 i_257_2_110 (.A1(n_257_2_109), .A2(n_257_2_5), .ZN(n_257_2_110));
   NAND2_X1 i_257_2_111 (.A1(CPU_Bus[17]), .A2(n_257_2_110), .ZN(n_257_2_111));
   NAND2_X1 i_257_2_112 (.A1(n_257_2_108), .A2(n_257_2_111), .ZN(n_257_2_112));
   NOR2_X1 i_257_2_113 (.A1(n_257_2_105), .A2(n_257_2_112), .ZN(n_257_2_113));
   NOR2_X1 i_257_2_114 (.A1(n_257_2_98), .A2(n_258), .ZN(n_257_2_114));
   NAND2_X1 i_257_2_115 (.A1(CPU_Bus[13]), .A2(n_257_2_114), .ZN(n_257_2_115));
   NOR2_X1 i_257_2_116 (.A1(n_257_2_102), .A2(n_258), .ZN(n_257_2_116));
   NAND2_X1 i_257_2_117 (.A1(CPU_Bus[9]), .A2(n_257_2_116), .ZN(n_257_2_117));
   NAND2_X1 i_257_2_118 (.A1(n_257_2_115), .A2(n_257_2_117), .ZN(n_257_2_118));
   NOR2_X1 i_257_2_119 (.A1(n_257_2_106), .A2(n_258), .ZN(n_257_2_119));
   NAND2_X1 i_257_2_120 (.A1(CPU_Bus[5]), .A2(n_257_2_119), .ZN(n_257_2_120));
   NOR2_X1 i_257_2_121 (.A1(n_257_2_109), .A2(n_258), .ZN(n_257_2_121));
   NAND2_X1 i_257_2_122 (.A1(CPU_Bus[1]), .A2(n_257_2_121), .ZN(n_257_2_122));
   NAND2_X1 i_257_2_123 (.A1(n_257_2_120), .A2(n_257_2_122), .ZN(n_257_2_123));
   NOR2_X1 i_257_2_124 (.A1(n_257_2_118), .A2(n_257_2_123), .ZN(n_257_2_124));
   NAND2_X1 i_257_2_125 (.A1(n_257_2_113), .A2(n_257_2_124), .ZN(n_257_2_125));
   NOR2_X1 i_257_2_126 (.A1(n_257_2_95), .A2(n_257_2_125), .ZN(n_257_2_126));
   NAND2_X1 i_257_2_127 (.A1(n_257_2_65), .A2(n_257_2_126), .ZN(n_257_14));
   NAND2_X1 i_257_4_0 (.A1(n_257_4_49), .A2(n_257_4_0), .ZN(n_257_15));
   NAND2_X1 i_257_4_1 (.A1(n_257_4_1), .A2(n_257_4_48), .ZN(n_257_4_0));
   NAND2_X1 i_257_4_2 (.A1(n_257_4_25), .A2(n_257_4_2), .ZN(n_257_4_1));
   NAND3_X1 i_257_4_3 (.A1(n_257_4_14), .A2(n_257_4_3), .A3(n_257), .ZN(
      n_257_4_2));
   NAND3_X1 i_257_4_4 (.A1(n_257_4_9), .A2(n_257_4_4), .A3(n_256), .ZN(n_257_4_3));
   NAND3_X1 i_257_4_5 (.A1(n_257_4_7), .A2(n_257_4_5), .A3(n_255), .ZN(n_257_4_4));
   NAND2_X1 i_257_4_6 (.A1(n_257_4_6), .A2(n_257_4_95), .ZN(n_257_4_5));
   INV_X1 i_257_4_7 (.A(CPU_Bus[11]), .ZN(n_257_4_6));
   NAND2_X1 i_257_4_8 (.A1(n_257_4_8), .A2(n_254), .ZN(n_257_4_7));
   INV_X1 i_257_4_9 (.A(CPU_Bus[12]), .ZN(n_257_4_8));
   NAND3_X1 i_257_4_10 (.A1(n_257_4_12), .A2(n_257_4_10), .A3(n_257_4_96), 
      .ZN(n_257_4_9));
   NAND2_X1 i_257_4_11 (.A1(n_257_4_11), .A2(n_254), .ZN(n_257_4_10));
   INV_X1 i_257_4_12 (.A(CPU_Bus[10]), .ZN(n_257_4_11));
   NAND2_X1 i_257_4_13 (.A1(n_257_4_13), .A2(n_257_4_95), .ZN(n_257_4_12));
   INV_X1 i_257_4_14 (.A(CPU_Bus[9]), .ZN(n_257_4_13));
   NAND3_X1 i_257_4_15 (.A1(n_257_4_20), .A2(n_257_4_15), .A3(n_257_4_97), 
      .ZN(n_257_4_14));
   NAND3_X1 i_257_4_16 (.A1(n_257_4_18), .A2(n_257_4_16), .A3(n_257_4_96), 
      .ZN(n_257_4_15));
   NAND2_X1 i_257_4_17 (.A1(n_257_4_17), .A2(n_257_4_95), .ZN(n_257_4_16));
   INV_X1 i_257_4_18 (.A(CPU_Bus[5]), .ZN(n_257_4_17));
   NAND2_X1 i_257_4_19 (.A1(n_257_4_19), .A2(n_254), .ZN(n_257_4_18));
   INV_X1 i_257_4_20 (.A(CPU_Bus[6]), .ZN(n_257_4_19));
   NAND3_X1 i_257_4_21 (.A1(n_257_4_23), .A2(n_257_4_21), .A3(n_255), .ZN(
      n_257_4_20));
   NAND2_X1 i_257_4_22 (.A1(n_257_4_22), .A2(n_254), .ZN(n_257_4_21));
   INV_X1 i_257_4_23 (.A(CPU_Bus[8]), .ZN(n_257_4_22));
   NAND2_X1 i_257_4_24 (.A1(n_257_4_24), .A2(n_257_4_95), .ZN(n_257_4_23));
   INV_X1 i_257_4_25 (.A(CPU_Bus[7]), .ZN(n_257_4_24));
   NAND3_X1 i_257_4_26 (.A1(n_257_4_37), .A2(n_257_4_26), .A3(n_257_4_98), 
      .ZN(n_257_4_25));
   NAND3_X1 i_257_4_27 (.A1(n_257_4_32), .A2(n_257_4_27), .A3(n_256), .ZN(
      n_257_4_26));
   NAND3_X1 i_257_4_28 (.A1(n_257_4_30), .A2(n_257_4_28), .A3(n_255), .ZN(
      n_257_4_27));
   NAND2_X1 i_257_4_29 (.A1(n_257_4_29), .A2(n_257_4_95), .ZN(n_257_4_28));
   INV_X1 i_257_4_30 (.A(CPU_Bus[3]), .ZN(n_257_4_29));
   NAND2_X1 i_257_4_31 (.A1(n_257_4_31), .A2(n_254), .ZN(n_257_4_30));
   INV_X1 i_257_4_32 (.A(CPU_Bus[4]), .ZN(n_257_4_31));
   NAND3_X1 i_257_4_33 (.A1(n_257_4_35), .A2(n_257_4_33), .A3(n_257_4_96), 
      .ZN(n_257_4_32));
   NAND2_X1 i_257_4_34 (.A1(n_257_4_34), .A2(n_254), .ZN(n_257_4_33));
   INV_X1 i_257_4_35 (.A(CPU_Bus[2]), .ZN(n_257_4_34));
   NAND2_X1 i_257_4_36 (.A1(n_257_4_36), .A2(n_257_4_95), .ZN(n_257_4_35));
   INV_X1 i_257_4_37 (.A(CPU_Bus[1]), .ZN(n_257_4_36));
   NAND3_X1 i_257_4_38 (.A1(n_257_4_43), .A2(n_257_4_38), .A3(n_257_4_97), 
      .ZN(n_257_4_37));
   NAND3_X1 i_257_4_39 (.A1(n_257_4_41), .A2(n_257_4_39), .A3(n_257_4_96), 
      .ZN(n_257_4_38));
   NAND2_X1 i_257_4_40 (.A1(n_257_4_40), .A2(n_257_4_95), .ZN(n_257_4_39));
   INV_X1 i_257_4_41 (.A(CPU_Bus[29]), .ZN(n_257_4_40));
   NAND2_X1 i_257_4_42 (.A1(n_257_4_42), .A2(n_254), .ZN(n_257_4_41));
   INV_X1 i_257_4_43 (.A(CPU_Bus[30]), .ZN(n_257_4_42));
   NAND3_X1 i_257_4_44 (.A1(n_257_4_46), .A2(n_257_4_44), .A3(n_255), .ZN(
      n_257_4_43));
   NAND2_X1 i_257_4_45 (.A1(n_257_4_45), .A2(n_254), .ZN(n_257_4_44));
   INV_X1 i_257_4_46 (.A(CPU_Bus[0]), .ZN(n_257_4_45));
   NAND2_X1 i_257_4_47 (.A1(n_257_4_47), .A2(n_257_4_95), .ZN(n_257_4_46));
   INV_X1 i_257_4_48 (.A(CPU_Bus[31]), .ZN(n_257_4_47));
   INV_X1 i_257_4_49 (.A(n_258), .ZN(n_257_4_48));
   NAND2_X1 i_257_4_50 (.A1(n_257_4_50), .A2(n_258), .ZN(n_257_4_49));
   NAND2_X1 i_257_4_51 (.A1(n_257_4_74), .A2(n_257_4_51), .ZN(n_257_4_50));
   NAND3_X1 i_257_4_52 (.A1(n_257_4_63), .A2(n_257_4_52), .A3(n_257), .ZN(
      n_257_4_51));
   NAND3_X1 i_257_4_53 (.A1(n_257_4_58), .A2(n_257_4_53), .A3(n_256), .ZN(
      n_257_4_52));
   NAND3_X1 i_257_4_54 (.A1(n_257_4_56), .A2(n_257_4_54), .A3(n_257_4_96), 
      .ZN(n_257_4_53));
   NAND2_X1 i_257_4_55 (.A1(n_257_4_55), .A2(n_254), .ZN(n_257_4_54));
   INV_X1 i_257_4_56 (.A(CPU_Bus[26]), .ZN(n_257_4_55));
   NAND2_X1 i_257_4_57 (.A1(n_257_4_57), .A2(n_257_4_95), .ZN(n_257_4_56));
   INV_X1 i_257_4_58 (.A(CPU_Bus[25]), .ZN(n_257_4_57));
   NAND3_X1 i_257_4_59 (.A1(n_257_4_61), .A2(n_257_4_59), .A3(n_255), .ZN(
      n_257_4_58));
   NAND2_X1 i_257_4_60 (.A1(n_257_4_60), .A2(n_254), .ZN(n_257_4_59));
   INV_X1 i_257_4_61 (.A(CPU_Bus[28]), .ZN(n_257_4_60));
   NAND2_X1 i_257_4_62 (.A1(n_257_4_62), .A2(n_257_4_95), .ZN(n_257_4_61));
   INV_X1 i_257_4_63 (.A(CPU_Bus[27]), .ZN(n_257_4_62));
   NAND3_X1 i_257_4_64 (.A1(n_257_4_69), .A2(n_257_4_64), .A3(n_257_4_97), 
      .ZN(n_257_4_63));
   NAND3_X1 i_257_4_65 (.A1(n_257_4_67), .A2(n_257_4_65), .A3(n_255), .ZN(
      n_257_4_64));
   NAND2_X1 i_257_4_66 (.A1(n_257_4_66), .A2(n_254), .ZN(n_257_4_65));
   INV_X1 i_257_4_67 (.A(CPU_Bus[24]), .ZN(n_257_4_66));
   NAND2_X1 i_257_4_68 (.A1(n_257_4_68), .A2(n_257_4_95), .ZN(n_257_4_67));
   INV_X1 i_257_4_69 (.A(CPU_Bus[23]), .ZN(n_257_4_68));
   NAND3_X1 i_257_4_70 (.A1(n_257_4_72), .A2(n_257_4_70), .A3(n_257_4_96), 
      .ZN(n_257_4_69));
   NAND2_X1 i_257_4_71 (.A1(n_257_4_71), .A2(n_254), .ZN(n_257_4_70));
   INV_X1 i_257_4_72 (.A(CPU_Bus[22]), .ZN(n_257_4_71));
   NAND2_X1 i_257_4_73 (.A1(n_257_4_73), .A2(n_257_4_95), .ZN(n_257_4_72));
   INV_X1 i_257_4_74 (.A(CPU_Bus[21]), .ZN(n_257_4_73));
   NAND3_X1 i_257_4_75 (.A1(n_257_4_86), .A2(n_257_4_98), .A3(n_257_4_75), 
      .ZN(n_257_4_74));
   NAND3_X1 i_257_4_76 (.A1(n_257_4_81), .A2(n_257_4_76), .A3(n_256), .ZN(
      n_257_4_75));
   NAND3_X1 i_257_4_77 (.A1(n_257_4_79), .A2(n_257_4_77), .A3(n_257_4_96), 
      .ZN(n_257_4_76));
   NAND2_X1 i_257_4_78 (.A1(n_257_4_78), .A2(n_254), .ZN(n_257_4_77));
   INV_X1 i_257_4_79 (.A(CPU_Bus[18]), .ZN(n_257_4_78));
   NAND2_X1 i_257_4_80 (.A1(n_257_4_80), .A2(n_257_4_95), .ZN(n_257_4_79));
   INV_X1 i_257_4_81 (.A(CPU_Bus[17]), .ZN(n_257_4_80));
   NAND3_X1 i_257_4_82 (.A1(n_257_4_84), .A2(n_257_4_82), .A3(n_255), .ZN(
      n_257_4_81));
   NAND2_X1 i_257_4_83 (.A1(n_257_4_83), .A2(n_254), .ZN(n_257_4_82));
   INV_X1 i_257_4_84 (.A(CPU_Bus[20]), .ZN(n_257_4_83));
   NAND2_X1 i_257_4_85 (.A1(n_257_4_85), .A2(n_257_4_95), .ZN(n_257_4_84));
   INV_X1 i_257_4_86 (.A(CPU_Bus[19]), .ZN(n_257_4_85));
   NAND3_X1 i_257_4_87 (.A1(n_257_4_92), .A2(n_257_4_97), .A3(n_257_4_87), 
      .ZN(n_257_4_86));
   NAND3_X1 i_257_4_88 (.A1(n_257_4_90), .A2(n_257_4_88), .A3(n_255), .ZN(
      n_257_4_87));
   NAND2_X1 i_257_4_89 (.A1(n_257_4_89), .A2(n_254), .ZN(n_257_4_88));
   INV_X1 i_257_4_90 (.A(CPU_Bus[16]), .ZN(n_257_4_89));
   NAND2_X1 i_257_4_91 (.A1(n_257_4_91), .A2(n_257_4_95), .ZN(n_257_4_90));
   INV_X1 i_257_4_92 (.A(CPU_Bus[15]), .ZN(n_257_4_91));
   OAI211_X1 i_257_4_93 (.A(n_257_4_93), .B(n_257_4_96), .C1(n_257_4_95), 
      .C2(CPU_Bus[14]), .ZN(n_257_4_92));
   NAND2_X1 i_257_4_94 (.A1(n_257_4_94), .A2(n_257_4_95), .ZN(n_257_4_93));
   INV_X1 i_257_4_95 (.A(CPU_Bus[13]), .ZN(n_257_4_94));
   INV_X1 i_257_4_96 (.A(n_254), .ZN(n_257_4_95));
   INV_X1 i_257_4_97 (.A(n_255), .ZN(n_257_4_96));
   INV_X1 i_257_4_98 (.A(n_256), .ZN(n_257_4_97));
   INV_X1 i_257_4_99 (.A(n_257), .ZN(n_257_4_98));
   NAND2_X1 i_257_5_0 (.A1(n_257_5_49), .A2(n_257_5_0), .ZN(n_257_16));
   NAND2_X1 i_257_5_1 (.A1(n_257_5_1), .A2(n_257_5_48), .ZN(n_257_5_0));
   NAND2_X1 i_257_5_2 (.A1(n_257_5_25), .A2(n_257_5_2), .ZN(n_257_5_1));
   NAND3_X1 i_257_5_3 (.A1(n_257_5_14), .A2(n_257_5_3), .A3(n_257), .ZN(
      n_257_5_2));
   NAND3_X1 i_257_5_4 (.A1(n_257_5_9), .A2(n_257_5_4), .A3(n_256), .ZN(n_257_5_3));
   NAND3_X1 i_257_5_5 (.A1(n_257_5_7), .A2(n_257_5_5), .A3(n_255), .ZN(n_257_5_4));
   NAND2_X1 i_257_5_6 (.A1(n_257_5_6), .A2(n_257_5_95), .ZN(n_257_5_5));
   INV_X1 i_257_5_7 (.A(CPU_Bus[10]), .ZN(n_257_5_6));
   NAND2_X1 i_257_5_8 (.A1(n_257_5_8), .A2(n_254), .ZN(n_257_5_7));
   INV_X1 i_257_5_9 (.A(CPU_Bus[11]), .ZN(n_257_5_8));
   NAND3_X1 i_257_5_10 (.A1(n_257_5_12), .A2(n_257_5_10), .A3(n_257_5_96), 
      .ZN(n_257_5_9));
   NAND2_X1 i_257_5_11 (.A1(n_257_5_11), .A2(n_254), .ZN(n_257_5_10));
   INV_X1 i_257_5_12 (.A(CPU_Bus[9]), .ZN(n_257_5_11));
   NAND2_X1 i_257_5_13 (.A1(n_257_5_13), .A2(n_257_5_95), .ZN(n_257_5_12));
   INV_X1 i_257_5_14 (.A(CPU_Bus[8]), .ZN(n_257_5_13));
   NAND3_X1 i_257_5_15 (.A1(n_257_5_20), .A2(n_257_5_15), .A3(n_257_5_97), 
      .ZN(n_257_5_14));
   NAND3_X1 i_257_5_16 (.A1(n_257_5_18), .A2(n_257_5_16), .A3(n_257_5_96), 
      .ZN(n_257_5_15));
   NAND2_X1 i_257_5_17 (.A1(n_257_5_17), .A2(n_257_5_95), .ZN(n_257_5_16));
   INV_X1 i_257_5_18 (.A(CPU_Bus[4]), .ZN(n_257_5_17));
   NAND2_X1 i_257_5_19 (.A1(n_257_5_19), .A2(n_254), .ZN(n_257_5_18));
   INV_X1 i_257_5_20 (.A(CPU_Bus[5]), .ZN(n_257_5_19));
   NAND3_X1 i_257_5_21 (.A1(n_257_5_23), .A2(n_257_5_21), .A3(n_255), .ZN(
      n_257_5_20));
   NAND2_X1 i_257_5_22 (.A1(n_257_5_22), .A2(n_254), .ZN(n_257_5_21));
   INV_X1 i_257_5_23 (.A(CPU_Bus[7]), .ZN(n_257_5_22));
   NAND2_X1 i_257_5_24 (.A1(n_257_5_24), .A2(n_257_5_95), .ZN(n_257_5_23));
   INV_X1 i_257_5_25 (.A(CPU_Bus[6]), .ZN(n_257_5_24));
   NAND3_X1 i_257_5_26 (.A1(n_257_5_37), .A2(n_257_5_26), .A3(n_257_5_98), 
      .ZN(n_257_5_25));
   NAND3_X1 i_257_5_27 (.A1(n_257_5_32), .A2(n_257_5_27), .A3(n_256), .ZN(
      n_257_5_26));
   NAND3_X1 i_257_5_28 (.A1(n_257_5_30), .A2(n_257_5_28), .A3(n_255), .ZN(
      n_257_5_27));
   NAND2_X1 i_257_5_29 (.A1(n_257_5_29), .A2(n_257_5_95), .ZN(n_257_5_28));
   INV_X1 i_257_5_30 (.A(CPU_Bus[2]), .ZN(n_257_5_29));
   NAND2_X1 i_257_5_31 (.A1(n_257_5_31), .A2(n_254), .ZN(n_257_5_30));
   INV_X1 i_257_5_32 (.A(CPU_Bus[3]), .ZN(n_257_5_31));
   NAND3_X1 i_257_5_33 (.A1(n_257_5_35), .A2(n_257_5_33), .A3(n_257_5_96), 
      .ZN(n_257_5_32));
   NAND2_X1 i_257_5_34 (.A1(n_257_5_34), .A2(n_254), .ZN(n_257_5_33));
   INV_X1 i_257_5_35 (.A(CPU_Bus[1]), .ZN(n_257_5_34));
   NAND2_X1 i_257_5_36 (.A1(n_257_5_36), .A2(n_257_5_95), .ZN(n_257_5_35));
   INV_X1 i_257_5_37 (.A(CPU_Bus[0]), .ZN(n_257_5_36));
   NAND3_X1 i_257_5_38 (.A1(n_257_5_43), .A2(n_257_5_38), .A3(n_257_5_97), 
      .ZN(n_257_5_37));
   NAND3_X1 i_257_5_39 (.A1(n_257_5_41), .A2(n_257_5_39), .A3(n_257_5_96), 
      .ZN(n_257_5_38));
   NAND2_X1 i_257_5_40 (.A1(n_257_5_40), .A2(n_257_5_95), .ZN(n_257_5_39));
   INV_X1 i_257_5_41 (.A(CPU_Bus[28]), .ZN(n_257_5_40));
   NAND2_X1 i_257_5_42 (.A1(n_257_5_42), .A2(n_254), .ZN(n_257_5_41));
   INV_X1 i_257_5_43 (.A(CPU_Bus[29]), .ZN(n_257_5_42));
   NAND3_X1 i_257_5_44 (.A1(n_257_5_46), .A2(n_257_5_44), .A3(n_255), .ZN(
      n_257_5_43));
   NAND2_X1 i_257_5_45 (.A1(n_257_5_45), .A2(n_254), .ZN(n_257_5_44));
   INV_X1 i_257_5_46 (.A(CPU_Bus[31]), .ZN(n_257_5_45));
   NAND2_X1 i_257_5_47 (.A1(n_257_5_47), .A2(n_257_5_95), .ZN(n_257_5_46));
   INV_X1 i_257_5_48 (.A(CPU_Bus[30]), .ZN(n_257_5_47));
   INV_X1 i_257_5_49 (.A(n_258), .ZN(n_257_5_48));
   NAND2_X1 i_257_5_50 (.A1(n_257_5_50), .A2(n_258), .ZN(n_257_5_49));
   NAND2_X1 i_257_5_51 (.A1(n_257_5_74), .A2(n_257_5_51), .ZN(n_257_5_50));
   NAND3_X1 i_257_5_52 (.A1(n_257_5_63), .A2(n_257_5_52), .A3(n_257), .ZN(
      n_257_5_51));
   NAND3_X1 i_257_5_53 (.A1(n_257_5_58), .A2(n_257_5_53), .A3(n_256), .ZN(
      n_257_5_52));
   NAND3_X1 i_257_5_54 (.A1(n_257_5_56), .A2(n_257_5_54), .A3(n_257_5_96), 
      .ZN(n_257_5_53));
   NAND2_X1 i_257_5_55 (.A1(n_257_5_55), .A2(n_254), .ZN(n_257_5_54));
   INV_X1 i_257_5_56 (.A(CPU_Bus[25]), .ZN(n_257_5_55));
   NAND2_X1 i_257_5_57 (.A1(n_257_5_57), .A2(n_257_5_95), .ZN(n_257_5_56));
   INV_X1 i_257_5_58 (.A(CPU_Bus[24]), .ZN(n_257_5_57));
   NAND3_X1 i_257_5_59 (.A1(n_257_5_61), .A2(n_257_5_59), .A3(n_255), .ZN(
      n_257_5_58));
   NAND2_X1 i_257_5_60 (.A1(n_257_5_60), .A2(n_254), .ZN(n_257_5_59));
   INV_X1 i_257_5_61 (.A(CPU_Bus[27]), .ZN(n_257_5_60));
   NAND2_X1 i_257_5_62 (.A1(n_257_5_62), .A2(n_257_5_95), .ZN(n_257_5_61));
   INV_X1 i_257_5_63 (.A(CPU_Bus[26]), .ZN(n_257_5_62));
   NAND3_X1 i_257_5_64 (.A1(n_257_5_69), .A2(n_257_5_64), .A3(n_257_5_97), 
      .ZN(n_257_5_63));
   NAND3_X1 i_257_5_65 (.A1(n_257_5_67), .A2(n_257_5_65), .A3(n_255), .ZN(
      n_257_5_64));
   NAND2_X1 i_257_5_66 (.A1(n_257_5_66), .A2(n_254), .ZN(n_257_5_65));
   INV_X1 i_257_5_67 (.A(CPU_Bus[23]), .ZN(n_257_5_66));
   NAND2_X1 i_257_5_68 (.A1(n_257_5_68), .A2(n_257_5_95), .ZN(n_257_5_67));
   INV_X1 i_257_5_69 (.A(CPU_Bus[22]), .ZN(n_257_5_68));
   NAND3_X1 i_257_5_70 (.A1(n_257_5_72), .A2(n_257_5_70), .A3(n_257_5_96), 
      .ZN(n_257_5_69));
   NAND2_X1 i_257_5_71 (.A1(n_257_5_71), .A2(n_254), .ZN(n_257_5_70));
   INV_X1 i_257_5_72 (.A(CPU_Bus[21]), .ZN(n_257_5_71));
   NAND2_X1 i_257_5_73 (.A1(n_257_5_73), .A2(n_257_5_95), .ZN(n_257_5_72));
   INV_X1 i_257_5_74 (.A(CPU_Bus[20]), .ZN(n_257_5_73));
   NAND3_X1 i_257_5_75 (.A1(n_257_5_86), .A2(n_257_5_98), .A3(n_257_5_75), 
      .ZN(n_257_5_74));
   NAND3_X1 i_257_5_76 (.A1(n_257_5_81), .A2(n_257_5_76), .A3(n_256), .ZN(
      n_257_5_75));
   NAND3_X1 i_257_5_77 (.A1(n_257_5_79), .A2(n_257_5_77), .A3(n_257_5_96), 
      .ZN(n_257_5_76));
   NAND2_X1 i_257_5_78 (.A1(n_257_5_78), .A2(n_254), .ZN(n_257_5_77));
   INV_X1 i_257_5_79 (.A(CPU_Bus[17]), .ZN(n_257_5_78));
   NAND2_X1 i_257_5_80 (.A1(n_257_5_80), .A2(n_257_5_95), .ZN(n_257_5_79));
   INV_X1 i_257_5_81 (.A(CPU_Bus[16]), .ZN(n_257_5_80));
   NAND3_X1 i_257_5_82 (.A1(n_257_5_84), .A2(n_257_5_82), .A3(n_255), .ZN(
      n_257_5_81));
   NAND2_X1 i_257_5_83 (.A1(n_257_5_83), .A2(n_254), .ZN(n_257_5_82));
   INV_X1 i_257_5_84 (.A(CPU_Bus[19]), .ZN(n_257_5_83));
   NAND2_X1 i_257_5_85 (.A1(n_257_5_85), .A2(n_257_5_95), .ZN(n_257_5_84));
   INV_X1 i_257_5_86 (.A(CPU_Bus[18]), .ZN(n_257_5_85));
   NAND3_X1 i_257_5_87 (.A1(n_257_5_92), .A2(n_257_5_97), .A3(n_257_5_87), 
      .ZN(n_257_5_86));
   NAND3_X1 i_257_5_88 (.A1(n_257_5_90), .A2(n_257_5_88), .A3(n_255), .ZN(
      n_257_5_87));
   NAND2_X1 i_257_5_89 (.A1(n_257_5_89), .A2(n_254), .ZN(n_257_5_88));
   INV_X1 i_257_5_90 (.A(CPU_Bus[15]), .ZN(n_257_5_89));
   NAND2_X1 i_257_5_91 (.A1(n_257_5_91), .A2(n_257_5_95), .ZN(n_257_5_90));
   INV_X1 i_257_5_92 (.A(CPU_Bus[14]), .ZN(n_257_5_91));
   OAI211_X1 i_257_5_93 (.A(n_257_5_93), .B(n_257_5_96), .C1(n_257_5_95), 
      .C2(CPU_Bus[13]), .ZN(n_257_5_92));
   NAND2_X1 i_257_5_94 (.A1(n_257_5_94), .A2(n_257_5_95), .ZN(n_257_5_93));
   INV_X1 i_257_5_95 (.A(CPU_Bus[12]), .ZN(n_257_5_94));
   INV_X1 i_257_5_96 (.A(n_254), .ZN(n_257_5_95));
   INV_X1 i_257_5_97 (.A(n_255), .ZN(n_257_5_96));
   INV_X1 i_257_5_98 (.A(n_256), .ZN(n_257_5_97));
   INV_X1 i_257_5_99 (.A(n_257), .ZN(n_257_5_98));
   INV_X1 i_257_7_0 (.A(n_257_7_0), .ZN(n_257_17));
   NAND2_X1 i_257_7_1 (.A1(n_257_7_49), .A2(n_257_7_1), .ZN(n_257_7_0));
   NAND3_X1 i_257_7_2 (.A1(n_257_7_25), .A2(n_257_7_2), .A3(n_257_7_48), 
      .ZN(n_257_7_1));
   NAND3_X1 i_257_7_3 (.A1(n_257_7_14), .A2(n_257_7_3), .A3(n_257), .ZN(
      n_257_7_2));
   NAND3_X1 i_257_7_4 (.A1(n_257_7_9), .A2(n_257_7_4), .A3(n_257_7_85), .ZN(
      n_257_7_3));
   NAND3_X1 i_257_7_5 (.A1(n_257_7_7), .A2(n_257_7_5), .A3(n_257_7_96), .ZN(
      n_257_7_4));
   NAND2_X1 i_257_7_6 (.A1(n_257_7_6), .A2(n_257_7_95), .ZN(n_257_7_5));
   INV_X1 i_257_7_7 (.A(CPU_Bus[3]), .ZN(n_257_7_6));
   NAND2_X1 i_257_7_8 (.A1(n_257_7_8), .A2(n_254), .ZN(n_257_7_7));
   INV_X1 i_257_7_9 (.A(CPU_Bus[4]), .ZN(n_257_7_8));
   NAND3_X1 i_257_7_10 (.A1(n_257_7_12), .A2(n_257_7_10), .A3(n_255), .ZN(
      n_257_7_9));
   NAND2_X1 i_257_7_11 (.A1(n_257_7_11), .A2(n_257_7_95), .ZN(n_257_7_10));
   INV_X1 i_257_7_12 (.A(CPU_Bus[5]), .ZN(n_257_7_11));
   NAND2_X1 i_257_7_13 (.A1(n_257_7_13), .A2(n_254), .ZN(n_257_7_12));
   INV_X1 i_257_7_14 (.A(CPU_Bus[6]), .ZN(n_257_7_13));
   NAND3_X1 i_257_7_15 (.A1(n_257_7_20), .A2(n_257_7_15), .A3(n_256), .ZN(
      n_257_7_14));
   NAND3_X1 i_257_7_16 (.A1(n_257_7_18), .A2(n_257_7_16), .A3(n_257_7_96), 
      .ZN(n_257_7_15));
   NAND2_X1 i_257_7_17 (.A1(n_257_7_17), .A2(n_257_7_95), .ZN(n_257_7_16));
   INV_X1 i_257_7_18 (.A(CPU_Bus[7]), .ZN(n_257_7_17));
   NAND2_X1 i_257_7_19 (.A1(n_257_7_19), .A2(n_254), .ZN(n_257_7_18));
   INV_X1 i_257_7_20 (.A(CPU_Bus[8]), .ZN(n_257_7_19));
   NAND3_X1 i_257_7_21 (.A1(n_257_7_23), .A2(n_257_7_21), .A3(n_255), .ZN(
      n_257_7_20));
   NAND2_X1 i_257_7_22 (.A1(n_257_7_22), .A2(n_257_7_95), .ZN(n_257_7_21));
   INV_X1 i_257_7_23 (.A(CPU_Bus[9]), .ZN(n_257_7_22));
   NAND2_X1 i_257_7_24 (.A1(n_257_7_24), .A2(n_254), .ZN(n_257_7_23));
   INV_X1 i_257_7_25 (.A(CPU_Bus[10]), .ZN(n_257_7_24));
   NAND3_X1 i_257_7_26 (.A1(n_257_7_37), .A2(n_257_7_26), .A3(n_257_7_97), 
      .ZN(n_257_7_25));
   NAND3_X1 i_257_7_27 (.A1(n_257_7_32), .A2(n_257_7_27), .A3(n_256), .ZN(
      n_257_7_26));
   NAND3_X1 i_257_7_28 (.A1(n_257_7_30), .A2(n_257_7_28), .A3(n_255), .ZN(
      n_257_7_27));
   NAND2_X1 i_257_7_29 (.A1(n_257_7_29), .A2(n_254), .ZN(n_257_7_28));
   INV_X1 i_257_7_30 (.A(CPU_Bus[2]), .ZN(n_257_7_29));
   NAND2_X1 i_257_7_31 (.A1(n_257_7_31), .A2(n_257_7_95), .ZN(n_257_7_30));
   INV_X1 i_257_7_32 (.A(CPU_Bus[1]), .ZN(n_257_7_31));
   NAND3_X1 i_257_7_33 (.A1(n_257_7_35), .A2(n_257_7_33), .A3(n_257_7_96), 
      .ZN(n_257_7_32));
   NAND2_X1 i_257_7_34 (.A1(n_257_7_34), .A2(n_257_7_95), .ZN(n_257_7_33));
   INV_X1 i_257_7_35 (.A(CPU_Bus[31]), .ZN(n_257_7_34));
   NAND2_X1 i_257_7_36 (.A1(n_257_7_36), .A2(n_254), .ZN(n_257_7_35));
   INV_X1 i_257_7_37 (.A(CPU_Bus[0]), .ZN(n_257_7_36));
   NAND3_X1 i_257_7_38 (.A1(n_257_7_43), .A2(n_257_7_38), .A3(n_257_7_85), 
      .ZN(n_257_7_37));
   NAND3_X1 i_257_7_39 (.A1(n_257_7_41), .A2(n_257_7_39), .A3(n_255), .ZN(
      n_257_7_38));
   NAND2_X1 i_257_7_40 (.A1(n_257_7_40), .A2(n_254), .ZN(n_257_7_39));
   INV_X1 i_257_7_41 (.A(CPU_Bus[30]), .ZN(n_257_7_40));
   NAND2_X1 i_257_7_42 (.A1(n_257_7_42), .A2(n_257_7_95), .ZN(n_257_7_41));
   INV_X1 i_257_7_43 (.A(CPU_Bus[29]), .ZN(n_257_7_42));
   NAND3_X1 i_257_7_44 (.A1(n_257_7_46), .A2(n_257_7_44), .A3(n_257_7_96), 
      .ZN(n_257_7_43));
   NAND2_X1 i_257_7_45 (.A1(n_257_7_45), .A2(n_257_7_95), .ZN(n_257_7_44));
   INV_X1 i_257_7_46 (.A(CPU_Bus[27]), .ZN(n_257_7_45));
   NAND2_X1 i_257_7_47 (.A1(n_257_7_47), .A2(n_254), .ZN(n_257_7_46));
   INV_X1 i_257_7_48 (.A(CPU_Bus[28]), .ZN(n_257_7_47));
   INV_X1 i_257_7_49 (.A(n_258), .ZN(n_257_7_48));
   NAND3_X1 i_257_7_50 (.A1(n_257_7_73), .A2(n_257_7_50), .A3(n_258), .ZN(
      n_257_7_49));
   NAND3_X1 i_257_7_51 (.A1(n_257_7_62), .A2(n_257_7_51), .A3(n_257), .ZN(
      n_257_7_50));
   NAND3_X1 i_257_7_52 (.A1(n_257_7_57), .A2(n_257_7_52), .A3(n_257_7_85), 
      .ZN(n_257_7_51));
   NAND3_X1 i_257_7_53 (.A1(n_257_7_55), .A2(n_257_7_53), .A3(n_257_7_96), 
      .ZN(n_257_7_52));
   NAND2_X1 i_257_7_54 (.A1(n_257_7_54), .A2(n_257_7_95), .ZN(n_257_7_53));
   INV_X1 i_257_7_55 (.A(CPU_Bus[19]), .ZN(n_257_7_54));
   NAND2_X1 i_257_7_56 (.A1(n_257_7_56), .A2(n_254), .ZN(n_257_7_55));
   INV_X1 i_257_7_57 (.A(CPU_Bus[20]), .ZN(n_257_7_56));
   NAND3_X1 i_257_7_58 (.A1(n_257_7_60), .A2(n_257_7_58), .A3(n_255), .ZN(
      n_257_7_57));
   NAND2_X1 i_257_7_59 (.A1(n_257_7_59), .A2(n_254), .ZN(n_257_7_58));
   INV_X1 i_257_7_60 (.A(CPU_Bus[22]), .ZN(n_257_7_59));
   NAND2_X1 i_257_7_61 (.A1(n_257_7_61), .A2(n_257_7_95), .ZN(n_257_7_60));
   INV_X1 i_257_7_62 (.A(CPU_Bus[21]), .ZN(n_257_7_61));
   NAND3_X1 i_257_7_63 (.A1(n_257_7_68), .A2(n_257_7_63), .A3(n_256), .ZN(
      n_257_7_62));
   NAND3_X1 i_257_7_64 (.A1(n_257_7_66), .A2(n_257_7_64), .A3(n_257_7_96), 
      .ZN(n_257_7_63));
   NAND2_X1 i_257_7_65 (.A1(n_257_7_65), .A2(n_254), .ZN(n_257_7_64));
   INV_X1 i_257_7_66 (.A(CPU_Bus[24]), .ZN(n_257_7_65));
   NAND2_X1 i_257_7_67 (.A1(n_257_7_67), .A2(n_257_7_95), .ZN(n_257_7_66));
   INV_X1 i_257_7_68 (.A(CPU_Bus[23]), .ZN(n_257_7_67));
   NAND3_X1 i_257_7_69 (.A1(n_257_7_71), .A2(n_257_7_69), .A3(n_255), .ZN(
      n_257_7_68));
   NAND2_X1 i_257_7_70 (.A1(n_257_7_70), .A2(n_257_7_95), .ZN(n_257_7_69));
   INV_X1 i_257_7_71 (.A(CPU_Bus[25]), .ZN(n_257_7_70));
   NAND2_X1 i_257_7_72 (.A1(n_257_7_72), .A2(n_254), .ZN(n_257_7_71));
   INV_X1 i_257_7_73 (.A(CPU_Bus[26]), .ZN(n_257_7_72));
   NAND3_X1 i_257_7_74 (.A1(n_257_7_86), .A2(n_257_7_74), .A3(n_257_7_97), 
      .ZN(n_257_7_73));
   NAND3_X1 i_257_7_75 (.A1(n_257_7_80), .A2(n_257_7_75), .A3(n_257_7_85), 
      .ZN(n_257_7_74));
   NAND3_X1 i_257_7_76 (.A1(n_257_7_78), .A2(n_257_7_76), .A3(n_257_7_96), 
      .ZN(n_257_7_75));
   NAND2_X1 i_257_7_77 (.A1(n_257_7_77), .A2(n_254), .ZN(n_257_7_76));
   INV_X1 i_257_7_78 (.A(CPU_Bus[12]), .ZN(n_257_7_77));
   NAND2_X1 i_257_7_79 (.A1(n_257_7_79), .A2(n_257_7_95), .ZN(n_257_7_78));
   INV_X1 i_257_7_80 (.A(CPU_Bus[11]), .ZN(n_257_7_79));
   NAND3_X1 i_257_7_81 (.A1(n_257_7_83), .A2(n_257_7_81), .A3(n_255), .ZN(
      n_257_7_80));
   NAND2_X1 i_257_7_82 (.A1(n_257_7_82), .A2(n_254), .ZN(n_257_7_81));
   INV_X1 i_257_7_83 (.A(CPU_Bus[14]), .ZN(n_257_7_82));
   NAND2_X1 i_257_7_84 (.A1(n_257_7_84), .A2(n_257_7_95), .ZN(n_257_7_83));
   INV_X1 i_257_7_85 (.A(CPU_Bus[13]), .ZN(n_257_7_84));
   INV_X1 i_257_7_86 (.A(n_256), .ZN(n_257_7_85));
   NAND3_X1 i_257_7_87 (.A1(n_257_7_92), .A2(n_257_7_87), .A3(n_256), .ZN(
      n_257_7_86));
   NAND3_X1 i_257_7_88 (.A1(n_257_7_90), .A2(n_257_7_88), .A3(n_255), .ZN(
      n_257_7_87));
   NAND2_X1 i_257_7_89 (.A1(n_257_7_89), .A2(n_257_7_95), .ZN(n_257_7_88));
   INV_X1 i_257_7_90 (.A(CPU_Bus[17]), .ZN(n_257_7_89));
   NAND2_X1 i_257_7_91 (.A1(n_257_7_91), .A2(n_254), .ZN(n_257_7_90));
   INV_X1 i_257_7_92 (.A(CPU_Bus[18]), .ZN(n_257_7_91));
   OAI211_X1 i_257_7_93 (.A(n_257_7_93), .B(n_257_7_96), .C1(n_257_7_95), 
      .C2(CPU_Bus[16]), .ZN(n_257_7_92));
   NAND2_X1 i_257_7_94 (.A1(n_257_7_94), .A2(n_257_7_95), .ZN(n_257_7_93));
   INV_X1 i_257_7_95 (.A(CPU_Bus[15]), .ZN(n_257_7_94));
   INV_X1 i_257_7_96 (.A(n_254), .ZN(n_257_7_95));
   INV_X1 i_257_7_97 (.A(n_255), .ZN(n_257_7_96));
   INV_X1 i_257_7_98 (.A(n_257), .ZN(n_257_7_97));
   INV_X1 i_257_8_0 (.A(n_257_8_0), .ZN(n_257_18));
   NAND2_X1 i_257_8_1 (.A1(n_257_8_49), .A2(n_257_8_1), .ZN(n_257_8_0));
   NAND3_X1 i_257_8_2 (.A1(n_257_8_25), .A2(n_257_8_2), .A3(n_257_8_48), 
      .ZN(n_257_8_1));
   NAND3_X1 i_257_8_3 (.A1(n_257_8_14), .A2(n_257_8_3), .A3(n_257), .ZN(
      n_257_8_2));
   NAND3_X1 i_257_8_4 (.A1(n_257_8_9), .A2(n_257_8_4), .A3(n_257_8_85), .ZN(
      n_257_8_3));
   NAND3_X1 i_257_8_5 (.A1(n_257_8_7), .A2(n_257_8_5), .A3(n_257_8_96), .ZN(
      n_257_8_4));
   NAND2_X1 i_257_8_6 (.A1(n_257_8_6), .A2(n_257_8_95), .ZN(n_257_8_5));
   INV_X1 i_257_8_7 (.A(CPU_Bus[2]), .ZN(n_257_8_6));
   NAND2_X1 i_257_8_8 (.A1(n_257_8_8), .A2(n_254), .ZN(n_257_8_7));
   INV_X1 i_257_8_9 (.A(CPU_Bus[3]), .ZN(n_257_8_8));
   NAND3_X1 i_257_8_10 (.A1(n_257_8_12), .A2(n_257_8_10), .A3(n_255), .ZN(
      n_257_8_9));
   NAND2_X1 i_257_8_11 (.A1(n_257_8_11), .A2(n_257_8_95), .ZN(n_257_8_10));
   INV_X1 i_257_8_12 (.A(CPU_Bus[4]), .ZN(n_257_8_11));
   NAND2_X1 i_257_8_13 (.A1(n_257_8_13), .A2(n_254), .ZN(n_257_8_12));
   INV_X1 i_257_8_14 (.A(CPU_Bus[5]), .ZN(n_257_8_13));
   NAND3_X1 i_257_8_15 (.A1(n_257_8_20), .A2(n_257_8_15), .A3(n_256), .ZN(
      n_257_8_14));
   NAND3_X1 i_257_8_16 (.A1(n_257_8_18), .A2(n_257_8_16), .A3(n_257_8_96), 
      .ZN(n_257_8_15));
   NAND2_X1 i_257_8_17 (.A1(n_257_8_17), .A2(n_257_8_95), .ZN(n_257_8_16));
   INV_X1 i_257_8_18 (.A(CPU_Bus[6]), .ZN(n_257_8_17));
   NAND2_X1 i_257_8_19 (.A1(n_257_8_19), .A2(n_254), .ZN(n_257_8_18));
   INV_X1 i_257_8_20 (.A(CPU_Bus[7]), .ZN(n_257_8_19));
   NAND3_X1 i_257_8_21 (.A1(n_257_8_23), .A2(n_257_8_21), .A3(n_255), .ZN(
      n_257_8_20));
   NAND2_X1 i_257_8_22 (.A1(n_257_8_22), .A2(n_257_8_95), .ZN(n_257_8_21));
   INV_X1 i_257_8_23 (.A(CPU_Bus[8]), .ZN(n_257_8_22));
   NAND2_X1 i_257_8_24 (.A1(n_257_8_24), .A2(n_254), .ZN(n_257_8_23));
   INV_X1 i_257_8_25 (.A(CPU_Bus[9]), .ZN(n_257_8_24));
   NAND3_X1 i_257_8_26 (.A1(n_257_8_37), .A2(n_257_8_26), .A3(n_257_8_97), 
      .ZN(n_257_8_25));
   NAND3_X1 i_257_8_27 (.A1(n_257_8_32), .A2(n_257_8_27), .A3(n_256), .ZN(
      n_257_8_26));
   NAND3_X1 i_257_8_28 (.A1(n_257_8_30), .A2(n_257_8_28), .A3(n_255), .ZN(
      n_257_8_27));
   NAND2_X1 i_257_8_29 (.A1(n_257_8_29), .A2(n_254), .ZN(n_257_8_28));
   INV_X1 i_257_8_30 (.A(CPU_Bus[1]), .ZN(n_257_8_29));
   NAND2_X1 i_257_8_31 (.A1(n_257_8_31), .A2(n_257_8_95), .ZN(n_257_8_30));
   INV_X1 i_257_8_32 (.A(CPU_Bus[0]), .ZN(n_257_8_31));
   NAND3_X1 i_257_8_33 (.A1(n_257_8_35), .A2(n_257_8_33), .A3(n_257_8_96), 
      .ZN(n_257_8_32));
   NAND2_X1 i_257_8_34 (.A1(n_257_8_34), .A2(n_257_8_95), .ZN(n_257_8_33));
   INV_X1 i_257_8_35 (.A(CPU_Bus[30]), .ZN(n_257_8_34));
   NAND2_X1 i_257_8_36 (.A1(n_257_8_36), .A2(n_254), .ZN(n_257_8_35));
   INV_X1 i_257_8_37 (.A(CPU_Bus[31]), .ZN(n_257_8_36));
   NAND3_X1 i_257_8_38 (.A1(n_257_8_43), .A2(n_257_8_38), .A3(n_257_8_85), 
      .ZN(n_257_8_37));
   NAND3_X1 i_257_8_39 (.A1(n_257_8_41), .A2(n_257_8_39), .A3(n_255), .ZN(
      n_257_8_38));
   NAND2_X1 i_257_8_40 (.A1(n_257_8_40), .A2(n_254), .ZN(n_257_8_39));
   INV_X1 i_257_8_41 (.A(CPU_Bus[29]), .ZN(n_257_8_40));
   NAND2_X1 i_257_8_42 (.A1(n_257_8_42), .A2(n_257_8_95), .ZN(n_257_8_41));
   INV_X1 i_257_8_43 (.A(CPU_Bus[28]), .ZN(n_257_8_42));
   NAND3_X1 i_257_8_44 (.A1(n_257_8_46), .A2(n_257_8_44), .A3(n_257_8_96), 
      .ZN(n_257_8_43));
   NAND2_X1 i_257_8_45 (.A1(n_257_8_45), .A2(n_257_8_95), .ZN(n_257_8_44));
   INV_X1 i_257_8_46 (.A(CPU_Bus[26]), .ZN(n_257_8_45));
   NAND2_X1 i_257_8_47 (.A1(n_257_8_47), .A2(n_254), .ZN(n_257_8_46));
   INV_X1 i_257_8_48 (.A(CPU_Bus[27]), .ZN(n_257_8_47));
   INV_X1 i_257_8_49 (.A(n_258), .ZN(n_257_8_48));
   NAND3_X1 i_257_8_50 (.A1(n_257_8_73), .A2(n_257_8_50), .A3(n_258), .ZN(
      n_257_8_49));
   NAND3_X1 i_257_8_51 (.A1(n_257_8_62), .A2(n_257_8_51), .A3(n_257), .ZN(
      n_257_8_50));
   NAND3_X1 i_257_8_52 (.A1(n_257_8_57), .A2(n_257_8_52), .A3(n_257_8_85), 
      .ZN(n_257_8_51));
   NAND3_X1 i_257_8_53 (.A1(n_257_8_55), .A2(n_257_8_53), .A3(n_257_8_96), 
      .ZN(n_257_8_52));
   NAND2_X1 i_257_8_54 (.A1(n_257_8_54), .A2(n_257_8_95), .ZN(n_257_8_53));
   INV_X1 i_257_8_55 (.A(CPU_Bus[18]), .ZN(n_257_8_54));
   NAND2_X1 i_257_8_56 (.A1(n_257_8_56), .A2(n_254), .ZN(n_257_8_55));
   INV_X1 i_257_8_57 (.A(CPU_Bus[19]), .ZN(n_257_8_56));
   NAND3_X1 i_257_8_58 (.A1(n_257_8_60), .A2(n_257_8_58), .A3(n_255), .ZN(
      n_257_8_57));
   NAND2_X1 i_257_8_59 (.A1(n_257_8_59), .A2(n_254), .ZN(n_257_8_58));
   INV_X1 i_257_8_60 (.A(CPU_Bus[21]), .ZN(n_257_8_59));
   NAND2_X1 i_257_8_61 (.A1(n_257_8_61), .A2(n_257_8_95), .ZN(n_257_8_60));
   INV_X1 i_257_8_62 (.A(CPU_Bus[20]), .ZN(n_257_8_61));
   NAND3_X1 i_257_8_63 (.A1(n_257_8_68), .A2(n_257_8_63), .A3(n_256), .ZN(
      n_257_8_62));
   NAND3_X1 i_257_8_64 (.A1(n_257_8_66), .A2(n_257_8_64), .A3(n_257_8_96), 
      .ZN(n_257_8_63));
   NAND2_X1 i_257_8_65 (.A1(n_257_8_65), .A2(n_254), .ZN(n_257_8_64));
   INV_X1 i_257_8_66 (.A(CPU_Bus[23]), .ZN(n_257_8_65));
   NAND2_X1 i_257_8_67 (.A1(n_257_8_67), .A2(n_257_8_95), .ZN(n_257_8_66));
   INV_X1 i_257_8_68 (.A(CPU_Bus[22]), .ZN(n_257_8_67));
   NAND3_X1 i_257_8_69 (.A1(n_257_8_71), .A2(n_257_8_69), .A3(n_255), .ZN(
      n_257_8_68));
   NAND2_X1 i_257_8_70 (.A1(n_257_8_70), .A2(n_257_8_95), .ZN(n_257_8_69));
   INV_X1 i_257_8_71 (.A(CPU_Bus[24]), .ZN(n_257_8_70));
   NAND2_X1 i_257_8_72 (.A1(n_257_8_72), .A2(n_254), .ZN(n_257_8_71));
   INV_X1 i_257_8_73 (.A(CPU_Bus[25]), .ZN(n_257_8_72));
   NAND3_X1 i_257_8_74 (.A1(n_257_8_86), .A2(n_257_8_74), .A3(n_257_8_97), 
      .ZN(n_257_8_73));
   NAND3_X1 i_257_8_75 (.A1(n_257_8_80), .A2(n_257_8_75), .A3(n_257_8_85), 
      .ZN(n_257_8_74));
   NAND3_X1 i_257_8_76 (.A1(n_257_8_78), .A2(n_257_8_76), .A3(n_257_8_96), 
      .ZN(n_257_8_75));
   NAND2_X1 i_257_8_77 (.A1(n_257_8_77), .A2(n_254), .ZN(n_257_8_76));
   INV_X1 i_257_8_78 (.A(CPU_Bus[11]), .ZN(n_257_8_77));
   NAND2_X1 i_257_8_79 (.A1(n_257_8_79), .A2(n_257_8_95), .ZN(n_257_8_78));
   INV_X1 i_257_8_80 (.A(CPU_Bus[10]), .ZN(n_257_8_79));
   NAND3_X1 i_257_8_81 (.A1(n_257_8_83), .A2(n_257_8_81), .A3(n_255), .ZN(
      n_257_8_80));
   NAND2_X1 i_257_8_82 (.A1(n_257_8_82), .A2(n_254), .ZN(n_257_8_81));
   INV_X1 i_257_8_83 (.A(CPU_Bus[13]), .ZN(n_257_8_82));
   NAND2_X1 i_257_8_84 (.A1(n_257_8_84), .A2(n_257_8_95), .ZN(n_257_8_83));
   INV_X1 i_257_8_85 (.A(CPU_Bus[12]), .ZN(n_257_8_84));
   INV_X1 i_257_8_86 (.A(n_256), .ZN(n_257_8_85));
   NAND3_X1 i_257_8_87 (.A1(n_257_8_92), .A2(n_257_8_87), .A3(n_256), .ZN(
      n_257_8_86));
   NAND3_X1 i_257_8_88 (.A1(n_257_8_90), .A2(n_257_8_88), .A3(n_255), .ZN(
      n_257_8_87));
   NAND2_X1 i_257_8_89 (.A1(n_257_8_89), .A2(n_257_8_95), .ZN(n_257_8_88));
   INV_X1 i_257_8_90 (.A(CPU_Bus[16]), .ZN(n_257_8_89));
   NAND2_X1 i_257_8_91 (.A1(n_257_8_91), .A2(n_254), .ZN(n_257_8_90));
   INV_X1 i_257_8_92 (.A(CPU_Bus[17]), .ZN(n_257_8_91));
   OAI211_X1 i_257_8_93 (.A(n_257_8_93), .B(n_257_8_96), .C1(n_257_8_95), 
      .C2(CPU_Bus[15]), .ZN(n_257_8_92));
   NAND2_X1 i_257_8_94 (.A1(n_257_8_94), .A2(n_257_8_95), .ZN(n_257_8_93));
   INV_X1 i_257_8_95 (.A(CPU_Bus[14]), .ZN(n_257_8_94));
   INV_X1 i_257_8_96 (.A(n_254), .ZN(n_257_8_95));
   INV_X1 i_257_8_97 (.A(n_255), .ZN(n_257_8_96));
   INV_X1 i_257_8_98 (.A(n_257), .ZN(n_257_8_97));
   NAND2_X1 i_257_9_0 (.A1(n_257_9_49), .A2(n_257_9_0), .ZN(n_257_19));
   NAND2_X1 i_257_9_1 (.A1(n_257_9_1), .A2(n_257_9_48), .ZN(n_257_9_0));
   NAND2_X1 i_257_9_2 (.A1(n_257_9_25), .A2(n_257_9_2), .ZN(n_257_9_1));
   NAND3_X1 i_257_9_3 (.A1(n_257_9_14), .A2(n_257_9_3), .A3(n_257), .ZN(
      n_257_9_2));
   NAND3_X1 i_257_9_4 (.A1(n_257_9_9), .A2(n_257_9_4), .A3(n_256), .ZN(n_257_9_3));
   NAND3_X1 i_257_9_5 (.A1(n_257_9_7), .A2(n_257_9_5), .A3(n_255), .ZN(n_257_9_4));
   NAND2_X1 i_257_9_6 (.A1(n_257_9_6), .A2(n_257_9_95), .ZN(n_257_9_5));
   INV_X1 i_257_9_7 (.A(CPU_Bus[7]), .ZN(n_257_9_6));
   NAND2_X1 i_257_9_8 (.A1(n_257_9_8), .A2(n_254), .ZN(n_257_9_7));
   INV_X1 i_257_9_9 (.A(CPU_Bus[8]), .ZN(n_257_9_8));
   NAND3_X1 i_257_9_10 (.A1(n_257_9_12), .A2(n_257_9_10), .A3(n_257_9_96), 
      .ZN(n_257_9_9));
   NAND2_X1 i_257_9_11 (.A1(n_257_9_11), .A2(n_254), .ZN(n_257_9_10));
   INV_X1 i_257_9_12 (.A(CPU_Bus[6]), .ZN(n_257_9_11));
   NAND2_X1 i_257_9_13 (.A1(n_257_9_13), .A2(n_257_9_95), .ZN(n_257_9_12));
   INV_X1 i_257_9_14 (.A(CPU_Bus[5]), .ZN(n_257_9_13));
   NAND3_X1 i_257_9_15 (.A1(n_257_9_20), .A2(n_257_9_15), .A3(n_257_9_97), 
      .ZN(n_257_9_14));
   NAND3_X1 i_257_9_16 (.A1(n_257_9_18), .A2(n_257_9_16), .A3(n_257_9_96), 
      .ZN(n_257_9_15));
   NAND2_X1 i_257_9_17 (.A1(n_257_9_17), .A2(n_257_9_95), .ZN(n_257_9_16));
   INV_X1 i_257_9_18 (.A(CPU_Bus[1]), .ZN(n_257_9_17));
   NAND2_X1 i_257_9_19 (.A1(n_257_9_19), .A2(n_254), .ZN(n_257_9_18));
   INV_X1 i_257_9_20 (.A(CPU_Bus[2]), .ZN(n_257_9_19));
   NAND3_X1 i_257_9_21 (.A1(n_257_9_23), .A2(n_257_9_21), .A3(n_255), .ZN(
      n_257_9_20));
   NAND2_X1 i_257_9_22 (.A1(n_257_9_22), .A2(n_254), .ZN(n_257_9_21));
   INV_X1 i_257_9_23 (.A(CPU_Bus[4]), .ZN(n_257_9_22));
   NAND2_X1 i_257_9_24 (.A1(n_257_9_24), .A2(n_257_9_95), .ZN(n_257_9_23));
   INV_X1 i_257_9_25 (.A(CPU_Bus[3]), .ZN(n_257_9_24));
   NAND3_X1 i_257_9_26 (.A1(n_257_9_37), .A2(n_257_9_26), .A3(n_257_9_98), 
      .ZN(n_257_9_25));
   NAND3_X1 i_257_9_27 (.A1(n_257_9_32), .A2(n_257_9_27), .A3(n_256), .ZN(
      n_257_9_26));
   NAND3_X1 i_257_9_28 (.A1(n_257_9_30), .A2(n_257_9_28), .A3(n_255), .ZN(
      n_257_9_27));
   NAND2_X1 i_257_9_29 (.A1(n_257_9_29), .A2(n_257_9_95), .ZN(n_257_9_28));
   INV_X1 i_257_9_30 (.A(CPU_Bus[31]), .ZN(n_257_9_29));
   NAND2_X1 i_257_9_31 (.A1(n_257_9_31), .A2(n_254), .ZN(n_257_9_30));
   INV_X1 i_257_9_32 (.A(CPU_Bus[0]), .ZN(n_257_9_31));
   NAND3_X1 i_257_9_33 (.A1(n_257_9_35), .A2(n_257_9_33), .A3(n_257_9_96), 
      .ZN(n_257_9_32));
   NAND2_X1 i_257_9_34 (.A1(n_257_9_34), .A2(n_254), .ZN(n_257_9_33));
   INV_X1 i_257_9_35 (.A(CPU_Bus[30]), .ZN(n_257_9_34));
   NAND2_X1 i_257_9_36 (.A1(n_257_9_36), .A2(n_257_9_95), .ZN(n_257_9_35));
   INV_X1 i_257_9_37 (.A(CPU_Bus[29]), .ZN(n_257_9_36));
   NAND3_X1 i_257_9_38 (.A1(n_257_9_43), .A2(n_257_9_38), .A3(n_257_9_97), 
      .ZN(n_257_9_37));
   NAND3_X1 i_257_9_39 (.A1(n_257_9_41), .A2(n_257_9_39), .A3(n_257_9_96), 
      .ZN(n_257_9_38));
   NAND2_X1 i_257_9_40 (.A1(n_257_9_40), .A2(n_257_9_95), .ZN(n_257_9_39));
   INV_X1 i_257_9_41 (.A(CPU_Bus[25]), .ZN(n_257_9_40));
   NAND2_X1 i_257_9_42 (.A1(n_257_9_42), .A2(n_254), .ZN(n_257_9_41));
   INV_X1 i_257_9_43 (.A(CPU_Bus[26]), .ZN(n_257_9_42));
   NAND3_X1 i_257_9_44 (.A1(n_257_9_46), .A2(n_257_9_44), .A3(n_255), .ZN(
      n_257_9_43));
   NAND2_X1 i_257_9_45 (.A1(n_257_9_45), .A2(n_254), .ZN(n_257_9_44));
   INV_X1 i_257_9_46 (.A(CPU_Bus[28]), .ZN(n_257_9_45));
   NAND2_X1 i_257_9_47 (.A1(n_257_9_47), .A2(n_257_9_95), .ZN(n_257_9_46));
   INV_X1 i_257_9_48 (.A(CPU_Bus[27]), .ZN(n_257_9_47));
   INV_X1 i_257_9_49 (.A(n_258), .ZN(n_257_9_48));
   NAND2_X1 i_257_9_50 (.A1(n_257_9_50), .A2(n_258), .ZN(n_257_9_49));
   NAND2_X1 i_257_9_51 (.A1(n_257_9_74), .A2(n_257_9_51), .ZN(n_257_9_50));
   NAND3_X1 i_257_9_52 (.A1(n_257_9_63), .A2(n_257_9_52), .A3(n_257), .ZN(
      n_257_9_51));
   NAND3_X1 i_257_9_53 (.A1(n_257_9_58), .A2(n_257_9_53), .A3(n_256), .ZN(
      n_257_9_52));
   NAND3_X1 i_257_9_54 (.A1(n_257_9_56), .A2(n_257_9_54), .A3(n_257_9_96), 
      .ZN(n_257_9_53));
   NAND2_X1 i_257_9_55 (.A1(n_257_9_55), .A2(n_254), .ZN(n_257_9_54));
   INV_X1 i_257_9_56 (.A(CPU_Bus[22]), .ZN(n_257_9_55));
   NAND2_X1 i_257_9_57 (.A1(n_257_9_57), .A2(n_257_9_95), .ZN(n_257_9_56));
   INV_X1 i_257_9_58 (.A(CPU_Bus[21]), .ZN(n_257_9_57));
   NAND3_X1 i_257_9_59 (.A1(n_257_9_61), .A2(n_257_9_59), .A3(n_255), .ZN(
      n_257_9_58));
   NAND2_X1 i_257_9_60 (.A1(n_257_9_60), .A2(n_254), .ZN(n_257_9_59));
   INV_X1 i_257_9_61 (.A(CPU_Bus[24]), .ZN(n_257_9_60));
   NAND2_X1 i_257_9_62 (.A1(n_257_9_62), .A2(n_257_9_95), .ZN(n_257_9_61));
   INV_X1 i_257_9_63 (.A(CPU_Bus[23]), .ZN(n_257_9_62));
   NAND3_X1 i_257_9_64 (.A1(n_257_9_69), .A2(n_257_9_64), .A3(n_257_9_97), 
      .ZN(n_257_9_63));
   NAND3_X1 i_257_9_65 (.A1(n_257_9_67), .A2(n_257_9_65), .A3(n_255), .ZN(
      n_257_9_64));
   NAND2_X1 i_257_9_66 (.A1(n_257_9_66), .A2(n_254), .ZN(n_257_9_65));
   INV_X1 i_257_9_67 (.A(CPU_Bus[20]), .ZN(n_257_9_66));
   NAND2_X1 i_257_9_68 (.A1(n_257_9_68), .A2(n_257_9_95), .ZN(n_257_9_67));
   INV_X1 i_257_9_69 (.A(CPU_Bus[19]), .ZN(n_257_9_68));
   NAND3_X1 i_257_9_70 (.A1(n_257_9_72), .A2(n_257_9_70), .A3(n_257_9_96), 
      .ZN(n_257_9_69));
   NAND2_X1 i_257_9_71 (.A1(n_257_9_71), .A2(n_254), .ZN(n_257_9_70));
   INV_X1 i_257_9_72 (.A(CPU_Bus[18]), .ZN(n_257_9_71));
   NAND2_X1 i_257_9_73 (.A1(n_257_9_73), .A2(n_257_9_95), .ZN(n_257_9_72));
   INV_X1 i_257_9_74 (.A(CPU_Bus[17]), .ZN(n_257_9_73));
   NAND3_X1 i_257_9_75 (.A1(n_257_9_86), .A2(n_257_9_98), .A3(n_257_9_75), 
      .ZN(n_257_9_74));
   NAND3_X1 i_257_9_76 (.A1(n_257_9_81), .A2(n_257_9_76), .A3(n_256), .ZN(
      n_257_9_75));
   NAND3_X1 i_257_9_77 (.A1(n_257_9_79), .A2(n_257_9_77), .A3(n_257_9_96), 
      .ZN(n_257_9_76));
   NAND2_X1 i_257_9_78 (.A1(n_257_9_78), .A2(n_254), .ZN(n_257_9_77));
   INV_X1 i_257_9_79 (.A(CPU_Bus[14]), .ZN(n_257_9_78));
   NAND2_X1 i_257_9_80 (.A1(n_257_9_80), .A2(n_257_9_95), .ZN(n_257_9_79));
   INV_X1 i_257_9_81 (.A(CPU_Bus[13]), .ZN(n_257_9_80));
   NAND3_X1 i_257_9_82 (.A1(n_257_9_84), .A2(n_257_9_82), .A3(n_255), .ZN(
      n_257_9_81));
   NAND2_X1 i_257_9_83 (.A1(n_257_9_83), .A2(n_254), .ZN(n_257_9_82));
   INV_X1 i_257_9_84 (.A(CPU_Bus[16]), .ZN(n_257_9_83));
   NAND2_X1 i_257_9_85 (.A1(n_257_9_85), .A2(n_257_9_95), .ZN(n_257_9_84));
   INV_X1 i_257_9_86 (.A(CPU_Bus[15]), .ZN(n_257_9_85));
   NAND3_X1 i_257_9_87 (.A1(n_257_9_92), .A2(n_257_9_97), .A3(n_257_9_87), 
      .ZN(n_257_9_86));
   NAND3_X1 i_257_9_88 (.A1(n_257_9_90), .A2(n_257_9_88), .A3(n_255), .ZN(
      n_257_9_87));
   NAND2_X1 i_257_9_89 (.A1(n_257_9_89), .A2(n_254), .ZN(n_257_9_88));
   INV_X1 i_257_9_90 (.A(CPU_Bus[12]), .ZN(n_257_9_89));
   NAND2_X1 i_257_9_91 (.A1(n_257_9_91), .A2(n_257_9_95), .ZN(n_257_9_90));
   INV_X1 i_257_9_92 (.A(CPU_Bus[11]), .ZN(n_257_9_91));
   OAI211_X1 i_257_9_93 (.A(n_257_9_93), .B(n_257_9_96), .C1(n_257_9_95), 
      .C2(CPU_Bus[10]), .ZN(n_257_9_92));
   NAND2_X1 i_257_9_94 (.A1(n_257_9_94), .A2(n_257_9_95), .ZN(n_257_9_93));
   INV_X1 i_257_9_95 (.A(CPU_Bus[9]), .ZN(n_257_9_94));
   INV_X1 i_257_9_96 (.A(n_254), .ZN(n_257_9_95));
   INV_X1 i_257_9_97 (.A(n_255), .ZN(n_257_9_96));
   INV_X1 i_257_9_98 (.A(n_256), .ZN(n_257_9_97));
   INV_X1 i_257_9_99 (.A(n_257), .ZN(n_257_9_98));
   NAND2_X1 i_257_10_0 (.A1(n_257_10_49), .A2(n_257_10_0), .ZN(n_257_20));
   NAND2_X1 i_257_10_1 (.A1(n_257_10_1), .A2(n_257_10_48), .ZN(n_257_10_0));
   NAND2_X1 i_257_10_2 (.A1(n_257_10_25), .A2(n_257_10_2), .ZN(n_257_10_1));
   NAND3_X1 i_257_10_3 (.A1(n_257_10_14), .A2(n_257_10_3), .A3(n_257), .ZN(
      n_257_10_2));
   NAND3_X1 i_257_10_4 (.A1(n_257_10_9), .A2(n_257_10_4), .A3(n_256), .ZN(
      n_257_10_3));
   NAND3_X1 i_257_10_5 (.A1(n_257_10_7), .A2(n_257_10_5), .A3(n_255), .ZN(
      n_257_10_4));
   NAND2_X1 i_257_10_6 (.A1(n_257_10_6), .A2(n_257_10_95), .ZN(n_257_10_5));
   INV_X1 i_257_10_7 (.A(CPU_Bus[6]), .ZN(n_257_10_6));
   NAND2_X1 i_257_10_8 (.A1(n_257_10_8), .A2(n_254), .ZN(n_257_10_7));
   INV_X1 i_257_10_9 (.A(CPU_Bus[7]), .ZN(n_257_10_8));
   NAND3_X1 i_257_10_10 (.A1(n_257_10_12), .A2(n_257_10_10), .A3(n_257_10_96), 
      .ZN(n_257_10_9));
   NAND2_X1 i_257_10_11 (.A1(n_257_10_11), .A2(n_254), .ZN(n_257_10_10));
   INV_X1 i_257_10_12 (.A(CPU_Bus[5]), .ZN(n_257_10_11));
   NAND2_X1 i_257_10_13 (.A1(n_257_10_13), .A2(n_257_10_95), .ZN(n_257_10_12));
   INV_X1 i_257_10_14 (.A(CPU_Bus[4]), .ZN(n_257_10_13));
   NAND3_X1 i_257_10_15 (.A1(n_257_10_20), .A2(n_257_10_15), .A3(n_257_10_97), 
      .ZN(n_257_10_14));
   NAND3_X1 i_257_10_16 (.A1(n_257_10_18), .A2(n_257_10_16), .A3(n_257_10_96), 
      .ZN(n_257_10_15));
   NAND2_X1 i_257_10_17 (.A1(n_257_10_17), .A2(n_257_10_95), .ZN(n_257_10_16));
   INV_X1 i_257_10_18 (.A(CPU_Bus[0]), .ZN(n_257_10_17));
   NAND2_X1 i_257_10_19 (.A1(n_257_10_19), .A2(n_254), .ZN(n_257_10_18));
   INV_X1 i_257_10_20 (.A(CPU_Bus[1]), .ZN(n_257_10_19));
   NAND3_X1 i_257_10_21 (.A1(n_257_10_23), .A2(n_257_10_21), .A3(n_255), 
      .ZN(n_257_10_20));
   NAND2_X1 i_257_10_22 (.A1(n_257_10_22), .A2(n_254), .ZN(n_257_10_21));
   INV_X1 i_257_10_23 (.A(CPU_Bus[3]), .ZN(n_257_10_22));
   NAND2_X1 i_257_10_24 (.A1(n_257_10_24), .A2(n_257_10_95), .ZN(n_257_10_23));
   INV_X1 i_257_10_25 (.A(CPU_Bus[2]), .ZN(n_257_10_24));
   NAND3_X1 i_257_10_26 (.A1(n_257_10_37), .A2(n_257_10_26), .A3(n_257_10_98), 
      .ZN(n_257_10_25));
   NAND3_X1 i_257_10_27 (.A1(n_257_10_32), .A2(n_257_10_27), .A3(n_256), 
      .ZN(n_257_10_26));
   NAND3_X1 i_257_10_28 (.A1(n_257_10_30), .A2(n_257_10_28), .A3(n_255), 
      .ZN(n_257_10_27));
   NAND2_X1 i_257_10_29 (.A1(n_257_10_29), .A2(n_257_10_95), .ZN(n_257_10_28));
   INV_X1 i_257_10_30 (.A(CPU_Bus[30]), .ZN(n_257_10_29));
   NAND2_X1 i_257_10_31 (.A1(n_257_10_31), .A2(n_254), .ZN(n_257_10_30));
   INV_X1 i_257_10_32 (.A(CPU_Bus[31]), .ZN(n_257_10_31));
   NAND3_X1 i_257_10_33 (.A1(n_257_10_35), .A2(n_257_10_33), .A3(n_257_10_96), 
      .ZN(n_257_10_32));
   NAND2_X1 i_257_10_34 (.A1(n_257_10_34), .A2(n_254), .ZN(n_257_10_33));
   INV_X1 i_257_10_35 (.A(CPU_Bus[29]), .ZN(n_257_10_34));
   NAND2_X1 i_257_10_36 (.A1(n_257_10_36), .A2(n_257_10_95), .ZN(n_257_10_35));
   INV_X1 i_257_10_37 (.A(CPU_Bus[28]), .ZN(n_257_10_36));
   NAND3_X1 i_257_10_38 (.A1(n_257_10_43), .A2(n_257_10_38), .A3(n_257_10_97), 
      .ZN(n_257_10_37));
   NAND3_X1 i_257_10_39 (.A1(n_257_10_41), .A2(n_257_10_39), .A3(n_257_10_96), 
      .ZN(n_257_10_38));
   NAND2_X1 i_257_10_40 (.A1(n_257_10_40), .A2(n_257_10_95), .ZN(n_257_10_39));
   INV_X1 i_257_10_41 (.A(CPU_Bus[24]), .ZN(n_257_10_40));
   NAND2_X1 i_257_10_42 (.A1(n_257_10_42), .A2(n_254), .ZN(n_257_10_41));
   INV_X1 i_257_10_43 (.A(CPU_Bus[25]), .ZN(n_257_10_42));
   NAND3_X1 i_257_10_44 (.A1(n_257_10_46), .A2(n_257_10_44), .A3(n_255), 
      .ZN(n_257_10_43));
   NAND2_X1 i_257_10_45 (.A1(n_257_10_45), .A2(n_254), .ZN(n_257_10_44));
   INV_X1 i_257_10_46 (.A(CPU_Bus[27]), .ZN(n_257_10_45));
   NAND2_X1 i_257_10_47 (.A1(n_257_10_47), .A2(n_257_10_95), .ZN(n_257_10_46));
   INV_X1 i_257_10_48 (.A(CPU_Bus[26]), .ZN(n_257_10_47));
   INV_X1 i_257_10_49 (.A(n_258), .ZN(n_257_10_48));
   NAND2_X1 i_257_10_50 (.A1(n_257_10_50), .A2(n_258), .ZN(n_257_10_49));
   NAND2_X1 i_257_10_51 (.A1(n_257_10_74), .A2(n_257_10_51), .ZN(n_257_10_50));
   NAND3_X1 i_257_10_52 (.A1(n_257_10_63), .A2(n_257_10_52), .A3(n_257), 
      .ZN(n_257_10_51));
   NAND3_X1 i_257_10_53 (.A1(n_257_10_58), .A2(n_257_10_53), .A3(n_256), 
      .ZN(n_257_10_52));
   NAND3_X1 i_257_10_54 (.A1(n_257_10_56), .A2(n_257_10_54), .A3(n_257_10_96), 
      .ZN(n_257_10_53));
   NAND2_X1 i_257_10_55 (.A1(n_257_10_55), .A2(n_254), .ZN(n_257_10_54));
   INV_X1 i_257_10_56 (.A(CPU_Bus[21]), .ZN(n_257_10_55));
   NAND2_X1 i_257_10_57 (.A1(n_257_10_57), .A2(n_257_10_95), .ZN(n_257_10_56));
   INV_X1 i_257_10_58 (.A(CPU_Bus[20]), .ZN(n_257_10_57));
   NAND3_X1 i_257_10_59 (.A1(n_257_10_61), .A2(n_257_10_59), .A3(n_255), 
      .ZN(n_257_10_58));
   NAND2_X1 i_257_10_60 (.A1(n_257_10_60), .A2(n_254), .ZN(n_257_10_59));
   INV_X1 i_257_10_61 (.A(CPU_Bus[23]), .ZN(n_257_10_60));
   NAND2_X1 i_257_10_62 (.A1(n_257_10_62), .A2(n_257_10_95), .ZN(n_257_10_61));
   INV_X1 i_257_10_63 (.A(CPU_Bus[22]), .ZN(n_257_10_62));
   NAND3_X1 i_257_10_64 (.A1(n_257_10_69), .A2(n_257_10_64), .A3(n_257_10_97), 
      .ZN(n_257_10_63));
   NAND3_X1 i_257_10_65 (.A1(n_257_10_67), .A2(n_257_10_65), .A3(n_255), 
      .ZN(n_257_10_64));
   NAND2_X1 i_257_10_66 (.A1(n_257_10_66), .A2(n_254), .ZN(n_257_10_65));
   INV_X1 i_257_10_67 (.A(CPU_Bus[19]), .ZN(n_257_10_66));
   NAND2_X1 i_257_10_68 (.A1(n_257_10_68), .A2(n_257_10_95), .ZN(n_257_10_67));
   INV_X1 i_257_10_69 (.A(CPU_Bus[18]), .ZN(n_257_10_68));
   NAND3_X1 i_257_10_70 (.A1(n_257_10_72), .A2(n_257_10_70), .A3(n_257_10_96), 
      .ZN(n_257_10_69));
   NAND2_X1 i_257_10_71 (.A1(n_257_10_71), .A2(n_254), .ZN(n_257_10_70));
   INV_X1 i_257_10_72 (.A(CPU_Bus[17]), .ZN(n_257_10_71));
   NAND2_X1 i_257_10_73 (.A1(n_257_10_73), .A2(n_257_10_95), .ZN(n_257_10_72));
   INV_X1 i_257_10_74 (.A(CPU_Bus[16]), .ZN(n_257_10_73));
   NAND3_X1 i_257_10_75 (.A1(n_257_10_86), .A2(n_257_10_98), .A3(n_257_10_75), 
      .ZN(n_257_10_74));
   NAND3_X1 i_257_10_76 (.A1(n_257_10_81), .A2(n_257_10_76), .A3(n_256), 
      .ZN(n_257_10_75));
   NAND3_X1 i_257_10_77 (.A1(n_257_10_79), .A2(n_257_10_77), .A3(n_257_10_96), 
      .ZN(n_257_10_76));
   NAND2_X1 i_257_10_78 (.A1(n_257_10_78), .A2(n_254), .ZN(n_257_10_77));
   INV_X1 i_257_10_79 (.A(CPU_Bus[13]), .ZN(n_257_10_78));
   NAND2_X1 i_257_10_80 (.A1(n_257_10_80), .A2(n_257_10_95), .ZN(n_257_10_79));
   INV_X1 i_257_10_81 (.A(CPU_Bus[12]), .ZN(n_257_10_80));
   NAND3_X1 i_257_10_82 (.A1(n_257_10_84), .A2(n_257_10_82), .A3(n_255), 
      .ZN(n_257_10_81));
   NAND2_X1 i_257_10_83 (.A1(n_257_10_83), .A2(n_254), .ZN(n_257_10_82));
   INV_X1 i_257_10_84 (.A(CPU_Bus[15]), .ZN(n_257_10_83));
   NAND2_X1 i_257_10_85 (.A1(n_257_10_85), .A2(n_257_10_95), .ZN(n_257_10_84));
   INV_X1 i_257_10_86 (.A(CPU_Bus[14]), .ZN(n_257_10_85));
   NAND3_X1 i_257_10_87 (.A1(n_257_10_92), .A2(n_257_10_97), .A3(n_257_10_87), 
      .ZN(n_257_10_86));
   NAND3_X1 i_257_10_88 (.A1(n_257_10_90), .A2(n_257_10_88), .A3(n_255), 
      .ZN(n_257_10_87));
   NAND2_X1 i_257_10_89 (.A1(n_257_10_89), .A2(n_254), .ZN(n_257_10_88));
   INV_X1 i_257_10_90 (.A(CPU_Bus[11]), .ZN(n_257_10_89));
   NAND2_X1 i_257_10_91 (.A1(n_257_10_91), .A2(n_257_10_95), .ZN(n_257_10_90));
   INV_X1 i_257_10_92 (.A(CPU_Bus[10]), .ZN(n_257_10_91));
   OAI211_X1 i_257_10_93 (.A(n_257_10_93), .B(n_257_10_96), .C1(n_257_10_95), 
      .C2(CPU_Bus[9]), .ZN(n_257_10_92));
   NAND2_X1 i_257_10_94 (.A1(n_257_10_94), .A2(n_257_10_95), .ZN(n_257_10_93));
   INV_X1 i_257_10_95 (.A(CPU_Bus[8]), .ZN(n_257_10_94));
   INV_X1 i_257_10_96 (.A(n_254), .ZN(n_257_10_95));
   INV_X1 i_257_10_97 (.A(n_255), .ZN(n_257_10_96));
   INV_X1 i_257_10_98 (.A(n_256), .ZN(n_257_10_97));
   INV_X1 i_257_10_99 (.A(n_257), .ZN(n_257_10_98));
   INV_X1 i_257_11_0 (.A(n_254), .ZN(n_257_11_0));
   NAND2_X1 i_257_11_1 (.A1(n_257_11_0), .A2(n_255), .ZN(n_257_11_1));
   INV_X1 i_257_11_2 (.A(n_256), .ZN(n_257_11_2));
   NOR2_X1 i_257_11_3 (.A1(n_257_11_1), .A2(n_257_11_2), .ZN(n_257_11_3));
   NAND2_X1 i_257_11_4 (.A1(n_257_11_3), .A2(n_257), .ZN(n_257_11_4));
   INV_X1 i_257_11_5 (.A(n_258), .ZN(n_257_11_5));
   NOR2_X1 i_257_11_6 (.A1(n_257_11_4), .A2(n_257_11_5), .ZN(n_257_11_6));
   NAND2_X1 i_257_11_7 (.A1(CPU_Bus[21]), .A2(n_257_11_6), .ZN(n_257_11_7));
   INV_X1 i_257_11_8 (.A(n_255), .ZN(n_257_11_8));
   NAND2_X1 i_257_11_9 (.A1(n_257_11_0), .A2(n_257_11_8), .ZN(n_257_11_9));
   NOR2_X1 i_257_11_10 (.A1(n_257_11_9), .A2(n_257_11_2), .ZN(n_257_11_10));
   NAND2_X1 i_257_11_11 (.A1(n_257_11_10), .A2(n_257), .ZN(n_257_11_11));
   NOR2_X1 i_257_11_12 (.A1(n_257_11_11), .A2(n_257_11_5), .ZN(n_257_11_12));
   NAND2_X1 i_257_11_13 (.A1(CPU_Bus[19]), .A2(n_257_11_12), .ZN(n_257_11_13));
   NAND2_X1 i_257_11_14 (.A1(n_257_11_7), .A2(n_257_11_13), .ZN(n_257_11_14));
   NOR2_X1 i_257_11_15 (.A1(n_257_11_1), .A2(n_256), .ZN(n_257_11_15));
   NAND2_X1 i_257_11_16 (.A1(n_257_11_15), .A2(n_257), .ZN(n_257_11_16));
   NOR2_X1 i_257_11_17 (.A1(n_257_11_16), .A2(n_257_11_5), .ZN(n_257_11_17));
   NAND2_X1 i_257_11_18 (.A1(CPU_Bus[17]), .A2(n_257_11_17), .ZN(n_257_11_18));
   NOR2_X1 i_257_11_19 (.A1(n_257_11_9), .A2(n_256), .ZN(n_257_11_19));
   NAND2_X1 i_257_11_20 (.A1(n_257_11_19), .A2(n_257), .ZN(n_257_11_20));
   NOR2_X1 i_257_11_21 (.A1(n_257_11_20), .A2(n_257_11_5), .ZN(n_257_11_21));
   NAND2_X1 i_257_11_22 (.A1(CPU_Bus[15]), .A2(n_257_11_21), .ZN(n_257_11_22));
   NAND2_X1 i_257_11_23 (.A1(n_257_11_18), .A2(n_257_11_22), .ZN(n_257_11_23));
   NOR2_X1 i_257_11_24 (.A1(n_257_11_14), .A2(n_257_11_23), .ZN(n_257_11_24));
   INV_X1 i_257_11_25 (.A(n_257), .ZN(n_257_11_25));
   NAND2_X1 i_257_11_26 (.A1(n_257_11_3), .A2(n_257_11_25), .ZN(n_257_11_26));
   NOR2_X1 i_257_11_27 (.A1(n_257_11_26), .A2(n_257_11_5), .ZN(n_257_11_27));
   NAND2_X1 i_257_11_28 (.A1(CPU_Bus[13]), .A2(n_257_11_27), .ZN(n_257_11_28));
   NAND2_X1 i_257_11_29 (.A1(n_257_11_10), .A2(n_257_11_25), .ZN(n_257_11_29));
   NOR2_X1 i_257_11_30 (.A1(n_257_11_29), .A2(n_257_11_5), .ZN(n_257_11_30));
   NAND2_X1 i_257_11_31 (.A1(CPU_Bus[11]), .A2(n_257_11_30), .ZN(n_257_11_31));
   NAND2_X1 i_257_11_32 (.A1(n_257_11_28), .A2(n_257_11_31), .ZN(n_257_11_32));
   NAND2_X1 i_257_11_33 (.A1(n_257_11_15), .A2(n_257_11_25), .ZN(n_257_11_33));
   NOR2_X1 i_257_11_34 (.A1(n_257_11_33), .A2(n_257_11_5), .ZN(n_257_11_34));
   NAND2_X1 i_257_11_35 (.A1(CPU_Bus[9]), .A2(n_257_11_34), .ZN(n_257_11_35));
   NAND2_X1 i_257_11_36 (.A1(n_257_11_19), .A2(n_257_11_25), .ZN(n_257_11_36));
   NOR2_X1 i_257_11_37 (.A1(n_257_11_36), .A2(n_257_11_5), .ZN(n_257_11_37));
   NAND2_X1 i_257_11_38 (.A1(CPU_Bus[7]), .A2(n_257_11_37), .ZN(n_257_11_38));
   NAND2_X1 i_257_11_39 (.A1(n_257_11_35), .A2(n_257_11_38), .ZN(n_257_11_39));
   NOR2_X1 i_257_11_40 (.A1(n_257_11_32), .A2(n_257_11_39), .ZN(n_257_11_40));
   NAND2_X1 i_257_11_41 (.A1(n_257_11_24), .A2(n_257_11_40), .ZN(n_257_11_41));
   NOR2_X1 i_257_11_42 (.A1(n_257_11_4), .A2(n_258), .ZN(n_257_11_42));
   NAND2_X1 i_257_11_43 (.A1(CPU_Bus[5]), .A2(n_257_11_42), .ZN(n_257_11_43));
   NOR2_X1 i_257_11_44 (.A1(n_257_11_11), .A2(n_258), .ZN(n_257_11_44));
   NAND2_X1 i_257_11_45 (.A1(CPU_Bus[3]), .A2(n_257_11_44), .ZN(n_257_11_45));
   NAND2_X1 i_257_11_46 (.A1(n_257_11_43), .A2(n_257_11_45), .ZN(n_257_11_46));
   NOR2_X1 i_257_11_47 (.A1(n_257_11_16), .A2(n_258), .ZN(n_257_11_47));
   NAND2_X1 i_257_11_48 (.A1(CPU_Bus[1]), .A2(n_257_11_47), .ZN(n_257_11_48));
   NOR2_X1 i_257_11_49 (.A1(n_257_11_20), .A2(n_258), .ZN(n_257_11_49));
   NAND2_X1 i_257_11_50 (.A1(CPU_Bus[31]), .A2(n_257_11_49), .ZN(n_257_11_50));
   NAND2_X1 i_257_11_51 (.A1(n_257_11_48), .A2(n_257_11_50), .ZN(n_257_11_51));
   NOR2_X1 i_257_11_52 (.A1(n_257_11_46), .A2(n_257_11_51), .ZN(n_257_11_52));
   NOR2_X1 i_257_11_53 (.A1(n_257_11_26), .A2(n_258), .ZN(n_257_11_53));
   NAND2_X1 i_257_11_54 (.A1(CPU_Bus[29]), .A2(n_257_11_53), .ZN(n_257_11_54));
   NOR2_X1 i_257_11_55 (.A1(n_257_11_29), .A2(n_258), .ZN(n_257_11_55));
   NAND2_X1 i_257_11_56 (.A1(CPU_Bus[27]), .A2(n_257_11_55), .ZN(n_257_11_56));
   NAND2_X1 i_257_11_57 (.A1(n_257_11_54), .A2(n_257_11_56), .ZN(n_257_11_57));
   NOR2_X1 i_257_11_58 (.A1(n_257_11_33), .A2(n_258), .ZN(n_257_11_58));
   NAND2_X1 i_257_11_59 (.A1(CPU_Bus[25]), .A2(n_257_11_58), .ZN(n_257_11_59));
   NOR2_X1 i_257_11_60 (.A1(n_257_11_36), .A2(n_258), .ZN(n_257_11_60));
   NAND2_X1 i_257_11_61 (.A1(CPU_Bus[23]), .A2(n_257_11_60), .ZN(n_257_11_61));
   NAND2_X1 i_257_11_62 (.A1(n_257_11_59), .A2(n_257_11_61), .ZN(n_257_11_62));
   NOR2_X1 i_257_11_63 (.A1(n_257_11_57), .A2(n_257_11_62), .ZN(n_257_11_63));
   NAND2_X1 i_257_11_64 (.A1(n_257_11_52), .A2(n_257_11_63), .ZN(n_257_11_64));
   NOR2_X1 i_257_11_65 (.A1(n_257_11_41), .A2(n_257_11_64), .ZN(n_257_11_65));
   NAND2_X1 i_257_11_66 (.A1(n_257_11_8), .A2(n_254), .ZN(n_257_11_66));
   NOR2_X1 i_257_11_67 (.A1(n_257_11_66), .A2(n_257_11_2), .ZN(n_257_11_67));
   NAND2_X1 i_257_11_68 (.A1(n_257_11_67), .A2(n_257), .ZN(n_257_11_68));
   NOR2_X1 i_257_11_69 (.A1(n_257_11_68), .A2(n_257_11_5), .ZN(n_257_11_69));
   NAND2_X1 i_257_11_70 (.A1(CPU_Bus[20]), .A2(n_257_11_69), .ZN(n_257_11_70));
   NOR2_X1 i_257_11_71 (.A1(n_257_11_66), .A2(n_256), .ZN(n_257_11_71));
   NAND2_X1 i_257_11_72 (.A1(n_257_11_71), .A2(n_257), .ZN(n_257_11_72));
   NOR2_X1 i_257_11_73 (.A1(n_257_11_72), .A2(n_257_11_5), .ZN(n_257_11_73));
   NAND2_X1 i_257_11_74 (.A1(CPU_Bus[16]), .A2(n_257_11_73), .ZN(n_257_11_74));
   NAND2_X1 i_257_11_75 (.A1(n_257_11_70), .A2(n_257_11_74), .ZN(n_257_11_75));
   NAND2_X1 i_257_11_76 (.A1(n_257_11_67), .A2(n_257_11_25), .ZN(n_257_11_76));
   NOR2_X1 i_257_11_77 (.A1(n_257_11_76), .A2(n_257_11_5), .ZN(n_257_11_77));
   NAND2_X1 i_257_11_78 (.A1(CPU_Bus[12]), .A2(n_257_11_77), .ZN(n_257_11_78));
   NAND2_X1 i_257_11_79 (.A1(n_257_11_71), .A2(n_257_11_25), .ZN(n_257_11_79));
   NOR2_X1 i_257_11_80 (.A1(n_257_11_79), .A2(n_257_11_5), .ZN(n_257_11_80));
   NAND2_X1 i_257_11_81 (.A1(CPU_Bus[8]), .A2(n_257_11_80), .ZN(n_257_11_81));
   NAND2_X1 i_257_11_82 (.A1(n_257_11_78), .A2(n_257_11_81), .ZN(n_257_11_82));
   NOR2_X1 i_257_11_83 (.A1(n_257_11_75), .A2(n_257_11_82), .ZN(n_257_11_83));
   NOR2_X1 i_257_11_84 (.A1(n_257_11_68), .A2(n_258), .ZN(n_257_11_84));
   NAND2_X1 i_257_11_85 (.A1(CPU_Bus[4]), .A2(n_257_11_84), .ZN(n_257_11_85));
   NOR2_X1 i_257_11_86 (.A1(n_257_11_72), .A2(n_258), .ZN(n_257_11_86));
   NAND2_X1 i_257_11_87 (.A1(CPU_Bus[0]), .A2(n_257_11_86), .ZN(n_257_11_87));
   NAND2_X1 i_257_11_88 (.A1(n_257_11_85), .A2(n_257_11_87), .ZN(n_257_11_88));
   NOR2_X1 i_257_11_89 (.A1(n_257_11_76), .A2(n_258), .ZN(n_257_11_89));
   NAND2_X1 i_257_11_90 (.A1(CPU_Bus[28]), .A2(n_257_11_89), .ZN(n_257_11_90));
   NOR2_X1 i_257_11_91 (.A1(n_257_11_79), .A2(n_258), .ZN(n_257_11_91));
   NAND2_X1 i_257_11_92 (.A1(CPU_Bus[24]), .A2(n_257_11_91), .ZN(n_257_11_92));
   NAND2_X1 i_257_11_93 (.A1(n_257_11_90), .A2(n_257_11_92), .ZN(n_257_11_93));
   NOR2_X1 i_257_11_94 (.A1(n_257_11_88), .A2(n_257_11_93), .ZN(n_257_11_94));
   NAND2_X1 i_257_11_95 (.A1(n_257_11_83), .A2(n_257_11_94), .ZN(n_257_11_95));
   NAND2_X1 i_257_11_96 (.A1(n_254), .A2(n_255), .ZN(n_257_11_96));
   NOR2_X1 i_257_11_97 (.A1(n_257_11_96), .A2(n_257_11_2), .ZN(n_257_11_97));
   NAND2_X1 i_257_11_98 (.A1(n_257_11_97), .A2(n_257), .ZN(n_257_11_98));
   NOR2_X1 i_257_11_99 (.A1(n_257_11_98), .A2(n_257_11_5), .ZN(n_257_11_99));
   NAND2_X1 i_257_11_100 (.A1(CPU_Bus[22]), .A2(n_257_11_99), .ZN(n_257_11_100));
   NOR2_X1 i_257_11_101 (.A1(n_257_11_96), .A2(n_256), .ZN(n_257_11_101));
   NAND2_X1 i_257_11_102 (.A1(n_257_11_101), .A2(n_257), .ZN(n_257_11_102));
   NOR2_X1 i_257_11_103 (.A1(n_257_11_102), .A2(n_257_11_5), .ZN(n_257_11_103));
   NAND2_X1 i_257_11_104 (.A1(CPU_Bus[18]), .A2(n_257_11_103), .ZN(n_257_11_104));
   NAND2_X1 i_257_11_105 (.A1(n_257_11_100), .A2(n_257_11_104), .ZN(n_257_11_105));
   NAND2_X1 i_257_11_106 (.A1(n_257_11_97), .A2(n_257_11_25), .ZN(n_257_11_106));
   NOR2_X1 i_257_11_107 (.A1(n_257_11_106), .A2(n_257_11_5), .ZN(n_257_11_107));
   NAND2_X1 i_257_11_108 (.A1(CPU_Bus[14]), .A2(n_257_11_107), .ZN(n_257_11_108));
   NAND2_X1 i_257_11_109 (.A1(n_257_11_101), .A2(n_257_11_25), .ZN(n_257_11_109));
   NOR2_X1 i_257_11_110 (.A1(n_257_11_109), .A2(n_257_11_5), .ZN(n_257_11_110));
   NAND2_X1 i_257_11_111 (.A1(CPU_Bus[10]), .A2(n_257_11_110), .ZN(n_257_11_111));
   NAND2_X1 i_257_11_112 (.A1(n_257_11_108), .A2(n_257_11_111), .ZN(n_257_11_112));
   NOR2_X1 i_257_11_113 (.A1(n_257_11_105), .A2(n_257_11_112), .ZN(n_257_11_113));
   NOR2_X1 i_257_11_114 (.A1(n_257_11_98), .A2(n_258), .ZN(n_257_11_114));
   NAND2_X1 i_257_11_115 (.A1(CPU_Bus[6]), .A2(n_257_11_114), .ZN(n_257_11_115));
   NOR2_X1 i_257_11_116 (.A1(n_257_11_102), .A2(n_258), .ZN(n_257_11_116));
   NAND2_X1 i_257_11_117 (.A1(CPU_Bus[2]), .A2(n_257_11_116), .ZN(n_257_11_117));
   NAND2_X1 i_257_11_118 (.A1(n_257_11_115), .A2(n_257_11_117), .ZN(n_257_11_118));
   NOR2_X1 i_257_11_119 (.A1(n_257_11_106), .A2(n_258), .ZN(n_257_11_119));
   NAND2_X1 i_257_11_120 (.A1(CPU_Bus[30]), .A2(n_257_11_119), .ZN(n_257_11_120));
   NOR2_X1 i_257_11_121 (.A1(n_257_11_109), .A2(n_258), .ZN(n_257_11_121));
   NAND2_X1 i_257_11_122 (.A1(CPU_Bus[26]), .A2(n_257_11_121), .ZN(n_257_11_122));
   NAND2_X1 i_257_11_123 (.A1(n_257_11_120), .A2(n_257_11_122), .ZN(n_257_11_123));
   NOR2_X1 i_257_11_124 (.A1(n_257_11_118), .A2(n_257_11_123), .ZN(n_257_11_124));
   NAND2_X1 i_257_11_125 (.A1(n_257_11_113), .A2(n_257_11_124), .ZN(n_257_11_125));
   NOR2_X1 i_257_11_126 (.A1(n_257_11_95), .A2(n_257_11_125), .ZN(n_257_11_126));
   NAND2_X1 i_257_11_127 (.A1(n_257_11_65), .A2(n_257_11_126), .ZN(n_257_21));
   INV_X1 i_257_12_0 (.A(n_257_12_0), .ZN(n_257_22));
   NAND2_X1 i_257_12_1 (.A1(n_257_12_49), .A2(n_257_12_1), .ZN(n_257_12_0));
   NAND3_X1 i_257_12_2 (.A1(n_257_12_25), .A2(n_257_12_2), .A3(n_257_12_48), 
      .ZN(n_257_12_1));
   NAND3_X1 i_257_12_3 (.A1(n_257_12_14), .A2(n_257_12_3), .A3(n_257), .ZN(
      n_257_12_2));
   NAND3_X1 i_257_12_4 (.A1(n_257_12_9), .A2(n_257_12_4), .A3(n_257_12_85), 
      .ZN(n_257_12_3));
   NAND3_X1 i_257_12_5 (.A1(n_257_12_7), .A2(n_257_12_5), .A3(n_257_12_96), 
      .ZN(n_257_12_4));
   NAND2_X1 i_257_12_6 (.A1(n_257_12_6), .A2(n_257_12_95), .ZN(n_257_12_5));
   INV_X1 i_257_12_7 (.A(CPU_Bus[30]), .ZN(n_257_12_6));
   NAND2_X1 i_257_12_8 (.A1(n_257_12_8), .A2(n_254), .ZN(n_257_12_7));
   INV_X1 i_257_12_9 (.A(CPU_Bus[31]), .ZN(n_257_12_8));
   NAND3_X1 i_257_12_10 (.A1(n_257_12_12), .A2(n_257_12_10), .A3(n_255), 
      .ZN(n_257_12_9));
   NAND2_X1 i_257_12_11 (.A1(n_257_12_11), .A2(n_257_12_95), .ZN(n_257_12_10));
   INV_X1 i_257_12_12 (.A(CPU_Bus[0]), .ZN(n_257_12_11));
   NAND2_X1 i_257_12_13 (.A1(n_257_12_13), .A2(n_254), .ZN(n_257_12_12));
   INV_X1 i_257_12_14 (.A(CPU_Bus[1]), .ZN(n_257_12_13));
   NAND3_X1 i_257_12_15 (.A1(n_257_12_20), .A2(n_257_12_15), .A3(n_256), 
      .ZN(n_257_12_14));
   NAND3_X1 i_257_12_16 (.A1(n_257_12_18), .A2(n_257_12_16), .A3(n_257_12_96), 
      .ZN(n_257_12_15));
   NAND2_X1 i_257_12_17 (.A1(n_257_12_17), .A2(n_257_12_95), .ZN(n_257_12_16));
   INV_X1 i_257_12_18 (.A(CPU_Bus[2]), .ZN(n_257_12_17));
   NAND2_X1 i_257_12_19 (.A1(n_257_12_19), .A2(n_254), .ZN(n_257_12_18));
   INV_X1 i_257_12_20 (.A(CPU_Bus[3]), .ZN(n_257_12_19));
   NAND3_X1 i_257_12_21 (.A1(n_257_12_23), .A2(n_257_12_21), .A3(n_255), 
      .ZN(n_257_12_20));
   NAND2_X1 i_257_12_22 (.A1(n_257_12_22), .A2(n_257_12_95), .ZN(n_257_12_21));
   INV_X1 i_257_12_23 (.A(CPU_Bus[4]), .ZN(n_257_12_22));
   NAND2_X1 i_257_12_24 (.A1(n_257_12_24), .A2(n_254), .ZN(n_257_12_23));
   INV_X1 i_257_12_25 (.A(CPU_Bus[5]), .ZN(n_257_12_24));
   NAND3_X1 i_257_12_26 (.A1(n_257_12_37), .A2(n_257_12_26), .A3(n_257_12_97), 
      .ZN(n_257_12_25));
   NAND3_X1 i_257_12_27 (.A1(n_257_12_32), .A2(n_257_12_27), .A3(n_256), 
      .ZN(n_257_12_26));
   NAND3_X1 i_257_12_28 (.A1(n_257_12_30), .A2(n_257_12_28), .A3(n_255), 
      .ZN(n_257_12_27));
   NAND2_X1 i_257_12_29 (.A1(n_257_12_29), .A2(n_254), .ZN(n_257_12_28));
   INV_X1 i_257_12_30 (.A(CPU_Bus[29]), .ZN(n_257_12_29));
   NAND2_X1 i_257_12_31 (.A1(n_257_12_31), .A2(n_257_12_95), .ZN(n_257_12_30));
   INV_X1 i_257_12_32 (.A(CPU_Bus[28]), .ZN(n_257_12_31));
   NAND3_X1 i_257_12_33 (.A1(n_257_12_35), .A2(n_257_12_33), .A3(n_257_12_96), 
      .ZN(n_257_12_32));
   NAND2_X1 i_257_12_34 (.A1(n_257_12_34), .A2(n_257_12_95), .ZN(n_257_12_33));
   INV_X1 i_257_12_35 (.A(CPU_Bus[26]), .ZN(n_257_12_34));
   NAND2_X1 i_257_12_36 (.A1(n_257_12_36), .A2(n_254), .ZN(n_257_12_35));
   INV_X1 i_257_12_37 (.A(CPU_Bus[27]), .ZN(n_257_12_36));
   NAND3_X1 i_257_12_38 (.A1(n_257_12_43), .A2(n_257_12_38), .A3(n_257_12_85), 
      .ZN(n_257_12_37));
   NAND3_X1 i_257_12_39 (.A1(n_257_12_41), .A2(n_257_12_39), .A3(n_255), 
      .ZN(n_257_12_38));
   NAND2_X1 i_257_12_40 (.A1(n_257_12_40), .A2(n_254), .ZN(n_257_12_39));
   INV_X1 i_257_12_41 (.A(CPU_Bus[25]), .ZN(n_257_12_40));
   NAND2_X1 i_257_12_42 (.A1(n_257_12_42), .A2(n_257_12_95), .ZN(n_257_12_41));
   INV_X1 i_257_12_43 (.A(CPU_Bus[24]), .ZN(n_257_12_42));
   NAND3_X1 i_257_12_44 (.A1(n_257_12_46), .A2(n_257_12_44), .A3(n_257_12_96), 
      .ZN(n_257_12_43));
   NAND2_X1 i_257_12_45 (.A1(n_257_12_45), .A2(n_257_12_95), .ZN(n_257_12_44));
   INV_X1 i_257_12_46 (.A(CPU_Bus[22]), .ZN(n_257_12_45));
   NAND2_X1 i_257_12_47 (.A1(n_257_12_47), .A2(n_254), .ZN(n_257_12_46));
   INV_X1 i_257_12_48 (.A(CPU_Bus[23]), .ZN(n_257_12_47));
   INV_X1 i_257_12_49 (.A(n_258), .ZN(n_257_12_48));
   NAND3_X1 i_257_12_50 (.A1(n_257_12_73), .A2(n_257_12_50), .A3(n_258), 
      .ZN(n_257_12_49));
   NAND3_X1 i_257_12_51 (.A1(n_257_12_62), .A2(n_257_12_51), .A3(n_257), 
      .ZN(n_257_12_50));
   NAND3_X1 i_257_12_52 (.A1(n_257_12_57), .A2(n_257_12_52), .A3(n_257_12_85), 
      .ZN(n_257_12_51));
   NAND3_X1 i_257_12_53 (.A1(n_257_12_55), .A2(n_257_12_53), .A3(n_257_12_96), 
      .ZN(n_257_12_52));
   NAND2_X1 i_257_12_54 (.A1(n_257_12_54), .A2(n_257_12_95), .ZN(n_257_12_53));
   INV_X1 i_257_12_55 (.A(CPU_Bus[14]), .ZN(n_257_12_54));
   NAND2_X1 i_257_12_56 (.A1(n_257_12_56), .A2(n_254), .ZN(n_257_12_55));
   INV_X1 i_257_12_57 (.A(CPU_Bus[15]), .ZN(n_257_12_56));
   NAND3_X1 i_257_12_58 (.A1(n_257_12_60), .A2(n_257_12_58), .A3(n_255), 
      .ZN(n_257_12_57));
   NAND2_X1 i_257_12_59 (.A1(n_257_12_59), .A2(n_254), .ZN(n_257_12_58));
   INV_X1 i_257_12_60 (.A(CPU_Bus[17]), .ZN(n_257_12_59));
   NAND2_X1 i_257_12_61 (.A1(n_257_12_61), .A2(n_257_12_95), .ZN(n_257_12_60));
   INV_X1 i_257_12_62 (.A(CPU_Bus[16]), .ZN(n_257_12_61));
   NAND3_X1 i_257_12_63 (.A1(n_257_12_68), .A2(n_257_12_63), .A3(n_256), 
      .ZN(n_257_12_62));
   NAND3_X1 i_257_12_64 (.A1(n_257_12_66), .A2(n_257_12_64), .A3(n_257_12_96), 
      .ZN(n_257_12_63));
   NAND2_X1 i_257_12_65 (.A1(n_257_12_65), .A2(n_254), .ZN(n_257_12_64));
   INV_X1 i_257_12_66 (.A(CPU_Bus[19]), .ZN(n_257_12_65));
   NAND2_X1 i_257_12_67 (.A1(n_257_12_67), .A2(n_257_12_95), .ZN(n_257_12_66));
   INV_X1 i_257_12_68 (.A(CPU_Bus[18]), .ZN(n_257_12_67));
   NAND3_X1 i_257_12_69 (.A1(n_257_12_71), .A2(n_257_12_69), .A3(n_255), 
      .ZN(n_257_12_68));
   NAND2_X1 i_257_12_70 (.A1(n_257_12_70), .A2(n_257_12_95), .ZN(n_257_12_69));
   INV_X1 i_257_12_71 (.A(CPU_Bus[20]), .ZN(n_257_12_70));
   NAND2_X1 i_257_12_72 (.A1(n_257_12_72), .A2(n_254), .ZN(n_257_12_71));
   INV_X1 i_257_12_73 (.A(CPU_Bus[21]), .ZN(n_257_12_72));
   NAND3_X1 i_257_12_74 (.A1(n_257_12_86), .A2(n_257_12_74), .A3(n_257_12_97), 
      .ZN(n_257_12_73));
   NAND3_X1 i_257_12_75 (.A1(n_257_12_80), .A2(n_257_12_75), .A3(n_257_12_85), 
      .ZN(n_257_12_74));
   NAND3_X1 i_257_12_76 (.A1(n_257_12_78), .A2(n_257_12_76), .A3(n_257_12_96), 
      .ZN(n_257_12_75));
   NAND2_X1 i_257_12_77 (.A1(n_257_12_77), .A2(n_254), .ZN(n_257_12_76));
   INV_X1 i_257_12_78 (.A(CPU_Bus[7]), .ZN(n_257_12_77));
   NAND2_X1 i_257_12_79 (.A1(n_257_12_79), .A2(n_257_12_95), .ZN(n_257_12_78));
   INV_X1 i_257_12_80 (.A(CPU_Bus[6]), .ZN(n_257_12_79));
   NAND3_X1 i_257_12_81 (.A1(n_257_12_83), .A2(n_257_12_81), .A3(n_255), 
      .ZN(n_257_12_80));
   NAND2_X1 i_257_12_82 (.A1(n_257_12_82), .A2(n_254), .ZN(n_257_12_81));
   INV_X1 i_257_12_83 (.A(CPU_Bus[9]), .ZN(n_257_12_82));
   NAND2_X1 i_257_12_84 (.A1(n_257_12_84), .A2(n_257_12_95), .ZN(n_257_12_83));
   INV_X1 i_257_12_85 (.A(CPU_Bus[8]), .ZN(n_257_12_84));
   INV_X1 i_257_12_86 (.A(n_256), .ZN(n_257_12_85));
   NAND3_X1 i_257_12_87 (.A1(n_257_12_92), .A2(n_257_12_87), .A3(n_256), 
      .ZN(n_257_12_86));
   NAND3_X1 i_257_12_88 (.A1(n_257_12_90), .A2(n_257_12_88), .A3(n_255), 
      .ZN(n_257_12_87));
   NAND2_X1 i_257_12_89 (.A1(n_257_12_89), .A2(n_257_12_95), .ZN(n_257_12_88));
   INV_X1 i_257_12_90 (.A(CPU_Bus[12]), .ZN(n_257_12_89));
   NAND2_X1 i_257_12_91 (.A1(n_257_12_91), .A2(n_254), .ZN(n_257_12_90));
   INV_X1 i_257_12_92 (.A(CPU_Bus[13]), .ZN(n_257_12_91));
   OAI211_X1 i_257_12_93 (.A(n_257_12_93), .B(n_257_12_96), .C1(n_257_12_95), 
      .C2(CPU_Bus[11]), .ZN(n_257_12_92));
   NAND2_X1 i_257_12_94 (.A1(n_257_12_94), .A2(n_257_12_95), .ZN(n_257_12_93));
   INV_X1 i_257_12_95 (.A(CPU_Bus[10]), .ZN(n_257_12_94));
   INV_X1 i_257_12_96 (.A(n_254), .ZN(n_257_12_95));
   INV_X1 i_257_12_97 (.A(n_255), .ZN(n_257_12_96));
   INV_X1 i_257_12_98 (.A(n_257), .ZN(n_257_12_97));
   NAND2_X1 i_257_13_0 (.A1(n_257_13_0), .A2(n_257_13_36), .ZN(n_257_23));
   NAND2_X1 i_257_13_1 (.A1(n_257_13_1), .A2(n_258), .ZN(n_257_13_0));
   NAND2_X1 i_257_13_2 (.A1(n_257_13_19), .A2(n_257_13_2), .ZN(n_257_13_1));
   NAND3_X1 i_257_13_3 (.A1(n_257_13_11), .A2(n_257_13_3), .A3(n_257_13_87), 
      .ZN(n_257_13_2));
   NAND2_X1 i_257_13_4 (.A1(n_257_13_4), .A2(n_257_13_86), .ZN(n_257_13_3));
   NAND2_X1 i_257_13_5 (.A1(n_257_13_8), .A2(n_257_13_5), .ZN(n_257_13_4));
   NAND3_X1 i_257_13_6 (.A1(n_257_13_7), .A2(n_257_13_6), .A3(n_255), .ZN(
      n_257_13_5));
   NAND2_X1 i_257_13_7 (.A1(CPU_Bus[7]), .A2(n_257_13_82), .ZN(n_257_13_6));
   NAND2_X1 i_257_13_8 (.A1(CPU_Bus[8]), .A2(n_254), .ZN(n_257_13_7));
   NAND3_X1 i_257_13_9 (.A1(n_257_13_10), .A2(n_257_13_9), .A3(n_257_13_85), 
      .ZN(n_257_13_8));
   NAND2_X1 i_257_13_10 (.A1(CPU_Bus[5]), .A2(n_257_13_82), .ZN(n_257_13_9));
   NAND2_X1 i_257_13_11 (.A1(CPU_Bus[6]), .A2(n_254), .ZN(n_257_13_10));
   NAND2_X1 i_257_13_12 (.A1(n_257_13_12), .A2(n_256), .ZN(n_257_13_11));
   NAND2_X1 i_257_13_13 (.A1(n_257_13_16), .A2(n_257_13_13), .ZN(n_257_13_12));
   NAND3_X1 i_257_13_14 (.A1(n_257_13_15), .A2(n_257_13_14), .A3(n_255), 
      .ZN(n_257_13_13));
   NAND2_X1 i_257_13_15 (.A1(CPU_Bus[11]), .A2(n_257_13_82), .ZN(n_257_13_14));
   NAND2_X1 i_257_13_16 (.A1(CPU_Bus[12]), .A2(n_254), .ZN(n_257_13_15));
   NAND3_X1 i_257_13_17 (.A1(n_257_13_18), .A2(n_257_13_17), .A3(n_257_13_85), 
      .ZN(n_257_13_16));
   NAND2_X1 i_257_13_18 (.A1(CPU_Bus[9]), .A2(n_257_13_82), .ZN(n_257_13_17));
   NAND2_X1 i_257_13_19 (.A1(CPU_Bus[10]), .A2(n_254), .ZN(n_257_13_18));
   NAND3_X1 i_257_13_20 (.A1(n_257_13_28), .A2(n_257_13_20), .A3(n_257), 
      .ZN(n_257_13_19));
   NAND2_X1 i_257_13_21 (.A1(n_257_13_21), .A2(n_257_13_86), .ZN(n_257_13_20));
   NAND2_X1 i_257_13_22 (.A1(n_257_13_25), .A2(n_257_13_22), .ZN(n_257_13_21));
   NAND3_X1 i_257_13_23 (.A1(n_257_13_24), .A2(n_257_13_23), .A3(n_255), 
      .ZN(n_257_13_22));
   NAND2_X1 i_257_13_24 (.A1(CPU_Bus[15]), .A2(n_257_13_82), .ZN(n_257_13_23));
   NAND2_X1 i_257_13_25 (.A1(CPU_Bus[16]), .A2(n_254), .ZN(n_257_13_24));
   NAND3_X1 i_257_13_26 (.A1(n_257_13_27), .A2(n_257_13_26), .A3(n_257_13_85), 
      .ZN(n_257_13_25));
   NAND2_X1 i_257_13_27 (.A1(CPU_Bus[13]), .A2(n_257_13_82), .ZN(n_257_13_26));
   NAND2_X1 i_257_13_28 (.A1(CPU_Bus[14]), .A2(n_254), .ZN(n_257_13_27));
   NAND2_X1 i_257_13_29 (.A1(n_257_13_29), .A2(n_256), .ZN(n_257_13_28));
   NAND2_X1 i_257_13_30 (.A1(n_257_13_33), .A2(n_257_13_30), .ZN(n_257_13_29));
   NAND3_X1 i_257_13_31 (.A1(n_257_13_32), .A2(n_257_13_31), .A3(n_255), 
      .ZN(n_257_13_30));
   NAND2_X1 i_257_13_32 (.A1(CPU_Bus[19]), .A2(n_257_13_82), .ZN(n_257_13_31));
   NAND2_X1 i_257_13_33 (.A1(CPU_Bus[20]), .A2(n_254), .ZN(n_257_13_32));
   NAND3_X1 i_257_13_34 (.A1(n_257_13_35), .A2(n_257_13_34), .A3(n_257_13_85), 
      .ZN(n_257_13_33));
   NAND2_X1 i_257_13_35 (.A1(CPU_Bus[17]), .A2(n_257_13_82), .ZN(n_257_13_34));
   NAND2_X1 i_257_13_36 (.A1(CPU_Bus[18]), .A2(n_254), .ZN(n_257_13_35));
   NAND2_X1 i_257_13_37 (.A1(n_257_13_37), .A2(n_257_13_88), .ZN(n_257_13_36));
   NAND2_X1 i_257_13_38 (.A1(n_257_13_61), .A2(n_257_13_38), .ZN(n_257_13_37));
   NAND3_X1 i_257_13_39 (.A1(n_257_13_50), .A2(n_257_13_39), .A3(n_257), 
      .ZN(n_257_13_38));
   NAND3_X1 i_257_13_40 (.A1(n_257_13_45), .A2(n_257_13_40), .A3(n_257_13_86), 
      .ZN(n_257_13_39));
   NAND3_X1 i_257_13_41 (.A1(n_257_13_43), .A2(n_257_13_41), .A3(n_255), 
      .ZN(n_257_13_40));
   NAND2_X1 i_257_13_42 (.A1(n_257_13_42), .A2(n_257_13_82), .ZN(n_257_13_41));
   INV_X1 i_257_13_43 (.A(CPU_Bus[31]), .ZN(n_257_13_42));
   NAND2_X1 i_257_13_44 (.A1(n_257_13_44), .A2(n_254), .ZN(n_257_13_43));
   INV_X1 i_257_13_45 (.A(CPU_Bus[0]), .ZN(n_257_13_44));
   NAND3_X1 i_257_13_46 (.A1(n_257_13_48), .A2(n_257_13_46), .A3(n_257_13_85), 
      .ZN(n_257_13_45));
   NAND2_X1 i_257_13_47 (.A1(n_257_13_47), .A2(n_257_13_82), .ZN(n_257_13_46));
   INV_X1 i_257_13_48 (.A(CPU_Bus[29]), .ZN(n_257_13_47));
   NAND2_X1 i_257_13_49 (.A1(n_257_13_49), .A2(n_254), .ZN(n_257_13_48));
   INV_X1 i_257_13_50 (.A(CPU_Bus[30]), .ZN(n_257_13_49));
   NAND3_X1 i_257_13_51 (.A1(n_257_13_56), .A2(n_257_13_51), .A3(n_256), 
      .ZN(n_257_13_50));
   NAND3_X1 i_257_13_52 (.A1(n_257_13_54), .A2(n_257_13_52), .A3(n_257_13_85), 
      .ZN(n_257_13_51));
   NAND2_X1 i_257_13_53 (.A1(n_257_13_53), .A2(n_257_13_82), .ZN(n_257_13_52));
   INV_X1 i_257_13_54 (.A(CPU_Bus[1]), .ZN(n_257_13_53));
   NAND2_X1 i_257_13_55 (.A1(n_257_13_55), .A2(n_254), .ZN(n_257_13_54));
   INV_X1 i_257_13_56 (.A(CPU_Bus[2]), .ZN(n_257_13_55));
   NAND3_X1 i_257_13_57 (.A1(n_257_13_59), .A2(n_257_13_57), .A3(n_255), 
      .ZN(n_257_13_56));
   NAND2_X1 i_257_13_58 (.A1(n_257_13_58), .A2(n_257_13_82), .ZN(n_257_13_57));
   INV_X1 i_257_13_59 (.A(CPU_Bus[3]), .ZN(n_257_13_58));
   NAND2_X1 i_257_13_60 (.A1(n_257_13_60), .A2(n_254), .ZN(n_257_13_59));
   INV_X1 i_257_13_61 (.A(CPU_Bus[4]), .ZN(n_257_13_60));
   NAND3_X1 i_257_13_62 (.A1(n_257_13_73), .A2(n_257_13_62), .A3(n_257_13_87), 
      .ZN(n_257_13_61));
   NAND3_X1 i_257_13_63 (.A1(n_257_13_68), .A2(n_257_13_63), .A3(n_256), 
      .ZN(n_257_13_62));
   NAND3_X1 i_257_13_64 (.A1(n_257_13_66), .A2(n_257_13_64), .A3(n_257_13_85), 
      .ZN(n_257_13_63));
   NAND2_X1 i_257_13_65 (.A1(n_257_13_65), .A2(n_257_13_82), .ZN(n_257_13_64));
   INV_X1 i_257_13_66 (.A(CPU_Bus[25]), .ZN(n_257_13_65));
   NAND2_X1 i_257_13_67 (.A1(n_257_13_67), .A2(n_254), .ZN(n_257_13_66));
   INV_X1 i_257_13_68 (.A(CPU_Bus[26]), .ZN(n_257_13_67));
   NAND3_X1 i_257_13_69 (.A1(n_257_13_71), .A2(n_257_13_69), .A3(n_255), 
      .ZN(n_257_13_68));
   NAND2_X1 i_257_13_70 (.A1(n_257_13_70), .A2(n_257_13_82), .ZN(n_257_13_69));
   INV_X1 i_257_13_71 (.A(CPU_Bus[27]), .ZN(n_257_13_70));
   NAND2_X1 i_257_13_72 (.A1(n_257_13_72), .A2(n_254), .ZN(n_257_13_71));
   INV_X1 i_257_13_73 (.A(CPU_Bus[28]), .ZN(n_257_13_72));
   NAND3_X1 i_257_13_74 (.A1(n_257_13_79), .A2(n_257_13_74), .A3(n_257_13_86), 
      .ZN(n_257_13_73));
   NAND3_X1 i_257_13_75 (.A1(n_257_13_77), .A2(n_257_13_75), .A3(n_255), 
      .ZN(n_257_13_74));
   NAND2_X1 i_257_13_76 (.A1(n_257_13_76), .A2(n_257_13_82), .ZN(n_257_13_75));
   INV_X1 i_257_13_77 (.A(CPU_Bus[23]), .ZN(n_257_13_76));
   NAND2_X1 i_257_13_78 (.A1(n_257_13_78), .A2(n_254), .ZN(n_257_13_77));
   INV_X1 i_257_13_79 (.A(CPU_Bus[24]), .ZN(n_257_13_78));
   NAND3_X1 i_257_13_80 (.A1(n_257_13_83), .A2(n_257_13_80), .A3(n_257_13_85), 
      .ZN(n_257_13_79));
   NAND2_X1 i_257_13_81 (.A1(n_257_13_81), .A2(n_257_13_82), .ZN(n_257_13_80));
   INV_X1 i_257_13_82 (.A(CPU_Bus[21]), .ZN(n_257_13_81));
   INV_X1 i_257_13_83 (.A(n_254), .ZN(n_257_13_82));
   NAND2_X1 i_257_13_84 (.A1(n_257_13_84), .A2(n_254), .ZN(n_257_13_83));
   INV_X1 i_257_13_85 (.A(CPU_Bus[22]), .ZN(n_257_13_84));
   INV_X1 i_257_13_86 (.A(n_255), .ZN(n_257_13_85));
   INV_X1 i_257_13_87 (.A(n_256), .ZN(n_257_13_86));
   INV_X1 i_257_13_88 (.A(n_257), .ZN(n_257_13_87));
   INV_X1 i_257_13_89 (.A(n_258), .ZN(n_257_13_88));
   NAND2_X1 i_257_14_0 (.A1(n_257_14_49), .A2(n_257_14_0), .ZN(n_257_24));
   NAND2_X1 i_257_14_1 (.A1(n_257_14_1), .A2(n_257_14_48), .ZN(n_257_14_0));
   NAND2_X1 i_257_14_2 (.A1(n_257_14_25), .A2(n_257_14_2), .ZN(n_257_14_1));
   NAND3_X1 i_257_14_3 (.A1(n_257_14_14), .A2(n_257_14_3), .A3(n_257), .ZN(
      n_257_14_2));
   NAND3_X1 i_257_14_4 (.A1(n_257_14_9), .A2(n_257_14_4), .A3(n_256), .ZN(
      n_257_14_3));
   NAND3_X1 i_257_14_5 (.A1(n_257_14_7), .A2(n_257_14_5), .A3(n_255), .ZN(
      n_257_14_4));
   NAND2_X1 i_257_14_6 (.A1(n_257_14_6), .A2(n_257_14_95), .ZN(n_257_14_5));
   INV_X1 i_257_14_7 (.A(CPU_Bus[2]), .ZN(n_257_14_6));
   NAND2_X1 i_257_14_8 (.A1(n_257_14_8), .A2(n_254), .ZN(n_257_14_7));
   INV_X1 i_257_14_9 (.A(CPU_Bus[3]), .ZN(n_257_14_8));
   NAND3_X1 i_257_14_10 (.A1(n_257_14_12), .A2(n_257_14_10), .A3(n_257_14_96), 
      .ZN(n_257_14_9));
   NAND2_X1 i_257_14_11 (.A1(n_257_14_11), .A2(n_254), .ZN(n_257_14_10));
   INV_X1 i_257_14_12 (.A(CPU_Bus[1]), .ZN(n_257_14_11));
   NAND2_X1 i_257_14_13 (.A1(n_257_14_13), .A2(n_257_14_95), .ZN(n_257_14_12));
   INV_X1 i_257_14_14 (.A(CPU_Bus[0]), .ZN(n_257_14_13));
   NAND3_X1 i_257_14_15 (.A1(n_257_14_20), .A2(n_257_14_15), .A3(n_257_14_97), 
      .ZN(n_257_14_14));
   NAND3_X1 i_257_14_16 (.A1(n_257_14_18), .A2(n_257_14_16), .A3(n_257_14_96), 
      .ZN(n_257_14_15));
   NAND2_X1 i_257_14_17 (.A1(n_257_14_17), .A2(n_257_14_95), .ZN(n_257_14_16));
   INV_X1 i_257_14_18 (.A(CPU_Bus[28]), .ZN(n_257_14_17));
   NAND2_X1 i_257_14_19 (.A1(n_257_14_19), .A2(n_254), .ZN(n_257_14_18));
   INV_X1 i_257_14_20 (.A(CPU_Bus[29]), .ZN(n_257_14_19));
   NAND3_X1 i_257_14_21 (.A1(n_257_14_23), .A2(n_257_14_21), .A3(n_255), 
      .ZN(n_257_14_20));
   NAND2_X1 i_257_14_22 (.A1(n_257_14_22), .A2(n_254), .ZN(n_257_14_21));
   INV_X1 i_257_14_23 (.A(CPU_Bus[31]), .ZN(n_257_14_22));
   NAND2_X1 i_257_14_24 (.A1(n_257_14_24), .A2(n_257_14_95), .ZN(n_257_14_23));
   INV_X1 i_257_14_25 (.A(CPU_Bus[30]), .ZN(n_257_14_24));
   NAND3_X1 i_257_14_26 (.A1(n_257_14_37), .A2(n_257_14_26), .A3(n_257_14_98), 
      .ZN(n_257_14_25));
   NAND3_X1 i_257_14_27 (.A1(n_257_14_32), .A2(n_257_14_27), .A3(n_256), 
      .ZN(n_257_14_26));
   NAND3_X1 i_257_14_28 (.A1(n_257_14_30), .A2(n_257_14_28), .A3(n_255), 
      .ZN(n_257_14_27));
   NAND2_X1 i_257_14_29 (.A1(n_257_14_29), .A2(n_257_14_95), .ZN(n_257_14_28));
   INV_X1 i_257_14_30 (.A(CPU_Bus[26]), .ZN(n_257_14_29));
   NAND2_X1 i_257_14_31 (.A1(n_257_14_31), .A2(n_254), .ZN(n_257_14_30));
   INV_X1 i_257_14_32 (.A(CPU_Bus[27]), .ZN(n_257_14_31));
   NAND3_X1 i_257_14_33 (.A1(n_257_14_35), .A2(n_257_14_33), .A3(n_257_14_96), 
      .ZN(n_257_14_32));
   NAND2_X1 i_257_14_34 (.A1(n_257_14_34), .A2(n_254), .ZN(n_257_14_33));
   INV_X1 i_257_14_35 (.A(CPU_Bus[25]), .ZN(n_257_14_34));
   NAND2_X1 i_257_14_36 (.A1(n_257_14_36), .A2(n_257_14_95), .ZN(n_257_14_35));
   INV_X1 i_257_14_37 (.A(CPU_Bus[24]), .ZN(n_257_14_36));
   NAND3_X1 i_257_14_38 (.A1(n_257_14_43), .A2(n_257_14_38), .A3(n_257_14_97), 
      .ZN(n_257_14_37));
   NAND3_X1 i_257_14_39 (.A1(n_257_14_41), .A2(n_257_14_39), .A3(n_257_14_96), 
      .ZN(n_257_14_38));
   NAND2_X1 i_257_14_40 (.A1(n_257_14_40), .A2(n_257_14_95), .ZN(n_257_14_39));
   INV_X1 i_257_14_41 (.A(CPU_Bus[20]), .ZN(n_257_14_40));
   NAND2_X1 i_257_14_42 (.A1(n_257_14_42), .A2(n_254), .ZN(n_257_14_41));
   INV_X1 i_257_14_43 (.A(CPU_Bus[21]), .ZN(n_257_14_42));
   NAND3_X1 i_257_14_44 (.A1(n_257_14_46), .A2(n_257_14_44), .A3(n_255), 
      .ZN(n_257_14_43));
   NAND2_X1 i_257_14_45 (.A1(n_257_14_45), .A2(n_254), .ZN(n_257_14_44));
   INV_X1 i_257_14_46 (.A(CPU_Bus[23]), .ZN(n_257_14_45));
   NAND2_X1 i_257_14_47 (.A1(n_257_14_47), .A2(n_257_14_95), .ZN(n_257_14_46));
   INV_X1 i_257_14_48 (.A(CPU_Bus[22]), .ZN(n_257_14_47));
   INV_X1 i_257_14_49 (.A(n_258), .ZN(n_257_14_48));
   NAND2_X1 i_257_14_50 (.A1(n_257_14_50), .A2(n_258), .ZN(n_257_14_49));
   NAND2_X1 i_257_14_51 (.A1(n_257_14_74), .A2(n_257_14_51), .ZN(n_257_14_50));
   NAND3_X1 i_257_14_52 (.A1(n_257_14_63), .A2(n_257_14_52), .A3(n_257), 
      .ZN(n_257_14_51));
   NAND3_X1 i_257_14_53 (.A1(n_257_14_58), .A2(n_257_14_53), .A3(n_256), 
      .ZN(n_257_14_52));
   NAND3_X1 i_257_14_54 (.A1(n_257_14_56), .A2(n_257_14_54), .A3(n_257_14_96), 
      .ZN(n_257_14_53));
   NAND2_X1 i_257_14_55 (.A1(n_257_14_55), .A2(n_254), .ZN(n_257_14_54));
   INV_X1 i_257_14_56 (.A(CPU_Bus[17]), .ZN(n_257_14_55));
   NAND2_X1 i_257_14_57 (.A1(n_257_14_57), .A2(n_257_14_95), .ZN(n_257_14_56));
   INV_X1 i_257_14_58 (.A(CPU_Bus[16]), .ZN(n_257_14_57));
   NAND3_X1 i_257_14_59 (.A1(n_257_14_61), .A2(n_257_14_59), .A3(n_255), 
      .ZN(n_257_14_58));
   NAND2_X1 i_257_14_60 (.A1(n_257_14_60), .A2(n_254), .ZN(n_257_14_59));
   INV_X1 i_257_14_61 (.A(CPU_Bus[19]), .ZN(n_257_14_60));
   NAND2_X1 i_257_14_62 (.A1(n_257_14_62), .A2(n_257_14_95), .ZN(n_257_14_61));
   INV_X1 i_257_14_63 (.A(CPU_Bus[18]), .ZN(n_257_14_62));
   NAND3_X1 i_257_14_64 (.A1(n_257_14_69), .A2(n_257_14_64), .A3(n_257_14_97), 
      .ZN(n_257_14_63));
   NAND3_X1 i_257_14_65 (.A1(n_257_14_67), .A2(n_257_14_65), .A3(n_255), 
      .ZN(n_257_14_64));
   NAND2_X1 i_257_14_66 (.A1(n_257_14_66), .A2(n_254), .ZN(n_257_14_65));
   INV_X1 i_257_14_67 (.A(CPU_Bus[15]), .ZN(n_257_14_66));
   NAND2_X1 i_257_14_68 (.A1(n_257_14_68), .A2(n_257_14_95), .ZN(n_257_14_67));
   INV_X1 i_257_14_69 (.A(CPU_Bus[14]), .ZN(n_257_14_68));
   NAND3_X1 i_257_14_70 (.A1(n_257_14_72), .A2(n_257_14_70), .A3(n_257_14_96), 
      .ZN(n_257_14_69));
   NAND2_X1 i_257_14_71 (.A1(n_257_14_71), .A2(n_254), .ZN(n_257_14_70));
   INV_X1 i_257_14_72 (.A(CPU_Bus[13]), .ZN(n_257_14_71));
   NAND2_X1 i_257_14_73 (.A1(n_257_14_73), .A2(n_257_14_95), .ZN(n_257_14_72));
   INV_X1 i_257_14_74 (.A(CPU_Bus[12]), .ZN(n_257_14_73));
   NAND3_X1 i_257_14_75 (.A1(n_257_14_86), .A2(n_257_14_98), .A3(n_257_14_75), 
      .ZN(n_257_14_74));
   NAND3_X1 i_257_14_76 (.A1(n_257_14_81), .A2(n_257_14_76), .A3(n_256), 
      .ZN(n_257_14_75));
   NAND3_X1 i_257_14_77 (.A1(n_257_14_79), .A2(n_257_14_77), .A3(n_257_14_96), 
      .ZN(n_257_14_76));
   NAND2_X1 i_257_14_78 (.A1(n_257_14_78), .A2(n_254), .ZN(n_257_14_77));
   INV_X1 i_257_14_79 (.A(CPU_Bus[9]), .ZN(n_257_14_78));
   NAND2_X1 i_257_14_80 (.A1(n_257_14_80), .A2(n_257_14_95), .ZN(n_257_14_79));
   INV_X1 i_257_14_81 (.A(CPU_Bus[8]), .ZN(n_257_14_80));
   NAND3_X1 i_257_14_82 (.A1(n_257_14_84), .A2(n_257_14_82), .A3(n_255), 
      .ZN(n_257_14_81));
   NAND2_X1 i_257_14_83 (.A1(n_257_14_83), .A2(n_254), .ZN(n_257_14_82));
   INV_X1 i_257_14_84 (.A(CPU_Bus[11]), .ZN(n_257_14_83));
   NAND2_X1 i_257_14_85 (.A1(n_257_14_85), .A2(n_257_14_95), .ZN(n_257_14_84));
   INV_X1 i_257_14_86 (.A(CPU_Bus[10]), .ZN(n_257_14_85));
   NAND3_X1 i_257_14_87 (.A1(n_257_14_92), .A2(n_257_14_97), .A3(n_257_14_87), 
      .ZN(n_257_14_86));
   NAND3_X1 i_257_14_88 (.A1(n_257_14_90), .A2(n_257_14_88), .A3(n_255), 
      .ZN(n_257_14_87));
   NAND2_X1 i_257_14_89 (.A1(n_257_14_89), .A2(n_254), .ZN(n_257_14_88));
   INV_X1 i_257_14_90 (.A(CPU_Bus[7]), .ZN(n_257_14_89));
   NAND2_X1 i_257_14_91 (.A1(n_257_14_91), .A2(n_257_14_95), .ZN(n_257_14_90));
   INV_X1 i_257_14_92 (.A(CPU_Bus[6]), .ZN(n_257_14_91));
   OAI211_X1 i_257_14_93 (.A(n_257_14_93), .B(n_257_14_96), .C1(n_257_14_95), 
      .C2(CPU_Bus[5]), .ZN(n_257_14_92));
   NAND2_X1 i_257_14_94 (.A1(n_257_14_94), .A2(n_257_14_95), .ZN(n_257_14_93));
   INV_X1 i_257_14_95 (.A(CPU_Bus[4]), .ZN(n_257_14_94));
   INV_X1 i_257_14_96 (.A(n_254), .ZN(n_257_14_95));
   INV_X1 i_257_14_97 (.A(n_255), .ZN(n_257_14_96));
   INV_X1 i_257_14_98 (.A(n_256), .ZN(n_257_14_97));
   INV_X1 i_257_14_99 (.A(n_257), .ZN(n_257_14_98));
   INV_X1 i_257_15_0 (.A(n_254), .ZN(n_257_15_0));
   NAND2_X1 i_257_15_1 (.A1(n_257_15_0), .A2(n_255), .ZN(n_257_15_1));
   INV_X1 i_257_15_2 (.A(n_256), .ZN(n_257_15_2));
   NOR2_X1 i_257_15_3 (.A1(n_257_15_1), .A2(n_257_15_2), .ZN(n_257_15_3));
   NAND2_X1 i_257_15_4 (.A1(n_257_15_3), .A2(n_257), .ZN(n_257_15_4));
   INV_X1 i_257_15_5 (.A(n_258), .ZN(n_257_15_5));
   NOR2_X1 i_257_15_6 (.A1(n_257_15_4), .A2(n_257_15_5), .ZN(n_257_15_6));
   NAND2_X1 i_257_15_7 (.A1(CPU_Bus[17]), .A2(n_257_15_6), .ZN(n_257_15_7));
   INV_X1 i_257_15_8 (.A(n_255), .ZN(n_257_15_8));
   NAND2_X1 i_257_15_9 (.A1(n_257_15_0), .A2(n_257_15_8), .ZN(n_257_15_9));
   NOR2_X1 i_257_15_10 (.A1(n_257_15_9), .A2(n_257_15_2), .ZN(n_257_15_10));
   NAND2_X1 i_257_15_11 (.A1(n_257_15_10), .A2(n_257), .ZN(n_257_15_11));
   NOR2_X1 i_257_15_12 (.A1(n_257_15_11), .A2(n_257_15_5), .ZN(n_257_15_12));
   NAND2_X1 i_257_15_13 (.A1(CPU_Bus[15]), .A2(n_257_15_12), .ZN(n_257_15_13));
   NAND2_X1 i_257_15_14 (.A1(n_257_15_7), .A2(n_257_15_13), .ZN(n_257_15_14));
   NOR2_X1 i_257_15_15 (.A1(n_257_15_1), .A2(n_256), .ZN(n_257_15_15));
   NAND2_X1 i_257_15_16 (.A1(n_257_15_15), .A2(n_257), .ZN(n_257_15_16));
   NOR2_X1 i_257_15_17 (.A1(n_257_15_16), .A2(n_257_15_5), .ZN(n_257_15_17));
   NAND2_X1 i_257_15_18 (.A1(CPU_Bus[13]), .A2(n_257_15_17), .ZN(n_257_15_18));
   NOR2_X1 i_257_15_19 (.A1(n_257_15_9), .A2(n_256), .ZN(n_257_15_19));
   NAND2_X1 i_257_15_20 (.A1(n_257_15_19), .A2(n_257), .ZN(n_257_15_20));
   NOR2_X1 i_257_15_21 (.A1(n_257_15_20), .A2(n_257_15_5), .ZN(n_257_15_21));
   NAND2_X1 i_257_15_22 (.A1(CPU_Bus[11]), .A2(n_257_15_21), .ZN(n_257_15_22));
   NAND2_X1 i_257_15_23 (.A1(n_257_15_18), .A2(n_257_15_22), .ZN(n_257_15_23));
   NOR2_X1 i_257_15_24 (.A1(n_257_15_14), .A2(n_257_15_23), .ZN(n_257_15_24));
   INV_X1 i_257_15_25 (.A(n_257), .ZN(n_257_15_25));
   NAND2_X1 i_257_15_26 (.A1(n_257_15_3), .A2(n_257_15_25), .ZN(n_257_15_26));
   NOR2_X1 i_257_15_27 (.A1(n_257_15_26), .A2(n_257_15_5), .ZN(n_257_15_27));
   NAND2_X1 i_257_15_28 (.A1(CPU_Bus[9]), .A2(n_257_15_27), .ZN(n_257_15_28));
   NAND2_X1 i_257_15_29 (.A1(n_257_15_10), .A2(n_257_15_25), .ZN(n_257_15_29));
   NOR2_X1 i_257_15_30 (.A1(n_257_15_29), .A2(n_257_15_5), .ZN(n_257_15_30));
   NAND2_X1 i_257_15_31 (.A1(CPU_Bus[7]), .A2(n_257_15_30), .ZN(n_257_15_31));
   NAND2_X1 i_257_15_32 (.A1(n_257_15_28), .A2(n_257_15_31), .ZN(n_257_15_32));
   NAND2_X1 i_257_15_33 (.A1(n_257_15_15), .A2(n_257_15_25), .ZN(n_257_15_33));
   NOR2_X1 i_257_15_34 (.A1(n_257_15_33), .A2(n_257_15_5), .ZN(n_257_15_34));
   NAND2_X1 i_257_15_35 (.A1(CPU_Bus[5]), .A2(n_257_15_34), .ZN(n_257_15_35));
   NAND2_X1 i_257_15_36 (.A1(n_257_15_19), .A2(n_257_15_25), .ZN(n_257_15_36));
   NOR2_X1 i_257_15_37 (.A1(n_257_15_36), .A2(n_257_15_5), .ZN(n_257_15_37));
   NAND2_X1 i_257_15_38 (.A1(CPU_Bus[3]), .A2(n_257_15_37), .ZN(n_257_15_38));
   NAND2_X1 i_257_15_39 (.A1(n_257_15_35), .A2(n_257_15_38), .ZN(n_257_15_39));
   NOR2_X1 i_257_15_40 (.A1(n_257_15_32), .A2(n_257_15_39), .ZN(n_257_15_40));
   NAND2_X1 i_257_15_41 (.A1(n_257_15_24), .A2(n_257_15_40), .ZN(n_257_15_41));
   NOR2_X1 i_257_15_42 (.A1(n_257_15_4), .A2(n_258), .ZN(n_257_15_42));
   NAND2_X1 i_257_15_43 (.A1(CPU_Bus[1]), .A2(n_257_15_42), .ZN(n_257_15_43));
   NOR2_X1 i_257_15_44 (.A1(n_257_15_11), .A2(n_258), .ZN(n_257_15_44));
   NAND2_X1 i_257_15_45 (.A1(CPU_Bus[31]), .A2(n_257_15_44), .ZN(n_257_15_45));
   NAND2_X1 i_257_15_46 (.A1(n_257_15_43), .A2(n_257_15_45), .ZN(n_257_15_46));
   NOR2_X1 i_257_15_47 (.A1(n_257_15_16), .A2(n_258), .ZN(n_257_15_47));
   NAND2_X1 i_257_15_48 (.A1(CPU_Bus[29]), .A2(n_257_15_47), .ZN(n_257_15_48));
   NOR2_X1 i_257_15_49 (.A1(n_257_15_20), .A2(n_258), .ZN(n_257_15_49));
   NAND2_X1 i_257_15_50 (.A1(CPU_Bus[27]), .A2(n_257_15_49), .ZN(n_257_15_50));
   NAND2_X1 i_257_15_51 (.A1(n_257_15_48), .A2(n_257_15_50), .ZN(n_257_15_51));
   NOR2_X1 i_257_15_52 (.A1(n_257_15_46), .A2(n_257_15_51), .ZN(n_257_15_52));
   NOR2_X1 i_257_15_53 (.A1(n_257_15_26), .A2(n_258), .ZN(n_257_15_53));
   NAND2_X1 i_257_15_54 (.A1(CPU_Bus[25]), .A2(n_257_15_53), .ZN(n_257_15_54));
   NOR2_X1 i_257_15_55 (.A1(n_257_15_29), .A2(n_258), .ZN(n_257_15_55));
   NAND2_X1 i_257_15_56 (.A1(CPU_Bus[23]), .A2(n_257_15_55), .ZN(n_257_15_56));
   NAND2_X1 i_257_15_57 (.A1(n_257_15_54), .A2(n_257_15_56), .ZN(n_257_15_57));
   NOR2_X1 i_257_15_58 (.A1(n_257_15_33), .A2(n_258), .ZN(n_257_15_58));
   NAND2_X1 i_257_15_59 (.A1(CPU_Bus[21]), .A2(n_257_15_58), .ZN(n_257_15_59));
   NOR2_X1 i_257_15_60 (.A1(n_257_15_36), .A2(n_258), .ZN(n_257_15_60));
   NAND2_X1 i_257_15_61 (.A1(CPU_Bus[19]), .A2(n_257_15_60), .ZN(n_257_15_61));
   NAND2_X1 i_257_15_62 (.A1(n_257_15_59), .A2(n_257_15_61), .ZN(n_257_15_62));
   NOR2_X1 i_257_15_63 (.A1(n_257_15_57), .A2(n_257_15_62), .ZN(n_257_15_63));
   NAND2_X1 i_257_15_64 (.A1(n_257_15_52), .A2(n_257_15_63), .ZN(n_257_15_64));
   NOR2_X1 i_257_15_65 (.A1(n_257_15_41), .A2(n_257_15_64), .ZN(n_257_15_65));
   NAND2_X1 i_257_15_66 (.A1(n_257_15_8), .A2(n_254), .ZN(n_257_15_66));
   NOR2_X1 i_257_15_67 (.A1(n_257_15_66), .A2(n_257_15_2), .ZN(n_257_15_67));
   NAND2_X1 i_257_15_68 (.A1(n_257_15_67), .A2(n_257), .ZN(n_257_15_68));
   NOR2_X1 i_257_15_69 (.A1(n_257_15_68), .A2(n_257_15_5), .ZN(n_257_15_69));
   NAND2_X1 i_257_15_70 (.A1(CPU_Bus[16]), .A2(n_257_15_69), .ZN(n_257_15_70));
   NOR2_X1 i_257_15_71 (.A1(n_257_15_66), .A2(n_256), .ZN(n_257_15_71));
   NAND2_X1 i_257_15_72 (.A1(n_257_15_71), .A2(n_257), .ZN(n_257_15_72));
   NOR2_X1 i_257_15_73 (.A1(n_257_15_72), .A2(n_257_15_5), .ZN(n_257_15_73));
   NAND2_X1 i_257_15_74 (.A1(CPU_Bus[12]), .A2(n_257_15_73), .ZN(n_257_15_74));
   NAND2_X1 i_257_15_75 (.A1(n_257_15_70), .A2(n_257_15_74), .ZN(n_257_15_75));
   NAND2_X1 i_257_15_76 (.A1(n_257_15_67), .A2(n_257_15_25), .ZN(n_257_15_76));
   NOR2_X1 i_257_15_77 (.A1(n_257_15_76), .A2(n_257_15_5), .ZN(n_257_15_77));
   NAND2_X1 i_257_15_78 (.A1(CPU_Bus[8]), .A2(n_257_15_77), .ZN(n_257_15_78));
   NAND2_X1 i_257_15_79 (.A1(n_257_15_71), .A2(n_257_15_25), .ZN(n_257_15_79));
   NOR2_X1 i_257_15_80 (.A1(n_257_15_79), .A2(n_257_15_5), .ZN(n_257_15_80));
   NAND2_X1 i_257_15_81 (.A1(CPU_Bus[4]), .A2(n_257_15_80), .ZN(n_257_15_81));
   NAND2_X1 i_257_15_82 (.A1(n_257_15_78), .A2(n_257_15_81), .ZN(n_257_15_82));
   NOR2_X1 i_257_15_83 (.A1(n_257_15_75), .A2(n_257_15_82), .ZN(n_257_15_83));
   NOR2_X1 i_257_15_84 (.A1(n_257_15_68), .A2(n_258), .ZN(n_257_15_84));
   NAND2_X1 i_257_15_85 (.A1(CPU_Bus[0]), .A2(n_257_15_84), .ZN(n_257_15_85));
   NOR2_X1 i_257_15_86 (.A1(n_257_15_72), .A2(n_258), .ZN(n_257_15_86));
   NAND2_X1 i_257_15_87 (.A1(CPU_Bus[28]), .A2(n_257_15_86), .ZN(n_257_15_87));
   NAND2_X1 i_257_15_88 (.A1(n_257_15_85), .A2(n_257_15_87), .ZN(n_257_15_88));
   NOR2_X1 i_257_15_89 (.A1(n_257_15_76), .A2(n_258), .ZN(n_257_15_89));
   NAND2_X1 i_257_15_90 (.A1(CPU_Bus[24]), .A2(n_257_15_89), .ZN(n_257_15_90));
   NOR2_X1 i_257_15_91 (.A1(n_257_15_79), .A2(n_258), .ZN(n_257_15_91));
   NAND2_X1 i_257_15_92 (.A1(CPU_Bus[20]), .A2(n_257_15_91), .ZN(n_257_15_92));
   NAND2_X1 i_257_15_93 (.A1(n_257_15_90), .A2(n_257_15_92), .ZN(n_257_15_93));
   NOR2_X1 i_257_15_94 (.A1(n_257_15_88), .A2(n_257_15_93), .ZN(n_257_15_94));
   NAND2_X1 i_257_15_95 (.A1(n_257_15_83), .A2(n_257_15_94), .ZN(n_257_15_95));
   NAND2_X1 i_257_15_96 (.A1(n_254), .A2(n_255), .ZN(n_257_15_96));
   NOR2_X1 i_257_15_97 (.A1(n_257_15_96), .A2(n_257_15_2), .ZN(n_257_15_97));
   NAND2_X1 i_257_15_98 (.A1(n_257_15_97), .A2(n_257), .ZN(n_257_15_98));
   NOR2_X1 i_257_15_99 (.A1(n_257_15_98), .A2(n_257_15_5), .ZN(n_257_15_99));
   NAND2_X1 i_257_15_100 (.A1(CPU_Bus[18]), .A2(n_257_15_99), .ZN(n_257_15_100));
   NOR2_X1 i_257_15_101 (.A1(n_257_15_96), .A2(n_256), .ZN(n_257_15_101));
   NAND2_X1 i_257_15_102 (.A1(n_257_15_101), .A2(n_257), .ZN(n_257_15_102));
   NOR2_X1 i_257_15_103 (.A1(n_257_15_102), .A2(n_257_15_5), .ZN(n_257_15_103));
   NAND2_X1 i_257_15_104 (.A1(CPU_Bus[14]), .A2(n_257_15_103), .ZN(n_257_15_104));
   NAND2_X1 i_257_15_105 (.A1(n_257_15_100), .A2(n_257_15_104), .ZN(n_257_15_105));
   NAND2_X1 i_257_15_106 (.A1(n_257_15_97), .A2(n_257_15_25), .ZN(n_257_15_106));
   NOR2_X1 i_257_15_107 (.A1(n_257_15_106), .A2(n_257_15_5), .ZN(n_257_15_107));
   NAND2_X1 i_257_15_108 (.A1(CPU_Bus[10]), .A2(n_257_15_107), .ZN(n_257_15_108));
   NAND2_X1 i_257_15_109 (.A1(n_257_15_101), .A2(n_257_15_25), .ZN(n_257_15_109));
   NOR2_X1 i_257_15_110 (.A1(n_257_15_109), .A2(n_257_15_5), .ZN(n_257_15_110));
   NAND2_X1 i_257_15_111 (.A1(CPU_Bus[6]), .A2(n_257_15_110), .ZN(n_257_15_111));
   NAND2_X1 i_257_15_112 (.A1(n_257_15_108), .A2(n_257_15_111), .ZN(n_257_15_112));
   NOR2_X1 i_257_15_113 (.A1(n_257_15_105), .A2(n_257_15_112), .ZN(n_257_15_113));
   NOR2_X1 i_257_15_114 (.A1(n_257_15_98), .A2(n_258), .ZN(n_257_15_114));
   NAND2_X1 i_257_15_115 (.A1(CPU_Bus[2]), .A2(n_257_15_114), .ZN(n_257_15_115));
   NOR2_X1 i_257_15_116 (.A1(n_257_15_102), .A2(n_258), .ZN(n_257_15_116));
   NAND2_X1 i_257_15_117 (.A1(CPU_Bus[30]), .A2(n_257_15_116), .ZN(n_257_15_117));
   NAND2_X1 i_257_15_118 (.A1(n_257_15_115), .A2(n_257_15_117), .ZN(n_257_15_118));
   NOR2_X1 i_257_15_119 (.A1(n_257_15_106), .A2(n_258), .ZN(n_257_15_119));
   NAND2_X1 i_257_15_120 (.A1(CPU_Bus[26]), .A2(n_257_15_119), .ZN(n_257_15_120));
   NOR2_X1 i_257_15_121 (.A1(n_257_15_109), .A2(n_258), .ZN(n_257_15_121));
   NAND2_X1 i_257_15_122 (.A1(CPU_Bus[22]), .A2(n_257_15_121), .ZN(n_257_15_122));
   NAND2_X1 i_257_15_123 (.A1(n_257_15_120), .A2(n_257_15_122), .ZN(n_257_15_123));
   NOR2_X1 i_257_15_124 (.A1(n_257_15_118), .A2(n_257_15_123), .ZN(n_257_15_124));
   NAND2_X1 i_257_15_125 (.A1(n_257_15_113), .A2(n_257_15_124), .ZN(n_257_15_125));
   NOR2_X1 i_257_15_126 (.A1(n_257_15_95), .A2(n_257_15_125), .ZN(n_257_15_126));
   NAND2_X1 i_257_15_127 (.A1(n_257_15_65), .A2(n_257_15_126), .ZN(n_257_25));
   INV_X1 i_257_16_0 (.A(n_254), .ZN(n_257_16_0));
   NAND2_X1 i_257_16_1 (.A1(n_257_16_0), .A2(n_255), .ZN(n_257_16_1));
   INV_X1 i_257_16_2 (.A(n_256), .ZN(n_257_16_2));
   NOR2_X1 i_257_16_3 (.A1(n_257_16_1), .A2(n_257_16_2), .ZN(n_257_16_3));
   NAND2_X1 i_257_16_4 (.A1(n_257_16_3), .A2(n_257), .ZN(n_257_16_4));
   INV_X1 i_257_16_5 (.A(n_258), .ZN(n_257_16_5));
   NOR2_X1 i_257_16_6 (.A1(n_257_16_4), .A2(n_257_16_5), .ZN(n_257_16_6));
   NAND2_X1 i_257_16_7 (.A1(CPU_Bus[16]), .A2(n_257_16_6), .ZN(n_257_16_7));
   INV_X1 i_257_16_8 (.A(n_255), .ZN(n_257_16_8));
   NAND2_X1 i_257_16_9 (.A1(n_257_16_0), .A2(n_257_16_8), .ZN(n_257_16_9));
   NOR2_X1 i_257_16_10 (.A1(n_257_16_9), .A2(n_257_16_2), .ZN(n_257_16_10));
   NAND2_X1 i_257_16_11 (.A1(n_257_16_10), .A2(n_257), .ZN(n_257_16_11));
   NOR2_X1 i_257_16_12 (.A1(n_257_16_11), .A2(n_257_16_5), .ZN(n_257_16_12));
   NAND2_X1 i_257_16_13 (.A1(CPU_Bus[14]), .A2(n_257_16_12), .ZN(n_257_16_13));
   NAND2_X1 i_257_16_14 (.A1(n_257_16_7), .A2(n_257_16_13), .ZN(n_257_16_14));
   NOR2_X1 i_257_16_15 (.A1(n_257_16_1), .A2(n_256), .ZN(n_257_16_15));
   NAND2_X1 i_257_16_16 (.A1(n_257_16_15), .A2(n_257), .ZN(n_257_16_16));
   NOR2_X1 i_257_16_17 (.A1(n_257_16_16), .A2(n_257_16_5), .ZN(n_257_16_17));
   NAND2_X1 i_257_16_18 (.A1(CPU_Bus[12]), .A2(n_257_16_17), .ZN(n_257_16_18));
   NOR2_X1 i_257_16_19 (.A1(n_257_16_9), .A2(n_256), .ZN(n_257_16_19));
   NAND2_X1 i_257_16_20 (.A1(n_257_16_19), .A2(n_257), .ZN(n_257_16_20));
   NOR2_X1 i_257_16_21 (.A1(n_257_16_20), .A2(n_257_16_5), .ZN(n_257_16_21));
   NAND2_X1 i_257_16_22 (.A1(CPU_Bus[10]), .A2(n_257_16_21), .ZN(n_257_16_22));
   NAND2_X1 i_257_16_23 (.A1(n_257_16_18), .A2(n_257_16_22), .ZN(n_257_16_23));
   NOR2_X1 i_257_16_24 (.A1(n_257_16_14), .A2(n_257_16_23), .ZN(n_257_16_24));
   INV_X1 i_257_16_25 (.A(n_257), .ZN(n_257_16_25));
   NAND2_X1 i_257_16_26 (.A1(n_257_16_3), .A2(n_257_16_25), .ZN(n_257_16_26));
   NOR2_X1 i_257_16_27 (.A1(n_257_16_26), .A2(n_257_16_5), .ZN(n_257_16_27));
   NAND2_X1 i_257_16_28 (.A1(CPU_Bus[8]), .A2(n_257_16_27), .ZN(n_257_16_28));
   NAND2_X1 i_257_16_29 (.A1(n_257_16_10), .A2(n_257_16_25), .ZN(n_257_16_29));
   NOR2_X1 i_257_16_30 (.A1(n_257_16_29), .A2(n_257_16_5), .ZN(n_257_16_30));
   NAND2_X1 i_257_16_31 (.A1(CPU_Bus[6]), .A2(n_257_16_30), .ZN(n_257_16_31));
   NAND2_X1 i_257_16_32 (.A1(n_257_16_28), .A2(n_257_16_31), .ZN(n_257_16_32));
   NAND2_X1 i_257_16_33 (.A1(n_257_16_15), .A2(n_257_16_25), .ZN(n_257_16_33));
   NOR2_X1 i_257_16_34 (.A1(n_257_16_33), .A2(n_257_16_5), .ZN(n_257_16_34));
   NAND2_X1 i_257_16_35 (.A1(CPU_Bus[4]), .A2(n_257_16_34), .ZN(n_257_16_35));
   NAND2_X1 i_257_16_36 (.A1(n_257_16_19), .A2(n_257_16_25), .ZN(n_257_16_36));
   NOR2_X1 i_257_16_37 (.A1(n_257_16_36), .A2(n_257_16_5), .ZN(n_257_16_37));
   NAND2_X1 i_257_16_38 (.A1(CPU_Bus[2]), .A2(n_257_16_37), .ZN(n_257_16_38));
   NAND2_X1 i_257_16_39 (.A1(n_257_16_35), .A2(n_257_16_38), .ZN(n_257_16_39));
   NOR2_X1 i_257_16_40 (.A1(n_257_16_32), .A2(n_257_16_39), .ZN(n_257_16_40));
   NAND2_X1 i_257_16_41 (.A1(n_257_16_24), .A2(n_257_16_40), .ZN(n_257_16_41));
   NOR2_X1 i_257_16_42 (.A1(n_257_16_4), .A2(n_258), .ZN(n_257_16_42));
   NAND2_X1 i_257_16_43 (.A1(CPU_Bus[0]), .A2(n_257_16_42), .ZN(n_257_16_43));
   NOR2_X1 i_257_16_44 (.A1(n_257_16_11), .A2(n_258), .ZN(n_257_16_44));
   NAND2_X1 i_257_16_45 (.A1(CPU_Bus[30]), .A2(n_257_16_44), .ZN(n_257_16_45));
   NAND2_X1 i_257_16_46 (.A1(n_257_16_43), .A2(n_257_16_45), .ZN(n_257_16_46));
   NOR2_X1 i_257_16_47 (.A1(n_257_16_16), .A2(n_258), .ZN(n_257_16_47));
   NAND2_X1 i_257_16_48 (.A1(CPU_Bus[28]), .A2(n_257_16_47), .ZN(n_257_16_48));
   NOR2_X1 i_257_16_49 (.A1(n_257_16_20), .A2(n_258), .ZN(n_257_16_49));
   NAND2_X1 i_257_16_50 (.A1(CPU_Bus[26]), .A2(n_257_16_49), .ZN(n_257_16_50));
   NAND2_X1 i_257_16_51 (.A1(n_257_16_48), .A2(n_257_16_50), .ZN(n_257_16_51));
   NOR2_X1 i_257_16_52 (.A1(n_257_16_46), .A2(n_257_16_51), .ZN(n_257_16_52));
   NOR2_X1 i_257_16_53 (.A1(n_257_16_26), .A2(n_258), .ZN(n_257_16_53));
   NAND2_X1 i_257_16_54 (.A1(CPU_Bus[24]), .A2(n_257_16_53), .ZN(n_257_16_54));
   NOR2_X1 i_257_16_55 (.A1(n_257_16_29), .A2(n_258), .ZN(n_257_16_55));
   NAND2_X1 i_257_16_56 (.A1(CPU_Bus[22]), .A2(n_257_16_55), .ZN(n_257_16_56));
   NAND2_X1 i_257_16_57 (.A1(n_257_16_54), .A2(n_257_16_56), .ZN(n_257_16_57));
   NOR2_X1 i_257_16_58 (.A1(n_257_16_33), .A2(n_258), .ZN(n_257_16_58));
   NAND2_X1 i_257_16_59 (.A1(CPU_Bus[20]), .A2(n_257_16_58), .ZN(n_257_16_59));
   NOR2_X1 i_257_16_60 (.A1(n_257_16_36), .A2(n_258), .ZN(n_257_16_60));
   NAND2_X1 i_257_16_61 (.A1(CPU_Bus[18]), .A2(n_257_16_60), .ZN(n_257_16_61));
   NAND2_X1 i_257_16_62 (.A1(n_257_16_59), .A2(n_257_16_61), .ZN(n_257_16_62));
   NOR2_X1 i_257_16_63 (.A1(n_257_16_57), .A2(n_257_16_62), .ZN(n_257_16_63));
   NAND2_X1 i_257_16_64 (.A1(n_257_16_52), .A2(n_257_16_63), .ZN(n_257_16_64));
   NOR2_X1 i_257_16_65 (.A1(n_257_16_41), .A2(n_257_16_64), .ZN(n_257_16_65));
   NAND2_X1 i_257_16_66 (.A1(n_257_16_8), .A2(n_254), .ZN(n_257_16_66));
   NOR2_X1 i_257_16_67 (.A1(n_257_16_66), .A2(n_257_16_2), .ZN(n_257_16_67));
   NAND2_X1 i_257_16_68 (.A1(n_257_16_67), .A2(n_257), .ZN(n_257_16_68));
   NOR2_X1 i_257_16_69 (.A1(n_257_16_68), .A2(n_257_16_5), .ZN(n_257_16_69));
   NAND2_X1 i_257_16_70 (.A1(CPU_Bus[15]), .A2(n_257_16_69), .ZN(n_257_16_70));
   NOR2_X1 i_257_16_71 (.A1(n_257_16_66), .A2(n_256), .ZN(n_257_16_71));
   NAND2_X1 i_257_16_72 (.A1(n_257_16_71), .A2(n_257), .ZN(n_257_16_72));
   NOR2_X1 i_257_16_73 (.A1(n_257_16_72), .A2(n_257_16_5), .ZN(n_257_16_73));
   NAND2_X1 i_257_16_74 (.A1(CPU_Bus[11]), .A2(n_257_16_73), .ZN(n_257_16_74));
   NAND2_X1 i_257_16_75 (.A1(n_257_16_70), .A2(n_257_16_74), .ZN(n_257_16_75));
   NAND2_X1 i_257_16_76 (.A1(n_257_16_67), .A2(n_257_16_25), .ZN(n_257_16_76));
   NOR2_X1 i_257_16_77 (.A1(n_257_16_76), .A2(n_257_16_5), .ZN(n_257_16_77));
   NAND2_X1 i_257_16_78 (.A1(CPU_Bus[7]), .A2(n_257_16_77), .ZN(n_257_16_78));
   NAND2_X1 i_257_16_79 (.A1(n_257_16_71), .A2(n_257_16_25), .ZN(n_257_16_79));
   NOR2_X1 i_257_16_80 (.A1(n_257_16_79), .A2(n_257_16_5), .ZN(n_257_16_80));
   NAND2_X1 i_257_16_81 (.A1(CPU_Bus[3]), .A2(n_257_16_80), .ZN(n_257_16_81));
   NAND2_X1 i_257_16_82 (.A1(n_257_16_78), .A2(n_257_16_81), .ZN(n_257_16_82));
   NOR2_X1 i_257_16_83 (.A1(n_257_16_75), .A2(n_257_16_82), .ZN(n_257_16_83));
   NOR2_X1 i_257_16_84 (.A1(n_257_16_68), .A2(n_258), .ZN(n_257_16_84));
   NAND2_X1 i_257_16_85 (.A1(CPU_Bus[31]), .A2(n_257_16_84), .ZN(n_257_16_85));
   NOR2_X1 i_257_16_86 (.A1(n_257_16_72), .A2(n_258), .ZN(n_257_16_86));
   NAND2_X1 i_257_16_87 (.A1(CPU_Bus[27]), .A2(n_257_16_86), .ZN(n_257_16_87));
   NAND2_X1 i_257_16_88 (.A1(n_257_16_85), .A2(n_257_16_87), .ZN(n_257_16_88));
   NOR2_X1 i_257_16_89 (.A1(n_257_16_76), .A2(n_258), .ZN(n_257_16_89));
   NAND2_X1 i_257_16_90 (.A1(CPU_Bus[23]), .A2(n_257_16_89), .ZN(n_257_16_90));
   NOR2_X1 i_257_16_91 (.A1(n_257_16_79), .A2(n_258), .ZN(n_257_16_91));
   NAND2_X1 i_257_16_92 (.A1(CPU_Bus[19]), .A2(n_257_16_91), .ZN(n_257_16_92));
   NAND2_X1 i_257_16_93 (.A1(n_257_16_90), .A2(n_257_16_92), .ZN(n_257_16_93));
   NOR2_X1 i_257_16_94 (.A1(n_257_16_88), .A2(n_257_16_93), .ZN(n_257_16_94));
   NAND2_X1 i_257_16_95 (.A1(n_257_16_83), .A2(n_257_16_94), .ZN(n_257_16_95));
   NAND2_X1 i_257_16_96 (.A1(n_254), .A2(n_255), .ZN(n_257_16_96));
   NOR2_X1 i_257_16_97 (.A1(n_257_16_96), .A2(n_257_16_2), .ZN(n_257_16_97));
   NAND2_X1 i_257_16_98 (.A1(n_257_16_97), .A2(n_257), .ZN(n_257_16_98));
   NOR2_X1 i_257_16_99 (.A1(n_257_16_98), .A2(n_257_16_5), .ZN(n_257_16_99));
   NAND2_X1 i_257_16_100 (.A1(CPU_Bus[17]), .A2(n_257_16_99), .ZN(n_257_16_100));
   NOR2_X1 i_257_16_101 (.A1(n_257_16_96), .A2(n_256), .ZN(n_257_16_101));
   NAND2_X1 i_257_16_102 (.A1(n_257_16_101), .A2(n_257), .ZN(n_257_16_102));
   NOR2_X1 i_257_16_103 (.A1(n_257_16_102), .A2(n_257_16_5), .ZN(n_257_16_103));
   NAND2_X1 i_257_16_104 (.A1(CPU_Bus[13]), .A2(n_257_16_103), .ZN(n_257_16_104));
   NAND2_X1 i_257_16_105 (.A1(n_257_16_100), .A2(n_257_16_104), .ZN(n_257_16_105));
   NAND2_X1 i_257_16_106 (.A1(n_257_16_97), .A2(n_257_16_25), .ZN(n_257_16_106));
   NOR2_X1 i_257_16_107 (.A1(n_257_16_106), .A2(n_257_16_5), .ZN(n_257_16_107));
   NAND2_X1 i_257_16_108 (.A1(CPU_Bus[9]), .A2(n_257_16_107), .ZN(n_257_16_108));
   NAND2_X1 i_257_16_109 (.A1(n_257_16_101), .A2(n_257_16_25), .ZN(n_257_16_109));
   NOR2_X1 i_257_16_110 (.A1(n_257_16_109), .A2(n_257_16_5), .ZN(n_257_16_110));
   NAND2_X1 i_257_16_111 (.A1(CPU_Bus[5]), .A2(n_257_16_110), .ZN(n_257_16_111));
   NAND2_X1 i_257_16_112 (.A1(n_257_16_108), .A2(n_257_16_111), .ZN(n_257_16_112));
   NOR2_X1 i_257_16_113 (.A1(n_257_16_105), .A2(n_257_16_112), .ZN(n_257_16_113));
   NOR2_X1 i_257_16_114 (.A1(n_257_16_98), .A2(n_258), .ZN(n_257_16_114));
   NAND2_X1 i_257_16_115 (.A1(CPU_Bus[1]), .A2(n_257_16_114), .ZN(n_257_16_115));
   NOR2_X1 i_257_16_116 (.A1(n_257_16_102), .A2(n_258), .ZN(n_257_16_116));
   NAND2_X1 i_257_16_117 (.A1(CPU_Bus[29]), .A2(n_257_16_116), .ZN(n_257_16_117));
   NAND2_X1 i_257_16_118 (.A1(n_257_16_115), .A2(n_257_16_117), .ZN(n_257_16_118));
   NOR2_X1 i_257_16_119 (.A1(n_257_16_106), .A2(n_258), .ZN(n_257_16_119));
   NAND2_X1 i_257_16_120 (.A1(CPU_Bus[25]), .A2(n_257_16_119), .ZN(n_257_16_120));
   NOR2_X1 i_257_16_121 (.A1(n_257_16_109), .A2(n_258), .ZN(n_257_16_121));
   NAND2_X1 i_257_16_122 (.A1(CPU_Bus[21]), .A2(n_257_16_121), .ZN(n_257_16_122));
   NAND2_X1 i_257_16_123 (.A1(n_257_16_120), .A2(n_257_16_122), .ZN(n_257_16_123));
   NOR2_X1 i_257_16_124 (.A1(n_257_16_118), .A2(n_257_16_123), .ZN(n_257_16_124));
   NAND2_X1 i_257_16_125 (.A1(n_257_16_113), .A2(n_257_16_124), .ZN(n_257_16_125));
   NOR2_X1 i_257_16_126 (.A1(n_257_16_95), .A2(n_257_16_125), .ZN(n_257_16_126));
   NAND2_X1 i_257_16_127 (.A1(n_257_16_65), .A2(n_257_16_126), .ZN(n_257_26));
   NAND2_X1 i_257_17_0 (.A1(n_257_17_49), .A2(n_257_17_0), .ZN(n_257_27));
   NAND2_X1 i_257_17_1 (.A1(n_257_17_1), .A2(n_257_17_48), .ZN(n_257_17_0));
   NAND2_X1 i_257_17_2 (.A1(n_257_17_25), .A2(n_257_17_2), .ZN(n_257_17_1));
   NAND3_X1 i_257_17_3 (.A1(n_257_17_14), .A2(n_257_17_3), .A3(n_257), .ZN(
      n_257_17_2));
   NAND3_X1 i_257_17_4 (.A1(n_257_17_9), .A2(n_257_17_4), .A3(n_256), .ZN(
      n_257_17_3));
   NAND3_X1 i_257_17_5 (.A1(n_257_17_7), .A2(n_257_17_5), .A3(n_255), .ZN(
      n_257_17_4));
   NAND2_X1 i_257_17_6 (.A1(n_257_17_6), .A2(n_257_17_95), .ZN(n_257_17_5));
   INV_X1 i_257_17_7 (.A(CPU_Bus[31]), .ZN(n_257_17_6));
   NAND2_X1 i_257_17_8 (.A1(n_257_17_8), .A2(n_254), .ZN(n_257_17_7));
   INV_X1 i_257_17_9 (.A(CPU_Bus[0]), .ZN(n_257_17_8));
   NAND3_X1 i_257_17_10 (.A1(n_257_17_12), .A2(n_257_17_10), .A3(n_257_17_96), 
      .ZN(n_257_17_9));
   NAND2_X1 i_257_17_11 (.A1(n_257_17_11), .A2(n_254), .ZN(n_257_17_10));
   INV_X1 i_257_17_12 (.A(CPU_Bus[30]), .ZN(n_257_17_11));
   NAND2_X1 i_257_17_13 (.A1(n_257_17_13), .A2(n_257_17_95), .ZN(n_257_17_12));
   INV_X1 i_257_17_14 (.A(CPU_Bus[29]), .ZN(n_257_17_13));
   NAND3_X1 i_257_17_15 (.A1(n_257_17_20), .A2(n_257_17_15), .A3(n_257_17_97), 
      .ZN(n_257_17_14));
   NAND3_X1 i_257_17_16 (.A1(n_257_17_18), .A2(n_257_17_16), .A3(n_257_17_96), 
      .ZN(n_257_17_15));
   NAND2_X1 i_257_17_17 (.A1(n_257_17_17), .A2(n_257_17_95), .ZN(n_257_17_16));
   INV_X1 i_257_17_18 (.A(CPU_Bus[25]), .ZN(n_257_17_17));
   NAND2_X1 i_257_17_19 (.A1(n_257_17_19), .A2(n_254), .ZN(n_257_17_18));
   INV_X1 i_257_17_20 (.A(CPU_Bus[26]), .ZN(n_257_17_19));
   NAND3_X1 i_257_17_21 (.A1(n_257_17_23), .A2(n_257_17_21), .A3(n_255), 
      .ZN(n_257_17_20));
   NAND2_X1 i_257_17_22 (.A1(n_257_17_22), .A2(n_254), .ZN(n_257_17_21));
   INV_X1 i_257_17_23 (.A(CPU_Bus[28]), .ZN(n_257_17_22));
   NAND2_X1 i_257_17_24 (.A1(n_257_17_24), .A2(n_257_17_95), .ZN(n_257_17_23));
   INV_X1 i_257_17_25 (.A(CPU_Bus[27]), .ZN(n_257_17_24));
   NAND3_X1 i_257_17_26 (.A1(n_257_17_37), .A2(n_257_17_26), .A3(n_257_17_98), 
      .ZN(n_257_17_25));
   NAND3_X1 i_257_17_27 (.A1(n_257_17_32), .A2(n_257_17_27), .A3(n_256), 
      .ZN(n_257_17_26));
   NAND3_X1 i_257_17_28 (.A1(n_257_17_30), .A2(n_257_17_28), .A3(n_255), 
      .ZN(n_257_17_27));
   NAND2_X1 i_257_17_29 (.A1(n_257_17_29), .A2(n_257_17_95), .ZN(n_257_17_28));
   INV_X1 i_257_17_30 (.A(CPU_Bus[23]), .ZN(n_257_17_29));
   NAND2_X1 i_257_17_31 (.A1(n_257_17_31), .A2(n_254), .ZN(n_257_17_30));
   INV_X1 i_257_17_32 (.A(CPU_Bus[24]), .ZN(n_257_17_31));
   NAND3_X1 i_257_17_33 (.A1(n_257_17_35), .A2(n_257_17_33), .A3(n_257_17_96), 
      .ZN(n_257_17_32));
   NAND2_X1 i_257_17_34 (.A1(n_257_17_34), .A2(n_254), .ZN(n_257_17_33));
   INV_X1 i_257_17_35 (.A(CPU_Bus[22]), .ZN(n_257_17_34));
   NAND2_X1 i_257_17_36 (.A1(n_257_17_36), .A2(n_257_17_95), .ZN(n_257_17_35));
   INV_X1 i_257_17_37 (.A(CPU_Bus[21]), .ZN(n_257_17_36));
   NAND3_X1 i_257_17_38 (.A1(n_257_17_43), .A2(n_257_17_38), .A3(n_257_17_97), 
      .ZN(n_257_17_37));
   NAND3_X1 i_257_17_39 (.A1(n_257_17_41), .A2(n_257_17_39), .A3(n_257_17_96), 
      .ZN(n_257_17_38));
   NAND2_X1 i_257_17_40 (.A1(n_257_17_40), .A2(n_257_17_95), .ZN(n_257_17_39));
   INV_X1 i_257_17_41 (.A(CPU_Bus[17]), .ZN(n_257_17_40));
   NAND2_X1 i_257_17_42 (.A1(n_257_17_42), .A2(n_254), .ZN(n_257_17_41));
   INV_X1 i_257_17_43 (.A(CPU_Bus[18]), .ZN(n_257_17_42));
   NAND3_X1 i_257_17_44 (.A1(n_257_17_46), .A2(n_257_17_44), .A3(n_255), 
      .ZN(n_257_17_43));
   NAND2_X1 i_257_17_45 (.A1(n_257_17_45), .A2(n_254), .ZN(n_257_17_44));
   INV_X1 i_257_17_46 (.A(CPU_Bus[20]), .ZN(n_257_17_45));
   NAND2_X1 i_257_17_47 (.A1(n_257_17_47), .A2(n_257_17_95), .ZN(n_257_17_46));
   INV_X1 i_257_17_48 (.A(CPU_Bus[19]), .ZN(n_257_17_47));
   INV_X1 i_257_17_49 (.A(n_258), .ZN(n_257_17_48));
   NAND2_X1 i_257_17_50 (.A1(n_257_17_50), .A2(n_258), .ZN(n_257_17_49));
   NAND2_X1 i_257_17_51 (.A1(n_257_17_74), .A2(n_257_17_51), .ZN(n_257_17_50));
   NAND3_X1 i_257_17_52 (.A1(n_257_17_63), .A2(n_257_17_52), .A3(n_257), 
      .ZN(n_257_17_51));
   NAND3_X1 i_257_17_53 (.A1(n_257_17_58), .A2(n_257_17_53), .A3(n_256), 
      .ZN(n_257_17_52));
   NAND3_X1 i_257_17_54 (.A1(n_257_17_56), .A2(n_257_17_54), .A3(n_257_17_96), 
      .ZN(n_257_17_53));
   NAND2_X1 i_257_17_55 (.A1(n_257_17_55), .A2(n_254), .ZN(n_257_17_54));
   INV_X1 i_257_17_56 (.A(CPU_Bus[14]), .ZN(n_257_17_55));
   NAND2_X1 i_257_17_57 (.A1(n_257_17_57), .A2(n_257_17_95), .ZN(n_257_17_56));
   INV_X1 i_257_17_58 (.A(CPU_Bus[13]), .ZN(n_257_17_57));
   NAND3_X1 i_257_17_59 (.A1(n_257_17_61), .A2(n_257_17_59), .A3(n_255), 
      .ZN(n_257_17_58));
   NAND2_X1 i_257_17_60 (.A1(n_257_17_60), .A2(n_254), .ZN(n_257_17_59));
   INV_X1 i_257_17_61 (.A(CPU_Bus[16]), .ZN(n_257_17_60));
   NAND2_X1 i_257_17_62 (.A1(n_257_17_62), .A2(n_257_17_95), .ZN(n_257_17_61));
   INV_X1 i_257_17_63 (.A(CPU_Bus[15]), .ZN(n_257_17_62));
   NAND3_X1 i_257_17_64 (.A1(n_257_17_69), .A2(n_257_17_64), .A3(n_257_17_97), 
      .ZN(n_257_17_63));
   NAND3_X1 i_257_17_65 (.A1(n_257_17_67), .A2(n_257_17_65), .A3(n_255), 
      .ZN(n_257_17_64));
   NAND2_X1 i_257_17_66 (.A1(n_257_17_66), .A2(n_254), .ZN(n_257_17_65));
   INV_X1 i_257_17_67 (.A(CPU_Bus[12]), .ZN(n_257_17_66));
   NAND2_X1 i_257_17_68 (.A1(n_257_17_68), .A2(n_257_17_95), .ZN(n_257_17_67));
   INV_X1 i_257_17_69 (.A(CPU_Bus[11]), .ZN(n_257_17_68));
   NAND3_X1 i_257_17_70 (.A1(n_257_17_72), .A2(n_257_17_70), .A3(n_257_17_96), 
      .ZN(n_257_17_69));
   NAND2_X1 i_257_17_71 (.A1(n_257_17_71), .A2(n_254), .ZN(n_257_17_70));
   INV_X1 i_257_17_72 (.A(CPU_Bus[10]), .ZN(n_257_17_71));
   NAND2_X1 i_257_17_73 (.A1(n_257_17_73), .A2(n_257_17_95), .ZN(n_257_17_72));
   INV_X1 i_257_17_74 (.A(CPU_Bus[9]), .ZN(n_257_17_73));
   NAND3_X1 i_257_17_75 (.A1(n_257_17_86), .A2(n_257_17_98), .A3(n_257_17_75), 
      .ZN(n_257_17_74));
   NAND3_X1 i_257_17_76 (.A1(n_257_17_81), .A2(n_257_17_76), .A3(n_256), 
      .ZN(n_257_17_75));
   NAND3_X1 i_257_17_77 (.A1(n_257_17_79), .A2(n_257_17_77), .A3(n_257_17_96), 
      .ZN(n_257_17_76));
   NAND2_X1 i_257_17_78 (.A1(n_257_17_78), .A2(n_254), .ZN(n_257_17_77));
   INV_X1 i_257_17_79 (.A(CPU_Bus[6]), .ZN(n_257_17_78));
   NAND2_X1 i_257_17_80 (.A1(n_257_17_80), .A2(n_257_17_95), .ZN(n_257_17_79));
   INV_X1 i_257_17_81 (.A(CPU_Bus[5]), .ZN(n_257_17_80));
   NAND3_X1 i_257_17_82 (.A1(n_257_17_84), .A2(n_257_17_82), .A3(n_255), 
      .ZN(n_257_17_81));
   NAND2_X1 i_257_17_83 (.A1(n_257_17_83), .A2(n_254), .ZN(n_257_17_82));
   INV_X1 i_257_17_84 (.A(CPU_Bus[8]), .ZN(n_257_17_83));
   NAND2_X1 i_257_17_85 (.A1(n_257_17_85), .A2(n_257_17_95), .ZN(n_257_17_84));
   INV_X1 i_257_17_86 (.A(CPU_Bus[7]), .ZN(n_257_17_85));
   NAND3_X1 i_257_17_87 (.A1(n_257_17_92), .A2(n_257_17_97), .A3(n_257_17_87), 
      .ZN(n_257_17_86));
   NAND3_X1 i_257_17_88 (.A1(n_257_17_90), .A2(n_257_17_88), .A3(n_255), 
      .ZN(n_257_17_87));
   NAND2_X1 i_257_17_89 (.A1(n_257_17_89), .A2(n_254), .ZN(n_257_17_88));
   INV_X1 i_257_17_90 (.A(CPU_Bus[4]), .ZN(n_257_17_89));
   NAND2_X1 i_257_17_91 (.A1(n_257_17_91), .A2(n_257_17_95), .ZN(n_257_17_90));
   INV_X1 i_257_17_92 (.A(CPU_Bus[3]), .ZN(n_257_17_91));
   OAI211_X1 i_257_17_93 (.A(n_257_17_93), .B(n_257_17_96), .C1(n_257_17_95), 
      .C2(CPU_Bus[2]), .ZN(n_257_17_92));
   NAND2_X1 i_257_17_94 (.A1(n_257_17_94), .A2(n_257_17_95), .ZN(n_257_17_93));
   INV_X1 i_257_17_95 (.A(CPU_Bus[1]), .ZN(n_257_17_94));
   INV_X1 i_257_17_96 (.A(n_254), .ZN(n_257_17_95));
   INV_X1 i_257_17_97 (.A(n_255), .ZN(n_257_17_96));
   INV_X1 i_257_17_98 (.A(n_256), .ZN(n_257_17_97));
   INV_X1 i_257_17_99 (.A(n_257), .ZN(n_257_17_98));
   INV_X1 i_257_18_0 (.A(n_257_18_0), .ZN(n_257_28));
   NAND2_X1 i_257_18_1 (.A1(n_257_18_49), .A2(n_257_18_1), .ZN(n_257_18_0));
   NAND3_X1 i_257_18_2 (.A1(n_257_18_25), .A2(n_257_18_2), .A3(n_257_18_48), 
      .ZN(n_257_18_1));
   NAND3_X1 i_257_18_3 (.A1(n_257_18_14), .A2(n_257_18_3), .A3(n_257), .ZN(
      n_257_18_2));
   NAND3_X1 i_257_18_4 (.A1(n_257_18_9), .A2(n_257_18_4), .A3(n_257_18_85), 
      .ZN(n_257_18_3));
   NAND3_X1 i_257_18_5 (.A1(n_257_18_7), .A2(n_257_18_5), .A3(n_257_18_96), 
      .ZN(n_257_18_4));
   NAND2_X1 i_257_18_6 (.A1(n_257_18_6), .A2(n_257_18_95), .ZN(n_257_18_5));
   INV_X1 i_257_18_7 (.A(CPU_Bus[24]), .ZN(n_257_18_6));
   NAND2_X1 i_257_18_8 (.A1(n_257_18_8), .A2(n_254), .ZN(n_257_18_7));
   INV_X1 i_257_18_9 (.A(CPU_Bus[25]), .ZN(n_257_18_8));
   NAND3_X1 i_257_18_10 (.A1(n_257_18_12), .A2(n_257_18_10), .A3(n_255), 
      .ZN(n_257_18_9));
   NAND2_X1 i_257_18_11 (.A1(n_257_18_11), .A2(n_257_18_95), .ZN(n_257_18_10));
   INV_X1 i_257_18_12 (.A(CPU_Bus[26]), .ZN(n_257_18_11));
   NAND2_X1 i_257_18_13 (.A1(n_257_18_13), .A2(n_254), .ZN(n_257_18_12));
   INV_X1 i_257_18_14 (.A(CPU_Bus[27]), .ZN(n_257_18_13));
   NAND3_X1 i_257_18_15 (.A1(n_257_18_20), .A2(n_257_18_15), .A3(n_256), 
      .ZN(n_257_18_14));
   NAND3_X1 i_257_18_16 (.A1(n_257_18_18), .A2(n_257_18_16), .A3(n_257_18_96), 
      .ZN(n_257_18_15));
   NAND2_X1 i_257_18_17 (.A1(n_257_18_17), .A2(n_257_18_95), .ZN(n_257_18_16));
   INV_X1 i_257_18_18 (.A(CPU_Bus[28]), .ZN(n_257_18_17));
   NAND2_X1 i_257_18_19 (.A1(n_257_18_19), .A2(n_254), .ZN(n_257_18_18));
   INV_X1 i_257_18_20 (.A(CPU_Bus[29]), .ZN(n_257_18_19));
   NAND3_X1 i_257_18_21 (.A1(n_257_18_23), .A2(n_257_18_21), .A3(n_255), 
      .ZN(n_257_18_20));
   NAND2_X1 i_257_18_22 (.A1(n_257_18_22), .A2(n_257_18_95), .ZN(n_257_18_21));
   INV_X1 i_257_18_23 (.A(CPU_Bus[30]), .ZN(n_257_18_22));
   NAND2_X1 i_257_18_24 (.A1(n_257_18_24), .A2(n_254), .ZN(n_257_18_23));
   INV_X1 i_257_18_25 (.A(CPU_Bus[31]), .ZN(n_257_18_24));
   NAND3_X1 i_257_18_26 (.A1(n_257_18_37), .A2(n_257_18_26), .A3(n_257_18_97), 
      .ZN(n_257_18_25));
   NAND3_X1 i_257_18_27 (.A1(n_257_18_32), .A2(n_257_18_27), .A3(n_256), 
      .ZN(n_257_18_26));
   NAND3_X1 i_257_18_28 (.A1(n_257_18_30), .A2(n_257_18_28), .A3(n_255), 
      .ZN(n_257_18_27));
   NAND2_X1 i_257_18_29 (.A1(n_257_18_29), .A2(n_254), .ZN(n_257_18_28));
   INV_X1 i_257_18_30 (.A(CPU_Bus[23]), .ZN(n_257_18_29));
   NAND2_X1 i_257_18_31 (.A1(n_257_18_31), .A2(n_257_18_95), .ZN(n_257_18_30));
   INV_X1 i_257_18_32 (.A(CPU_Bus[22]), .ZN(n_257_18_31));
   NAND3_X1 i_257_18_33 (.A1(n_257_18_35), .A2(n_257_18_33), .A3(n_257_18_96), 
      .ZN(n_257_18_32));
   NAND2_X1 i_257_18_34 (.A1(n_257_18_34), .A2(n_257_18_95), .ZN(n_257_18_33));
   INV_X1 i_257_18_35 (.A(CPU_Bus[20]), .ZN(n_257_18_34));
   NAND2_X1 i_257_18_36 (.A1(n_257_18_36), .A2(n_254), .ZN(n_257_18_35));
   INV_X1 i_257_18_37 (.A(CPU_Bus[21]), .ZN(n_257_18_36));
   NAND3_X1 i_257_18_38 (.A1(n_257_18_43), .A2(n_257_18_38), .A3(n_257_18_85), 
      .ZN(n_257_18_37));
   NAND3_X1 i_257_18_39 (.A1(n_257_18_41), .A2(n_257_18_39), .A3(n_255), 
      .ZN(n_257_18_38));
   NAND2_X1 i_257_18_40 (.A1(n_257_18_40), .A2(n_254), .ZN(n_257_18_39));
   INV_X1 i_257_18_41 (.A(CPU_Bus[19]), .ZN(n_257_18_40));
   NAND2_X1 i_257_18_42 (.A1(n_257_18_42), .A2(n_257_18_95), .ZN(n_257_18_41));
   INV_X1 i_257_18_43 (.A(CPU_Bus[18]), .ZN(n_257_18_42));
   NAND3_X1 i_257_18_44 (.A1(n_257_18_46), .A2(n_257_18_44), .A3(n_257_18_96), 
      .ZN(n_257_18_43));
   NAND2_X1 i_257_18_45 (.A1(n_257_18_45), .A2(n_257_18_95), .ZN(n_257_18_44));
   INV_X1 i_257_18_46 (.A(CPU_Bus[16]), .ZN(n_257_18_45));
   NAND2_X1 i_257_18_47 (.A1(n_257_18_47), .A2(n_254), .ZN(n_257_18_46));
   INV_X1 i_257_18_48 (.A(CPU_Bus[17]), .ZN(n_257_18_47));
   INV_X1 i_257_18_49 (.A(n_258), .ZN(n_257_18_48));
   NAND3_X1 i_257_18_50 (.A1(n_257_18_73), .A2(n_257_18_50), .A3(n_258), 
      .ZN(n_257_18_49));
   NAND3_X1 i_257_18_51 (.A1(n_257_18_62), .A2(n_257_18_51), .A3(n_257), 
      .ZN(n_257_18_50));
   NAND3_X1 i_257_18_52 (.A1(n_257_18_57), .A2(n_257_18_52), .A3(n_257_18_85), 
      .ZN(n_257_18_51));
   NAND3_X1 i_257_18_53 (.A1(n_257_18_55), .A2(n_257_18_53), .A3(n_257_18_96), 
      .ZN(n_257_18_52));
   NAND2_X1 i_257_18_54 (.A1(n_257_18_54), .A2(n_257_18_95), .ZN(n_257_18_53));
   INV_X1 i_257_18_55 (.A(CPU_Bus[8]), .ZN(n_257_18_54));
   NAND2_X1 i_257_18_56 (.A1(n_257_18_56), .A2(n_254), .ZN(n_257_18_55));
   INV_X1 i_257_18_57 (.A(CPU_Bus[9]), .ZN(n_257_18_56));
   NAND3_X1 i_257_18_58 (.A1(n_257_18_60), .A2(n_257_18_58), .A3(n_255), 
      .ZN(n_257_18_57));
   NAND2_X1 i_257_18_59 (.A1(n_257_18_59), .A2(n_254), .ZN(n_257_18_58));
   INV_X1 i_257_18_60 (.A(CPU_Bus[11]), .ZN(n_257_18_59));
   NAND2_X1 i_257_18_61 (.A1(n_257_18_61), .A2(n_257_18_95), .ZN(n_257_18_60));
   INV_X1 i_257_18_62 (.A(CPU_Bus[10]), .ZN(n_257_18_61));
   NAND3_X1 i_257_18_63 (.A1(n_257_18_68), .A2(n_257_18_63), .A3(n_256), 
      .ZN(n_257_18_62));
   NAND3_X1 i_257_18_64 (.A1(n_257_18_66), .A2(n_257_18_64), .A3(n_257_18_96), 
      .ZN(n_257_18_63));
   NAND2_X1 i_257_18_65 (.A1(n_257_18_65), .A2(n_254), .ZN(n_257_18_64));
   INV_X1 i_257_18_66 (.A(CPU_Bus[13]), .ZN(n_257_18_65));
   NAND2_X1 i_257_18_67 (.A1(n_257_18_67), .A2(n_257_18_95), .ZN(n_257_18_66));
   INV_X1 i_257_18_68 (.A(CPU_Bus[12]), .ZN(n_257_18_67));
   NAND3_X1 i_257_18_69 (.A1(n_257_18_71), .A2(n_257_18_69), .A3(n_255), 
      .ZN(n_257_18_68));
   NAND2_X1 i_257_18_70 (.A1(n_257_18_70), .A2(n_257_18_95), .ZN(n_257_18_69));
   INV_X1 i_257_18_71 (.A(CPU_Bus[14]), .ZN(n_257_18_70));
   NAND2_X1 i_257_18_72 (.A1(n_257_18_72), .A2(n_254), .ZN(n_257_18_71));
   INV_X1 i_257_18_73 (.A(CPU_Bus[15]), .ZN(n_257_18_72));
   NAND3_X1 i_257_18_74 (.A1(n_257_18_86), .A2(n_257_18_74), .A3(n_257_18_97), 
      .ZN(n_257_18_73));
   NAND3_X1 i_257_18_75 (.A1(n_257_18_80), .A2(n_257_18_75), .A3(n_257_18_85), 
      .ZN(n_257_18_74));
   NAND3_X1 i_257_18_76 (.A1(n_257_18_78), .A2(n_257_18_76), .A3(n_257_18_96), 
      .ZN(n_257_18_75));
   NAND2_X1 i_257_18_77 (.A1(n_257_18_77), .A2(n_254), .ZN(n_257_18_76));
   INV_X1 i_257_18_78 (.A(CPU_Bus[1]), .ZN(n_257_18_77));
   NAND2_X1 i_257_18_79 (.A1(n_257_18_79), .A2(n_257_18_95), .ZN(n_257_18_78));
   INV_X1 i_257_18_80 (.A(CPU_Bus[0]), .ZN(n_257_18_79));
   NAND3_X1 i_257_18_81 (.A1(n_257_18_83), .A2(n_257_18_81), .A3(n_255), 
      .ZN(n_257_18_80));
   NAND2_X1 i_257_18_82 (.A1(n_257_18_82), .A2(n_254), .ZN(n_257_18_81));
   INV_X1 i_257_18_83 (.A(CPU_Bus[3]), .ZN(n_257_18_82));
   NAND2_X1 i_257_18_84 (.A1(n_257_18_84), .A2(n_257_18_95), .ZN(n_257_18_83));
   INV_X1 i_257_18_85 (.A(CPU_Bus[2]), .ZN(n_257_18_84));
   INV_X1 i_257_18_86 (.A(n_256), .ZN(n_257_18_85));
   NAND3_X1 i_257_18_87 (.A1(n_257_18_92), .A2(n_257_18_87), .A3(n_256), 
      .ZN(n_257_18_86));
   NAND3_X1 i_257_18_88 (.A1(n_257_18_90), .A2(n_257_18_88), .A3(n_255), 
      .ZN(n_257_18_87));
   NAND2_X1 i_257_18_89 (.A1(n_257_18_89), .A2(n_257_18_95), .ZN(n_257_18_88));
   INV_X1 i_257_18_90 (.A(CPU_Bus[6]), .ZN(n_257_18_89));
   NAND2_X1 i_257_18_91 (.A1(n_257_18_91), .A2(n_254), .ZN(n_257_18_90));
   INV_X1 i_257_18_92 (.A(CPU_Bus[7]), .ZN(n_257_18_91));
   OAI211_X1 i_257_18_93 (.A(n_257_18_93), .B(n_257_18_96), .C1(n_257_18_95), 
      .C2(CPU_Bus[5]), .ZN(n_257_18_92));
   NAND2_X1 i_257_18_94 (.A1(n_257_18_94), .A2(n_257_18_95), .ZN(n_257_18_93));
   INV_X1 i_257_18_95 (.A(CPU_Bus[4]), .ZN(n_257_18_94));
   INV_X1 i_257_18_96 (.A(n_254), .ZN(n_257_18_95));
   INV_X1 i_257_18_97 (.A(n_255), .ZN(n_257_18_96));
   INV_X1 i_257_18_98 (.A(n_257), .ZN(n_257_18_97));
   datapath__1_338 i_257_19 (.PacketSize(PacketSize), .p_0({n_257_34, uc_104, 
      uc_105, uc_106, uc_107, uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, 
      uc_114, uc_115, uc_116, uc_117, uc_118, uc_119, uc_120, uc_121, uc_122, 
      uc_123, uc_124, uc_125, uc_126, uc_127, uc_128, n_257_33, n_257_32, 
      n_257_31, n_257_30, n_257_29, uc_129}));
   datapath__1_339 i_257_20 (.p_0({uc_130, uc_131, uc_132, uc_133, uc_134, 
      uc_135, uc_136, uc_137, uc_138, uc_139, uc_140, uc_141, uc_142, uc_143, 
      uc_144, uc_145, uc_146, uc_147, uc_148, uc_149, uc_150, uc_151, uc_152, 
      uc_153, uc_154, n_257_34, n_257_33, n_257_32, n_257_31, n_257_30, n_257_29, 
      n_151}), .p_1({n_257_66, n_257_65, n_257_64, n_257_63, n_257_62, n_257_61, 
      n_257_60, n_257_59, n_257_58, n_257_57, n_257_56, n_257_55, n_257_54, 
      n_257_53, n_257_52, n_257_51, n_257_50, n_257_49, n_257_48, n_257_47, 
      n_257_46, n_257_45, n_257_44, n_257_43, n_257_42, n_257_41, n_257_40, 
      n_257_39, n_257_38, n_257_37, n_257_36, n_257_35}));
   NAND2_X1 i_257_21_0 (.A1(n_257_21_49), .A2(n_257_21_0), .ZN(n_257_67));
   NAND2_X1 i_257_21_1 (.A1(n_257_21_1), .A2(n_257_21_48), .ZN(n_257_21_0));
   NAND2_X1 i_257_21_2 (.A1(n_257_21_25), .A2(n_257_21_2), .ZN(n_257_21_1));
   NAND3_X1 i_257_21_3 (.A1(n_257_21_14), .A2(n_257_21_3), .A3(n_257), .ZN(
      n_257_21_2));
   NAND3_X1 i_257_21_4 (.A1(n_257_21_9), .A2(n_257_21_4), .A3(n_256), .ZN(
      n_257_21_3));
   NAND3_X1 i_257_21_5 (.A1(n_257_21_7), .A2(n_257_21_5), .A3(n_255), .ZN(
      n_257_21_4));
   NAND2_X1 i_257_21_6 (.A1(n_257_21_6), .A2(n_257_21_95), .ZN(n_257_21_5));
   INV_X1 i_257_21_7 (.A(CPU_Bus[28]), .ZN(n_257_21_6));
   NAND2_X1 i_257_21_8 (.A1(n_257_21_8), .A2(n_254), .ZN(n_257_21_7));
   INV_X1 i_257_21_9 (.A(CPU_Bus[29]), .ZN(n_257_21_8));
   NAND3_X1 i_257_21_10 (.A1(n_257_21_12), .A2(n_257_21_10), .A3(n_257_21_96), 
      .ZN(n_257_21_9));
   NAND2_X1 i_257_21_11 (.A1(n_257_21_11), .A2(n_254), .ZN(n_257_21_10));
   INV_X1 i_257_21_12 (.A(CPU_Bus[27]), .ZN(n_257_21_11));
   NAND2_X1 i_257_21_13 (.A1(n_257_21_13), .A2(n_257_21_95), .ZN(n_257_21_12));
   INV_X1 i_257_21_14 (.A(CPU_Bus[26]), .ZN(n_257_21_13));
   NAND3_X1 i_257_21_15 (.A1(n_257_21_20), .A2(n_257_21_15), .A3(n_257_21_97), 
      .ZN(n_257_21_14));
   NAND3_X1 i_257_21_16 (.A1(n_257_21_18), .A2(n_257_21_16), .A3(n_257_21_96), 
      .ZN(n_257_21_15));
   NAND2_X1 i_257_21_17 (.A1(n_257_21_17), .A2(n_257_21_95), .ZN(n_257_21_16));
   INV_X1 i_257_21_18 (.A(CPU_Bus[22]), .ZN(n_257_21_17));
   NAND2_X1 i_257_21_19 (.A1(n_257_21_19), .A2(n_254), .ZN(n_257_21_18));
   INV_X1 i_257_21_20 (.A(CPU_Bus[23]), .ZN(n_257_21_19));
   NAND3_X1 i_257_21_21 (.A1(n_257_21_23), .A2(n_257_21_21), .A3(n_255), 
      .ZN(n_257_21_20));
   NAND2_X1 i_257_21_22 (.A1(n_257_21_22), .A2(n_254), .ZN(n_257_21_21));
   INV_X1 i_257_21_23 (.A(CPU_Bus[25]), .ZN(n_257_21_22));
   NAND2_X1 i_257_21_24 (.A1(n_257_21_24), .A2(n_257_21_95), .ZN(n_257_21_23));
   INV_X1 i_257_21_25 (.A(CPU_Bus[24]), .ZN(n_257_21_24));
   NAND3_X1 i_257_21_26 (.A1(n_257_21_37), .A2(n_257_21_26), .A3(n_257_21_98), 
      .ZN(n_257_21_25));
   NAND3_X1 i_257_21_27 (.A1(n_257_21_32), .A2(n_257_21_27), .A3(n_256), 
      .ZN(n_257_21_26));
   NAND3_X1 i_257_21_28 (.A1(n_257_21_30), .A2(n_257_21_28), .A3(n_255), 
      .ZN(n_257_21_27));
   NAND2_X1 i_257_21_29 (.A1(n_257_21_29), .A2(n_257_21_95), .ZN(n_257_21_28));
   INV_X1 i_257_21_30 (.A(CPU_Bus[20]), .ZN(n_257_21_29));
   NAND2_X1 i_257_21_31 (.A1(n_257_21_31), .A2(n_254), .ZN(n_257_21_30));
   INV_X1 i_257_21_32 (.A(CPU_Bus[21]), .ZN(n_257_21_31));
   NAND3_X1 i_257_21_33 (.A1(n_257_21_35), .A2(n_257_21_33), .A3(n_257_21_96), 
      .ZN(n_257_21_32));
   NAND2_X1 i_257_21_34 (.A1(n_257_21_34), .A2(n_254), .ZN(n_257_21_33));
   INV_X1 i_257_21_35 (.A(CPU_Bus[19]), .ZN(n_257_21_34));
   NAND2_X1 i_257_21_36 (.A1(n_257_21_36), .A2(n_257_21_95), .ZN(n_257_21_35));
   INV_X1 i_257_21_37 (.A(CPU_Bus[18]), .ZN(n_257_21_36));
   NAND3_X1 i_257_21_38 (.A1(n_257_21_43), .A2(n_257_21_38), .A3(n_257_21_97), 
      .ZN(n_257_21_37));
   NAND3_X1 i_257_21_39 (.A1(n_257_21_41), .A2(n_257_21_39), .A3(n_257_21_96), 
      .ZN(n_257_21_38));
   NAND2_X1 i_257_21_40 (.A1(n_257_21_40), .A2(n_257_21_95), .ZN(n_257_21_39));
   INV_X1 i_257_21_41 (.A(CPU_Bus[14]), .ZN(n_257_21_40));
   NAND2_X1 i_257_21_42 (.A1(n_257_21_42), .A2(n_254), .ZN(n_257_21_41));
   INV_X1 i_257_21_43 (.A(CPU_Bus[15]), .ZN(n_257_21_42));
   NAND3_X1 i_257_21_44 (.A1(n_257_21_46), .A2(n_257_21_44), .A3(n_255), 
      .ZN(n_257_21_43));
   NAND2_X1 i_257_21_45 (.A1(n_257_21_45), .A2(n_254), .ZN(n_257_21_44));
   INV_X1 i_257_21_46 (.A(CPU_Bus[17]), .ZN(n_257_21_45));
   NAND2_X1 i_257_21_47 (.A1(n_257_21_47), .A2(n_257_21_95), .ZN(n_257_21_46));
   INV_X1 i_257_21_48 (.A(CPU_Bus[16]), .ZN(n_257_21_47));
   INV_X1 i_257_21_49 (.A(n_258), .ZN(n_257_21_48));
   NAND2_X1 i_257_21_50 (.A1(n_257_21_50), .A2(n_258), .ZN(n_257_21_49));
   NAND2_X1 i_257_21_51 (.A1(n_257_21_74), .A2(n_257_21_51), .ZN(n_257_21_50));
   NAND3_X1 i_257_21_52 (.A1(n_257_21_63), .A2(n_257_21_52), .A3(n_257), 
      .ZN(n_257_21_51));
   NAND3_X1 i_257_21_53 (.A1(n_257_21_58), .A2(n_257_21_53), .A3(n_256), 
      .ZN(n_257_21_52));
   NAND3_X1 i_257_21_54 (.A1(n_257_21_56), .A2(n_257_21_54), .A3(n_257_21_96), 
      .ZN(n_257_21_53));
   NAND2_X1 i_257_21_55 (.A1(n_257_21_55), .A2(n_254), .ZN(n_257_21_54));
   INV_X1 i_257_21_56 (.A(CPU_Bus[11]), .ZN(n_257_21_55));
   NAND2_X1 i_257_21_57 (.A1(n_257_21_57), .A2(n_257_21_95), .ZN(n_257_21_56));
   INV_X1 i_257_21_58 (.A(CPU_Bus[10]), .ZN(n_257_21_57));
   NAND3_X1 i_257_21_59 (.A1(n_257_21_61), .A2(n_257_21_59), .A3(n_255), 
      .ZN(n_257_21_58));
   NAND2_X1 i_257_21_60 (.A1(n_257_21_60), .A2(n_254), .ZN(n_257_21_59));
   INV_X1 i_257_21_61 (.A(CPU_Bus[13]), .ZN(n_257_21_60));
   NAND2_X1 i_257_21_62 (.A1(n_257_21_62), .A2(n_257_21_95), .ZN(n_257_21_61));
   INV_X1 i_257_21_63 (.A(CPU_Bus[12]), .ZN(n_257_21_62));
   NAND3_X1 i_257_21_64 (.A1(n_257_21_69), .A2(n_257_21_64), .A3(n_257_21_97), 
      .ZN(n_257_21_63));
   NAND3_X1 i_257_21_65 (.A1(n_257_21_67), .A2(n_257_21_65), .A3(n_255), 
      .ZN(n_257_21_64));
   NAND2_X1 i_257_21_66 (.A1(n_257_21_66), .A2(n_254), .ZN(n_257_21_65));
   INV_X1 i_257_21_67 (.A(CPU_Bus[9]), .ZN(n_257_21_66));
   NAND2_X1 i_257_21_68 (.A1(n_257_21_68), .A2(n_257_21_95), .ZN(n_257_21_67));
   INV_X1 i_257_21_69 (.A(CPU_Bus[8]), .ZN(n_257_21_68));
   NAND3_X1 i_257_21_70 (.A1(n_257_21_72), .A2(n_257_21_70), .A3(n_257_21_96), 
      .ZN(n_257_21_69));
   NAND2_X1 i_257_21_71 (.A1(n_257_21_71), .A2(n_254), .ZN(n_257_21_70));
   INV_X1 i_257_21_72 (.A(CPU_Bus[7]), .ZN(n_257_21_71));
   NAND2_X1 i_257_21_73 (.A1(n_257_21_73), .A2(n_257_21_95), .ZN(n_257_21_72));
   INV_X1 i_257_21_74 (.A(CPU_Bus[6]), .ZN(n_257_21_73));
   NAND3_X1 i_257_21_75 (.A1(n_257_21_86), .A2(n_257_21_98), .A3(n_257_21_75), 
      .ZN(n_257_21_74));
   NAND3_X1 i_257_21_76 (.A1(n_257_21_81), .A2(n_257_21_76), .A3(n_256), 
      .ZN(n_257_21_75));
   NAND3_X1 i_257_21_77 (.A1(n_257_21_79), .A2(n_257_21_77), .A3(n_257_21_96), 
      .ZN(n_257_21_76));
   NAND2_X1 i_257_21_78 (.A1(n_257_21_78), .A2(n_254), .ZN(n_257_21_77));
   INV_X1 i_257_21_79 (.A(CPU_Bus[3]), .ZN(n_257_21_78));
   NAND2_X1 i_257_21_80 (.A1(n_257_21_80), .A2(n_257_21_95), .ZN(n_257_21_79));
   INV_X1 i_257_21_81 (.A(CPU_Bus[2]), .ZN(n_257_21_80));
   NAND3_X1 i_257_21_82 (.A1(n_257_21_84), .A2(n_257_21_82), .A3(n_255), 
      .ZN(n_257_21_81));
   NAND2_X1 i_257_21_83 (.A1(n_257_21_83), .A2(n_254), .ZN(n_257_21_82));
   INV_X1 i_257_21_84 (.A(CPU_Bus[5]), .ZN(n_257_21_83));
   NAND2_X1 i_257_21_85 (.A1(n_257_21_85), .A2(n_257_21_95), .ZN(n_257_21_84));
   INV_X1 i_257_21_86 (.A(CPU_Bus[4]), .ZN(n_257_21_85));
   NAND3_X1 i_257_21_87 (.A1(n_257_21_92), .A2(n_257_21_97), .A3(n_257_21_87), 
      .ZN(n_257_21_86));
   NAND3_X1 i_257_21_88 (.A1(n_257_21_90), .A2(n_257_21_88), .A3(n_255), 
      .ZN(n_257_21_87));
   NAND2_X1 i_257_21_89 (.A1(n_257_21_89), .A2(n_254), .ZN(n_257_21_88));
   INV_X1 i_257_21_90 (.A(CPU_Bus[1]), .ZN(n_257_21_89));
   NAND2_X1 i_257_21_91 (.A1(n_257_21_91), .A2(n_257_21_95), .ZN(n_257_21_90));
   INV_X1 i_257_21_92 (.A(CPU_Bus[0]), .ZN(n_257_21_91));
   OAI211_X1 i_257_21_93 (.A(n_257_21_93), .B(n_257_21_96), .C1(n_257_21_95), 
      .C2(CPU_Bus[31]), .ZN(n_257_21_92));
   NAND2_X1 i_257_21_94 (.A1(n_257_21_94), .A2(n_257_21_95), .ZN(n_257_21_93));
   INV_X1 i_257_21_95 (.A(CPU_Bus[30]), .ZN(n_257_21_94));
   INV_X1 i_257_21_96 (.A(n_254), .ZN(n_257_21_95));
   INV_X1 i_257_21_97 (.A(n_255), .ZN(n_257_21_96));
   INV_X1 i_257_21_98 (.A(n_256), .ZN(n_257_21_97));
   INV_X1 i_257_21_99 (.A(n_257), .ZN(n_257_21_98));
   INV_X1 i_257_22_0 (.A(n_257_22_0), .ZN(n_257_68));
   NAND2_X1 i_257_22_1 (.A1(n_257_22_49), .A2(n_257_22_1), .ZN(n_257_22_0));
   NAND3_X1 i_257_22_2 (.A1(n_257_22_25), .A2(n_257_22_2), .A3(n_257_22_48), 
      .ZN(n_257_22_1));
   NAND3_X1 i_257_22_3 (.A1(n_257_22_14), .A2(n_257_22_3), .A3(n_257), .ZN(
      n_257_22_2));
   NAND3_X1 i_257_22_4 (.A1(n_257_22_9), .A2(n_257_22_4), .A3(n_257_22_85), 
      .ZN(n_257_22_3));
   NAND3_X1 i_257_22_5 (.A1(n_257_22_7), .A2(n_257_22_5), .A3(n_257_22_96), 
      .ZN(n_257_22_4));
   NAND2_X1 i_257_22_6 (.A1(n_257_22_6), .A2(n_257_22_95), .ZN(n_257_22_5));
   INV_X1 i_257_22_7 (.A(CPU_Bus[21]), .ZN(n_257_22_6));
   NAND2_X1 i_257_22_8 (.A1(n_257_22_8), .A2(n_254), .ZN(n_257_22_7));
   INV_X1 i_257_22_9 (.A(CPU_Bus[22]), .ZN(n_257_22_8));
   NAND3_X1 i_257_22_10 (.A1(n_257_22_12), .A2(n_257_22_10), .A3(n_255), 
      .ZN(n_257_22_9));
   NAND2_X1 i_257_22_11 (.A1(n_257_22_11), .A2(n_257_22_95), .ZN(n_257_22_10));
   INV_X1 i_257_22_12 (.A(CPU_Bus[23]), .ZN(n_257_22_11));
   NAND2_X1 i_257_22_13 (.A1(n_257_22_13), .A2(n_254), .ZN(n_257_22_12));
   INV_X1 i_257_22_14 (.A(CPU_Bus[24]), .ZN(n_257_22_13));
   NAND3_X1 i_257_22_15 (.A1(n_257_22_20), .A2(n_257_22_15), .A3(n_256), 
      .ZN(n_257_22_14));
   NAND3_X1 i_257_22_16 (.A1(n_257_22_18), .A2(n_257_22_16), .A3(n_257_22_96), 
      .ZN(n_257_22_15));
   NAND2_X1 i_257_22_17 (.A1(n_257_22_17), .A2(n_257_22_95), .ZN(n_257_22_16));
   INV_X1 i_257_22_18 (.A(CPU_Bus[25]), .ZN(n_257_22_17));
   NAND2_X1 i_257_22_19 (.A1(n_257_22_19), .A2(n_254), .ZN(n_257_22_18));
   INV_X1 i_257_22_20 (.A(CPU_Bus[26]), .ZN(n_257_22_19));
   NAND3_X1 i_257_22_21 (.A1(n_257_22_23), .A2(n_257_22_21), .A3(n_255), 
      .ZN(n_257_22_20));
   NAND2_X1 i_257_22_22 (.A1(n_257_22_22), .A2(n_257_22_95), .ZN(n_257_22_21));
   INV_X1 i_257_22_23 (.A(CPU_Bus[27]), .ZN(n_257_22_22));
   NAND2_X1 i_257_22_24 (.A1(n_257_22_24), .A2(n_254), .ZN(n_257_22_23));
   INV_X1 i_257_22_25 (.A(CPU_Bus[28]), .ZN(n_257_22_24));
   NAND3_X1 i_257_22_26 (.A1(n_257_22_37), .A2(n_257_22_26), .A3(n_257_22_97), 
      .ZN(n_257_22_25));
   NAND3_X1 i_257_22_27 (.A1(n_257_22_32), .A2(n_257_22_27), .A3(n_256), 
      .ZN(n_257_22_26));
   NAND3_X1 i_257_22_28 (.A1(n_257_22_30), .A2(n_257_22_28), .A3(n_255), 
      .ZN(n_257_22_27));
   NAND2_X1 i_257_22_29 (.A1(n_257_22_29), .A2(n_254), .ZN(n_257_22_28));
   INV_X1 i_257_22_30 (.A(CPU_Bus[20]), .ZN(n_257_22_29));
   NAND2_X1 i_257_22_31 (.A1(n_257_22_31), .A2(n_257_22_95), .ZN(n_257_22_30));
   INV_X1 i_257_22_32 (.A(CPU_Bus[19]), .ZN(n_257_22_31));
   NAND3_X1 i_257_22_33 (.A1(n_257_22_35), .A2(n_257_22_33), .A3(n_257_22_96), 
      .ZN(n_257_22_32));
   NAND2_X1 i_257_22_34 (.A1(n_257_22_34), .A2(n_257_22_95), .ZN(n_257_22_33));
   INV_X1 i_257_22_35 (.A(CPU_Bus[17]), .ZN(n_257_22_34));
   NAND2_X1 i_257_22_36 (.A1(n_257_22_36), .A2(n_254), .ZN(n_257_22_35));
   INV_X1 i_257_22_37 (.A(CPU_Bus[18]), .ZN(n_257_22_36));
   NAND3_X1 i_257_22_38 (.A1(n_257_22_43), .A2(n_257_22_38), .A3(n_257_22_85), 
      .ZN(n_257_22_37));
   NAND3_X1 i_257_22_39 (.A1(n_257_22_41), .A2(n_257_22_39), .A3(n_255), 
      .ZN(n_257_22_38));
   NAND2_X1 i_257_22_40 (.A1(n_257_22_40), .A2(n_254), .ZN(n_257_22_39));
   INV_X1 i_257_22_41 (.A(CPU_Bus[16]), .ZN(n_257_22_40));
   NAND2_X1 i_257_22_42 (.A1(n_257_22_42), .A2(n_257_22_95), .ZN(n_257_22_41));
   INV_X1 i_257_22_43 (.A(CPU_Bus[15]), .ZN(n_257_22_42));
   NAND3_X1 i_257_22_44 (.A1(n_257_22_46), .A2(n_257_22_44), .A3(n_257_22_96), 
      .ZN(n_257_22_43));
   NAND2_X1 i_257_22_45 (.A1(n_257_22_45), .A2(n_257_22_95), .ZN(n_257_22_44));
   INV_X1 i_257_22_46 (.A(CPU_Bus[13]), .ZN(n_257_22_45));
   NAND2_X1 i_257_22_47 (.A1(n_257_22_47), .A2(n_254), .ZN(n_257_22_46));
   INV_X1 i_257_22_48 (.A(CPU_Bus[14]), .ZN(n_257_22_47));
   INV_X1 i_257_22_49 (.A(n_258), .ZN(n_257_22_48));
   NAND3_X1 i_257_22_50 (.A1(n_257_22_73), .A2(n_257_22_50), .A3(n_258), 
      .ZN(n_257_22_49));
   NAND3_X1 i_257_22_51 (.A1(n_257_22_62), .A2(n_257_22_51), .A3(n_257), 
      .ZN(n_257_22_50));
   NAND3_X1 i_257_22_52 (.A1(n_257_22_57), .A2(n_257_22_52), .A3(n_257_22_85), 
      .ZN(n_257_22_51));
   NAND3_X1 i_257_22_53 (.A1(n_257_22_55), .A2(n_257_22_53), .A3(n_257_22_96), 
      .ZN(n_257_22_52));
   NAND2_X1 i_257_22_54 (.A1(n_257_22_54), .A2(n_257_22_95), .ZN(n_257_22_53));
   INV_X1 i_257_22_55 (.A(CPU_Bus[5]), .ZN(n_257_22_54));
   NAND2_X1 i_257_22_56 (.A1(n_257_22_56), .A2(n_254), .ZN(n_257_22_55));
   INV_X1 i_257_22_57 (.A(CPU_Bus[6]), .ZN(n_257_22_56));
   NAND3_X1 i_257_22_58 (.A1(n_257_22_60), .A2(n_257_22_58), .A3(n_255), 
      .ZN(n_257_22_57));
   NAND2_X1 i_257_22_59 (.A1(n_257_22_59), .A2(n_254), .ZN(n_257_22_58));
   INV_X1 i_257_22_60 (.A(CPU_Bus[8]), .ZN(n_257_22_59));
   NAND2_X1 i_257_22_61 (.A1(n_257_22_61), .A2(n_257_22_95), .ZN(n_257_22_60));
   INV_X1 i_257_22_62 (.A(CPU_Bus[7]), .ZN(n_257_22_61));
   NAND3_X1 i_257_22_63 (.A1(n_257_22_68), .A2(n_257_22_63), .A3(n_256), 
      .ZN(n_257_22_62));
   NAND3_X1 i_257_22_64 (.A1(n_257_22_66), .A2(n_257_22_64), .A3(n_257_22_96), 
      .ZN(n_257_22_63));
   NAND2_X1 i_257_22_65 (.A1(n_257_22_65), .A2(n_254), .ZN(n_257_22_64));
   INV_X1 i_257_22_66 (.A(CPU_Bus[10]), .ZN(n_257_22_65));
   NAND2_X1 i_257_22_67 (.A1(n_257_22_67), .A2(n_257_22_95), .ZN(n_257_22_66));
   INV_X1 i_257_22_68 (.A(CPU_Bus[9]), .ZN(n_257_22_67));
   NAND3_X1 i_257_22_69 (.A1(n_257_22_71), .A2(n_257_22_69), .A3(n_255), 
      .ZN(n_257_22_68));
   NAND2_X1 i_257_22_70 (.A1(n_257_22_70), .A2(n_257_22_95), .ZN(n_257_22_69));
   INV_X1 i_257_22_71 (.A(CPU_Bus[11]), .ZN(n_257_22_70));
   NAND2_X1 i_257_22_72 (.A1(n_257_22_72), .A2(n_254), .ZN(n_257_22_71));
   INV_X1 i_257_22_73 (.A(CPU_Bus[12]), .ZN(n_257_22_72));
   NAND3_X1 i_257_22_74 (.A1(n_257_22_86), .A2(n_257_22_74), .A3(n_257_22_97), 
      .ZN(n_257_22_73));
   NAND3_X1 i_257_22_75 (.A1(n_257_22_80), .A2(n_257_22_75), .A3(n_257_22_85), 
      .ZN(n_257_22_74));
   NAND3_X1 i_257_22_76 (.A1(n_257_22_78), .A2(n_257_22_76), .A3(n_257_22_96), 
      .ZN(n_257_22_75));
   NAND2_X1 i_257_22_77 (.A1(n_257_22_77), .A2(n_254), .ZN(n_257_22_76));
   INV_X1 i_257_22_78 (.A(CPU_Bus[30]), .ZN(n_257_22_77));
   NAND2_X1 i_257_22_79 (.A1(n_257_22_79), .A2(n_257_22_95), .ZN(n_257_22_78));
   INV_X1 i_257_22_80 (.A(CPU_Bus[29]), .ZN(n_257_22_79));
   NAND3_X1 i_257_22_81 (.A1(n_257_22_83), .A2(n_257_22_81), .A3(n_255), 
      .ZN(n_257_22_80));
   NAND2_X1 i_257_22_82 (.A1(n_257_22_82), .A2(n_254), .ZN(n_257_22_81));
   INV_X1 i_257_22_83 (.A(CPU_Bus[0]), .ZN(n_257_22_82));
   NAND2_X1 i_257_22_84 (.A1(n_257_22_84), .A2(n_257_22_95), .ZN(n_257_22_83));
   INV_X1 i_257_22_85 (.A(CPU_Bus[31]), .ZN(n_257_22_84));
   INV_X1 i_257_22_86 (.A(n_256), .ZN(n_257_22_85));
   NAND3_X1 i_257_22_87 (.A1(n_257_22_92), .A2(n_257_22_87), .A3(n_256), 
      .ZN(n_257_22_86));
   NAND3_X1 i_257_22_88 (.A1(n_257_22_90), .A2(n_257_22_88), .A3(n_255), 
      .ZN(n_257_22_87));
   NAND2_X1 i_257_22_89 (.A1(n_257_22_89), .A2(n_257_22_95), .ZN(n_257_22_88));
   INV_X1 i_257_22_90 (.A(CPU_Bus[3]), .ZN(n_257_22_89));
   NAND2_X1 i_257_22_91 (.A1(n_257_22_91), .A2(n_254), .ZN(n_257_22_90));
   INV_X1 i_257_22_92 (.A(CPU_Bus[4]), .ZN(n_257_22_91));
   OAI211_X1 i_257_22_93 (.A(n_257_22_93), .B(n_257_22_96), .C1(n_257_22_95), 
      .C2(CPU_Bus[2]), .ZN(n_257_22_92));
   NAND2_X1 i_257_22_94 (.A1(n_257_22_94), .A2(n_257_22_95), .ZN(n_257_22_93));
   INV_X1 i_257_22_95 (.A(CPU_Bus[1]), .ZN(n_257_22_94));
   INV_X1 i_257_22_96 (.A(n_254), .ZN(n_257_22_95));
   INV_X1 i_257_22_97 (.A(n_255), .ZN(n_257_22_96));
   INV_X1 i_257_22_98 (.A(n_257), .ZN(n_257_22_97));
   datapath__1_344 i_257_23 (.PacketSize(PacketSize), .p_0({n_257_74, uc_155, 
      uc_156, uc_157, uc_158, uc_159, uc_160, uc_161, uc_162, uc_163, uc_164, 
      uc_165, uc_166, uc_167, uc_168, uc_169, uc_170, uc_171, uc_172, uc_173, 
      uc_174, uc_175, uc_176, uc_177, uc_178, uc_179, n_257_73, n_257_72, 
      n_257_71, n_257_70, n_257_69, uc_180}));
   datapath__1_345 i_257_24 (.p_0({uc_181, uc_182, uc_183, uc_184, uc_185, 
      uc_186, uc_187, uc_188, uc_189, uc_190, uc_191, uc_192, uc_193, uc_194, 
      uc_195, uc_196, uc_197, uc_198, uc_199, uc_200, uc_201, uc_202, uc_203, 
      uc_204, uc_205, n_257_74, n_257_73, n_257_72, n_257_71, n_257_70, n_257_69, 
      n_151}), .p_1({n_257_106, n_257_105, n_257_104, n_257_103, n_257_102, 
      n_257_101, n_257_100, n_257_99, n_257_98, n_257_97, n_257_96, n_257_95, 
      n_257_94, n_257_93, n_257_92, n_257_91, n_257_90, n_257_89, n_257_88, 
      n_257_87, n_257_86, n_257_85, n_257_84, n_257_83, n_257_82, n_257_81, 
      n_257_80, n_257_79, n_257_78, n_257_77, n_257_76, n_257_75}));
   INV_X1 i_257_25_0 (.A(n_254), .ZN(n_257_25_0));
   NAND2_X1 i_257_25_1 (.A1(n_257_25_0), .A2(n_255), .ZN(n_257_25_1));
   INV_X1 i_257_25_2 (.A(n_256), .ZN(n_257_25_2));
   NOR2_X1 i_257_25_3 (.A1(n_257_25_1), .A2(n_257_25_2), .ZN(n_257_25_3));
   NAND2_X1 i_257_25_4 (.A1(n_257_25_3), .A2(n_257), .ZN(n_257_25_4));
   INV_X1 i_257_25_5 (.A(n_258), .ZN(n_257_25_5));
   NOR2_X1 i_257_25_6 (.A1(n_257_25_4), .A2(n_257_25_5), .ZN(n_257_25_6));
   NAND2_X1 i_257_25_7 (.A1(CPU_Bus[10]), .A2(n_257_25_6), .ZN(n_257_25_7));
   INV_X1 i_257_25_8 (.A(n_255), .ZN(n_257_25_8));
   NAND2_X1 i_257_25_9 (.A1(n_257_25_0), .A2(n_257_25_8), .ZN(n_257_25_9));
   NOR2_X1 i_257_25_10 (.A1(n_257_25_9), .A2(n_257_25_2), .ZN(n_257_25_10));
   NAND2_X1 i_257_25_11 (.A1(n_257_25_10), .A2(n_257), .ZN(n_257_25_11));
   NOR2_X1 i_257_25_12 (.A1(n_257_25_11), .A2(n_257_25_5), .ZN(n_257_25_12));
   NAND2_X1 i_257_25_13 (.A1(CPU_Bus[8]), .A2(n_257_25_12), .ZN(n_257_25_13));
   NAND2_X1 i_257_25_14 (.A1(n_257_25_7), .A2(n_257_25_13), .ZN(n_257_25_14));
   NOR2_X1 i_257_25_15 (.A1(n_257_25_1), .A2(n_256), .ZN(n_257_25_15));
   NAND2_X1 i_257_25_16 (.A1(n_257_25_15), .A2(n_257), .ZN(n_257_25_16));
   NOR2_X1 i_257_25_17 (.A1(n_257_25_16), .A2(n_257_25_5), .ZN(n_257_25_17));
   NAND2_X1 i_257_25_18 (.A1(CPU_Bus[6]), .A2(n_257_25_17), .ZN(n_257_25_18));
   NOR2_X1 i_257_25_19 (.A1(n_257_25_9), .A2(n_256), .ZN(n_257_25_19));
   NAND2_X1 i_257_25_20 (.A1(n_257_25_19), .A2(n_257), .ZN(n_257_25_20));
   NOR2_X1 i_257_25_21 (.A1(n_257_25_20), .A2(n_257_25_5), .ZN(n_257_25_21));
   NAND2_X1 i_257_25_22 (.A1(CPU_Bus[4]), .A2(n_257_25_21), .ZN(n_257_25_22));
   NAND2_X1 i_257_25_23 (.A1(n_257_25_18), .A2(n_257_25_22), .ZN(n_257_25_23));
   NOR2_X1 i_257_25_24 (.A1(n_257_25_14), .A2(n_257_25_23), .ZN(n_257_25_24));
   INV_X1 i_257_25_25 (.A(n_257), .ZN(n_257_25_25));
   NAND2_X1 i_257_25_26 (.A1(n_257_25_3), .A2(n_257_25_25), .ZN(n_257_25_26));
   NOR2_X1 i_257_25_27 (.A1(n_257_25_26), .A2(n_257_25_5), .ZN(n_257_25_27));
   NAND2_X1 i_257_25_28 (.A1(CPU_Bus[2]), .A2(n_257_25_27), .ZN(n_257_25_28));
   NAND2_X1 i_257_25_29 (.A1(n_257_25_10), .A2(n_257_25_25), .ZN(n_257_25_29));
   NOR2_X1 i_257_25_30 (.A1(n_257_25_29), .A2(n_257_25_5), .ZN(n_257_25_30));
   NAND2_X1 i_257_25_31 (.A1(CPU_Bus[0]), .A2(n_257_25_30), .ZN(n_257_25_31));
   NAND2_X1 i_257_25_32 (.A1(n_257_25_28), .A2(n_257_25_31), .ZN(n_257_25_32));
   NAND2_X1 i_257_25_33 (.A1(n_257_25_15), .A2(n_257_25_25), .ZN(n_257_25_33));
   NOR2_X1 i_257_25_34 (.A1(n_257_25_33), .A2(n_257_25_5), .ZN(n_257_25_34));
   NAND2_X1 i_257_25_35 (.A1(CPU_Bus[30]), .A2(n_257_25_34), .ZN(n_257_25_35));
   NAND2_X1 i_257_25_36 (.A1(n_257_25_19), .A2(n_257_25_25), .ZN(n_257_25_36));
   NOR2_X1 i_257_25_37 (.A1(n_257_25_36), .A2(n_257_25_5), .ZN(n_257_25_37));
   NAND2_X1 i_257_25_38 (.A1(CPU_Bus[28]), .A2(n_257_25_37), .ZN(n_257_25_38));
   NAND2_X1 i_257_25_39 (.A1(n_257_25_35), .A2(n_257_25_38), .ZN(n_257_25_39));
   NOR2_X1 i_257_25_40 (.A1(n_257_25_32), .A2(n_257_25_39), .ZN(n_257_25_40));
   NAND2_X1 i_257_25_41 (.A1(n_257_25_24), .A2(n_257_25_40), .ZN(n_257_25_41));
   NOR2_X1 i_257_25_42 (.A1(n_257_25_4), .A2(n_258), .ZN(n_257_25_42));
   NAND2_X1 i_257_25_43 (.A1(CPU_Bus[26]), .A2(n_257_25_42), .ZN(n_257_25_43));
   NOR2_X1 i_257_25_44 (.A1(n_257_25_11), .A2(n_258), .ZN(n_257_25_44));
   NAND2_X1 i_257_25_45 (.A1(CPU_Bus[24]), .A2(n_257_25_44), .ZN(n_257_25_45));
   NAND2_X1 i_257_25_46 (.A1(n_257_25_43), .A2(n_257_25_45), .ZN(n_257_25_46));
   NOR2_X1 i_257_25_47 (.A1(n_257_25_16), .A2(n_258), .ZN(n_257_25_47));
   NAND2_X1 i_257_25_48 (.A1(CPU_Bus[22]), .A2(n_257_25_47), .ZN(n_257_25_48));
   NOR2_X1 i_257_25_49 (.A1(n_257_25_20), .A2(n_258), .ZN(n_257_25_49));
   NAND2_X1 i_257_25_50 (.A1(CPU_Bus[20]), .A2(n_257_25_49), .ZN(n_257_25_50));
   NAND2_X1 i_257_25_51 (.A1(n_257_25_48), .A2(n_257_25_50), .ZN(n_257_25_51));
   NOR2_X1 i_257_25_52 (.A1(n_257_25_46), .A2(n_257_25_51), .ZN(n_257_25_52));
   NOR2_X1 i_257_25_53 (.A1(n_257_25_26), .A2(n_258), .ZN(n_257_25_53));
   NAND2_X1 i_257_25_54 (.A1(CPU_Bus[18]), .A2(n_257_25_53), .ZN(n_257_25_54));
   NOR2_X1 i_257_25_55 (.A1(n_257_25_29), .A2(n_258), .ZN(n_257_25_55));
   NAND2_X1 i_257_25_56 (.A1(CPU_Bus[16]), .A2(n_257_25_55), .ZN(n_257_25_56));
   NAND2_X1 i_257_25_57 (.A1(n_257_25_54), .A2(n_257_25_56), .ZN(n_257_25_57));
   NOR2_X1 i_257_25_58 (.A1(n_257_25_33), .A2(n_258), .ZN(n_257_25_58));
   NAND2_X1 i_257_25_59 (.A1(CPU_Bus[14]), .A2(n_257_25_58), .ZN(n_257_25_59));
   NOR2_X1 i_257_25_60 (.A1(n_257_25_36), .A2(n_258), .ZN(n_257_25_60));
   NAND2_X1 i_257_25_61 (.A1(CPU_Bus[12]), .A2(n_257_25_60), .ZN(n_257_25_61));
   NAND2_X1 i_257_25_62 (.A1(n_257_25_59), .A2(n_257_25_61), .ZN(n_257_25_62));
   NOR2_X1 i_257_25_63 (.A1(n_257_25_57), .A2(n_257_25_62), .ZN(n_257_25_63));
   NAND2_X1 i_257_25_64 (.A1(n_257_25_52), .A2(n_257_25_63), .ZN(n_257_25_64));
   NOR2_X1 i_257_25_65 (.A1(n_257_25_41), .A2(n_257_25_64), .ZN(n_257_25_65));
   NAND2_X1 i_257_25_66 (.A1(n_257_25_8), .A2(n_254), .ZN(n_257_25_66));
   NOR2_X1 i_257_25_67 (.A1(n_257_25_66), .A2(n_257_25_2), .ZN(n_257_25_67));
   NAND2_X1 i_257_25_68 (.A1(n_257_25_67), .A2(n_257), .ZN(n_257_25_68));
   NOR2_X1 i_257_25_69 (.A1(n_257_25_68), .A2(n_257_25_5), .ZN(n_257_25_69));
   NAND2_X1 i_257_25_70 (.A1(CPU_Bus[9]), .A2(n_257_25_69), .ZN(n_257_25_70));
   NOR2_X1 i_257_25_71 (.A1(n_257_25_66), .A2(n_256), .ZN(n_257_25_71));
   NAND2_X1 i_257_25_72 (.A1(n_257_25_71), .A2(n_257), .ZN(n_257_25_72));
   NOR2_X1 i_257_25_73 (.A1(n_257_25_72), .A2(n_257_25_5), .ZN(n_257_25_73));
   NAND2_X1 i_257_25_74 (.A1(CPU_Bus[5]), .A2(n_257_25_73), .ZN(n_257_25_74));
   NAND2_X1 i_257_25_75 (.A1(n_257_25_70), .A2(n_257_25_74), .ZN(n_257_25_75));
   NAND2_X1 i_257_25_76 (.A1(n_257_25_67), .A2(n_257_25_25), .ZN(n_257_25_76));
   NOR2_X1 i_257_25_77 (.A1(n_257_25_76), .A2(n_257_25_5), .ZN(n_257_25_77));
   NAND2_X1 i_257_25_78 (.A1(CPU_Bus[1]), .A2(n_257_25_77), .ZN(n_257_25_78));
   NAND2_X1 i_257_25_79 (.A1(n_257_25_71), .A2(n_257_25_25), .ZN(n_257_25_79));
   NOR2_X1 i_257_25_80 (.A1(n_257_25_79), .A2(n_257_25_5), .ZN(n_257_25_80));
   NAND2_X1 i_257_25_81 (.A1(CPU_Bus[29]), .A2(n_257_25_80), .ZN(n_257_25_81));
   NAND2_X1 i_257_25_82 (.A1(n_257_25_78), .A2(n_257_25_81), .ZN(n_257_25_82));
   NOR2_X1 i_257_25_83 (.A1(n_257_25_75), .A2(n_257_25_82), .ZN(n_257_25_83));
   NOR2_X1 i_257_25_84 (.A1(n_257_25_68), .A2(n_258), .ZN(n_257_25_84));
   NAND2_X1 i_257_25_85 (.A1(CPU_Bus[25]), .A2(n_257_25_84), .ZN(n_257_25_85));
   NOR2_X1 i_257_25_86 (.A1(n_257_25_72), .A2(n_258), .ZN(n_257_25_86));
   NAND2_X1 i_257_25_87 (.A1(CPU_Bus[21]), .A2(n_257_25_86), .ZN(n_257_25_87));
   NAND2_X1 i_257_25_88 (.A1(n_257_25_85), .A2(n_257_25_87), .ZN(n_257_25_88));
   NOR2_X1 i_257_25_89 (.A1(n_257_25_76), .A2(n_258), .ZN(n_257_25_89));
   NAND2_X1 i_257_25_90 (.A1(CPU_Bus[17]), .A2(n_257_25_89), .ZN(n_257_25_90));
   NOR2_X1 i_257_25_91 (.A1(n_257_25_79), .A2(n_258), .ZN(n_257_25_91));
   NAND2_X1 i_257_25_92 (.A1(CPU_Bus[13]), .A2(n_257_25_91), .ZN(n_257_25_92));
   NAND2_X1 i_257_25_93 (.A1(n_257_25_90), .A2(n_257_25_92), .ZN(n_257_25_93));
   NOR2_X1 i_257_25_94 (.A1(n_257_25_88), .A2(n_257_25_93), .ZN(n_257_25_94));
   NAND2_X1 i_257_25_95 (.A1(n_257_25_83), .A2(n_257_25_94), .ZN(n_257_25_95));
   NAND2_X1 i_257_25_96 (.A1(n_254), .A2(n_255), .ZN(n_257_25_96));
   NOR2_X1 i_257_25_97 (.A1(n_257_25_96), .A2(n_257_25_2), .ZN(n_257_25_97));
   NAND2_X1 i_257_25_98 (.A1(n_257_25_97), .A2(n_257), .ZN(n_257_25_98));
   NOR2_X1 i_257_25_99 (.A1(n_257_25_98), .A2(n_257_25_5), .ZN(n_257_25_99));
   NAND2_X1 i_257_25_100 (.A1(CPU_Bus[11]), .A2(n_257_25_99), .ZN(n_257_25_100));
   NOR2_X1 i_257_25_101 (.A1(n_257_25_96), .A2(n_256), .ZN(n_257_25_101));
   NAND2_X1 i_257_25_102 (.A1(n_257_25_101), .A2(n_257), .ZN(n_257_25_102));
   NOR2_X1 i_257_25_103 (.A1(n_257_25_102), .A2(n_257_25_5), .ZN(n_257_25_103));
   NAND2_X1 i_257_25_104 (.A1(CPU_Bus[7]), .A2(n_257_25_103), .ZN(n_257_25_104));
   NAND2_X1 i_257_25_105 (.A1(n_257_25_100), .A2(n_257_25_104), .ZN(n_257_25_105));
   NAND2_X1 i_257_25_106 (.A1(n_257_25_97), .A2(n_257_25_25), .ZN(n_257_25_106));
   NOR2_X1 i_257_25_107 (.A1(n_257_25_106), .A2(n_257_25_5), .ZN(n_257_25_107));
   NAND2_X1 i_257_25_108 (.A1(CPU_Bus[3]), .A2(n_257_25_107), .ZN(n_257_25_108));
   NAND2_X1 i_257_25_109 (.A1(n_257_25_101), .A2(n_257_25_25), .ZN(n_257_25_109));
   NOR2_X1 i_257_25_110 (.A1(n_257_25_109), .A2(n_257_25_5), .ZN(n_257_25_110));
   NAND2_X1 i_257_25_111 (.A1(CPU_Bus[31]), .A2(n_257_25_110), .ZN(n_257_25_111));
   NAND2_X1 i_257_25_112 (.A1(n_257_25_108), .A2(n_257_25_111), .ZN(n_257_25_112));
   NOR2_X1 i_257_25_113 (.A1(n_257_25_105), .A2(n_257_25_112), .ZN(n_257_25_113));
   NOR2_X1 i_257_25_114 (.A1(n_257_25_98), .A2(n_258), .ZN(n_257_25_114));
   NAND2_X1 i_257_25_115 (.A1(CPU_Bus[27]), .A2(n_257_25_114), .ZN(n_257_25_115));
   NOR2_X1 i_257_25_116 (.A1(n_257_25_102), .A2(n_258), .ZN(n_257_25_116));
   NAND2_X1 i_257_25_117 (.A1(CPU_Bus[23]), .A2(n_257_25_116), .ZN(n_257_25_117));
   NAND2_X1 i_257_25_118 (.A1(n_257_25_115), .A2(n_257_25_117), .ZN(n_257_25_118));
   NOR2_X1 i_257_25_119 (.A1(n_257_25_106), .A2(n_258), .ZN(n_257_25_119));
   NAND2_X1 i_257_25_120 (.A1(CPU_Bus[19]), .A2(n_257_25_119), .ZN(n_257_25_120));
   NOR2_X1 i_257_25_121 (.A1(n_257_25_109), .A2(n_258), .ZN(n_257_25_121));
   NAND2_X1 i_257_25_122 (.A1(CPU_Bus[15]), .A2(n_257_25_121), .ZN(n_257_25_122));
   NAND2_X1 i_257_25_123 (.A1(n_257_25_120), .A2(n_257_25_122), .ZN(n_257_25_123));
   NOR2_X1 i_257_25_124 (.A1(n_257_25_118), .A2(n_257_25_123), .ZN(n_257_25_124));
   NAND2_X1 i_257_25_125 (.A1(n_257_25_113), .A2(n_257_25_124), .ZN(n_257_25_125));
   NOR2_X1 i_257_25_126 (.A1(n_257_25_95), .A2(n_257_25_125), .ZN(n_257_25_126));
   NAND2_X1 i_257_25_127 (.A1(n_257_25_65), .A2(n_257_25_126), .ZN(n_257_107));
   datapath__1_347 i_257_26 (.PacketSize({PacketSize[5], PacketSize[4], 
      PacketSize[3], PacketSize[2], PacketSize[1], 1'b0}), .p_0({n_257_112, 
      uc_206, uc_207, uc_208, uc_209, uc_210, uc_211, uc_212, uc_213, uc_214, 
      uc_215, uc_216, uc_217, uc_218, uc_219, uc_220, uc_221, uc_222, uc_223, 
      uc_224, uc_225, uc_226, uc_227, uc_228, uc_229, uc_230, n_257_111, 
      n_257_110, n_257_109, n_257_108, uc_231, uc_232}));
   datapath__1_348 i_257_27 (.p_0({uc_233, uc_234, uc_235, uc_236, uc_237, 
      uc_238, uc_239, uc_240, uc_241, uc_242, uc_243, uc_244, uc_245, uc_246, 
      uc_247, uc_248, uc_249, uc_250, uc_251, uc_252, uc_253, uc_254, uc_255, 
      uc_256, uc_257, n_257_112, n_257_111, n_257_110, n_257_109, n_257_108, 
      n_257_1091, PacketSize[0]}), .p_1({n_257_144, n_257_143, n_257_142, 
      n_257_141, n_257_140, n_257_139, n_257_138, n_257_137, n_257_136, 
      n_257_135, n_257_134, n_257_133, n_257_132, n_257_131, n_257_130, 
      n_257_129, n_257_128, n_257_127, n_257_126, n_257_125, n_257_124, 
      n_257_123, n_257_122, n_257_121, n_257_120, n_257_119, n_257_118, 
      n_257_117, n_257_116, n_257_115, n_257_114, n_257_113}));
   INV_X1 i_257_28_0 (.A(n_254), .ZN(n_257_28_0));
   NAND2_X1 i_257_28_1 (.A1(n_257_28_0), .A2(n_255), .ZN(n_257_28_1));
   INV_X1 i_257_28_2 (.A(n_256), .ZN(n_257_28_2));
   NOR2_X1 i_257_28_3 (.A1(n_257_28_1), .A2(n_257_28_2), .ZN(n_257_28_3));
   NAND2_X1 i_257_28_4 (.A1(n_257_28_3), .A2(n_257), .ZN(n_257_28_4));
   INV_X1 i_257_28_5 (.A(n_258), .ZN(n_257_28_5));
   NOR2_X1 i_257_28_6 (.A1(n_257_28_4), .A2(n_257_28_5), .ZN(n_257_28_6));
   NAND2_X1 i_257_28_7 (.A1(CPU_Bus[9]), .A2(n_257_28_6), .ZN(n_257_28_7));
   INV_X1 i_257_28_8 (.A(n_255), .ZN(n_257_28_8));
   NAND2_X1 i_257_28_9 (.A1(n_257_28_0), .A2(n_257_28_8), .ZN(n_257_28_9));
   NOR2_X1 i_257_28_10 (.A1(n_257_28_9), .A2(n_257_28_2), .ZN(n_257_28_10));
   NAND2_X1 i_257_28_11 (.A1(n_257_28_10), .A2(n_257), .ZN(n_257_28_11));
   NOR2_X1 i_257_28_12 (.A1(n_257_28_11), .A2(n_257_28_5), .ZN(n_257_28_12));
   NAND2_X1 i_257_28_13 (.A1(CPU_Bus[7]), .A2(n_257_28_12), .ZN(n_257_28_13));
   NAND2_X1 i_257_28_14 (.A1(n_257_28_7), .A2(n_257_28_13), .ZN(n_257_28_14));
   NOR2_X1 i_257_28_15 (.A1(n_257_28_1), .A2(n_256), .ZN(n_257_28_15));
   NAND2_X1 i_257_28_16 (.A1(n_257_28_15), .A2(n_257), .ZN(n_257_28_16));
   NOR2_X1 i_257_28_17 (.A1(n_257_28_16), .A2(n_257_28_5), .ZN(n_257_28_17));
   NAND2_X1 i_257_28_18 (.A1(CPU_Bus[5]), .A2(n_257_28_17), .ZN(n_257_28_18));
   NOR2_X1 i_257_28_19 (.A1(n_257_28_9), .A2(n_256), .ZN(n_257_28_19));
   NAND2_X1 i_257_28_20 (.A1(n_257_28_19), .A2(n_257), .ZN(n_257_28_20));
   NOR2_X1 i_257_28_21 (.A1(n_257_28_20), .A2(n_257_28_5), .ZN(n_257_28_21));
   NAND2_X1 i_257_28_22 (.A1(CPU_Bus[3]), .A2(n_257_28_21), .ZN(n_257_28_22));
   NAND2_X1 i_257_28_23 (.A1(n_257_28_18), .A2(n_257_28_22), .ZN(n_257_28_23));
   NOR2_X1 i_257_28_24 (.A1(n_257_28_14), .A2(n_257_28_23), .ZN(n_257_28_24));
   INV_X1 i_257_28_25 (.A(n_257), .ZN(n_257_28_25));
   NAND2_X1 i_257_28_26 (.A1(n_257_28_3), .A2(n_257_28_25), .ZN(n_257_28_26));
   NOR2_X1 i_257_28_27 (.A1(n_257_28_26), .A2(n_257_28_5), .ZN(n_257_28_27));
   NAND2_X1 i_257_28_28 (.A1(CPU_Bus[1]), .A2(n_257_28_27), .ZN(n_257_28_28));
   NAND2_X1 i_257_28_29 (.A1(n_257_28_10), .A2(n_257_28_25), .ZN(n_257_28_29));
   NOR2_X1 i_257_28_30 (.A1(n_257_28_29), .A2(n_257_28_5), .ZN(n_257_28_30));
   NAND2_X1 i_257_28_31 (.A1(CPU_Bus[31]), .A2(n_257_28_30), .ZN(n_257_28_31));
   NAND2_X1 i_257_28_32 (.A1(n_257_28_28), .A2(n_257_28_31), .ZN(n_257_28_32));
   NAND2_X1 i_257_28_33 (.A1(n_257_28_15), .A2(n_257_28_25), .ZN(n_257_28_33));
   NOR2_X1 i_257_28_34 (.A1(n_257_28_33), .A2(n_257_28_5), .ZN(n_257_28_34));
   NAND2_X1 i_257_28_35 (.A1(CPU_Bus[29]), .A2(n_257_28_34), .ZN(n_257_28_35));
   NAND2_X1 i_257_28_36 (.A1(n_257_28_19), .A2(n_257_28_25), .ZN(n_257_28_36));
   NOR2_X1 i_257_28_37 (.A1(n_257_28_36), .A2(n_257_28_5), .ZN(n_257_28_37));
   NAND2_X1 i_257_28_38 (.A1(CPU_Bus[27]), .A2(n_257_28_37), .ZN(n_257_28_38));
   NAND2_X1 i_257_28_39 (.A1(n_257_28_35), .A2(n_257_28_38), .ZN(n_257_28_39));
   NOR2_X1 i_257_28_40 (.A1(n_257_28_32), .A2(n_257_28_39), .ZN(n_257_28_40));
   NAND2_X1 i_257_28_41 (.A1(n_257_28_24), .A2(n_257_28_40), .ZN(n_257_28_41));
   NOR2_X1 i_257_28_42 (.A1(n_257_28_4), .A2(n_258), .ZN(n_257_28_42));
   NAND2_X1 i_257_28_43 (.A1(CPU_Bus[25]), .A2(n_257_28_42), .ZN(n_257_28_43));
   NOR2_X1 i_257_28_44 (.A1(n_257_28_11), .A2(n_258), .ZN(n_257_28_44));
   NAND2_X1 i_257_28_45 (.A1(CPU_Bus[23]), .A2(n_257_28_44), .ZN(n_257_28_45));
   NAND2_X1 i_257_28_46 (.A1(n_257_28_43), .A2(n_257_28_45), .ZN(n_257_28_46));
   NOR2_X1 i_257_28_47 (.A1(n_257_28_16), .A2(n_258), .ZN(n_257_28_47));
   NAND2_X1 i_257_28_48 (.A1(CPU_Bus[21]), .A2(n_257_28_47), .ZN(n_257_28_48));
   NOR2_X1 i_257_28_49 (.A1(n_257_28_20), .A2(n_258), .ZN(n_257_28_49));
   NAND2_X1 i_257_28_50 (.A1(CPU_Bus[19]), .A2(n_257_28_49), .ZN(n_257_28_50));
   NAND2_X1 i_257_28_51 (.A1(n_257_28_48), .A2(n_257_28_50), .ZN(n_257_28_51));
   NOR2_X1 i_257_28_52 (.A1(n_257_28_46), .A2(n_257_28_51), .ZN(n_257_28_52));
   NOR2_X1 i_257_28_53 (.A1(n_257_28_26), .A2(n_258), .ZN(n_257_28_53));
   NAND2_X1 i_257_28_54 (.A1(CPU_Bus[17]), .A2(n_257_28_53), .ZN(n_257_28_54));
   NOR2_X1 i_257_28_55 (.A1(n_257_28_29), .A2(n_258), .ZN(n_257_28_55));
   NAND2_X1 i_257_28_56 (.A1(CPU_Bus[15]), .A2(n_257_28_55), .ZN(n_257_28_56));
   NAND2_X1 i_257_28_57 (.A1(n_257_28_54), .A2(n_257_28_56), .ZN(n_257_28_57));
   NOR2_X1 i_257_28_58 (.A1(n_257_28_33), .A2(n_258), .ZN(n_257_28_58));
   NAND2_X1 i_257_28_59 (.A1(CPU_Bus[13]), .A2(n_257_28_58), .ZN(n_257_28_59));
   NOR2_X1 i_257_28_60 (.A1(n_257_28_36), .A2(n_258), .ZN(n_257_28_60));
   NAND2_X1 i_257_28_61 (.A1(CPU_Bus[11]), .A2(n_257_28_60), .ZN(n_257_28_61));
   NAND2_X1 i_257_28_62 (.A1(n_257_28_59), .A2(n_257_28_61), .ZN(n_257_28_62));
   NOR2_X1 i_257_28_63 (.A1(n_257_28_57), .A2(n_257_28_62), .ZN(n_257_28_63));
   NAND2_X1 i_257_28_64 (.A1(n_257_28_52), .A2(n_257_28_63), .ZN(n_257_28_64));
   NOR2_X1 i_257_28_65 (.A1(n_257_28_41), .A2(n_257_28_64), .ZN(n_257_28_65));
   NAND2_X1 i_257_28_66 (.A1(n_257_28_8), .A2(n_254), .ZN(n_257_28_66));
   NOR2_X1 i_257_28_67 (.A1(n_257_28_66), .A2(n_257_28_2), .ZN(n_257_28_67));
   NAND2_X1 i_257_28_68 (.A1(n_257_28_67), .A2(n_257), .ZN(n_257_28_68));
   NOR2_X1 i_257_28_69 (.A1(n_257_28_68), .A2(n_257_28_5), .ZN(n_257_28_69));
   NAND2_X1 i_257_28_70 (.A1(CPU_Bus[8]), .A2(n_257_28_69), .ZN(n_257_28_70));
   NOR2_X1 i_257_28_71 (.A1(n_257_28_66), .A2(n_256), .ZN(n_257_28_71));
   NAND2_X1 i_257_28_72 (.A1(n_257_28_71), .A2(n_257), .ZN(n_257_28_72));
   NOR2_X1 i_257_28_73 (.A1(n_257_28_72), .A2(n_257_28_5), .ZN(n_257_28_73));
   NAND2_X1 i_257_28_74 (.A1(CPU_Bus[4]), .A2(n_257_28_73), .ZN(n_257_28_74));
   NAND2_X1 i_257_28_75 (.A1(n_257_28_70), .A2(n_257_28_74), .ZN(n_257_28_75));
   NAND2_X1 i_257_28_76 (.A1(n_257_28_67), .A2(n_257_28_25), .ZN(n_257_28_76));
   NOR2_X1 i_257_28_77 (.A1(n_257_28_76), .A2(n_257_28_5), .ZN(n_257_28_77));
   NAND2_X1 i_257_28_78 (.A1(CPU_Bus[0]), .A2(n_257_28_77), .ZN(n_257_28_78));
   NAND2_X1 i_257_28_79 (.A1(n_257_28_71), .A2(n_257_28_25), .ZN(n_257_28_79));
   NOR2_X1 i_257_28_80 (.A1(n_257_28_79), .A2(n_257_28_5), .ZN(n_257_28_80));
   NAND2_X1 i_257_28_81 (.A1(CPU_Bus[28]), .A2(n_257_28_80), .ZN(n_257_28_81));
   NAND2_X1 i_257_28_82 (.A1(n_257_28_78), .A2(n_257_28_81), .ZN(n_257_28_82));
   NOR2_X1 i_257_28_83 (.A1(n_257_28_75), .A2(n_257_28_82), .ZN(n_257_28_83));
   NOR2_X1 i_257_28_84 (.A1(n_257_28_68), .A2(n_258), .ZN(n_257_28_84));
   NAND2_X1 i_257_28_85 (.A1(CPU_Bus[24]), .A2(n_257_28_84), .ZN(n_257_28_85));
   NOR2_X1 i_257_28_86 (.A1(n_257_28_72), .A2(n_258), .ZN(n_257_28_86));
   NAND2_X1 i_257_28_87 (.A1(CPU_Bus[20]), .A2(n_257_28_86), .ZN(n_257_28_87));
   NAND2_X1 i_257_28_88 (.A1(n_257_28_85), .A2(n_257_28_87), .ZN(n_257_28_88));
   NOR2_X1 i_257_28_89 (.A1(n_257_28_76), .A2(n_258), .ZN(n_257_28_89));
   NAND2_X1 i_257_28_90 (.A1(CPU_Bus[16]), .A2(n_257_28_89), .ZN(n_257_28_90));
   NOR2_X1 i_257_28_91 (.A1(n_257_28_79), .A2(n_258), .ZN(n_257_28_91));
   NAND2_X1 i_257_28_92 (.A1(CPU_Bus[12]), .A2(n_257_28_91), .ZN(n_257_28_92));
   NAND2_X1 i_257_28_93 (.A1(n_257_28_90), .A2(n_257_28_92), .ZN(n_257_28_93));
   NOR2_X1 i_257_28_94 (.A1(n_257_28_88), .A2(n_257_28_93), .ZN(n_257_28_94));
   NAND2_X1 i_257_28_95 (.A1(n_257_28_83), .A2(n_257_28_94), .ZN(n_257_28_95));
   NAND2_X1 i_257_28_96 (.A1(n_254), .A2(n_255), .ZN(n_257_28_96));
   NOR2_X1 i_257_28_97 (.A1(n_257_28_96), .A2(n_257_28_2), .ZN(n_257_28_97));
   NAND2_X1 i_257_28_98 (.A1(n_257_28_97), .A2(n_257), .ZN(n_257_28_98));
   NOR2_X1 i_257_28_99 (.A1(n_257_28_98), .A2(n_257_28_5), .ZN(n_257_28_99));
   NAND2_X1 i_257_28_100 (.A1(CPU_Bus[10]), .A2(n_257_28_99), .ZN(n_257_28_100));
   NOR2_X1 i_257_28_101 (.A1(n_257_28_96), .A2(n_256), .ZN(n_257_28_101));
   NAND2_X1 i_257_28_102 (.A1(n_257_28_101), .A2(n_257), .ZN(n_257_28_102));
   NOR2_X1 i_257_28_103 (.A1(n_257_28_102), .A2(n_257_28_5), .ZN(n_257_28_103));
   NAND2_X1 i_257_28_104 (.A1(CPU_Bus[6]), .A2(n_257_28_103), .ZN(n_257_28_104));
   NAND2_X1 i_257_28_105 (.A1(n_257_28_100), .A2(n_257_28_104), .ZN(n_257_28_105));
   NAND2_X1 i_257_28_106 (.A1(n_257_28_97), .A2(n_257_28_25), .ZN(n_257_28_106));
   NOR2_X1 i_257_28_107 (.A1(n_257_28_106), .A2(n_257_28_5), .ZN(n_257_28_107));
   NAND2_X1 i_257_28_108 (.A1(CPU_Bus[2]), .A2(n_257_28_107), .ZN(n_257_28_108));
   NAND2_X1 i_257_28_109 (.A1(n_257_28_101), .A2(n_257_28_25), .ZN(n_257_28_109));
   NOR2_X1 i_257_28_110 (.A1(n_257_28_109), .A2(n_257_28_5), .ZN(n_257_28_110));
   NAND2_X1 i_257_28_111 (.A1(CPU_Bus[30]), .A2(n_257_28_110), .ZN(n_257_28_111));
   NAND2_X1 i_257_28_112 (.A1(n_257_28_108), .A2(n_257_28_111), .ZN(n_257_28_112));
   NOR2_X1 i_257_28_113 (.A1(n_257_28_105), .A2(n_257_28_112), .ZN(n_257_28_113));
   NOR2_X1 i_257_28_114 (.A1(n_257_28_98), .A2(n_258), .ZN(n_257_28_114));
   NAND2_X1 i_257_28_115 (.A1(CPU_Bus[26]), .A2(n_257_28_114), .ZN(n_257_28_115));
   NOR2_X1 i_257_28_116 (.A1(n_257_28_102), .A2(n_258), .ZN(n_257_28_116));
   NAND2_X1 i_257_28_117 (.A1(CPU_Bus[22]), .A2(n_257_28_116), .ZN(n_257_28_117));
   NAND2_X1 i_257_28_118 (.A1(n_257_28_115), .A2(n_257_28_117), .ZN(n_257_28_118));
   NOR2_X1 i_257_28_119 (.A1(n_257_28_106), .A2(n_258), .ZN(n_257_28_119));
   NAND2_X1 i_257_28_120 (.A1(CPU_Bus[18]), .A2(n_257_28_119), .ZN(n_257_28_120));
   NOR2_X1 i_257_28_121 (.A1(n_257_28_109), .A2(n_258), .ZN(n_257_28_121));
   NAND2_X1 i_257_28_122 (.A1(CPU_Bus[14]), .A2(n_257_28_121), .ZN(n_257_28_122));
   NAND2_X1 i_257_28_123 (.A1(n_257_28_120), .A2(n_257_28_122), .ZN(n_257_28_123));
   NOR2_X1 i_257_28_124 (.A1(n_257_28_118), .A2(n_257_28_123), .ZN(n_257_28_124));
   NAND2_X1 i_257_28_125 (.A1(n_257_28_113), .A2(n_257_28_124), .ZN(n_257_28_125));
   NOR2_X1 i_257_28_126 (.A1(n_257_28_95), .A2(n_257_28_125), .ZN(n_257_28_126));
   NAND2_X1 i_257_28_127 (.A1(n_257_28_65), .A2(n_257_28_126), .ZN(n_257_145));
   datapath__1_350 i_257_29 (.PacketSize(PacketSize), .p_0({n_257_151, uc_258, 
      uc_259, uc_260, uc_261, uc_262, uc_263, uc_264, uc_265, uc_266, uc_267, 
      uc_268, uc_269, uc_270, uc_271, uc_272, uc_273, uc_274, uc_275, uc_276, 
      uc_277, uc_278, uc_279, uc_280, uc_281, uc_282, n_257_150, n_257_149, 
      n_257_148, n_257_147, n_257_146, uc_283}));
   datapath__1_351 i_257_30 (.p_0({uc_284, uc_285, uc_286, uc_287, uc_288, 
      uc_289, uc_290, uc_291, uc_292, uc_293, uc_294, uc_295, uc_296, uc_297, 
      uc_298, uc_299, uc_300, uc_301, uc_302, uc_303, uc_304, uc_305, uc_306, 
      uc_307, uc_308, n_257_151, n_257_150, n_257_149, n_257_148, n_257_147, 
      n_257_146, n_151}), .p_1({n_257_183, n_257_182, n_257_181, n_257_180, 
      n_257_179, n_257_178, n_257_177, n_257_176, n_257_175, n_257_174, 
      n_257_173, n_257_172, n_257_171, n_257_170, n_257_169, n_257_168, 
      n_257_167, n_257_166, n_257_165, n_257_164, n_257_163, n_257_162, 
      n_257_161, n_257_160, n_257_159, n_257_158, n_257_157, n_257_156, 
      n_257_155, n_257_154, n_257_153, n_257_152}));
   NAND2_X1 i_257_31_0 (.A1(n_257_31_0), .A2(n_257_31_36), .ZN(n_257_184));
   NAND2_X1 i_257_31_1 (.A1(n_257_31_1), .A2(n_258), .ZN(n_257_31_0));
   NAND2_X1 i_257_31_2 (.A1(n_257_31_19), .A2(n_257_31_2), .ZN(n_257_31_1));
   NAND3_X1 i_257_31_3 (.A1(n_257_31_11), .A2(n_257_31_3), .A3(n_257_31_87), 
      .ZN(n_257_31_2));
   NAND2_X1 i_257_31_4 (.A1(n_257_31_4), .A2(n_257_31_86), .ZN(n_257_31_3));
   NAND2_X1 i_257_31_5 (.A1(n_257_31_8), .A2(n_257_31_5), .ZN(n_257_31_4));
   NAND3_X1 i_257_31_6 (.A1(n_257_31_7), .A2(n_257_31_6), .A3(n_255), .ZN(
      n_257_31_5));
   NAND2_X1 i_257_31_7 (.A1(CPU_Bus[28]), .A2(n_257_31_82), .ZN(n_257_31_6));
   NAND2_X1 i_257_31_8 (.A1(CPU_Bus[29]), .A2(n_254), .ZN(n_257_31_7));
   NAND3_X1 i_257_31_9 (.A1(n_257_31_10), .A2(n_257_31_9), .A3(n_257_31_85), 
      .ZN(n_257_31_8));
   NAND2_X1 i_257_31_10 (.A1(CPU_Bus[26]), .A2(n_257_31_82), .ZN(n_257_31_9));
   NAND2_X1 i_257_31_11 (.A1(CPU_Bus[27]), .A2(n_254), .ZN(n_257_31_10));
   NAND2_X1 i_257_31_12 (.A1(n_257_31_12), .A2(n_256), .ZN(n_257_31_11));
   NAND2_X1 i_257_31_13 (.A1(n_257_31_16), .A2(n_257_31_13), .ZN(n_257_31_12));
   NAND3_X1 i_257_31_14 (.A1(n_257_31_15), .A2(n_257_31_14), .A3(n_255), 
      .ZN(n_257_31_13));
   NAND2_X1 i_257_31_15 (.A1(CPU_Bus[0]), .A2(n_257_31_82), .ZN(n_257_31_14));
   NAND2_X1 i_257_31_16 (.A1(CPU_Bus[1]), .A2(n_254), .ZN(n_257_31_15));
   NAND3_X1 i_257_31_17 (.A1(n_257_31_18), .A2(n_257_31_17), .A3(n_257_31_85), 
      .ZN(n_257_31_16));
   NAND2_X1 i_257_31_18 (.A1(CPU_Bus[30]), .A2(n_257_31_82), .ZN(n_257_31_17));
   NAND2_X1 i_257_31_19 (.A1(CPU_Bus[31]), .A2(n_254), .ZN(n_257_31_18));
   NAND3_X1 i_257_31_20 (.A1(n_257_31_28), .A2(n_257_31_20), .A3(n_257), 
      .ZN(n_257_31_19));
   NAND2_X1 i_257_31_21 (.A1(n_257_31_21), .A2(n_257_31_86), .ZN(n_257_31_20));
   NAND2_X1 i_257_31_22 (.A1(n_257_31_25), .A2(n_257_31_22), .ZN(n_257_31_21));
   NAND3_X1 i_257_31_23 (.A1(n_257_31_24), .A2(n_257_31_23), .A3(n_255), 
      .ZN(n_257_31_22));
   NAND2_X1 i_257_31_24 (.A1(CPU_Bus[4]), .A2(n_257_31_82), .ZN(n_257_31_23));
   NAND2_X1 i_257_31_25 (.A1(CPU_Bus[5]), .A2(n_254), .ZN(n_257_31_24));
   NAND3_X1 i_257_31_26 (.A1(n_257_31_27), .A2(n_257_31_26), .A3(n_257_31_85), 
      .ZN(n_257_31_25));
   NAND2_X1 i_257_31_27 (.A1(CPU_Bus[2]), .A2(n_257_31_82), .ZN(n_257_31_26));
   NAND2_X1 i_257_31_28 (.A1(CPU_Bus[3]), .A2(n_254), .ZN(n_257_31_27));
   NAND2_X1 i_257_31_29 (.A1(n_257_31_29), .A2(n_256), .ZN(n_257_31_28));
   NAND2_X1 i_257_31_30 (.A1(n_257_31_33), .A2(n_257_31_30), .ZN(n_257_31_29));
   NAND3_X1 i_257_31_31 (.A1(n_257_31_32), .A2(n_257_31_31), .A3(n_255), 
      .ZN(n_257_31_30));
   NAND2_X1 i_257_31_32 (.A1(CPU_Bus[8]), .A2(n_257_31_82), .ZN(n_257_31_31));
   NAND2_X1 i_257_31_33 (.A1(CPU_Bus[9]), .A2(n_254), .ZN(n_257_31_32));
   NAND3_X1 i_257_31_34 (.A1(n_257_31_35), .A2(n_257_31_34), .A3(n_257_31_85), 
      .ZN(n_257_31_33));
   NAND2_X1 i_257_31_35 (.A1(CPU_Bus[6]), .A2(n_257_31_82), .ZN(n_257_31_34));
   NAND2_X1 i_257_31_36 (.A1(CPU_Bus[7]), .A2(n_254), .ZN(n_257_31_35));
   NAND2_X1 i_257_31_37 (.A1(n_257_31_37), .A2(n_257_31_88), .ZN(n_257_31_36));
   NAND2_X1 i_257_31_38 (.A1(n_257_31_61), .A2(n_257_31_38), .ZN(n_257_31_37));
   NAND3_X1 i_257_31_39 (.A1(n_257_31_50), .A2(n_257_31_39), .A3(n_257), 
      .ZN(n_257_31_38));
   NAND3_X1 i_257_31_40 (.A1(n_257_31_45), .A2(n_257_31_40), .A3(n_257_31_86), 
      .ZN(n_257_31_39));
   NAND3_X1 i_257_31_41 (.A1(n_257_31_43), .A2(n_257_31_41), .A3(n_255), 
      .ZN(n_257_31_40));
   NAND2_X1 i_257_31_42 (.A1(n_257_31_42), .A2(n_257_31_82), .ZN(n_257_31_41));
   INV_X1 i_257_31_43 (.A(CPU_Bus[20]), .ZN(n_257_31_42));
   NAND2_X1 i_257_31_44 (.A1(n_257_31_44), .A2(n_254), .ZN(n_257_31_43));
   INV_X1 i_257_31_45 (.A(CPU_Bus[21]), .ZN(n_257_31_44));
   NAND3_X1 i_257_31_46 (.A1(n_257_31_48), .A2(n_257_31_46), .A3(n_257_31_85), 
      .ZN(n_257_31_45));
   NAND2_X1 i_257_31_47 (.A1(n_257_31_47), .A2(n_257_31_82), .ZN(n_257_31_46));
   INV_X1 i_257_31_48 (.A(CPU_Bus[18]), .ZN(n_257_31_47));
   NAND2_X1 i_257_31_49 (.A1(n_257_31_49), .A2(n_254), .ZN(n_257_31_48));
   INV_X1 i_257_31_50 (.A(CPU_Bus[19]), .ZN(n_257_31_49));
   NAND3_X1 i_257_31_51 (.A1(n_257_31_56), .A2(n_257_31_51), .A3(n_256), 
      .ZN(n_257_31_50));
   NAND3_X1 i_257_31_52 (.A1(n_257_31_54), .A2(n_257_31_52), .A3(n_257_31_85), 
      .ZN(n_257_31_51));
   NAND2_X1 i_257_31_53 (.A1(n_257_31_53), .A2(n_257_31_82), .ZN(n_257_31_52));
   INV_X1 i_257_31_54 (.A(CPU_Bus[22]), .ZN(n_257_31_53));
   NAND2_X1 i_257_31_55 (.A1(n_257_31_55), .A2(n_254), .ZN(n_257_31_54));
   INV_X1 i_257_31_56 (.A(CPU_Bus[23]), .ZN(n_257_31_55));
   NAND3_X1 i_257_31_57 (.A1(n_257_31_59), .A2(n_257_31_57), .A3(n_255), 
      .ZN(n_257_31_56));
   NAND2_X1 i_257_31_58 (.A1(n_257_31_58), .A2(n_257_31_82), .ZN(n_257_31_57));
   INV_X1 i_257_31_59 (.A(CPU_Bus[24]), .ZN(n_257_31_58));
   NAND2_X1 i_257_31_60 (.A1(n_257_31_60), .A2(n_254), .ZN(n_257_31_59));
   INV_X1 i_257_31_61 (.A(CPU_Bus[25]), .ZN(n_257_31_60));
   NAND3_X1 i_257_31_62 (.A1(n_257_31_73), .A2(n_257_31_62), .A3(n_257_31_87), 
      .ZN(n_257_31_61));
   NAND3_X1 i_257_31_63 (.A1(n_257_31_68), .A2(n_257_31_63), .A3(n_256), 
      .ZN(n_257_31_62));
   NAND3_X1 i_257_31_64 (.A1(n_257_31_66), .A2(n_257_31_64), .A3(n_257_31_85), 
      .ZN(n_257_31_63));
   NAND2_X1 i_257_31_65 (.A1(n_257_31_65), .A2(n_257_31_82), .ZN(n_257_31_64));
   INV_X1 i_257_31_66 (.A(CPU_Bus[14]), .ZN(n_257_31_65));
   NAND2_X1 i_257_31_67 (.A1(n_257_31_67), .A2(n_254), .ZN(n_257_31_66));
   INV_X1 i_257_31_68 (.A(CPU_Bus[15]), .ZN(n_257_31_67));
   NAND3_X1 i_257_31_69 (.A1(n_257_31_71), .A2(n_257_31_69), .A3(n_255), 
      .ZN(n_257_31_68));
   NAND2_X1 i_257_31_70 (.A1(n_257_31_70), .A2(n_257_31_82), .ZN(n_257_31_69));
   INV_X1 i_257_31_71 (.A(CPU_Bus[16]), .ZN(n_257_31_70));
   NAND2_X1 i_257_31_72 (.A1(n_257_31_72), .A2(n_254), .ZN(n_257_31_71));
   INV_X1 i_257_31_73 (.A(CPU_Bus[17]), .ZN(n_257_31_72));
   NAND3_X1 i_257_31_74 (.A1(n_257_31_79), .A2(n_257_31_74), .A3(n_257_31_86), 
      .ZN(n_257_31_73));
   NAND3_X1 i_257_31_75 (.A1(n_257_31_77), .A2(n_257_31_75), .A3(n_255), 
      .ZN(n_257_31_74));
   NAND2_X1 i_257_31_76 (.A1(n_257_31_76), .A2(n_257_31_82), .ZN(n_257_31_75));
   INV_X1 i_257_31_77 (.A(CPU_Bus[12]), .ZN(n_257_31_76));
   NAND2_X1 i_257_31_78 (.A1(n_257_31_78), .A2(n_254), .ZN(n_257_31_77));
   INV_X1 i_257_31_79 (.A(CPU_Bus[13]), .ZN(n_257_31_78));
   NAND3_X1 i_257_31_80 (.A1(n_257_31_83), .A2(n_257_31_80), .A3(n_257_31_85), 
      .ZN(n_257_31_79));
   NAND2_X1 i_257_31_81 (.A1(n_257_31_81), .A2(n_257_31_82), .ZN(n_257_31_80));
   INV_X1 i_257_31_82 (.A(CPU_Bus[10]), .ZN(n_257_31_81));
   INV_X1 i_257_31_83 (.A(n_254), .ZN(n_257_31_82));
   NAND2_X1 i_257_31_84 (.A1(n_257_31_84), .A2(n_254), .ZN(n_257_31_83));
   INV_X1 i_257_31_85 (.A(CPU_Bus[11]), .ZN(n_257_31_84));
   INV_X1 i_257_31_86 (.A(n_255), .ZN(n_257_31_85));
   INV_X1 i_257_31_87 (.A(n_256), .ZN(n_257_31_86));
   INV_X1 i_257_31_88 (.A(n_257), .ZN(n_257_31_87));
   INV_X1 i_257_31_89 (.A(n_258), .ZN(n_257_31_88));
   INV_X1 i_257_32_0 (.A(n_254), .ZN(n_257_32_0));
   NAND2_X1 i_257_32_1 (.A1(n_257_32_0), .A2(n_255), .ZN(n_257_32_1));
   INV_X1 i_257_32_2 (.A(n_256), .ZN(n_257_32_2));
   NOR2_X1 i_257_32_3 (.A1(n_257_32_1), .A2(n_257_32_2), .ZN(n_257_32_3));
   NAND2_X1 i_257_32_4 (.A1(n_257_32_3), .A2(n_257), .ZN(n_257_32_4));
   INV_X1 i_257_32_5 (.A(n_258), .ZN(n_257_32_5));
   NOR2_X1 i_257_32_6 (.A1(n_257_32_4), .A2(n_257_32_5), .ZN(n_257_32_6));
   NAND2_X1 i_257_32_7 (.A1(CPU_Bus[7]), .A2(n_257_32_6), .ZN(n_257_32_7));
   INV_X1 i_257_32_8 (.A(n_255), .ZN(n_257_32_8));
   NAND2_X1 i_257_32_9 (.A1(n_257_32_0), .A2(n_257_32_8), .ZN(n_257_32_9));
   NOR2_X1 i_257_32_10 (.A1(n_257_32_9), .A2(n_257_32_2), .ZN(n_257_32_10));
   NAND2_X1 i_257_32_11 (.A1(n_257_32_10), .A2(n_257), .ZN(n_257_32_11));
   NOR2_X1 i_257_32_12 (.A1(n_257_32_11), .A2(n_257_32_5), .ZN(n_257_32_12));
   NAND2_X1 i_257_32_13 (.A1(CPU_Bus[5]), .A2(n_257_32_12), .ZN(n_257_32_13));
   NAND2_X1 i_257_32_14 (.A1(n_257_32_7), .A2(n_257_32_13), .ZN(n_257_32_14));
   NOR2_X1 i_257_32_15 (.A1(n_257_32_1), .A2(n_256), .ZN(n_257_32_15));
   NAND2_X1 i_257_32_16 (.A1(n_257_32_15), .A2(n_257), .ZN(n_257_32_16));
   NOR2_X1 i_257_32_17 (.A1(n_257_32_16), .A2(n_257_32_5), .ZN(n_257_32_17));
   NAND2_X1 i_257_32_18 (.A1(CPU_Bus[3]), .A2(n_257_32_17), .ZN(n_257_32_18));
   NOR2_X1 i_257_32_19 (.A1(n_257_32_9), .A2(n_256), .ZN(n_257_32_19));
   NAND2_X1 i_257_32_20 (.A1(n_257_32_19), .A2(n_257), .ZN(n_257_32_20));
   NOR2_X1 i_257_32_21 (.A1(n_257_32_20), .A2(n_257_32_5), .ZN(n_257_32_21));
   NAND2_X1 i_257_32_22 (.A1(CPU_Bus[1]), .A2(n_257_32_21), .ZN(n_257_32_22));
   NAND2_X1 i_257_32_23 (.A1(n_257_32_18), .A2(n_257_32_22), .ZN(n_257_32_23));
   NOR2_X1 i_257_32_24 (.A1(n_257_32_14), .A2(n_257_32_23), .ZN(n_257_32_24));
   INV_X1 i_257_32_25 (.A(n_257), .ZN(n_257_32_25));
   NAND2_X1 i_257_32_26 (.A1(n_257_32_3), .A2(n_257_32_25), .ZN(n_257_32_26));
   NOR2_X1 i_257_32_27 (.A1(n_257_32_26), .A2(n_257_32_5), .ZN(n_257_32_27));
   NAND2_X1 i_257_32_28 (.A1(CPU_Bus[31]), .A2(n_257_32_27), .ZN(n_257_32_28));
   NAND2_X1 i_257_32_29 (.A1(n_257_32_10), .A2(n_257_32_25), .ZN(n_257_32_29));
   NOR2_X1 i_257_32_30 (.A1(n_257_32_29), .A2(n_257_32_5), .ZN(n_257_32_30));
   NAND2_X1 i_257_32_31 (.A1(CPU_Bus[29]), .A2(n_257_32_30), .ZN(n_257_32_31));
   NAND2_X1 i_257_32_32 (.A1(n_257_32_28), .A2(n_257_32_31), .ZN(n_257_32_32));
   NAND2_X1 i_257_32_33 (.A1(n_257_32_15), .A2(n_257_32_25), .ZN(n_257_32_33));
   NOR2_X1 i_257_32_34 (.A1(n_257_32_33), .A2(n_257_32_5), .ZN(n_257_32_34));
   NAND2_X1 i_257_32_35 (.A1(CPU_Bus[27]), .A2(n_257_32_34), .ZN(n_257_32_35));
   NAND2_X1 i_257_32_36 (.A1(n_257_32_19), .A2(n_257_32_25), .ZN(n_257_32_36));
   NOR2_X1 i_257_32_37 (.A1(n_257_32_36), .A2(n_257_32_5), .ZN(n_257_32_37));
   NAND2_X1 i_257_32_38 (.A1(CPU_Bus[25]), .A2(n_257_32_37), .ZN(n_257_32_38));
   NAND2_X1 i_257_32_39 (.A1(n_257_32_35), .A2(n_257_32_38), .ZN(n_257_32_39));
   NOR2_X1 i_257_32_40 (.A1(n_257_32_32), .A2(n_257_32_39), .ZN(n_257_32_40));
   NAND2_X1 i_257_32_41 (.A1(n_257_32_24), .A2(n_257_32_40), .ZN(n_257_32_41));
   NOR2_X1 i_257_32_42 (.A1(n_257_32_4), .A2(n_258), .ZN(n_257_32_42));
   NAND2_X1 i_257_32_43 (.A1(CPU_Bus[23]), .A2(n_257_32_42), .ZN(n_257_32_43));
   NOR2_X1 i_257_32_44 (.A1(n_257_32_11), .A2(n_258), .ZN(n_257_32_44));
   NAND2_X1 i_257_32_45 (.A1(CPU_Bus[21]), .A2(n_257_32_44), .ZN(n_257_32_45));
   NAND2_X1 i_257_32_46 (.A1(n_257_32_43), .A2(n_257_32_45), .ZN(n_257_32_46));
   NOR2_X1 i_257_32_47 (.A1(n_257_32_16), .A2(n_258), .ZN(n_257_32_47));
   NAND2_X1 i_257_32_48 (.A1(CPU_Bus[19]), .A2(n_257_32_47), .ZN(n_257_32_48));
   NOR2_X1 i_257_32_49 (.A1(n_257_32_20), .A2(n_258), .ZN(n_257_32_49));
   NAND2_X1 i_257_32_50 (.A1(CPU_Bus[17]), .A2(n_257_32_49), .ZN(n_257_32_50));
   NAND2_X1 i_257_32_51 (.A1(n_257_32_48), .A2(n_257_32_50), .ZN(n_257_32_51));
   NOR2_X1 i_257_32_52 (.A1(n_257_32_46), .A2(n_257_32_51), .ZN(n_257_32_52));
   NOR2_X1 i_257_32_53 (.A1(n_257_32_26), .A2(n_258), .ZN(n_257_32_53));
   NAND2_X1 i_257_32_54 (.A1(CPU_Bus[15]), .A2(n_257_32_53), .ZN(n_257_32_54));
   NOR2_X1 i_257_32_55 (.A1(n_257_32_29), .A2(n_258), .ZN(n_257_32_55));
   NAND2_X1 i_257_32_56 (.A1(CPU_Bus[13]), .A2(n_257_32_55), .ZN(n_257_32_56));
   NAND2_X1 i_257_32_57 (.A1(n_257_32_54), .A2(n_257_32_56), .ZN(n_257_32_57));
   NOR2_X1 i_257_32_58 (.A1(n_257_32_33), .A2(n_258), .ZN(n_257_32_58));
   NAND2_X1 i_257_32_59 (.A1(CPU_Bus[11]), .A2(n_257_32_58), .ZN(n_257_32_59));
   NOR2_X1 i_257_32_60 (.A1(n_257_32_36), .A2(n_258), .ZN(n_257_32_60));
   NAND2_X1 i_257_32_61 (.A1(CPU_Bus[9]), .A2(n_257_32_60), .ZN(n_257_32_61));
   NAND2_X1 i_257_32_62 (.A1(n_257_32_59), .A2(n_257_32_61), .ZN(n_257_32_62));
   NOR2_X1 i_257_32_63 (.A1(n_257_32_57), .A2(n_257_32_62), .ZN(n_257_32_63));
   NAND2_X1 i_257_32_64 (.A1(n_257_32_52), .A2(n_257_32_63), .ZN(n_257_32_64));
   NOR2_X1 i_257_32_65 (.A1(n_257_32_41), .A2(n_257_32_64), .ZN(n_257_32_65));
   NAND2_X1 i_257_32_66 (.A1(n_257_32_8), .A2(n_254), .ZN(n_257_32_66));
   NOR2_X1 i_257_32_67 (.A1(n_257_32_66), .A2(n_257_32_2), .ZN(n_257_32_67));
   NAND2_X1 i_257_32_68 (.A1(n_257_32_67), .A2(n_257), .ZN(n_257_32_68));
   NOR2_X1 i_257_32_69 (.A1(n_257_32_68), .A2(n_257_32_5), .ZN(n_257_32_69));
   NAND2_X1 i_257_32_70 (.A1(CPU_Bus[6]), .A2(n_257_32_69), .ZN(n_257_32_70));
   NOR2_X1 i_257_32_71 (.A1(n_257_32_66), .A2(n_256), .ZN(n_257_32_71));
   NAND2_X1 i_257_32_72 (.A1(n_257_32_71), .A2(n_257), .ZN(n_257_32_72));
   NOR2_X1 i_257_32_73 (.A1(n_257_32_72), .A2(n_257_32_5), .ZN(n_257_32_73));
   NAND2_X1 i_257_32_74 (.A1(CPU_Bus[2]), .A2(n_257_32_73), .ZN(n_257_32_74));
   NAND2_X1 i_257_32_75 (.A1(n_257_32_70), .A2(n_257_32_74), .ZN(n_257_32_75));
   NAND2_X1 i_257_32_76 (.A1(n_257_32_67), .A2(n_257_32_25), .ZN(n_257_32_76));
   NOR2_X1 i_257_32_77 (.A1(n_257_32_76), .A2(n_257_32_5), .ZN(n_257_32_77));
   NAND2_X1 i_257_32_78 (.A1(CPU_Bus[30]), .A2(n_257_32_77), .ZN(n_257_32_78));
   NAND2_X1 i_257_32_79 (.A1(n_257_32_71), .A2(n_257_32_25), .ZN(n_257_32_79));
   NOR2_X1 i_257_32_80 (.A1(n_257_32_79), .A2(n_257_32_5), .ZN(n_257_32_80));
   NAND2_X1 i_257_32_81 (.A1(CPU_Bus[26]), .A2(n_257_32_80), .ZN(n_257_32_81));
   NAND2_X1 i_257_32_82 (.A1(n_257_32_78), .A2(n_257_32_81), .ZN(n_257_32_82));
   NOR2_X1 i_257_32_83 (.A1(n_257_32_75), .A2(n_257_32_82), .ZN(n_257_32_83));
   NOR2_X1 i_257_32_84 (.A1(n_257_32_68), .A2(n_258), .ZN(n_257_32_84));
   NAND2_X1 i_257_32_85 (.A1(CPU_Bus[22]), .A2(n_257_32_84), .ZN(n_257_32_85));
   NOR2_X1 i_257_32_86 (.A1(n_257_32_72), .A2(n_258), .ZN(n_257_32_86));
   NAND2_X1 i_257_32_87 (.A1(CPU_Bus[18]), .A2(n_257_32_86), .ZN(n_257_32_87));
   NAND2_X1 i_257_32_88 (.A1(n_257_32_85), .A2(n_257_32_87), .ZN(n_257_32_88));
   NOR2_X1 i_257_32_89 (.A1(n_257_32_76), .A2(n_258), .ZN(n_257_32_89));
   NAND2_X1 i_257_32_90 (.A1(CPU_Bus[14]), .A2(n_257_32_89), .ZN(n_257_32_90));
   NOR2_X1 i_257_32_91 (.A1(n_257_32_79), .A2(n_258), .ZN(n_257_32_91));
   NAND2_X1 i_257_32_92 (.A1(CPU_Bus[10]), .A2(n_257_32_91), .ZN(n_257_32_92));
   NAND2_X1 i_257_32_93 (.A1(n_257_32_90), .A2(n_257_32_92), .ZN(n_257_32_93));
   NOR2_X1 i_257_32_94 (.A1(n_257_32_88), .A2(n_257_32_93), .ZN(n_257_32_94));
   NAND2_X1 i_257_32_95 (.A1(n_257_32_83), .A2(n_257_32_94), .ZN(n_257_32_95));
   NAND2_X1 i_257_32_96 (.A1(n_254), .A2(n_255), .ZN(n_257_32_96));
   NOR2_X1 i_257_32_97 (.A1(n_257_32_96), .A2(n_257_32_2), .ZN(n_257_32_97));
   NAND2_X1 i_257_32_98 (.A1(n_257_32_97), .A2(n_257), .ZN(n_257_32_98));
   NOR2_X1 i_257_32_99 (.A1(n_257_32_98), .A2(n_257_32_5), .ZN(n_257_32_99));
   NAND2_X1 i_257_32_100 (.A1(CPU_Bus[8]), .A2(n_257_32_99), .ZN(n_257_32_100));
   NOR2_X1 i_257_32_101 (.A1(n_257_32_96), .A2(n_256), .ZN(n_257_32_101));
   NAND2_X1 i_257_32_102 (.A1(n_257_32_101), .A2(n_257), .ZN(n_257_32_102));
   NOR2_X1 i_257_32_103 (.A1(n_257_32_102), .A2(n_257_32_5), .ZN(n_257_32_103));
   NAND2_X1 i_257_32_104 (.A1(CPU_Bus[4]), .A2(n_257_32_103), .ZN(n_257_32_104));
   NAND2_X1 i_257_32_105 (.A1(n_257_32_100), .A2(n_257_32_104), .ZN(n_257_32_105));
   NAND2_X1 i_257_32_106 (.A1(n_257_32_97), .A2(n_257_32_25), .ZN(n_257_32_106));
   NOR2_X1 i_257_32_107 (.A1(n_257_32_106), .A2(n_257_32_5), .ZN(n_257_32_107));
   NAND2_X1 i_257_32_108 (.A1(CPU_Bus[0]), .A2(n_257_32_107), .ZN(n_257_32_108));
   NAND2_X1 i_257_32_109 (.A1(n_257_32_101), .A2(n_257_32_25), .ZN(n_257_32_109));
   NOR2_X1 i_257_32_110 (.A1(n_257_32_109), .A2(n_257_32_5), .ZN(n_257_32_110));
   NAND2_X1 i_257_32_111 (.A1(CPU_Bus[28]), .A2(n_257_32_110), .ZN(n_257_32_111));
   NAND2_X1 i_257_32_112 (.A1(n_257_32_108), .A2(n_257_32_111), .ZN(n_257_32_112));
   NOR2_X1 i_257_32_113 (.A1(n_257_32_105), .A2(n_257_32_112), .ZN(n_257_32_113));
   NOR2_X1 i_257_32_114 (.A1(n_257_32_98), .A2(n_258), .ZN(n_257_32_114));
   NAND2_X1 i_257_32_115 (.A1(CPU_Bus[24]), .A2(n_257_32_114), .ZN(n_257_32_115));
   NOR2_X1 i_257_32_116 (.A1(n_257_32_102), .A2(n_258), .ZN(n_257_32_116));
   NAND2_X1 i_257_32_117 (.A1(CPU_Bus[20]), .A2(n_257_32_116), .ZN(n_257_32_117));
   NAND2_X1 i_257_32_118 (.A1(n_257_32_115), .A2(n_257_32_117), .ZN(n_257_32_118));
   NOR2_X1 i_257_32_119 (.A1(n_257_32_106), .A2(n_258), .ZN(n_257_32_119));
   NAND2_X1 i_257_32_120 (.A1(CPU_Bus[16]), .A2(n_257_32_119), .ZN(n_257_32_120));
   NOR2_X1 i_257_32_121 (.A1(n_257_32_109), .A2(n_258), .ZN(n_257_32_121));
   NAND2_X1 i_257_32_122 (.A1(CPU_Bus[12]), .A2(n_257_32_121), .ZN(n_257_32_122));
   NAND2_X1 i_257_32_123 (.A1(n_257_32_120), .A2(n_257_32_122), .ZN(n_257_32_123));
   NOR2_X1 i_257_32_124 (.A1(n_257_32_118), .A2(n_257_32_123), .ZN(n_257_32_124));
   NAND2_X1 i_257_32_125 (.A1(n_257_32_113), .A2(n_257_32_124), .ZN(n_257_32_125));
   NOR2_X1 i_257_32_126 (.A1(n_257_32_95), .A2(n_257_32_125), .ZN(n_257_32_126));
   NAND2_X1 i_257_32_127 (.A1(n_257_32_65), .A2(n_257_32_126), .ZN(n_257_185));
   datapath__1_355 i_257_33 (.PacketSize(PacketSize), .p_0({n_257_191, uc_309, 
      uc_310, uc_311, uc_312, uc_313, uc_314, uc_315, uc_316, uc_317, uc_318, 
      uc_319, uc_320, uc_321, uc_322, uc_323, uc_324, uc_325, uc_326, uc_327, 
      uc_328, uc_329, uc_330, uc_331, uc_332, uc_333, n_257_190, n_257_189, 
      n_257_188, n_257_187, n_257_186, uc_334}));
   datapath__1_356 i_257_34 (.p_0({uc_335, uc_336, uc_337, uc_338, uc_339, 
      uc_340, uc_341, uc_342, uc_343, uc_344, uc_345, uc_346, uc_347, uc_348, 
      uc_349, uc_350, uc_351, uc_352, uc_353, uc_354, uc_355, uc_356, uc_357, 
      uc_358, uc_359, n_257_191, n_257_190, n_257_189, n_257_188, n_257_187, 
      n_257_186, n_151}), .p_1({n_257_223, n_257_222, n_257_221, n_257_220, 
      n_257_219, n_257_218, n_257_217, n_257_216, n_257_215, n_257_214, 
      n_257_213, n_257_212, n_257_211, n_257_210, n_257_209, n_257_208, 
      n_257_207, n_257_206, n_257_205, n_257_204, n_257_203, n_257_202, 
      n_257_201, n_257_200, n_257_199, n_257_198, n_257_197, n_257_196, 
      n_257_195, n_257_194, n_257_193, n_257_192}));
   INV_X1 i_257_35_0 (.A(n_254), .ZN(n_257_35_0));
   NAND2_X1 i_257_35_1 (.A1(n_257_35_0), .A2(n_255), .ZN(n_257_35_1));
   INV_X1 i_257_35_2 (.A(n_256), .ZN(n_257_35_2));
   NOR2_X1 i_257_35_3 (.A1(n_257_35_1), .A2(n_257_35_2), .ZN(n_257_35_3));
   NAND2_X1 i_257_35_4 (.A1(n_257_35_3), .A2(n_257), .ZN(n_257_35_4));
   INV_X1 i_257_35_5 (.A(n_258), .ZN(n_257_35_5));
   NOR2_X1 i_257_35_6 (.A1(n_257_35_4), .A2(n_257_35_5), .ZN(n_257_35_6));
   NAND2_X1 i_257_35_7 (.A1(CPU_Bus[6]), .A2(n_257_35_6), .ZN(n_257_35_7));
   INV_X1 i_257_35_8 (.A(n_255), .ZN(n_257_35_8));
   NAND2_X1 i_257_35_9 (.A1(n_257_35_0), .A2(n_257_35_8), .ZN(n_257_35_9));
   NOR2_X1 i_257_35_10 (.A1(n_257_35_9), .A2(n_257_35_2), .ZN(n_257_35_10));
   NAND2_X1 i_257_35_11 (.A1(n_257_35_10), .A2(n_257), .ZN(n_257_35_11));
   NOR2_X1 i_257_35_12 (.A1(n_257_35_11), .A2(n_257_35_5), .ZN(n_257_35_12));
   NAND2_X1 i_257_35_13 (.A1(CPU_Bus[4]), .A2(n_257_35_12), .ZN(n_257_35_13));
   NAND2_X1 i_257_35_14 (.A1(n_257_35_7), .A2(n_257_35_13), .ZN(n_257_35_14));
   NOR2_X1 i_257_35_15 (.A1(n_257_35_1), .A2(n_256), .ZN(n_257_35_15));
   NAND2_X1 i_257_35_16 (.A1(n_257_35_15), .A2(n_257), .ZN(n_257_35_16));
   NOR2_X1 i_257_35_17 (.A1(n_257_35_16), .A2(n_257_35_5), .ZN(n_257_35_17));
   NAND2_X1 i_257_35_18 (.A1(CPU_Bus[2]), .A2(n_257_35_17), .ZN(n_257_35_18));
   NOR2_X1 i_257_35_19 (.A1(n_257_35_9), .A2(n_256), .ZN(n_257_35_19));
   NAND2_X1 i_257_35_20 (.A1(n_257_35_19), .A2(n_257), .ZN(n_257_35_20));
   NOR2_X1 i_257_35_21 (.A1(n_257_35_20), .A2(n_257_35_5), .ZN(n_257_35_21));
   NAND2_X1 i_257_35_22 (.A1(CPU_Bus[0]), .A2(n_257_35_21), .ZN(n_257_35_22));
   NAND2_X1 i_257_35_23 (.A1(n_257_35_18), .A2(n_257_35_22), .ZN(n_257_35_23));
   NOR2_X1 i_257_35_24 (.A1(n_257_35_14), .A2(n_257_35_23), .ZN(n_257_35_24));
   INV_X1 i_257_35_25 (.A(n_257), .ZN(n_257_35_25));
   NAND2_X1 i_257_35_26 (.A1(n_257_35_3), .A2(n_257_35_25), .ZN(n_257_35_26));
   NOR2_X1 i_257_35_27 (.A1(n_257_35_26), .A2(n_257_35_5), .ZN(n_257_35_27));
   NAND2_X1 i_257_35_28 (.A1(CPU_Bus[30]), .A2(n_257_35_27), .ZN(n_257_35_28));
   NAND2_X1 i_257_35_29 (.A1(n_257_35_10), .A2(n_257_35_25), .ZN(n_257_35_29));
   NOR2_X1 i_257_35_30 (.A1(n_257_35_29), .A2(n_257_35_5), .ZN(n_257_35_30));
   NAND2_X1 i_257_35_31 (.A1(CPU_Bus[28]), .A2(n_257_35_30), .ZN(n_257_35_31));
   NAND2_X1 i_257_35_32 (.A1(n_257_35_28), .A2(n_257_35_31), .ZN(n_257_35_32));
   NAND2_X1 i_257_35_33 (.A1(n_257_35_15), .A2(n_257_35_25), .ZN(n_257_35_33));
   NOR2_X1 i_257_35_34 (.A1(n_257_35_33), .A2(n_257_35_5), .ZN(n_257_35_34));
   NAND2_X1 i_257_35_35 (.A1(CPU_Bus[26]), .A2(n_257_35_34), .ZN(n_257_35_35));
   NAND2_X1 i_257_35_36 (.A1(n_257_35_19), .A2(n_257_35_25), .ZN(n_257_35_36));
   NOR2_X1 i_257_35_37 (.A1(n_257_35_36), .A2(n_257_35_5), .ZN(n_257_35_37));
   NAND2_X1 i_257_35_38 (.A1(CPU_Bus[24]), .A2(n_257_35_37), .ZN(n_257_35_38));
   NAND2_X1 i_257_35_39 (.A1(n_257_35_35), .A2(n_257_35_38), .ZN(n_257_35_39));
   NOR2_X1 i_257_35_40 (.A1(n_257_35_32), .A2(n_257_35_39), .ZN(n_257_35_40));
   NAND2_X1 i_257_35_41 (.A1(n_257_35_24), .A2(n_257_35_40), .ZN(n_257_35_41));
   NOR2_X1 i_257_35_42 (.A1(n_257_35_4), .A2(n_258), .ZN(n_257_35_42));
   NAND2_X1 i_257_35_43 (.A1(CPU_Bus[22]), .A2(n_257_35_42), .ZN(n_257_35_43));
   NOR2_X1 i_257_35_44 (.A1(n_257_35_11), .A2(n_258), .ZN(n_257_35_44));
   NAND2_X1 i_257_35_45 (.A1(CPU_Bus[20]), .A2(n_257_35_44), .ZN(n_257_35_45));
   NAND2_X1 i_257_35_46 (.A1(n_257_35_43), .A2(n_257_35_45), .ZN(n_257_35_46));
   NOR2_X1 i_257_35_47 (.A1(n_257_35_16), .A2(n_258), .ZN(n_257_35_47));
   NAND2_X1 i_257_35_48 (.A1(CPU_Bus[18]), .A2(n_257_35_47), .ZN(n_257_35_48));
   NOR2_X1 i_257_35_49 (.A1(n_257_35_20), .A2(n_258), .ZN(n_257_35_49));
   NAND2_X1 i_257_35_50 (.A1(CPU_Bus[16]), .A2(n_257_35_49), .ZN(n_257_35_50));
   NAND2_X1 i_257_35_51 (.A1(n_257_35_48), .A2(n_257_35_50), .ZN(n_257_35_51));
   NOR2_X1 i_257_35_52 (.A1(n_257_35_46), .A2(n_257_35_51), .ZN(n_257_35_52));
   NOR2_X1 i_257_35_53 (.A1(n_257_35_26), .A2(n_258), .ZN(n_257_35_53));
   NAND2_X1 i_257_35_54 (.A1(CPU_Bus[14]), .A2(n_257_35_53), .ZN(n_257_35_54));
   NOR2_X1 i_257_35_55 (.A1(n_257_35_29), .A2(n_258), .ZN(n_257_35_55));
   NAND2_X1 i_257_35_56 (.A1(CPU_Bus[12]), .A2(n_257_35_55), .ZN(n_257_35_56));
   NAND2_X1 i_257_35_57 (.A1(n_257_35_54), .A2(n_257_35_56), .ZN(n_257_35_57));
   NOR2_X1 i_257_35_58 (.A1(n_257_35_33), .A2(n_258), .ZN(n_257_35_58));
   NAND2_X1 i_257_35_59 (.A1(CPU_Bus[10]), .A2(n_257_35_58), .ZN(n_257_35_59));
   NOR2_X1 i_257_35_60 (.A1(n_257_35_36), .A2(n_258), .ZN(n_257_35_60));
   NAND2_X1 i_257_35_61 (.A1(CPU_Bus[8]), .A2(n_257_35_60), .ZN(n_257_35_61));
   NAND2_X1 i_257_35_62 (.A1(n_257_35_59), .A2(n_257_35_61), .ZN(n_257_35_62));
   NOR2_X1 i_257_35_63 (.A1(n_257_35_57), .A2(n_257_35_62), .ZN(n_257_35_63));
   NAND2_X1 i_257_35_64 (.A1(n_257_35_52), .A2(n_257_35_63), .ZN(n_257_35_64));
   NOR2_X1 i_257_35_65 (.A1(n_257_35_41), .A2(n_257_35_64), .ZN(n_257_35_65));
   NAND2_X1 i_257_35_66 (.A1(n_257_35_8), .A2(n_254), .ZN(n_257_35_66));
   NOR2_X1 i_257_35_67 (.A1(n_257_35_66), .A2(n_257_35_2), .ZN(n_257_35_67));
   NAND2_X1 i_257_35_68 (.A1(n_257_35_67), .A2(n_257), .ZN(n_257_35_68));
   NOR2_X1 i_257_35_69 (.A1(n_257_35_68), .A2(n_257_35_5), .ZN(n_257_35_69));
   NAND2_X1 i_257_35_70 (.A1(CPU_Bus[5]), .A2(n_257_35_69), .ZN(n_257_35_70));
   NOR2_X1 i_257_35_71 (.A1(n_257_35_66), .A2(n_256), .ZN(n_257_35_71));
   NAND2_X1 i_257_35_72 (.A1(n_257_35_71), .A2(n_257), .ZN(n_257_35_72));
   NOR2_X1 i_257_35_73 (.A1(n_257_35_72), .A2(n_257_35_5), .ZN(n_257_35_73));
   NAND2_X1 i_257_35_74 (.A1(CPU_Bus[1]), .A2(n_257_35_73), .ZN(n_257_35_74));
   NAND2_X1 i_257_35_75 (.A1(n_257_35_70), .A2(n_257_35_74), .ZN(n_257_35_75));
   NAND2_X1 i_257_35_76 (.A1(n_257_35_67), .A2(n_257_35_25), .ZN(n_257_35_76));
   NOR2_X1 i_257_35_77 (.A1(n_257_35_76), .A2(n_257_35_5), .ZN(n_257_35_77));
   NAND2_X1 i_257_35_78 (.A1(CPU_Bus[29]), .A2(n_257_35_77), .ZN(n_257_35_78));
   NAND2_X1 i_257_35_79 (.A1(n_257_35_71), .A2(n_257_35_25), .ZN(n_257_35_79));
   NOR2_X1 i_257_35_80 (.A1(n_257_35_79), .A2(n_257_35_5), .ZN(n_257_35_80));
   NAND2_X1 i_257_35_81 (.A1(CPU_Bus[25]), .A2(n_257_35_80), .ZN(n_257_35_81));
   NAND2_X1 i_257_35_82 (.A1(n_257_35_78), .A2(n_257_35_81), .ZN(n_257_35_82));
   NOR2_X1 i_257_35_83 (.A1(n_257_35_75), .A2(n_257_35_82), .ZN(n_257_35_83));
   NOR2_X1 i_257_35_84 (.A1(n_257_35_68), .A2(n_258), .ZN(n_257_35_84));
   NAND2_X1 i_257_35_85 (.A1(CPU_Bus[21]), .A2(n_257_35_84), .ZN(n_257_35_85));
   NOR2_X1 i_257_35_86 (.A1(n_257_35_72), .A2(n_258), .ZN(n_257_35_86));
   NAND2_X1 i_257_35_87 (.A1(CPU_Bus[17]), .A2(n_257_35_86), .ZN(n_257_35_87));
   NAND2_X1 i_257_35_88 (.A1(n_257_35_85), .A2(n_257_35_87), .ZN(n_257_35_88));
   NOR2_X1 i_257_35_89 (.A1(n_257_35_76), .A2(n_258), .ZN(n_257_35_89));
   NAND2_X1 i_257_35_90 (.A1(CPU_Bus[13]), .A2(n_257_35_89), .ZN(n_257_35_90));
   NOR2_X1 i_257_35_91 (.A1(n_257_35_79), .A2(n_258), .ZN(n_257_35_91));
   NAND2_X1 i_257_35_92 (.A1(CPU_Bus[9]), .A2(n_257_35_91), .ZN(n_257_35_92));
   NAND2_X1 i_257_35_93 (.A1(n_257_35_90), .A2(n_257_35_92), .ZN(n_257_35_93));
   NOR2_X1 i_257_35_94 (.A1(n_257_35_88), .A2(n_257_35_93), .ZN(n_257_35_94));
   NAND2_X1 i_257_35_95 (.A1(n_257_35_83), .A2(n_257_35_94), .ZN(n_257_35_95));
   NAND2_X1 i_257_35_96 (.A1(n_254), .A2(n_255), .ZN(n_257_35_96));
   NOR2_X1 i_257_35_97 (.A1(n_257_35_96), .A2(n_257_35_2), .ZN(n_257_35_97));
   NAND2_X1 i_257_35_98 (.A1(n_257_35_97), .A2(n_257), .ZN(n_257_35_98));
   NOR2_X1 i_257_35_99 (.A1(n_257_35_98), .A2(n_257_35_5), .ZN(n_257_35_99));
   NAND2_X1 i_257_35_100 (.A1(CPU_Bus[7]), .A2(n_257_35_99), .ZN(n_257_35_100));
   NOR2_X1 i_257_35_101 (.A1(n_257_35_96), .A2(n_256), .ZN(n_257_35_101));
   NAND2_X1 i_257_35_102 (.A1(n_257_35_101), .A2(n_257), .ZN(n_257_35_102));
   NOR2_X1 i_257_35_103 (.A1(n_257_35_102), .A2(n_257_35_5), .ZN(n_257_35_103));
   NAND2_X1 i_257_35_104 (.A1(CPU_Bus[3]), .A2(n_257_35_103), .ZN(n_257_35_104));
   NAND2_X1 i_257_35_105 (.A1(n_257_35_100), .A2(n_257_35_104), .ZN(n_257_35_105));
   NAND2_X1 i_257_35_106 (.A1(n_257_35_97), .A2(n_257_35_25), .ZN(n_257_35_106));
   NOR2_X1 i_257_35_107 (.A1(n_257_35_106), .A2(n_257_35_5), .ZN(n_257_35_107));
   NAND2_X1 i_257_35_108 (.A1(CPU_Bus[31]), .A2(n_257_35_107), .ZN(n_257_35_108));
   NAND2_X1 i_257_35_109 (.A1(n_257_35_101), .A2(n_257_35_25), .ZN(n_257_35_109));
   NOR2_X1 i_257_35_110 (.A1(n_257_35_109), .A2(n_257_35_5), .ZN(n_257_35_110));
   NAND2_X1 i_257_35_111 (.A1(CPU_Bus[27]), .A2(n_257_35_110), .ZN(n_257_35_111));
   NAND2_X1 i_257_35_112 (.A1(n_257_35_108), .A2(n_257_35_111), .ZN(n_257_35_112));
   NOR2_X1 i_257_35_113 (.A1(n_257_35_105), .A2(n_257_35_112), .ZN(n_257_35_113));
   NOR2_X1 i_257_35_114 (.A1(n_257_35_98), .A2(n_258), .ZN(n_257_35_114));
   NAND2_X1 i_257_35_115 (.A1(CPU_Bus[23]), .A2(n_257_35_114), .ZN(n_257_35_115));
   NOR2_X1 i_257_35_116 (.A1(n_257_35_102), .A2(n_258), .ZN(n_257_35_116));
   NAND2_X1 i_257_35_117 (.A1(CPU_Bus[19]), .A2(n_257_35_116), .ZN(n_257_35_117));
   NAND2_X1 i_257_35_118 (.A1(n_257_35_115), .A2(n_257_35_117), .ZN(n_257_35_118));
   NOR2_X1 i_257_35_119 (.A1(n_257_35_106), .A2(n_258), .ZN(n_257_35_119));
   NAND2_X1 i_257_35_120 (.A1(CPU_Bus[15]), .A2(n_257_35_119), .ZN(n_257_35_120));
   NOR2_X1 i_257_35_121 (.A1(n_257_35_109), .A2(n_258), .ZN(n_257_35_121));
   NAND2_X1 i_257_35_122 (.A1(CPU_Bus[11]), .A2(n_257_35_121), .ZN(n_257_35_122));
   NAND2_X1 i_257_35_123 (.A1(n_257_35_120), .A2(n_257_35_122), .ZN(n_257_35_123));
   NOR2_X1 i_257_35_124 (.A1(n_257_35_118), .A2(n_257_35_123), .ZN(n_257_35_124));
   NAND2_X1 i_257_35_125 (.A1(n_257_35_113), .A2(n_257_35_124), .ZN(n_257_35_125));
   NOR2_X1 i_257_35_126 (.A1(n_257_35_95), .A2(n_257_35_125), .ZN(n_257_35_126));
   NAND2_X1 i_257_35_127 (.A1(n_257_35_65), .A2(n_257_35_126), .ZN(n_257_224));
   INV_X1 i_257_36_0 (.A(n_254), .ZN(n_257_36_0));
   NAND2_X1 i_257_36_1 (.A1(n_257_36_0), .A2(n_255), .ZN(n_257_36_1));
   INV_X1 i_257_36_2 (.A(n_256), .ZN(n_257_36_2));
   NOR2_X1 i_257_36_3 (.A1(n_257_36_1), .A2(n_257_36_2), .ZN(n_257_36_3));
   NAND2_X1 i_257_36_4 (.A1(n_257_36_3), .A2(n_257), .ZN(n_257_36_4));
   INV_X1 i_257_36_5 (.A(n_258), .ZN(n_257_36_5));
   NOR2_X1 i_257_36_6 (.A1(n_257_36_4), .A2(n_257_36_5), .ZN(n_257_36_6));
   NAND2_X1 i_257_36_7 (.A1(CPU_Bus[5]), .A2(n_257_36_6), .ZN(n_257_36_7));
   INV_X1 i_257_36_8 (.A(n_255), .ZN(n_257_36_8));
   NAND2_X1 i_257_36_9 (.A1(n_257_36_0), .A2(n_257_36_8), .ZN(n_257_36_9));
   NOR2_X1 i_257_36_10 (.A1(n_257_36_9), .A2(n_257_36_2), .ZN(n_257_36_10));
   NAND2_X1 i_257_36_11 (.A1(n_257_36_10), .A2(n_257), .ZN(n_257_36_11));
   NOR2_X1 i_257_36_12 (.A1(n_257_36_11), .A2(n_257_36_5), .ZN(n_257_36_12));
   NAND2_X1 i_257_36_13 (.A1(CPU_Bus[3]), .A2(n_257_36_12), .ZN(n_257_36_13));
   NAND2_X1 i_257_36_14 (.A1(n_257_36_7), .A2(n_257_36_13), .ZN(n_257_36_14));
   NOR2_X1 i_257_36_15 (.A1(n_257_36_1), .A2(n_256), .ZN(n_257_36_15));
   NAND2_X1 i_257_36_16 (.A1(n_257_36_15), .A2(n_257), .ZN(n_257_36_16));
   NOR2_X1 i_257_36_17 (.A1(n_257_36_16), .A2(n_257_36_5), .ZN(n_257_36_17));
   NAND2_X1 i_257_36_18 (.A1(CPU_Bus[1]), .A2(n_257_36_17), .ZN(n_257_36_18));
   NOR2_X1 i_257_36_19 (.A1(n_257_36_9), .A2(n_256), .ZN(n_257_36_19));
   NAND2_X1 i_257_36_20 (.A1(n_257_36_19), .A2(n_257), .ZN(n_257_36_20));
   NOR2_X1 i_257_36_21 (.A1(n_257_36_20), .A2(n_257_36_5), .ZN(n_257_36_21));
   NAND2_X1 i_257_36_22 (.A1(CPU_Bus[31]), .A2(n_257_36_21), .ZN(n_257_36_22));
   NAND2_X1 i_257_36_23 (.A1(n_257_36_18), .A2(n_257_36_22), .ZN(n_257_36_23));
   NOR2_X1 i_257_36_24 (.A1(n_257_36_14), .A2(n_257_36_23), .ZN(n_257_36_24));
   INV_X1 i_257_36_25 (.A(n_257), .ZN(n_257_36_25));
   NAND2_X1 i_257_36_26 (.A1(n_257_36_3), .A2(n_257_36_25), .ZN(n_257_36_26));
   NOR2_X1 i_257_36_27 (.A1(n_257_36_26), .A2(n_257_36_5), .ZN(n_257_36_27));
   NAND2_X1 i_257_36_28 (.A1(CPU_Bus[29]), .A2(n_257_36_27), .ZN(n_257_36_28));
   NAND2_X1 i_257_36_29 (.A1(n_257_36_10), .A2(n_257_36_25), .ZN(n_257_36_29));
   NOR2_X1 i_257_36_30 (.A1(n_257_36_29), .A2(n_257_36_5), .ZN(n_257_36_30));
   NAND2_X1 i_257_36_31 (.A1(CPU_Bus[27]), .A2(n_257_36_30), .ZN(n_257_36_31));
   NAND2_X1 i_257_36_32 (.A1(n_257_36_28), .A2(n_257_36_31), .ZN(n_257_36_32));
   NAND2_X1 i_257_36_33 (.A1(n_257_36_15), .A2(n_257_36_25), .ZN(n_257_36_33));
   NOR2_X1 i_257_36_34 (.A1(n_257_36_33), .A2(n_257_36_5), .ZN(n_257_36_34));
   NAND2_X1 i_257_36_35 (.A1(CPU_Bus[25]), .A2(n_257_36_34), .ZN(n_257_36_35));
   NAND2_X1 i_257_36_36 (.A1(n_257_36_19), .A2(n_257_36_25), .ZN(n_257_36_36));
   NOR2_X1 i_257_36_37 (.A1(n_257_36_36), .A2(n_257_36_5), .ZN(n_257_36_37));
   NAND2_X1 i_257_36_38 (.A1(CPU_Bus[23]), .A2(n_257_36_37), .ZN(n_257_36_38));
   NAND2_X1 i_257_36_39 (.A1(n_257_36_35), .A2(n_257_36_38), .ZN(n_257_36_39));
   NOR2_X1 i_257_36_40 (.A1(n_257_36_32), .A2(n_257_36_39), .ZN(n_257_36_40));
   NAND2_X1 i_257_36_41 (.A1(n_257_36_24), .A2(n_257_36_40), .ZN(n_257_36_41));
   NOR2_X1 i_257_36_42 (.A1(n_257_36_4), .A2(n_258), .ZN(n_257_36_42));
   NAND2_X1 i_257_36_43 (.A1(CPU_Bus[21]), .A2(n_257_36_42), .ZN(n_257_36_43));
   NOR2_X1 i_257_36_44 (.A1(n_257_36_11), .A2(n_258), .ZN(n_257_36_44));
   NAND2_X1 i_257_36_45 (.A1(CPU_Bus[19]), .A2(n_257_36_44), .ZN(n_257_36_45));
   NAND2_X1 i_257_36_46 (.A1(n_257_36_43), .A2(n_257_36_45), .ZN(n_257_36_46));
   NOR2_X1 i_257_36_47 (.A1(n_257_36_16), .A2(n_258), .ZN(n_257_36_47));
   NAND2_X1 i_257_36_48 (.A1(CPU_Bus[17]), .A2(n_257_36_47), .ZN(n_257_36_48));
   NOR2_X1 i_257_36_49 (.A1(n_257_36_20), .A2(n_258), .ZN(n_257_36_49));
   NAND2_X1 i_257_36_50 (.A1(CPU_Bus[15]), .A2(n_257_36_49), .ZN(n_257_36_50));
   NAND2_X1 i_257_36_51 (.A1(n_257_36_48), .A2(n_257_36_50), .ZN(n_257_36_51));
   NOR2_X1 i_257_36_52 (.A1(n_257_36_46), .A2(n_257_36_51), .ZN(n_257_36_52));
   NOR2_X1 i_257_36_53 (.A1(n_257_36_26), .A2(n_258), .ZN(n_257_36_53));
   NAND2_X1 i_257_36_54 (.A1(CPU_Bus[13]), .A2(n_257_36_53), .ZN(n_257_36_54));
   NOR2_X1 i_257_36_55 (.A1(n_257_36_29), .A2(n_258), .ZN(n_257_36_55));
   NAND2_X1 i_257_36_56 (.A1(CPU_Bus[11]), .A2(n_257_36_55), .ZN(n_257_36_56));
   NAND2_X1 i_257_36_57 (.A1(n_257_36_54), .A2(n_257_36_56), .ZN(n_257_36_57));
   NOR2_X1 i_257_36_58 (.A1(n_257_36_33), .A2(n_258), .ZN(n_257_36_58));
   NAND2_X1 i_257_36_59 (.A1(CPU_Bus[9]), .A2(n_257_36_58), .ZN(n_257_36_59));
   NOR2_X1 i_257_36_60 (.A1(n_257_36_36), .A2(n_258), .ZN(n_257_36_60));
   NAND2_X1 i_257_36_61 (.A1(CPU_Bus[7]), .A2(n_257_36_60), .ZN(n_257_36_61));
   NAND2_X1 i_257_36_62 (.A1(n_257_36_59), .A2(n_257_36_61), .ZN(n_257_36_62));
   NOR2_X1 i_257_36_63 (.A1(n_257_36_57), .A2(n_257_36_62), .ZN(n_257_36_63));
   NAND2_X1 i_257_36_64 (.A1(n_257_36_52), .A2(n_257_36_63), .ZN(n_257_36_64));
   NOR2_X1 i_257_36_65 (.A1(n_257_36_41), .A2(n_257_36_64), .ZN(n_257_36_65));
   NAND2_X1 i_257_36_66 (.A1(n_257_36_8), .A2(n_254), .ZN(n_257_36_66));
   NOR2_X1 i_257_36_67 (.A1(n_257_36_66), .A2(n_257_36_2), .ZN(n_257_36_67));
   NAND2_X1 i_257_36_68 (.A1(n_257_36_67), .A2(n_257), .ZN(n_257_36_68));
   NOR2_X1 i_257_36_69 (.A1(n_257_36_68), .A2(n_257_36_5), .ZN(n_257_36_69));
   NAND2_X1 i_257_36_70 (.A1(CPU_Bus[4]), .A2(n_257_36_69), .ZN(n_257_36_70));
   NOR2_X1 i_257_36_71 (.A1(n_257_36_66), .A2(n_256), .ZN(n_257_36_71));
   NAND2_X1 i_257_36_72 (.A1(n_257_36_71), .A2(n_257), .ZN(n_257_36_72));
   NOR2_X1 i_257_36_73 (.A1(n_257_36_72), .A2(n_257_36_5), .ZN(n_257_36_73));
   NAND2_X1 i_257_36_74 (.A1(CPU_Bus[0]), .A2(n_257_36_73), .ZN(n_257_36_74));
   NAND2_X1 i_257_36_75 (.A1(n_257_36_70), .A2(n_257_36_74), .ZN(n_257_36_75));
   NAND2_X1 i_257_36_76 (.A1(n_257_36_67), .A2(n_257_36_25), .ZN(n_257_36_76));
   NOR2_X1 i_257_36_77 (.A1(n_257_36_76), .A2(n_257_36_5), .ZN(n_257_36_77));
   NAND2_X1 i_257_36_78 (.A1(CPU_Bus[28]), .A2(n_257_36_77), .ZN(n_257_36_78));
   NAND2_X1 i_257_36_79 (.A1(n_257_36_71), .A2(n_257_36_25), .ZN(n_257_36_79));
   NOR2_X1 i_257_36_80 (.A1(n_257_36_79), .A2(n_257_36_5), .ZN(n_257_36_80));
   NAND2_X1 i_257_36_81 (.A1(CPU_Bus[24]), .A2(n_257_36_80), .ZN(n_257_36_81));
   NAND2_X1 i_257_36_82 (.A1(n_257_36_78), .A2(n_257_36_81), .ZN(n_257_36_82));
   NOR2_X1 i_257_36_83 (.A1(n_257_36_75), .A2(n_257_36_82), .ZN(n_257_36_83));
   NOR2_X1 i_257_36_84 (.A1(n_257_36_68), .A2(n_258), .ZN(n_257_36_84));
   NAND2_X1 i_257_36_85 (.A1(CPU_Bus[20]), .A2(n_257_36_84), .ZN(n_257_36_85));
   NOR2_X1 i_257_36_86 (.A1(n_257_36_72), .A2(n_258), .ZN(n_257_36_86));
   NAND2_X1 i_257_36_87 (.A1(CPU_Bus[16]), .A2(n_257_36_86), .ZN(n_257_36_87));
   NAND2_X1 i_257_36_88 (.A1(n_257_36_85), .A2(n_257_36_87), .ZN(n_257_36_88));
   NOR2_X1 i_257_36_89 (.A1(n_257_36_76), .A2(n_258), .ZN(n_257_36_89));
   NAND2_X1 i_257_36_90 (.A1(CPU_Bus[12]), .A2(n_257_36_89), .ZN(n_257_36_90));
   NOR2_X1 i_257_36_91 (.A1(n_257_36_79), .A2(n_258), .ZN(n_257_36_91));
   NAND2_X1 i_257_36_92 (.A1(CPU_Bus[8]), .A2(n_257_36_91), .ZN(n_257_36_92));
   NAND2_X1 i_257_36_93 (.A1(n_257_36_90), .A2(n_257_36_92), .ZN(n_257_36_93));
   NOR2_X1 i_257_36_94 (.A1(n_257_36_88), .A2(n_257_36_93), .ZN(n_257_36_94));
   NAND2_X1 i_257_36_95 (.A1(n_257_36_83), .A2(n_257_36_94), .ZN(n_257_36_95));
   NAND2_X1 i_257_36_96 (.A1(n_254), .A2(n_255), .ZN(n_257_36_96));
   NOR2_X1 i_257_36_97 (.A1(n_257_36_96), .A2(n_257_36_2), .ZN(n_257_36_97));
   NAND2_X1 i_257_36_98 (.A1(n_257_36_97), .A2(n_257), .ZN(n_257_36_98));
   NOR2_X1 i_257_36_99 (.A1(n_257_36_98), .A2(n_257_36_5), .ZN(n_257_36_99));
   NAND2_X1 i_257_36_100 (.A1(CPU_Bus[6]), .A2(n_257_36_99), .ZN(n_257_36_100));
   NOR2_X1 i_257_36_101 (.A1(n_257_36_96), .A2(n_256), .ZN(n_257_36_101));
   NAND2_X1 i_257_36_102 (.A1(n_257_36_101), .A2(n_257), .ZN(n_257_36_102));
   NOR2_X1 i_257_36_103 (.A1(n_257_36_102), .A2(n_257_36_5), .ZN(n_257_36_103));
   NAND2_X1 i_257_36_104 (.A1(CPU_Bus[2]), .A2(n_257_36_103), .ZN(n_257_36_104));
   NAND2_X1 i_257_36_105 (.A1(n_257_36_100), .A2(n_257_36_104), .ZN(n_257_36_105));
   NAND2_X1 i_257_36_106 (.A1(n_257_36_97), .A2(n_257_36_25), .ZN(n_257_36_106));
   NOR2_X1 i_257_36_107 (.A1(n_257_36_106), .A2(n_257_36_5), .ZN(n_257_36_107));
   NAND2_X1 i_257_36_108 (.A1(CPU_Bus[30]), .A2(n_257_36_107), .ZN(n_257_36_108));
   NAND2_X1 i_257_36_109 (.A1(n_257_36_101), .A2(n_257_36_25), .ZN(n_257_36_109));
   NOR2_X1 i_257_36_110 (.A1(n_257_36_109), .A2(n_257_36_5), .ZN(n_257_36_110));
   NAND2_X1 i_257_36_111 (.A1(CPU_Bus[26]), .A2(n_257_36_110), .ZN(n_257_36_111));
   NAND2_X1 i_257_36_112 (.A1(n_257_36_108), .A2(n_257_36_111), .ZN(n_257_36_112));
   NOR2_X1 i_257_36_113 (.A1(n_257_36_105), .A2(n_257_36_112), .ZN(n_257_36_113));
   NOR2_X1 i_257_36_114 (.A1(n_257_36_98), .A2(n_258), .ZN(n_257_36_114));
   NAND2_X1 i_257_36_115 (.A1(CPU_Bus[22]), .A2(n_257_36_114), .ZN(n_257_36_115));
   NOR2_X1 i_257_36_116 (.A1(n_257_36_102), .A2(n_258), .ZN(n_257_36_116));
   NAND2_X1 i_257_36_117 (.A1(CPU_Bus[18]), .A2(n_257_36_116), .ZN(n_257_36_117));
   NAND2_X1 i_257_36_118 (.A1(n_257_36_115), .A2(n_257_36_117), .ZN(n_257_36_118));
   NOR2_X1 i_257_36_119 (.A1(n_257_36_106), .A2(n_258), .ZN(n_257_36_119));
   NAND2_X1 i_257_36_120 (.A1(CPU_Bus[14]), .A2(n_257_36_119), .ZN(n_257_36_120));
   NOR2_X1 i_257_36_121 (.A1(n_257_36_109), .A2(n_258), .ZN(n_257_36_121));
   NAND2_X1 i_257_36_122 (.A1(CPU_Bus[10]), .A2(n_257_36_121), .ZN(n_257_36_122));
   NAND2_X1 i_257_36_123 (.A1(n_257_36_120), .A2(n_257_36_122), .ZN(n_257_36_123));
   NOR2_X1 i_257_36_124 (.A1(n_257_36_118), .A2(n_257_36_123), .ZN(n_257_36_124));
   NAND2_X1 i_257_36_125 (.A1(n_257_36_113), .A2(n_257_36_124), .ZN(n_257_36_125));
   NOR2_X1 i_257_36_126 (.A1(n_257_36_95), .A2(n_257_36_125), .ZN(n_257_36_126));
   NAND2_X1 i_257_36_127 (.A1(n_257_36_65), .A2(n_257_36_126), .ZN(n_257_225));
   datapath__1_361 i_257_37 (.PacketSize(PacketSize), .p_0({n_257_231, uc_360, 
      uc_361, uc_362, uc_363, uc_364, uc_365, uc_366, uc_367, uc_368, uc_369, 
      uc_370, uc_371, uc_372, uc_373, uc_374, uc_375, uc_376, uc_377, uc_378, 
      uc_379, uc_380, uc_381, uc_382, uc_383, uc_384, n_257_230, n_257_229, 
      n_257_228, n_257_227, n_257_226, uc_385}));
   datapath__1_362 i_257_38 (.p_0({uc_386, uc_387, uc_388, uc_389, uc_390, 
      uc_391, uc_392, uc_393, uc_394, uc_395, uc_396, uc_397, uc_398, uc_399, 
      uc_400, uc_401, uc_402, uc_403, uc_404, uc_405, uc_406, uc_407, uc_408, 
      uc_409, uc_410, n_257_231, n_257_230, n_257_229, n_257_228, n_257_227, 
      n_257_226, n_151}), .p_1({n_257_263, n_257_262, n_257_261, n_257_260, 
      n_257_259, n_257_258, n_257_257, n_257_256, n_257_255, n_257_254, 
      n_257_253, n_257_252, n_257_251, n_257_250, n_257_249, n_257_248, 
      n_257_247, n_257_246, n_257_245, n_257_244, n_257_243, n_257_242, 
      n_257_241, n_257_240, n_257_239, n_257_238, n_257_237, n_257_236, 
      n_257_235, n_257_234, n_257_233, n_257_232}));
   INV_X1 i_257_39_0 (.A(n_254), .ZN(n_257_39_0));
   NAND2_X1 i_257_39_1 (.A1(n_257_39_0), .A2(n_255), .ZN(n_257_39_1));
   INV_X1 i_257_39_2 (.A(n_256), .ZN(n_257_39_2));
   NOR2_X1 i_257_39_3 (.A1(n_257_39_1), .A2(n_257_39_2), .ZN(n_257_39_3));
   NAND2_X1 i_257_39_4 (.A1(n_257_39_3), .A2(n_257), .ZN(n_257_39_4));
   INV_X1 i_257_39_5 (.A(n_258), .ZN(n_257_39_5));
   NOR2_X1 i_257_39_6 (.A1(n_257_39_4), .A2(n_257_39_5), .ZN(n_257_39_6));
   NAND2_X1 i_257_39_7 (.A1(CPU_Bus[4]), .A2(n_257_39_6), .ZN(n_257_39_7));
   INV_X1 i_257_39_8 (.A(n_255), .ZN(n_257_39_8));
   NAND2_X1 i_257_39_9 (.A1(n_257_39_0), .A2(n_257_39_8), .ZN(n_257_39_9));
   NOR2_X1 i_257_39_10 (.A1(n_257_39_9), .A2(n_257_39_2), .ZN(n_257_39_10));
   NAND2_X1 i_257_39_11 (.A1(n_257_39_10), .A2(n_257), .ZN(n_257_39_11));
   NOR2_X1 i_257_39_12 (.A1(n_257_39_11), .A2(n_257_39_5), .ZN(n_257_39_12));
   NAND2_X1 i_257_39_13 (.A1(CPU_Bus[2]), .A2(n_257_39_12), .ZN(n_257_39_13));
   NAND2_X1 i_257_39_14 (.A1(n_257_39_7), .A2(n_257_39_13), .ZN(n_257_39_14));
   NOR2_X1 i_257_39_15 (.A1(n_257_39_1), .A2(n_256), .ZN(n_257_39_15));
   NAND2_X1 i_257_39_16 (.A1(n_257_39_15), .A2(n_257), .ZN(n_257_39_16));
   NOR2_X1 i_257_39_17 (.A1(n_257_39_16), .A2(n_257_39_5), .ZN(n_257_39_17));
   NAND2_X1 i_257_39_18 (.A1(CPU_Bus[0]), .A2(n_257_39_17), .ZN(n_257_39_18));
   NOR2_X1 i_257_39_19 (.A1(n_257_39_9), .A2(n_256), .ZN(n_257_39_19));
   NAND2_X1 i_257_39_20 (.A1(n_257_39_19), .A2(n_257), .ZN(n_257_39_20));
   NOR2_X1 i_257_39_21 (.A1(n_257_39_20), .A2(n_257_39_5), .ZN(n_257_39_21));
   NAND2_X1 i_257_39_22 (.A1(CPU_Bus[30]), .A2(n_257_39_21), .ZN(n_257_39_22));
   NAND2_X1 i_257_39_23 (.A1(n_257_39_18), .A2(n_257_39_22), .ZN(n_257_39_23));
   NOR2_X1 i_257_39_24 (.A1(n_257_39_14), .A2(n_257_39_23), .ZN(n_257_39_24));
   INV_X1 i_257_39_25 (.A(n_257), .ZN(n_257_39_25));
   NAND2_X1 i_257_39_26 (.A1(n_257_39_3), .A2(n_257_39_25), .ZN(n_257_39_26));
   NOR2_X1 i_257_39_27 (.A1(n_257_39_26), .A2(n_257_39_5), .ZN(n_257_39_27));
   NAND2_X1 i_257_39_28 (.A1(CPU_Bus[28]), .A2(n_257_39_27), .ZN(n_257_39_28));
   NAND2_X1 i_257_39_29 (.A1(n_257_39_10), .A2(n_257_39_25), .ZN(n_257_39_29));
   NOR2_X1 i_257_39_30 (.A1(n_257_39_29), .A2(n_257_39_5), .ZN(n_257_39_30));
   NAND2_X1 i_257_39_31 (.A1(CPU_Bus[26]), .A2(n_257_39_30), .ZN(n_257_39_31));
   NAND2_X1 i_257_39_32 (.A1(n_257_39_28), .A2(n_257_39_31), .ZN(n_257_39_32));
   NAND2_X1 i_257_39_33 (.A1(n_257_39_15), .A2(n_257_39_25), .ZN(n_257_39_33));
   NOR2_X1 i_257_39_34 (.A1(n_257_39_33), .A2(n_257_39_5), .ZN(n_257_39_34));
   NAND2_X1 i_257_39_35 (.A1(CPU_Bus[24]), .A2(n_257_39_34), .ZN(n_257_39_35));
   NAND2_X1 i_257_39_36 (.A1(n_257_39_19), .A2(n_257_39_25), .ZN(n_257_39_36));
   NOR2_X1 i_257_39_37 (.A1(n_257_39_36), .A2(n_257_39_5), .ZN(n_257_39_37));
   NAND2_X1 i_257_39_38 (.A1(CPU_Bus[22]), .A2(n_257_39_37), .ZN(n_257_39_38));
   NAND2_X1 i_257_39_39 (.A1(n_257_39_35), .A2(n_257_39_38), .ZN(n_257_39_39));
   NOR2_X1 i_257_39_40 (.A1(n_257_39_32), .A2(n_257_39_39), .ZN(n_257_39_40));
   NAND2_X1 i_257_39_41 (.A1(n_257_39_24), .A2(n_257_39_40), .ZN(n_257_39_41));
   NOR2_X1 i_257_39_42 (.A1(n_257_39_4), .A2(n_258), .ZN(n_257_39_42));
   NAND2_X1 i_257_39_43 (.A1(CPU_Bus[20]), .A2(n_257_39_42), .ZN(n_257_39_43));
   NOR2_X1 i_257_39_44 (.A1(n_257_39_11), .A2(n_258), .ZN(n_257_39_44));
   NAND2_X1 i_257_39_45 (.A1(CPU_Bus[18]), .A2(n_257_39_44), .ZN(n_257_39_45));
   NAND2_X1 i_257_39_46 (.A1(n_257_39_43), .A2(n_257_39_45), .ZN(n_257_39_46));
   NOR2_X1 i_257_39_47 (.A1(n_257_39_16), .A2(n_258), .ZN(n_257_39_47));
   NAND2_X1 i_257_39_48 (.A1(CPU_Bus[16]), .A2(n_257_39_47), .ZN(n_257_39_48));
   NOR2_X1 i_257_39_49 (.A1(n_257_39_20), .A2(n_258), .ZN(n_257_39_49));
   NAND2_X1 i_257_39_50 (.A1(CPU_Bus[14]), .A2(n_257_39_49), .ZN(n_257_39_50));
   NAND2_X1 i_257_39_51 (.A1(n_257_39_48), .A2(n_257_39_50), .ZN(n_257_39_51));
   NOR2_X1 i_257_39_52 (.A1(n_257_39_46), .A2(n_257_39_51), .ZN(n_257_39_52));
   NOR2_X1 i_257_39_53 (.A1(n_257_39_26), .A2(n_258), .ZN(n_257_39_53));
   NAND2_X1 i_257_39_54 (.A1(CPU_Bus[12]), .A2(n_257_39_53), .ZN(n_257_39_54));
   NOR2_X1 i_257_39_55 (.A1(n_257_39_29), .A2(n_258), .ZN(n_257_39_55));
   NAND2_X1 i_257_39_56 (.A1(CPU_Bus[10]), .A2(n_257_39_55), .ZN(n_257_39_56));
   NAND2_X1 i_257_39_57 (.A1(n_257_39_54), .A2(n_257_39_56), .ZN(n_257_39_57));
   NOR2_X1 i_257_39_58 (.A1(n_257_39_33), .A2(n_258), .ZN(n_257_39_58));
   NAND2_X1 i_257_39_59 (.A1(CPU_Bus[8]), .A2(n_257_39_58), .ZN(n_257_39_59));
   NOR2_X1 i_257_39_60 (.A1(n_257_39_36), .A2(n_258), .ZN(n_257_39_60));
   NAND2_X1 i_257_39_61 (.A1(CPU_Bus[6]), .A2(n_257_39_60), .ZN(n_257_39_61));
   NAND2_X1 i_257_39_62 (.A1(n_257_39_59), .A2(n_257_39_61), .ZN(n_257_39_62));
   NOR2_X1 i_257_39_63 (.A1(n_257_39_57), .A2(n_257_39_62), .ZN(n_257_39_63));
   NAND2_X1 i_257_39_64 (.A1(n_257_39_52), .A2(n_257_39_63), .ZN(n_257_39_64));
   NOR2_X1 i_257_39_65 (.A1(n_257_39_41), .A2(n_257_39_64), .ZN(n_257_39_65));
   NAND2_X1 i_257_39_66 (.A1(n_257_39_8), .A2(n_254), .ZN(n_257_39_66));
   NOR2_X1 i_257_39_67 (.A1(n_257_39_66), .A2(n_257_39_2), .ZN(n_257_39_67));
   NAND2_X1 i_257_39_68 (.A1(n_257_39_67), .A2(n_257), .ZN(n_257_39_68));
   NOR2_X1 i_257_39_69 (.A1(n_257_39_68), .A2(n_257_39_5), .ZN(n_257_39_69));
   NAND2_X1 i_257_39_70 (.A1(CPU_Bus[3]), .A2(n_257_39_69), .ZN(n_257_39_70));
   NOR2_X1 i_257_39_71 (.A1(n_257_39_66), .A2(n_256), .ZN(n_257_39_71));
   NAND2_X1 i_257_39_72 (.A1(n_257_39_71), .A2(n_257), .ZN(n_257_39_72));
   NOR2_X1 i_257_39_73 (.A1(n_257_39_72), .A2(n_257_39_5), .ZN(n_257_39_73));
   NAND2_X1 i_257_39_74 (.A1(CPU_Bus[31]), .A2(n_257_39_73), .ZN(n_257_39_74));
   NAND2_X1 i_257_39_75 (.A1(n_257_39_70), .A2(n_257_39_74), .ZN(n_257_39_75));
   NAND2_X1 i_257_39_76 (.A1(n_257_39_67), .A2(n_257_39_25), .ZN(n_257_39_76));
   NOR2_X1 i_257_39_77 (.A1(n_257_39_76), .A2(n_257_39_5), .ZN(n_257_39_77));
   NAND2_X1 i_257_39_78 (.A1(CPU_Bus[27]), .A2(n_257_39_77), .ZN(n_257_39_78));
   NAND2_X1 i_257_39_79 (.A1(n_257_39_71), .A2(n_257_39_25), .ZN(n_257_39_79));
   NOR2_X1 i_257_39_80 (.A1(n_257_39_79), .A2(n_257_39_5), .ZN(n_257_39_80));
   NAND2_X1 i_257_39_81 (.A1(CPU_Bus[23]), .A2(n_257_39_80), .ZN(n_257_39_81));
   NAND2_X1 i_257_39_82 (.A1(n_257_39_78), .A2(n_257_39_81), .ZN(n_257_39_82));
   NOR2_X1 i_257_39_83 (.A1(n_257_39_75), .A2(n_257_39_82), .ZN(n_257_39_83));
   NOR2_X1 i_257_39_84 (.A1(n_257_39_68), .A2(n_258), .ZN(n_257_39_84));
   NAND2_X1 i_257_39_85 (.A1(CPU_Bus[19]), .A2(n_257_39_84), .ZN(n_257_39_85));
   NOR2_X1 i_257_39_86 (.A1(n_257_39_72), .A2(n_258), .ZN(n_257_39_86));
   NAND2_X1 i_257_39_87 (.A1(CPU_Bus[15]), .A2(n_257_39_86), .ZN(n_257_39_87));
   NAND2_X1 i_257_39_88 (.A1(n_257_39_85), .A2(n_257_39_87), .ZN(n_257_39_88));
   NOR2_X1 i_257_39_89 (.A1(n_257_39_76), .A2(n_258), .ZN(n_257_39_89));
   NAND2_X1 i_257_39_90 (.A1(CPU_Bus[11]), .A2(n_257_39_89), .ZN(n_257_39_90));
   NOR2_X1 i_257_39_91 (.A1(n_257_39_79), .A2(n_258), .ZN(n_257_39_91));
   NAND2_X1 i_257_39_92 (.A1(CPU_Bus[7]), .A2(n_257_39_91), .ZN(n_257_39_92));
   NAND2_X1 i_257_39_93 (.A1(n_257_39_90), .A2(n_257_39_92), .ZN(n_257_39_93));
   NOR2_X1 i_257_39_94 (.A1(n_257_39_88), .A2(n_257_39_93), .ZN(n_257_39_94));
   NAND2_X1 i_257_39_95 (.A1(n_257_39_83), .A2(n_257_39_94), .ZN(n_257_39_95));
   NAND2_X1 i_257_39_96 (.A1(n_254), .A2(n_255), .ZN(n_257_39_96));
   NOR2_X1 i_257_39_97 (.A1(n_257_39_96), .A2(n_257_39_2), .ZN(n_257_39_97));
   NAND2_X1 i_257_39_98 (.A1(n_257_39_97), .A2(n_257), .ZN(n_257_39_98));
   NOR2_X1 i_257_39_99 (.A1(n_257_39_98), .A2(n_257_39_5), .ZN(n_257_39_99));
   NAND2_X1 i_257_39_100 (.A1(CPU_Bus[5]), .A2(n_257_39_99), .ZN(n_257_39_100));
   NOR2_X1 i_257_39_101 (.A1(n_257_39_96), .A2(n_256), .ZN(n_257_39_101));
   NAND2_X1 i_257_39_102 (.A1(n_257_39_101), .A2(n_257), .ZN(n_257_39_102));
   NOR2_X1 i_257_39_103 (.A1(n_257_39_102), .A2(n_257_39_5), .ZN(n_257_39_103));
   NAND2_X1 i_257_39_104 (.A1(CPU_Bus[1]), .A2(n_257_39_103), .ZN(n_257_39_104));
   NAND2_X1 i_257_39_105 (.A1(n_257_39_100), .A2(n_257_39_104), .ZN(n_257_39_105));
   NAND2_X1 i_257_39_106 (.A1(n_257_39_97), .A2(n_257_39_25), .ZN(n_257_39_106));
   NOR2_X1 i_257_39_107 (.A1(n_257_39_106), .A2(n_257_39_5), .ZN(n_257_39_107));
   NAND2_X1 i_257_39_108 (.A1(CPU_Bus[29]), .A2(n_257_39_107), .ZN(n_257_39_108));
   NAND2_X1 i_257_39_109 (.A1(n_257_39_101), .A2(n_257_39_25), .ZN(n_257_39_109));
   NOR2_X1 i_257_39_110 (.A1(n_257_39_109), .A2(n_257_39_5), .ZN(n_257_39_110));
   NAND2_X1 i_257_39_111 (.A1(CPU_Bus[25]), .A2(n_257_39_110), .ZN(n_257_39_111));
   NAND2_X1 i_257_39_112 (.A1(n_257_39_108), .A2(n_257_39_111), .ZN(n_257_39_112));
   NOR2_X1 i_257_39_113 (.A1(n_257_39_105), .A2(n_257_39_112), .ZN(n_257_39_113));
   NOR2_X1 i_257_39_114 (.A1(n_257_39_98), .A2(n_258), .ZN(n_257_39_114));
   NAND2_X1 i_257_39_115 (.A1(CPU_Bus[21]), .A2(n_257_39_114), .ZN(n_257_39_115));
   NOR2_X1 i_257_39_116 (.A1(n_257_39_102), .A2(n_258), .ZN(n_257_39_116));
   NAND2_X1 i_257_39_117 (.A1(CPU_Bus[17]), .A2(n_257_39_116), .ZN(n_257_39_117));
   NAND2_X1 i_257_39_118 (.A1(n_257_39_115), .A2(n_257_39_117), .ZN(n_257_39_118));
   NOR2_X1 i_257_39_119 (.A1(n_257_39_106), .A2(n_258), .ZN(n_257_39_119));
   NAND2_X1 i_257_39_120 (.A1(CPU_Bus[13]), .A2(n_257_39_119), .ZN(n_257_39_120));
   NOR2_X1 i_257_39_121 (.A1(n_257_39_109), .A2(n_258), .ZN(n_257_39_121));
   NAND2_X1 i_257_39_122 (.A1(CPU_Bus[9]), .A2(n_257_39_121), .ZN(n_257_39_122));
   NAND2_X1 i_257_39_123 (.A1(n_257_39_120), .A2(n_257_39_122), .ZN(n_257_39_123));
   NOR2_X1 i_257_39_124 (.A1(n_257_39_118), .A2(n_257_39_123), .ZN(n_257_39_124));
   NAND2_X1 i_257_39_125 (.A1(n_257_39_113), .A2(n_257_39_124), .ZN(n_257_39_125));
   NOR2_X1 i_257_39_126 (.A1(n_257_39_95), .A2(n_257_39_125), .ZN(n_257_39_126));
   NAND2_X1 i_257_39_127 (.A1(n_257_39_65), .A2(n_257_39_126), .ZN(n_257_264));
   INV_X1 i_257_40_0 (.A(n_254), .ZN(n_257_40_0));
   NAND2_X1 i_257_40_1 (.A1(n_257_40_0), .A2(n_255), .ZN(n_257_40_1));
   INV_X1 i_257_40_2 (.A(n_256), .ZN(n_257_40_2));
   NOR2_X1 i_257_40_3 (.A1(n_257_40_1), .A2(n_257_40_2), .ZN(n_257_40_3));
   NAND2_X1 i_257_40_4 (.A1(n_257_40_3), .A2(n_257), .ZN(n_257_40_4));
   INV_X1 i_257_40_5 (.A(n_258), .ZN(n_257_40_5));
   NOR2_X1 i_257_40_6 (.A1(n_257_40_4), .A2(n_257_40_5), .ZN(n_257_40_6));
   NAND2_X1 i_257_40_7 (.A1(CPU_Bus[3]), .A2(n_257_40_6), .ZN(n_257_40_7));
   INV_X1 i_257_40_8 (.A(n_255), .ZN(n_257_40_8));
   NAND2_X1 i_257_40_9 (.A1(n_257_40_0), .A2(n_257_40_8), .ZN(n_257_40_9));
   NOR2_X1 i_257_40_10 (.A1(n_257_40_9), .A2(n_257_40_2), .ZN(n_257_40_10));
   NAND2_X1 i_257_40_11 (.A1(n_257_40_10), .A2(n_257), .ZN(n_257_40_11));
   NOR2_X1 i_257_40_12 (.A1(n_257_40_11), .A2(n_257_40_5), .ZN(n_257_40_12));
   NAND2_X1 i_257_40_13 (.A1(CPU_Bus[1]), .A2(n_257_40_12), .ZN(n_257_40_13));
   NAND2_X1 i_257_40_14 (.A1(n_257_40_7), .A2(n_257_40_13), .ZN(n_257_40_14));
   NOR2_X1 i_257_40_15 (.A1(n_257_40_1), .A2(n_256), .ZN(n_257_40_15));
   NAND2_X1 i_257_40_16 (.A1(n_257_40_15), .A2(n_257), .ZN(n_257_40_16));
   NOR2_X1 i_257_40_17 (.A1(n_257_40_16), .A2(n_257_40_5), .ZN(n_257_40_17));
   NAND2_X1 i_257_40_18 (.A1(CPU_Bus[31]), .A2(n_257_40_17), .ZN(n_257_40_18));
   NOR2_X1 i_257_40_19 (.A1(n_257_40_9), .A2(n_256), .ZN(n_257_40_19));
   NAND2_X1 i_257_40_20 (.A1(n_257_40_19), .A2(n_257), .ZN(n_257_40_20));
   NOR2_X1 i_257_40_21 (.A1(n_257_40_20), .A2(n_257_40_5), .ZN(n_257_40_21));
   NAND2_X1 i_257_40_22 (.A1(CPU_Bus[29]), .A2(n_257_40_21), .ZN(n_257_40_22));
   NAND2_X1 i_257_40_23 (.A1(n_257_40_18), .A2(n_257_40_22), .ZN(n_257_40_23));
   NOR2_X1 i_257_40_24 (.A1(n_257_40_14), .A2(n_257_40_23), .ZN(n_257_40_24));
   INV_X1 i_257_40_25 (.A(n_257), .ZN(n_257_40_25));
   NAND2_X1 i_257_40_26 (.A1(n_257_40_3), .A2(n_257_40_25), .ZN(n_257_40_26));
   NOR2_X1 i_257_40_27 (.A1(n_257_40_26), .A2(n_257_40_5), .ZN(n_257_40_27));
   NAND2_X1 i_257_40_28 (.A1(CPU_Bus[27]), .A2(n_257_40_27), .ZN(n_257_40_28));
   NAND2_X1 i_257_40_29 (.A1(n_257_40_10), .A2(n_257_40_25), .ZN(n_257_40_29));
   NOR2_X1 i_257_40_30 (.A1(n_257_40_29), .A2(n_257_40_5), .ZN(n_257_40_30));
   NAND2_X1 i_257_40_31 (.A1(CPU_Bus[25]), .A2(n_257_40_30), .ZN(n_257_40_31));
   NAND2_X1 i_257_40_32 (.A1(n_257_40_28), .A2(n_257_40_31), .ZN(n_257_40_32));
   NAND2_X1 i_257_40_33 (.A1(n_257_40_15), .A2(n_257_40_25), .ZN(n_257_40_33));
   NOR2_X1 i_257_40_34 (.A1(n_257_40_33), .A2(n_257_40_5), .ZN(n_257_40_34));
   NAND2_X1 i_257_40_35 (.A1(CPU_Bus[23]), .A2(n_257_40_34), .ZN(n_257_40_35));
   NAND2_X1 i_257_40_36 (.A1(n_257_40_19), .A2(n_257_40_25), .ZN(n_257_40_36));
   NOR2_X1 i_257_40_37 (.A1(n_257_40_36), .A2(n_257_40_5), .ZN(n_257_40_37));
   NAND2_X1 i_257_40_38 (.A1(CPU_Bus[21]), .A2(n_257_40_37), .ZN(n_257_40_38));
   NAND2_X1 i_257_40_39 (.A1(n_257_40_35), .A2(n_257_40_38), .ZN(n_257_40_39));
   NOR2_X1 i_257_40_40 (.A1(n_257_40_32), .A2(n_257_40_39), .ZN(n_257_40_40));
   NAND2_X1 i_257_40_41 (.A1(n_257_40_24), .A2(n_257_40_40), .ZN(n_257_40_41));
   NOR2_X1 i_257_40_42 (.A1(n_257_40_4), .A2(n_258), .ZN(n_257_40_42));
   NAND2_X1 i_257_40_43 (.A1(CPU_Bus[19]), .A2(n_257_40_42), .ZN(n_257_40_43));
   NOR2_X1 i_257_40_44 (.A1(n_257_40_11), .A2(n_258), .ZN(n_257_40_44));
   NAND2_X1 i_257_40_45 (.A1(CPU_Bus[17]), .A2(n_257_40_44), .ZN(n_257_40_45));
   NAND2_X1 i_257_40_46 (.A1(n_257_40_43), .A2(n_257_40_45), .ZN(n_257_40_46));
   NOR2_X1 i_257_40_47 (.A1(n_257_40_16), .A2(n_258), .ZN(n_257_40_47));
   NAND2_X1 i_257_40_48 (.A1(CPU_Bus[15]), .A2(n_257_40_47), .ZN(n_257_40_48));
   NOR2_X1 i_257_40_49 (.A1(n_257_40_20), .A2(n_258), .ZN(n_257_40_49));
   NAND2_X1 i_257_40_50 (.A1(CPU_Bus[13]), .A2(n_257_40_49), .ZN(n_257_40_50));
   NAND2_X1 i_257_40_51 (.A1(n_257_40_48), .A2(n_257_40_50), .ZN(n_257_40_51));
   NOR2_X1 i_257_40_52 (.A1(n_257_40_46), .A2(n_257_40_51), .ZN(n_257_40_52));
   NOR2_X1 i_257_40_53 (.A1(n_257_40_26), .A2(n_258), .ZN(n_257_40_53));
   NAND2_X1 i_257_40_54 (.A1(CPU_Bus[11]), .A2(n_257_40_53), .ZN(n_257_40_54));
   NOR2_X1 i_257_40_55 (.A1(n_257_40_29), .A2(n_258), .ZN(n_257_40_55));
   NAND2_X1 i_257_40_56 (.A1(CPU_Bus[9]), .A2(n_257_40_55), .ZN(n_257_40_56));
   NAND2_X1 i_257_40_57 (.A1(n_257_40_54), .A2(n_257_40_56), .ZN(n_257_40_57));
   NOR2_X1 i_257_40_58 (.A1(n_257_40_33), .A2(n_258), .ZN(n_257_40_58));
   NAND2_X1 i_257_40_59 (.A1(CPU_Bus[7]), .A2(n_257_40_58), .ZN(n_257_40_59));
   NOR2_X1 i_257_40_60 (.A1(n_257_40_36), .A2(n_258), .ZN(n_257_40_60));
   NAND2_X1 i_257_40_61 (.A1(CPU_Bus[5]), .A2(n_257_40_60), .ZN(n_257_40_61));
   NAND2_X1 i_257_40_62 (.A1(n_257_40_59), .A2(n_257_40_61), .ZN(n_257_40_62));
   NOR2_X1 i_257_40_63 (.A1(n_257_40_57), .A2(n_257_40_62), .ZN(n_257_40_63));
   NAND2_X1 i_257_40_64 (.A1(n_257_40_52), .A2(n_257_40_63), .ZN(n_257_40_64));
   NOR2_X1 i_257_40_65 (.A1(n_257_40_41), .A2(n_257_40_64), .ZN(n_257_40_65));
   NAND2_X1 i_257_40_66 (.A1(n_257_40_8), .A2(n_254), .ZN(n_257_40_66));
   NOR2_X1 i_257_40_67 (.A1(n_257_40_66), .A2(n_257_40_2), .ZN(n_257_40_67));
   NAND2_X1 i_257_40_68 (.A1(n_257_40_67), .A2(n_257), .ZN(n_257_40_68));
   NOR2_X1 i_257_40_69 (.A1(n_257_40_68), .A2(n_257_40_5), .ZN(n_257_40_69));
   NAND2_X1 i_257_40_70 (.A1(CPU_Bus[2]), .A2(n_257_40_69), .ZN(n_257_40_70));
   NOR2_X1 i_257_40_71 (.A1(n_257_40_66), .A2(n_256), .ZN(n_257_40_71));
   NAND2_X1 i_257_40_72 (.A1(n_257_40_71), .A2(n_257), .ZN(n_257_40_72));
   NOR2_X1 i_257_40_73 (.A1(n_257_40_72), .A2(n_257_40_5), .ZN(n_257_40_73));
   NAND2_X1 i_257_40_74 (.A1(CPU_Bus[30]), .A2(n_257_40_73), .ZN(n_257_40_74));
   NAND2_X1 i_257_40_75 (.A1(n_257_40_70), .A2(n_257_40_74), .ZN(n_257_40_75));
   NAND2_X1 i_257_40_76 (.A1(n_257_40_67), .A2(n_257_40_25), .ZN(n_257_40_76));
   NOR2_X1 i_257_40_77 (.A1(n_257_40_76), .A2(n_257_40_5), .ZN(n_257_40_77));
   NAND2_X1 i_257_40_78 (.A1(CPU_Bus[26]), .A2(n_257_40_77), .ZN(n_257_40_78));
   NAND2_X1 i_257_40_79 (.A1(n_257_40_71), .A2(n_257_40_25), .ZN(n_257_40_79));
   NOR2_X1 i_257_40_80 (.A1(n_257_40_79), .A2(n_257_40_5), .ZN(n_257_40_80));
   NAND2_X1 i_257_40_81 (.A1(CPU_Bus[22]), .A2(n_257_40_80), .ZN(n_257_40_81));
   NAND2_X1 i_257_40_82 (.A1(n_257_40_78), .A2(n_257_40_81), .ZN(n_257_40_82));
   NOR2_X1 i_257_40_83 (.A1(n_257_40_75), .A2(n_257_40_82), .ZN(n_257_40_83));
   NOR2_X1 i_257_40_84 (.A1(n_257_40_68), .A2(n_258), .ZN(n_257_40_84));
   NAND2_X1 i_257_40_85 (.A1(CPU_Bus[18]), .A2(n_257_40_84), .ZN(n_257_40_85));
   NOR2_X1 i_257_40_86 (.A1(n_257_40_72), .A2(n_258), .ZN(n_257_40_86));
   NAND2_X1 i_257_40_87 (.A1(CPU_Bus[14]), .A2(n_257_40_86), .ZN(n_257_40_87));
   NAND2_X1 i_257_40_88 (.A1(n_257_40_85), .A2(n_257_40_87), .ZN(n_257_40_88));
   NOR2_X1 i_257_40_89 (.A1(n_257_40_76), .A2(n_258), .ZN(n_257_40_89));
   NAND2_X1 i_257_40_90 (.A1(CPU_Bus[10]), .A2(n_257_40_89), .ZN(n_257_40_90));
   NOR2_X1 i_257_40_91 (.A1(n_257_40_79), .A2(n_258), .ZN(n_257_40_91));
   NAND2_X1 i_257_40_92 (.A1(CPU_Bus[6]), .A2(n_257_40_91), .ZN(n_257_40_92));
   NAND2_X1 i_257_40_93 (.A1(n_257_40_90), .A2(n_257_40_92), .ZN(n_257_40_93));
   NOR2_X1 i_257_40_94 (.A1(n_257_40_88), .A2(n_257_40_93), .ZN(n_257_40_94));
   NAND2_X1 i_257_40_95 (.A1(n_257_40_83), .A2(n_257_40_94), .ZN(n_257_40_95));
   NAND2_X1 i_257_40_96 (.A1(n_254), .A2(n_255), .ZN(n_257_40_96));
   NOR2_X1 i_257_40_97 (.A1(n_257_40_96), .A2(n_257_40_2), .ZN(n_257_40_97));
   NAND2_X1 i_257_40_98 (.A1(n_257_40_97), .A2(n_257), .ZN(n_257_40_98));
   NOR2_X1 i_257_40_99 (.A1(n_257_40_98), .A2(n_257_40_5), .ZN(n_257_40_99));
   NAND2_X1 i_257_40_100 (.A1(CPU_Bus[4]), .A2(n_257_40_99), .ZN(n_257_40_100));
   NOR2_X1 i_257_40_101 (.A1(n_257_40_96), .A2(n_256), .ZN(n_257_40_101));
   NAND2_X1 i_257_40_102 (.A1(n_257_40_101), .A2(n_257), .ZN(n_257_40_102));
   NOR2_X1 i_257_40_103 (.A1(n_257_40_102), .A2(n_257_40_5), .ZN(n_257_40_103));
   NAND2_X1 i_257_40_104 (.A1(CPU_Bus[0]), .A2(n_257_40_103), .ZN(n_257_40_104));
   NAND2_X1 i_257_40_105 (.A1(n_257_40_100), .A2(n_257_40_104), .ZN(n_257_40_105));
   NAND2_X1 i_257_40_106 (.A1(n_257_40_97), .A2(n_257_40_25), .ZN(n_257_40_106));
   NOR2_X1 i_257_40_107 (.A1(n_257_40_106), .A2(n_257_40_5), .ZN(n_257_40_107));
   NAND2_X1 i_257_40_108 (.A1(CPU_Bus[28]), .A2(n_257_40_107), .ZN(n_257_40_108));
   NAND2_X1 i_257_40_109 (.A1(n_257_40_101), .A2(n_257_40_25), .ZN(n_257_40_109));
   NOR2_X1 i_257_40_110 (.A1(n_257_40_109), .A2(n_257_40_5), .ZN(n_257_40_110));
   NAND2_X1 i_257_40_111 (.A1(CPU_Bus[24]), .A2(n_257_40_110), .ZN(n_257_40_111));
   NAND2_X1 i_257_40_112 (.A1(n_257_40_108), .A2(n_257_40_111), .ZN(n_257_40_112));
   NOR2_X1 i_257_40_113 (.A1(n_257_40_105), .A2(n_257_40_112), .ZN(n_257_40_113));
   NOR2_X1 i_257_40_114 (.A1(n_257_40_98), .A2(n_258), .ZN(n_257_40_114));
   NAND2_X1 i_257_40_115 (.A1(CPU_Bus[20]), .A2(n_257_40_114), .ZN(n_257_40_115));
   NOR2_X1 i_257_40_116 (.A1(n_257_40_102), .A2(n_258), .ZN(n_257_40_116));
   NAND2_X1 i_257_40_117 (.A1(CPU_Bus[16]), .A2(n_257_40_116), .ZN(n_257_40_117));
   NAND2_X1 i_257_40_118 (.A1(n_257_40_115), .A2(n_257_40_117), .ZN(n_257_40_118));
   NOR2_X1 i_257_40_119 (.A1(n_257_40_106), .A2(n_258), .ZN(n_257_40_119));
   NAND2_X1 i_257_40_120 (.A1(CPU_Bus[12]), .A2(n_257_40_119), .ZN(n_257_40_120));
   NOR2_X1 i_257_40_121 (.A1(n_257_40_109), .A2(n_258), .ZN(n_257_40_121));
   NAND2_X1 i_257_40_122 (.A1(CPU_Bus[8]), .A2(n_257_40_121), .ZN(n_257_40_122));
   NAND2_X1 i_257_40_123 (.A1(n_257_40_120), .A2(n_257_40_122), .ZN(n_257_40_123));
   NOR2_X1 i_257_40_124 (.A1(n_257_40_118), .A2(n_257_40_123), .ZN(n_257_40_124));
   NAND2_X1 i_257_40_125 (.A1(n_257_40_113), .A2(n_257_40_124), .ZN(n_257_40_125));
   NOR2_X1 i_257_40_126 (.A1(n_257_40_95), .A2(n_257_40_125), .ZN(n_257_40_126));
   NAND2_X1 i_257_40_127 (.A1(n_257_40_65), .A2(n_257_40_126), .ZN(n_257_265));
   datapath__1_366 i_257_41 (.PacketSize(PacketSize), .p_0({n_257_271, uc_411, 
      uc_412, uc_413, uc_414, uc_415, uc_416, uc_417, uc_418, uc_419, uc_420, 
      uc_421, uc_422, uc_423, uc_424, uc_425, uc_426, uc_427, uc_428, uc_429, 
      uc_430, uc_431, uc_432, uc_433, uc_434, uc_435, n_257_270, n_257_269, 
      n_257_268, n_257_267, n_257_266, uc_436}));
   datapath__1_367 i_257_42 (.p_0({uc_437, uc_438, uc_439, uc_440, uc_441, 
      uc_442, uc_443, uc_444, uc_445, uc_446, uc_447, uc_448, uc_449, uc_450, 
      uc_451, uc_452, uc_453, uc_454, uc_455, uc_456, uc_457, uc_458, uc_459, 
      uc_460, uc_461, n_257_271, n_257_270, n_257_269, n_257_268, n_257_267, 
      n_257_266, n_151}), .p_1({n_257_303, n_257_302, n_257_301, n_257_300, 
      n_257_299, n_257_298, n_257_297, n_257_296, n_257_295, n_257_294, 
      n_257_293, n_257_292, n_257_291, n_257_290, n_257_289, n_257_288, 
      n_257_287, n_257_286, n_257_285, n_257_284, n_257_283, n_257_282, 
      n_257_281, n_257_280, n_257_279, n_257_278, n_257_277, n_257_276, 
      n_257_275, n_257_274, n_257_273, n_257_272}));
   INV_X1 i_257_43_0 (.A(n_254), .ZN(n_257_43_0));
   NAND2_X1 i_257_43_1 (.A1(n_257_43_0), .A2(n_255), .ZN(n_257_43_1));
   INV_X1 i_257_43_2 (.A(n_256), .ZN(n_257_43_2));
   NOR2_X1 i_257_43_3 (.A1(n_257_43_1), .A2(n_257_43_2), .ZN(n_257_43_3));
   NAND2_X1 i_257_43_4 (.A1(n_257_43_3), .A2(n_257), .ZN(n_257_43_4));
   INV_X1 i_257_43_5 (.A(n_258), .ZN(n_257_43_5));
   NOR2_X1 i_257_43_6 (.A1(n_257_43_4), .A2(n_257_43_5), .ZN(n_257_43_6));
   NAND2_X1 i_257_43_7 (.A1(CPU_Bus[2]), .A2(n_257_43_6), .ZN(n_257_43_7));
   INV_X1 i_257_43_8 (.A(n_255), .ZN(n_257_43_8));
   NAND2_X1 i_257_43_9 (.A1(n_257_43_0), .A2(n_257_43_8), .ZN(n_257_43_9));
   NOR2_X1 i_257_43_10 (.A1(n_257_43_9), .A2(n_257_43_2), .ZN(n_257_43_10));
   NAND2_X1 i_257_43_11 (.A1(n_257_43_10), .A2(n_257), .ZN(n_257_43_11));
   NOR2_X1 i_257_43_12 (.A1(n_257_43_11), .A2(n_257_43_5), .ZN(n_257_43_12));
   NAND2_X1 i_257_43_13 (.A1(CPU_Bus[0]), .A2(n_257_43_12), .ZN(n_257_43_13));
   NAND2_X1 i_257_43_14 (.A1(n_257_43_7), .A2(n_257_43_13), .ZN(n_257_43_14));
   NOR2_X1 i_257_43_15 (.A1(n_257_43_1), .A2(n_256), .ZN(n_257_43_15));
   NAND2_X1 i_257_43_16 (.A1(n_257_43_15), .A2(n_257), .ZN(n_257_43_16));
   NOR2_X1 i_257_43_17 (.A1(n_257_43_16), .A2(n_257_43_5), .ZN(n_257_43_17));
   NAND2_X1 i_257_43_18 (.A1(CPU_Bus[30]), .A2(n_257_43_17), .ZN(n_257_43_18));
   NOR2_X1 i_257_43_19 (.A1(n_257_43_9), .A2(n_256), .ZN(n_257_43_19));
   NAND2_X1 i_257_43_20 (.A1(n_257_43_19), .A2(n_257), .ZN(n_257_43_20));
   NOR2_X1 i_257_43_21 (.A1(n_257_43_20), .A2(n_257_43_5), .ZN(n_257_43_21));
   NAND2_X1 i_257_43_22 (.A1(CPU_Bus[28]), .A2(n_257_43_21), .ZN(n_257_43_22));
   NAND2_X1 i_257_43_23 (.A1(n_257_43_18), .A2(n_257_43_22), .ZN(n_257_43_23));
   NOR2_X1 i_257_43_24 (.A1(n_257_43_14), .A2(n_257_43_23), .ZN(n_257_43_24));
   INV_X1 i_257_43_25 (.A(n_257), .ZN(n_257_43_25));
   NAND2_X1 i_257_43_26 (.A1(n_257_43_3), .A2(n_257_43_25), .ZN(n_257_43_26));
   NOR2_X1 i_257_43_27 (.A1(n_257_43_26), .A2(n_257_43_5), .ZN(n_257_43_27));
   NAND2_X1 i_257_43_28 (.A1(CPU_Bus[26]), .A2(n_257_43_27), .ZN(n_257_43_28));
   NAND2_X1 i_257_43_29 (.A1(n_257_43_10), .A2(n_257_43_25), .ZN(n_257_43_29));
   NOR2_X1 i_257_43_30 (.A1(n_257_43_29), .A2(n_257_43_5), .ZN(n_257_43_30));
   NAND2_X1 i_257_43_31 (.A1(CPU_Bus[24]), .A2(n_257_43_30), .ZN(n_257_43_31));
   NAND2_X1 i_257_43_32 (.A1(n_257_43_28), .A2(n_257_43_31), .ZN(n_257_43_32));
   NAND2_X1 i_257_43_33 (.A1(n_257_43_15), .A2(n_257_43_25), .ZN(n_257_43_33));
   NOR2_X1 i_257_43_34 (.A1(n_257_43_33), .A2(n_257_43_5), .ZN(n_257_43_34));
   NAND2_X1 i_257_43_35 (.A1(CPU_Bus[22]), .A2(n_257_43_34), .ZN(n_257_43_35));
   NAND2_X1 i_257_43_36 (.A1(n_257_43_19), .A2(n_257_43_25), .ZN(n_257_43_36));
   NOR2_X1 i_257_43_37 (.A1(n_257_43_36), .A2(n_257_43_5), .ZN(n_257_43_37));
   NAND2_X1 i_257_43_38 (.A1(CPU_Bus[20]), .A2(n_257_43_37), .ZN(n_257_43_38));
   NAND2_X1 i_257_43_39 (.A1(n_257_43_35), .A2(n_257_43_38), .ZN(n_257_43_39));
   NOR2_X1 i_257_43_40 (.A1(n_257_43_32), .A2(n_257_43_39), .ZN(n_257_43_40));
   NAND2_X1 i_257_43_41 (.A1(n_257_43_24), .A2(n_257_43_40), .ZN(n_257_43_41));
   NOR2_X1 i_257_43_42 (.A1(n_257_43_4), .A2(n_258), .ZN(n_257_43_42));
   NAND2_X1 i_257_43_43 (.A1(CPU_Bus[18]), .A2(n_257_43_42), .ZN(n_257_43_43));
   NOR2_X1 i_257_43_44 (.A1(n_257_43_11), .A2(n_258), .ZN(n_257_43_44));
   NAND2_X1 i_257_43_45 (.A1(CPU_Bus[16]), .A2(n_257_43_44), .ZN(n_257_43_45));
   NAND2_X1 i_257_43_46 (.A1(n_257_43_43), .A2(n_257_43_45), .ZN(n_257_43_46));
   NOR2_X1 i_257_43_47 (.A1(n_257_43_16), .A2(n_258), .ZN(n_257_43_47));
   NAND2_X1 i_257_43_48 (.A1(CPU_Bus[14]), .A2(n_257_43_47), .ZN(n_257_43_48));
   NOR2_X1 i_257_43_49 (.A1(n_257_43_20), .A2(n_258), .ZN(n_257_43_49));
   NAND2_X1 i_257_43_50 (.A1(CPU_Bus[12]), .A2(n_257_43_49), .ZN(n_257_43_50));
   NAND2_X1 i_257_43_51 (.A1(n_257_43_48), .A2(n_257_43_50), .ZN(n_257_43_51));
   NOR2_X1 i_257_43_52 (.A1(n_257_43_46), .A2(n_257_43_51), .ZN(n_257_43_52));
   NOR2_X1 i_257_43_53 (.A1(n_257_43_26), .A2(n_258), .ZN(n_257_43_53));
   NAND2_X1 i_257_43_54 (.A1(CPU_Bus[10]), .A2(n_257_43_53), .ZN(n_257_43_54));
   NOR2_X1 i_257_43_55 (.A1(n_257_43_29), .A2(n_258), .ZN(n_257_43_55));
   NAND2_X1 i_257_43_56 (.A1(CPU_Bus[8]), .A2(n_257_43_55), .ZN(n_257_43_56));
   NAND2_X1 i_257_43_57 (.A1(n_257_43_54), .A2(n_257_43_56), .ZN(n_257_43_57));
   NOR2_X1 i_257_43_58 (.A1(n_257_43_33), .A2(n_258), .ZN(n_257_43_58));
   NAND2_X1 i_257_43_59 (.A1(CPU_Bus[6]), .A2(n_257_43_58), .ZN(n_257_43_59));
   NOR2_X1 i_257_43_60 (.A1(n_257_43_36), .A2(n_258), .ZN(n_257_43_60));
   NAND2_X1 i_257_43_61 (.A1(CPU_Bus[4]), .A2(n_257_43_60), .ZN(n_257_43_61));
   NAND2_X1 i_257_43_62 (.A1(n_257_43_59), .A2(n_257_43_61), .ZN(n_257_43_62));
   NOR2_X1 i_257_43_63 (.A1(n_257_43_57), .A2(n_257_43_62), .ZN(n_257_43_63));
   NAND2_X1 i_257_43_64 (.A1(n_257_43_52), .A2(n_257_43_63), .ZN(n_257_43_64));
   NOR2_X1 i_257_43_65 (.A1(n_257_43_41), .A2(n_257_43_64), .ZN(n_257_43_65));
   NAND2_X1 i_257_43_66 (.A1(n_257_43_8), .A2(n_254), .ZN(n_257_43_66));
   NOR2_X1 i_257_43_67 (.A1(n_257_43_66), .A2(n_257_43_2), .ZN(n_257_43_67));
   NAND2_X1 i_257_43_68 (.A1(n_257_43_67), .A2(n_257), .ZN(n_257_43_68));
   NOR2_X1 i_257_43_69 (.A1(n_257_43_68), .A2(n_257_43_5), .ZN(n_257_43_69));
   NAND2_X1 i_257_43_70 (.A1(CPU_Bus[1]), .A2(n_257_43_69), .ZN(n_257_43_70));
   NOR2_X1 i_257_43_71 (.A1(n_257_43_66), .A2(n_256), .ZN(n_257_43_71));
   NAND2_X1 i_257_43_72 (.A1(n_257_43_71), .A2(n_257), .ZN(n_257_43_72));
   NOR2_X1 i_257_43_73 (.A1(n_257_43_72), .A2(n_257_43_5), .ZN(n_257_43_73));
   NAND2_X1 i_257_43_74 (.A1(CPU_Bus[29]), .A2(n_257_43_73), .ZN(n_257_43_74));
   NAND2_X1 i_257_43_75 (.A1(n_257_43_70), .A2(n_257_43_74), .ZN(n_257_43_75));
   NAND2_X1 i_257_43_76 (.A1(n_257_43_67), .A2(n_257_43_25), .ZN(n_257_43_76));
   NOR2_X1 i_257_43_77 (.A1(n_257_43_76), .A2(n_257_43_5), .ZN(n_257_43_77));
   NAND2_X1 i_257_43_78 (.A1(CPU_Bus[25]), .A2(n_257_43_77), .ZN(n_257_43_78));
   NAND2_X1 i_257_43_79 (.A1(n_257_43_71), .A2(n_257_43_25), .ZN(n_257_43_79));
   NOR2_X1 i_257_43_80 (.A1(n_257_43_79), .A2(n_257_43_5), .ZN(n_257_43_80));
   NAND2_X1 i_257_43_81 (.A1(CPU_Bus[21]), .A2(n_257_43_80), .ZN(n_257_43_81));
   NAND2_X1 i_257_43_82 (.A1(n_257_43_78), .A2(n_257_43_81), .ZN(n_257_43_82));
   NOR2_X1 i_257_43_83 (.A1(n_257_43_75), .A2(n_257_43_82), .ZN(n_257_43_83));
   NOR2_X1 i_257_43_84 (.A1(n_257_43_68), .A2(n_258), .ZN(n_257_43_84));
   NAND2_X1 i_257_43_85 (.A1(CPU_Bus[17]), .A2(n_257_43_84), .ZN(n_257_43_85));
   NOR2_X1 i_257_43_86 (.A1(n_257_43_72), .A2(n_258), .ZN(n_257_43_86));
   NAND2_X1 i_257_43_87 (.A1(CPU_Bus[13]), .A2(n_257_43_86), .ZN(n_257_43_87));
   NAND2_X1 i_257_43_88 (.A1(n_257_43_85), .A2(n_257_43_87), .ZN(n_257_43_88));
   NOR2_X1 i_257_43_89 (.A1(n_257_43_76), .A2(n_258), .ZN(n_257_43_89));
   NAND2_X1 i_257_43_90 (.A1(CPU_Bus[9]), .A2(n_257_43_89), .ZN(n_257_43_90));
   NOR2_X1 i_257_43_91 (.A1(n_257_43_79), .A2(n_258), .ZN(n_257_43_91));
   NAND2_X1 i_257_43_92 (.A1(CPU_Bus[5]), .A2(n_257_43_91), .ZN(n_257_43_92));
   NAND2_X1 i_257_43_93 (.A1(n_257_43_90), .A2(n_257_43_92), .ZN(n_257_43_93));
   NOR2_X1 i_257_43_94 (.A1(n_257_43_88), .A2(n_257_43_93), .ZN(n_257_43_94));
   NAND2_X1 i_257_43_95 (.A1(n_257_43_83), .A2(n_257_43_94), .ZN(n_257_43_95));
   NAND2_X1 i_257_43_96 (.A1(n_254), .A2(n_255), .ZN(n_257_43_96));
   NOR2_X1 i_257_43_97 (.A1(n_257_43_96), .A2(n_257_43_2), .ZN(n_257_43_97));
   NAND2_X1 i_257_43_98 (.A1(n_257_43_97), .A2(n_257), .ZN(n_257_43_98));
   NOR2_X1 i_257_43_99 (.A1(n_257_43_98), .A2(n_257_43_5), .ZN(n_257_43_99));
   NAND2_X1 i_257_43_100 (.A1(CPU_Bus[3]), .A2(n_257_43_99), .ZN(n_257_43_100));
   NOR2_X1 i_257_43_101 (.A1(n_257_43_96), .A2(n_256), .ZN(n_257_43_101));
   NAND2_X1 i_257_43_102 (.A1(n_257_43_101), .A2(n_257), .ZN(n_257_43_102));
   NOR2_X1 i_257_43_103 (.A1(n_257_43_102), .A2(n_257_43_5), .ZN(n_257_43_103));
   NAND2_X1 i_257_43_104 (.A1(CPU_Bus[31]), .A2(n_257_43_103), .ZN(n_257_43_104));
   NAND2_X1 i_257_43_105 (.A1(n_257_43_100), .A2(n_257_43_104), .ZN(n_257_43_105));
   NAND2_X1 i_257_43_106 (.A1(n_257_43_97), .A2(n_257_43_25), .ZN(n_257_43_106));
   NOR2_X1 i_257_43_107 (.A1(n_257_43_106), .A2(n_257_43_5), .ZN(n_257_43_107));
   NAND2_X1 i_257_43_108 (.A1(CPU_Bus[27]), .A2(n_257_43_107), .ZN(n_257_43_108));
   NAND2_X1 i_257_43_109 (.A1(n_257_43_101), .A2(n_257_43_25), .ZN(n_257_43_109));
   NOR2_X1 i_257_43_110 (.A1(n_257_43_109), .A2(n_257_43_5), .ZN(n_257_43_110));
   NAND2_X1 i_257_43_111 (.A1(CPU_Bus[23]), .A2(n_257_43_110), .ZN(n_257_43_111));
   NAND2_X1 i_257_43_112 (.A1(n_257_43_108), .A2(n_257_43_111), .ZN(n_257_43_112));
   NOR2_X1 i_257_43_113 (.A1(n_257_43_105), .A2(n_257_43_112), .ZN(n_257_43_113));
   NOR2_X1 i_257_43_114 (.A1(n_257_43_98), .A2(n_258), .ZN(n_257_43_114));
   NAND2_X1 i_257_43_115 (.A1(CPU_Bus[19]), .A2(n_257_43_114), .ZN(n_257_43_115));
   NOR2_X1 i_257_43_116 (.A1(n_257_43_102), .A2(n_258), .ZN(n_257_43_116));
   NAND2_X1 i_257_43_117 (.A1(CPU_Bus[15]), .A2(n_257_43_116), .ZN(n_257_43_117));
   NAND2_X1 i_257_43_118 (.A1(n_257_43_115), .A2(n_257_43_117), .ZN(n_257_43_118));
   NOR2_X1 i_257_43_119 (.A1(n_257_43_106), .A2(n_258), .ZN(n_257_43_119));
   NAND2_X1 i_257_43_120 (.A1(CPU_Bus[11]), .A2(n_257_43_119), .ZN(n_257_43_120));
   NOR2_X1 i_257_43_121 (.A1(n_257_43_109), .A2(n_258), .ZN(n_257_43_121));
   NAND2_X1 i_257_43_122 (.A1(CPU_Bus[7]), .A2(n_257_43_121), .ZN(n_257_43_122));
   NAND2_X1 i_257_43_123 (.A1(n_257_43_120), .A2(n_257_43_122), .ZN(n_257_43_123));
   NOR2_X1 i_257_43_124 (.A1(n_257_43_118), .A2(n_257_43_123), .ZN(n_257_43_124));
   NAND2_X1 i_257_43_125 (.A1(n_257_43_113), .A2(n_257_43_124), .ZN(n_257_43_125));
   NOR2_X1 i_257_43_126 (.A1(n_257_43_95), .A2(n_257_43_125), .ZN(n_257_43_126));
   NAND2_X1 i_257_43_127 (.A1(n_257_43_65), .A2(n_257_43_126), .ZN(n_257_304));
   datapath__1_369 i_257_44 (.PacketSize({PacketSize[5], PacketSize[4], 
      PacketSize[3], PacketSize[2], PacketSize[1], 1'b0}), .p_0({n_257_309, 
      uc_462, uc_463, uc_464, uc_465, uc_466, uc_467, uc_468, uc_469, uc_470, 
      uc_471, uc_472, uc_473, uc_474, uc_475, uc_476, uc_477, uc_478, uc_479, 
      uc_480, uc_481, uc_482, uc_483, uc_484, uc_485, uc_486, n_257_308, 
      n_257_307, n_257_306, n_257_305, uc_487, uc_488}));
   datapath__1_370 i_257_45 (.p_0({uc_489, uc_490, uc_491, uc_492, uc_493, 
      uc_494, uc_495, uc_496, uc_497, uc_498, uc_499, uc_500, uc_501, uc_502, 
      uc_503, uc_504, uc_505, uc_506, uc_507, uc_508, uc_509, uc_510, uc_511, 
      uc_512, uc_513, n_257_309, n_257_308, n_257_307, n_257_306, n_257_305, 
      n_257_1091, PacketSize[0]}), .p_1({n_257_341, n_257_340, n_257_339, 
      n_257_338, n_257_337, n_257_336, n_257_335, n_257_334, n_257_333, 
      n_257_332, n_257_331, n_257_330, n_257_329, n_257_328, n_257_327, 
      n_257_326, n_257_325, n_257_324, n_257_323, n_257_322, n_257_321, 
      n_257_320, n_257_319, n_257_318, n_257_317, n_257_316, n_257_315, 
      n_257_314, n_257_313, n_257_312, n_257_311, n_257_310}));
   INV_X1 i_257_46_0 (.A(n_257_46_0), .ZN(n_257_342));
   NAND2_X1 i_257_46_1 (.A1(n_257_46_49), .A2(n_257_46_1), .ZN(n_257_46_0));
   NAND3_X1 i_257_46_2 (.A1(n_257_46_25), .A2(n_257_46_2), .A3(n_257_46_48), 
      .ZN(n_257_46_1));
   NAND3_X1 i_257_46_3 (.A1(n_257_46_14), .A2(n_257_46_3), .A3(n_257), .ZN(
      n_257_46_2));
   NAND3_X1 i_257_46_4 (.A1(n_257_46_9), .A2(n_257_46_4), .A3(n_257_46_85), 
      .ZN(n_257_46_3));
   NAND3_X1 i_257_46_5 (.A1(n_257_46_7), .A2(n_257_46_5), .A3(n_257_46_96), 
      .ZN(n_257_46_4));
   NAND2_X1 i_257_46_6 (.A1(n_257_46_6), .A2(n_257_46_95), .ZN(n_257_46_5));
   INV_X1 i_257_46_7 (.A(CPU_Bus[11]), .ZN(n_257_46_6));
   NAND2_X1 i_257_46_8 (.A1(n_257_46_8), .A2(n_254), .ZN(n_257_46_7));
   INV_X1 i_257_46_9 (.A(CPU_Bus[12]), .ZN(n_257_46_8));
   NAND3_X1 i_257_46_10 (.A1(n_257_46_12), .A2(n_257_46_10), .A3(n_255), 
      .ZN(n_257_46_9));
   NAND2_X1 i_257_46_11 (.A1(n_257_46_11), .A2(n_257_46_95), .ZN(n_257_46_10));
   INV_X1 i_257_46_12 (.A(CPU_Bus[13]), .ZN(n_257_46_11));
   NAND2_X1 i_257_46_13 (.A1(n_257_46_13), .A2(n_254), .ZN(n_257_46_12));
   INV_X1 i_257_46_14 (.A(CPU_Bus[14]), .ZN(n_257_46_13));
   NAND3_X1 i_257_46_15 (.A1(n_257_46_20), .A2(n_257_46_15), .A3(n_256), 
      .ZN(n_257_46_14));
   NAND3_X1 i_257_46_16 (.A1(n_257_46_18), .A2(n_257_46_16), .A3(n_257_46_96), 
      .ZN(n_257_46_15));
   NAND2_X1 i_257_46_17 (.A1(n_257_46_17), .A2(n_257_46_95), .ZN(n_257_46_16));
   INV_X1 i_257_46_18 (.A(CPU_Bus[15]), .ZN(n_257_46_17));
   NAND2_X1 i_257_46_19 (.A1(n_257_46_19), .A2(n_254), .ZN(n_257_46_18));
   INV_X1 i_257_46_20 (.A(CPU_Bus[16]), .ZN(n_257_46_19));
   NAND3_X1 i_257_46_21 (.A1(n_257_46_23), .A2(n_257_46_21), .A3(n_255), 
      .ZN(n_257_46_20));
   NAND2_X1 i_257_46_22 (.A1(n_257_46_22), .A2(n_257_46_95), .ZN(n_257_46_21));
   INV_X1 i_257_46_23 (.A(CPU_Bus[17]), .ZN(n_257_46_22));
   NAND2_X1 i_257_46_24 (.A1(n_257_46_24), .A2(n_254), .ZN(n_257_46_23));
   INV_X1 i_257_46_25 (.A(CPU_Bus[18]), .ZN(n_257_46_24));
   NAND3_X1 i_257_46_26 (.A1(n_257_46_37), .A2(n_257_46_26), .A3(n_257_46_97), 
      .ZN(n_257_46_25));
   NAND3_X1 i_257_46_27 (.A1(n_257_46_32), .A2(n_257_46_27), .A3(n_256), 
      .ZN(n_257_46_26));
   NAND3_X1 i_257_46_28 (.A1(n_257_46_30), .A2(n_257_46_28), .A3(n_255), 
      .ZN(n_257_46_27));
   NAND2_X1 i_257_46_29 (.A1(n_257_46_29), .A2(n_254), .ZN(n_257_46_28));
   INV_X1 i_257_46_30 (.A(CPU_Bus[10]), .ZN(n_257_46_29));
   NAND2_X1 i_257_46_31 (.A1(n_257_46_31), .A2(n_257_46_95), .ZN(n_257_46_30));
   INV_X1 i_257_46_32 (.A(CPU_Bus[9]), .ZN(n_257_46_31));
   NAND3_X1 i_257_46_33 (.A1(n_257_46_35), .A2(n_257_46_33), .A3(n_257_46_96), 
      .ZN(n_257_46_32));
   NAND2_X1 i_257_46_34 (.A1(n_257_46_34), .A2(n_257_46_95), .ZN(n_257_46_33));
   INV_X1 i_257_46_35 (.A(CPU_Bus[7]), .ZN(n_257_46_34));
   NAND2_X1 i_257_46_36 (.A1(n_257_46_36), .A2(n_254), .ZN(n_257_46_35));
   INV_X1 i_257_46_37 (.A(CPU_Bus[8]), .ZN(n_257_46_36));
   NAND3_X1 i_257_46_38 (.A1(n_257_46_43), .A2(n_257_46_38), .A3(n_257_46_85), 
      .ZN(n_257_46_37));
   NAND3_X1 i_257_46_39 (.A1(n_257_46_41), .A2(n_257_46_39), .A3(n_255), 
      .ZN(n_257_46_38));
   NAND2_X1 i_257_46_40 (.A1(n_257_46_40), .A2(n_254), .ZN(n_257_46_39));
   INV_X1 i_257_46_41 (.A(CPU_Bus[6]), .ZN(n_257_46_40));
   NAND2_X1 i_257_46_42 (.A1(n_257_46_42), .A2(n_257_46_95), .ZN(n_257_46_41));
   INV_X1 i_257_46_43 (.A(CPU_Bus[5]), .ZN(n_257_46_42));
   NAND3_X1 i_257_46_44 (.A1(n_257_46_46), .A2(n_257_46_44), .A3(n_257_46_96), 
      .ZN(n_257_46_43));
   NAND2_X1 i_257_46_45 (.A1(n_257_46_45), .A2(n_257_46_95), .ZN(n_257_46_44));
   INV_X1 i_257_46_46 (.A(CPU_Bus[3]), .ZN(n_257_46_45));
   NAND2_X1 i_257_46_47 (.A1(n_257_46_47), .A2(n_254), .ZN(n_257_46_46));
   INV_X1 i_257_46_48 (.A(CPU_Bus[4]), .ZN(n_257_46_47));
   INV_X1 i_257_46_49 (.A(n_258), .ZN(n_257_46_48));
   NAND3_X1 i_257_46_50 (.A1(n_257_46_73), .A2(n_257_46_50), .A3(n_258), 
      .ZN(n_257_46_49));
   NAND3_X1 i_257_46_51 (.A1(n_257_46_62), .A2(n_257_46_51), .A3(n_257), 
      .ZN(n_257_46_50));
   NAND3_X1 i_257_46_52 (.A1(n_257_46_57), .A2(n_257_46_52), .A3(n_257_46_85), 
      .ZN(n_257_46_51));
   NAND3_X1 i_257_46_53 (.A1(n_257_46_55), .A2(n_257_46_53), .A3(n_257_46_96), 
      .ZN(n_257_46_52));
   NAND2_X1 i_257_46_54 (.A1(n_257_46_54), .A2(n_257_46_95), .ZN(n_257_46_53));
   INV_X1 i_257_46_55 (.A(CPU_Bus[27]), .ZN(n_257_46_54));
   NAND2_X1 i_257_46_56 (.A1(n_257_46_56), .A2(n_254), .ZN(n_257_46_55));
   INV_X1 i_257_46_57 (.A(CPU_Bus[28]), .ZN(n_257_46_56));
   NAND3_X1 i_257_46_58 (.A1(n_257_46_60), .A2(n_257_46_58), .A3(n_255), 
      .ZN(n_257_46_57));
   NAND2_X1 i_257_46_59 (.A1(n_257_46_59), .A2(n_254), .ZN(n_257_46_58));
   INV_X1 i_257_46_60 (.A(CPU_Bus[30]), .ZN(n_257_46_59));
   NAND2_X1 i_257_46_61 (.A1(n_257_46_61), .A2(n_257_46_95), .ZN(n_257_46_60));
   INV_X1 i_257_46_62 (.A(CPU_Bus[29]), .ZN(n_257_46_61));
   NAND3_X1 i_257_46_63 (.A1(n_257_46_68), .A2(n_257_46_63), .A3(n_256), 
      .ZN(n_257_46_62));
   NAND3_X1 i_257_46_64 (.A1(n_257_46_66), .A2(n_257_46_64), .A3(n_257_46_96), 
      .ZN(n_257_46_63));
   NAND2_X1 i_257_46_65 (.A1(n_257_46_65), .A2(n_254), .ZN(n_257_46_64));
   INV_X1 i_257_46_66 (.A(CPU_Bus[0]), .ZN(n_257_46_65));
   NAND2_X1 i_257_46_67 (.A1(n_257_46_67), .A2(n_257_46_95), .ZN(n_257_46_66));
   INV_X1 i_257_46_68 (.A(CPU_Bus[31]), .ZN(n_257_46_67));
   NAND3_X1 i_257_46_69 (.A1(n_257_46_71), .A2(n_257_46_69), .A3(n_255), 
      .ZN(n_257_46_68));
   NAND2_X1 i_257_46_70 (.A1(n_257_46_70), .A2(n_257_46_95), .ZN(n_257_46_69));
   INV_X1 i_257_46_71 (.A(CPU_Bus[1]), .ZN(n_257_46_70));
   NAND2_X1 i_257_46_72 (.A1(n_257_46_72), .A2(n_254), .ZN(n_257_46_71));
   INV_X1 i_257_46_73 (.A(CPU_Bus[2]), .ZN(n_257_46_72));
   NAND3_X1 i_257_46_74 (.A1(n_257_46_86), .A2(n_257_46_74), .A3(n_257_46_97), 
      .ZN(n_257_46_73));
   NAND3_X1 i_257_46_75 (.A1(n_257_46_80), .A2(n_257_46_75), .A3(n_257_46_85), 
      .ZN(n_257_46_74));
   NAND3_X1 i_257_46_76 (.A1(n_257_46_78), .A2(n_257_46_76), .A3(n_257_46_96), 
      .ZN(n_257_46_75));
   NAND2_X1 i_257_46_77 (.A1(n_257_46_77), .A2(n_254), .ZN(n_257_46_76));
   INV_X1 i_257_46_78 (.A(CPU_Bus[20]), .ZN(n_257_46_77));
   NAND2_X1 i_257_46_79 (.A1(n_257_46_79), .A2(n_257_46_95), .ZN(n_257_46_78));
   INV_X1 i_257_46_80 (.A(CPU_Bus[19]), .ZN(n_257_46_79));
   NAND3_X1 i_257_46_81 (.A1(n_257_46_83), .A2(n_257_46_81), .A3(n_255), 
      .ZN(n_257_46_80));
   NAND2_X1 i_257_46_82 (.A1(n_257_46_82), .A2(n_254), .ZN(n_257_46_81));
   INV_X1 i_257_46_83 (.A(CPU_Bus[22]), .ZN(n_257_46_82));
   NAND2_X1 i_257_46_84 (.A1(n_257_46_84), .A2(n_257_46_95), .ZN(n_257_46_83));
   INV_X1 i_257_46_85 (.A(CPU_Bus[21]), .ZN(n_257_46_84));
   INV_X1 i_257_46_86 (.A(n_256), .ZN(n_257_46_85));
   NAND3_X1 i_257_46_87 (.A1(n_257_46_92), .A2(n_257_46_87), .A3(n_256), 
      .ZN(n_257_46_86));
   NAND3_X1 i_257_46_88 (.A1(n_257_46_90), .A2(n_257_46_88), .A3(n_255), 
      .ZN(n_257_46_87));
   NAND2_X1 i_257_46_89 (.A1(n_257_46_89), .A2(n_257_46_95), .ZN(n_257_46_88));
   INV_X1 i_257_46_90 (.A(CPU_Bus[25]), .ZN(n_257_46_89));
   NAND2_X1 i_257_46_91 (.A1(n_257_46_91), .A2(n_254), .ZN(n_257_46_90));
   INV_X1 i_257_46_92 (.A(CPU_Bus[26]), .ZN(n_257_46_91));
   OAI211_X1 i_257_46_93 (.A(n_257_46_93), .B(n_257_46_96), .C1(n_257_46_95), 
      .C2(CPU_Bus[24]), .ZN(n_257_46_92));
   NAND2_X1 i_257_46_94 (.A1(n_257_46_94), .A2(n_257_46_95), .ZN(n_257_46_93));
   INV_X1 i_257_46_95 (.A(CPU_Bus[23]), .ZN(n_257_46_94));
   INV_X1 i_257_46_96 (.A(n_254), .ZN(n_257_46_95));
   INV_X1 i_257_46_97 (.A(n_255), .ZN(n_257_46_96));
   INV_X1 i_257_46_98 (.A(n_257), .ZN(n_257_46_97));
   datapath__1_372 i_257_47 (.PacketSize(PacketSize), .p_0({n_257_348, uc_514, 
      uc_515, uc_516, uc_517, uc_518, uc_519, uc_520, uc_521, uc_522, uc_523, 
      uc_524, uc_525, uc_526, uc_527, uc_528, uc_529, uc_530, uc_531, uc_532, 
      uc_533, uc_534, uc_535, uc_536, uc_537, uc_538, n_257_347, n_257_346, 
      n_257_345, n_257_344, n_257_343, uc_539}));
   datapath__1_373 i_257_48 (.p_0({uc_540, uc_541, uc_542, uc_543, uc_544, 
      uc_545, uc_546, uc_547, uc_548, uc_549, uc_550, uc_551, uc_552, uc_553, 
      uc_554, uc_555, uc_556, uc_557, uc_558, uc_559, uc_560, uc_561, uc_562, 
      uc_563, uc_564, n_257_348, n_257_347, n_257_346, n_257_345, n_257_344, 
      n_257_343, n_151}), .p_1({n_257_380, n_257_379, n_257_378, n_257_377, 
      n_257_376, n_257_375, n_257_374, n_257_373, n_257_372, n_257_371, 
      n_257_370, n_257_369, n_257_368, n_257_367, n_257_366, n_257_365, 
      n_257_364, n_257_363, n_257_362, n_257_361, n_257_360, n_257_359, 
      n_257_358, n_257_357, n_257_356, n_257_355, n_257_354, n_257_353, 
      n_257_352, n_257_351, n_257_350, n_257_349}));
   NAND2_X1 i_257_49_0 (.A1(n_257_49_49), .A2(n_257_49_0), .ZN(n_257_381));
   NAND2_X1 i_257_49_1 (.A1(n_257_49_1), .A2(n_257_49_48), .ZN(n_257_49_0));
   NAND2_X1 i_257_49_2 (.A1(n_257_49_25), .A2(n_257_49_2), .ZN(n_257_49_1));
   NAND3_X1 i_257_49_3 (.A1(n_257_49_14), .A2(n_257_49_3), .A3(n_257), .ZN(
      n_257_49_2));
   NAND3_X1 i_257_49_4 (.A1(n_257_49_9), .A2(n_257_49_4), .A3(n_257_49_97), 
      .ZN(n_257_49_3));
   NAND3_X1 i_257_49_5 (.A1(n_257_49_7), .A2(n_257_49_5), .A3(n_257_49_96), 
      .ZN(n_257_49_4));
   NAND2_X1 i_257_49_6 (.A1(n_257_49_6), .A2(n_254), .ZN(n_257_49_5));
   INV_X1 i_257_49_7 (.A(CPU_Bus[11]), .ZN(n_257_49_6));
   NAND2_X1 i_257_49_8 (.A1(n_257_49_8), .A2(n_257_49_92), .ZN(n_257_49_7));
   INV_X1 i_257_49_9 (.A(CPU_Bus[10]), .ZN(n_257_49_8));
   NAND3_X1 i_257_49_10 (.A1(n_257_49_12), .A2(n_257_49_10), .A3(n_255), 
      .ZN(n_257_49_9));
   NAND2_X1 i_257_49_11 (.A1(n_257_49_11), .A2(n_257_49_92), .ZN(n_257_49_10));
   INV_X1 i_257_49_12 (.A(CPU_Bus[12]), .ZN(n_257_49_11));
   NAND2_X1 i_257_49_13 (.A1(n_257_49_13), .A2(n_254), .ZN(n_257_49_12));
   INV_X1 i_257_49_14 (.A(CPU_Bus[13]), .ZN(n_257_49_13));
   NAND3_X1 i_257_49_15 (.A1(n_257_49_20), .A2(n_257_49_15), .A3(n_256), 
      .ZN(n_257_49_14));
   NAND3_X1 i_257_49_16 (.A1(n_257_49_18), .A2(n_257_49_16), .A3(n_255), 
      .ZN(n_257_49_15));
   NAND2_X1 i_257_49_17 (.A1(n_257_49_17), .A2(n_257_49_92), .ZN(n_257_49_16));
   INV_X1 i_257_49_18 (.A(CPU_Bus[16]), .ZN(n_257_49_17));
   NAND2_X1 i_257_49_19 (.A1(n_257_49_19), .A2(n_254), .ZN(n_257_49_18));
   INV_X1 i_257_49_20 (.A(CPU_Bus[17]), .ZN(n_257_49_19));
   NAND3_X1 i_257_49_21 (.A1(n_257_49_23), .A2(n_257_49_21), .A3(n_257_49_96), 
      .ZN(n_257_49_20));
   NAND2_X1 i_257_49_22 (.A1(n_257_49_22), .A2(n_254), .ZN(n_257_49_21));
   INV_X1 i_257_49_23 (.A(CPU_Bus[15]), .ZN(n_257_49_22));
   NAND2_X1 i_257_49_24 (.A1(n_257_49_24), .A2(n_257_49_92), .ZN(n_257_49_23));
   INV_X1 i_257_49_25 (.A(CPU_Bus[14]), .ZN(n_257_49_24));
   NAND3_X1 i_257_49_26 (.A1(n_257_49_37), .A2(n_257_49_26), .A3(n_257_49_98), 
      .ZN(n_257_49_25));
   NAND3_X1 i_257_49_27 (.A1(n_257_49_32), .A2(n_257_49_27), .A3(n_256), 
      .ZN(n_257_49_26));
   NAND3_X1 i_257_49_28 (.A1(n_257_49_30), .A2(n_257_49_28), .A3(n_255), 
      .ZN(n_257_49_27));
   NAND2_X1 i_257_49_29 (.A1(n_257_49_29), .A2(n_257_49_92), .ZN(n_257_49_28));
   INV_X1 i_257_49_30 (.A(CPU_Bus[8]), .ZN(n_257_49_29));
   NAND2_X1 i_257_49_31 (.A1(n_257_49_31), .A2(n_254), .ZN(n_257_49_30));
   INV_X1 i_257_49_32 (.A(CPU_Bus[9]), .ZN(n_257_49_31));
   NAND3_X1 i_257_49_33 (.A1(n_257_49_35), .A2(n_257_49_33), .A3(n_257_49_96), 
      .ZN(n_257_49_32));
   NAND2_X1 i_257_49_34 (.A1(n_257_49_34), .A2(n_257_49_92), .ZN(n_257_49_33));
   INV_X1 i_257_49_35 (.A(CPU_Bus[6]), .ZN(n_257_49_34));
   NAND2_X1 i_257_49_36 (.A1(n_257_49_36), .A2(n_254), .ZN(n_257_49_35));
   INV_X1 i_257_49_37 (.A(CPU_Bus[7]), .ZN(n_257_49_36));
   NAND3_X1 i_257_49_38 (.A1(n_257_49_43), .A2(n_257_49_38), .A3(n_257_49_97), 
      .ZN(n_257_49_37));
   NAND3_X1 i_257_49_39 (.A1(n_257_49_41), .A2(n_257_49_39), .A3(n_257_49_96), 
      .ZN(n_257_49_38));
   NAND2_X1 i_257_49_40 (.A1(n_257_49_40), .A2(n_257_49_92), .ZN(n_257_49_39));
   INV_X1 i_257_49_41 (.A(CPU_Bus[2]), .ZN(n_257_49_40));
   NAND2_X1 i_257_49_42 (.A1(n_257_49_42), .A2(n_254), .ZN(n_257_49_41));
   INV_X1 i_257_49_43 (.A(CPU_Bus[3]), .ZN(n_257_49_42));
   NAND3_X1 i_257_49_44 (.A1(n_257_49_46), .A2(n_257_49_44), .A3(n_255), 
      .ZN(n_257_49_43));
   NAND2_X1 i_257_49_45 (.A1(n_257_49_45), .A2(n_257_49_92), .ZN(n_257_49_44));
   INV_X1 i_257_49_46 (.A(CPU_Bus[4]), .ZN(n_257_49_45));
   NAND2_X1 i_257_49_47 (.A1(n_257_49_47), .A2(n_254), .ZN(n_257_49_46));
   INV_X1 i_257_49_48 (.A(CPU_Bus[5]), .ZN(n_257_49_47));
   INV_X1 i_257_49_49 (.A(n_258), .ZN(n_257_49_48));
   NAND2_X1 i_257_49_50 (.A1(n_257_49_50), .A2(n_258), .ZN(n_257_49_49));
   NAND2_X1 i_257_49_51 (.A1(n_257_49_74), .A2(n_257_49_51), .ZN(n_257_49_50));
   NAND3_X1 i_257_49_52 (.A1(n_257_49_63), .A2(n_257_49_52), .A3(n_257), 
      .ZN(n_257_49_51));
   NAND3_X1 i_257_49_53 (.A1(n_257_49_58), .A2(n_257_49_53), .A3(n_257_49_97), 
      .ZN(n_257_49_52));
   NAND3_X1 i_257_49_54 (.A1(n_257_49_56), .A2(n_257_49_54), .A3(n_257_49_96), 
      .ZN(n_257_49_53));
   NAND2_X1 i_257_49_55 (.A1(n_257_49_55), .A2(n_254), .ZN(n_257_49_54));
   INV_X1 i_257_49_56 (.A(CPU_Bus[27]), .ZN(n_257_49_55));
   NAND2_X1 i_257_49_57 (.A1(n_257_49_57), .A2(n_257_49_92), .ZN(n_257_49_56));
   INV_X1 i_257_49_58 (.A(CPU_Bus[26]), .ZN(n_257_49_57));
   NAND3_X1 i_257_49_59 (.A1(n_257_49_61), .A2(n_257_49_59), .A3(n_255), 
      .ZN(n_257_49_58));
   NAND2_X1 i_257_49_60 (.A1(n_257_49_60), .A2(n_254), .ZN(n_257_49_59));
   INV_X1 i_257_49_61 (.A(CPU_Bus[29]), .ZN(n_257_49_60));
   NAND2_X1 i_257_49_62 (.A1(n_257_49_62), .A2(n_257_49_92), .ZN(n_257_49_61));
   INV_X1 i_257_49_63 (.A(CPU_Bus[28]), .ZN(n_257_49_62));
   NAND3_X1 i_257_49_64 (.A1(n_257_49_69), .A2(n_257_49_64), .A3(n_256), 
      .ZN(n_257_49_63));
   NAND3_X1 i_257_49_65 (.A1(n_257_49_67), .A2(n_257_49_65), .A3(n_255), 
      .ZN(n_257_49_64));
   NAND2_X1 i_257_49_66 (.A1(n_257_49_66), .A2(n_257_49_92), .ZN(n_257_49_65));
   INV_X1 i_257_49_67 (.A(CPU_Bus[0]), .ZN(n_257_49_66));
   NAND2_X1 i_257_49_68 (.A1(n_257_49_68), .A2(n_254), .ZN(n_257_49_67));
   INV_X1 i_257_49_69 (.A(CPU_Bus[1]), .ZN(n_257_49_68));
   NAND3_X1 i_257_49_70 (.A1(n_257_49_72), .A2(n_257_49_70), .A3(n_257_49_96), 
      .ZN(n_257_49_69));
   NAND2_X1 i_257_49_71 (.A1(n_257_49_71), .A2(n_257_49_92), .ZN(n_257_49_70));
   INV_X1 i_257_49_72 (.A(CPU_Bus[30]), .ZN(n_257_49_71));
   NAND2_X1 i_257_49_73 (.A1(n_257_49_73), .A2(n_254), .ZN(n_257_49_72));
   INV_X1 i_257_49_74 (.A(CPU_Bus[31]), .ZN(n_257_49_73));
   NAND3_X1 i_257_49_75 (.A1(n_257_49_86), .A2(n_257_49_98), .A3(n_257_49_75), 
      .ZN(n_257_49_74));
   NAND3_X1 i_257_49_76 (.A1(n_257_49_81), .A2(n_257_49_76), .A3(n_256), 
      .ZN(n_257_49_75));
   NAND3_X1 i_257_49_77 (.A1(n_257_49_79), .A2(n_257_49_77), .A3(n_257_49_96), 
      .ZN(n_257_49_76));
   NAND2_X1 i_257_49_78 (.A1(n_257_49_78), .A2(n_254), .ZN(n_257_49_77));
   INV_X1 i_257_49_79 (.A(CPU_Bus[23]), .ZN(n_257_49_78));
   NAND2_X1 i_257_49_80 (.A1(n_257_49_80), .A2(n_257_49_92), .ZN(n_257_49_79));
   INV_X1 i_257_49_81 (.A(CPU_Bus[22]), .ZN(n_257_49_80));
   NAND3_X1 i_257_49_82 (.A1(n_257_49_84), .A2(n_257_49_82), .A3(n_255), 
      .ZN(n_257_49_81));
   NAND2_X1 i_257_49_83 (.A1(n_257_49_83), .A2(n_254), .ZN(n_257_49_82));
   INV_X1 i_257_49_84 (.A(CPU_Bus[25]), .ZN(n_257_49_83));
   NAND2_X1 i_257_49_85 (.A1(n_257_49_85), .A2(n_257_49_92), .ZN(n_257_49_84));
   INV_X1 i_257_49_86 (.A(CPU_Bus[24]), .ZN(n_257_49_85));
   NAND3_X1 i_257_49_87 (.A1(n_257_49_93), .A2(n_257_49_97), .A3(n_257_49_87), 
      .ZN(n_257_49_86));
   NAND3_X1 i_257_49_88 (.A1(n_257_49_90), .A2(n_257_49_88), .A3(n_255), 
      .ZN(n_257_49_87));
   NAND2_X1 i_257_49_89 (.A1(n_257_49_89), .A2(n_254), .ZN(n_257_49_88));
   INV_X1 i_257_49_90 (.A(CPU_Bus[21]), .ZN(n_257_49_89));
   NAND2_X1 i_257_49_91 (.A1(n_257_49_91), .A2(n_257_49_92), .ZN(n_257_49_90));
   INV_X1 i_257_49_92 (.A(CPU_Bus[20]), .ZN(n_257_49_91));
   INV_X1 i_257_49_93 (.A(n_254), .ZN(n_257_49_92));
   OAI211_X1 i_257_49_94 (.A(n_257_49_94), .B(n_257_49_96), .C1(n_254), .C2(
      CPU_Bus[18]), .ZN(n_257_49_93));
   NAND2_X1 i_257_49_95 (.A1(n_257_49_95), .A2(n_254), .ZN(n_257_49_94));
   INV_X1 i_257_49_96 (.A(CPU_Bus[19]), .ZN(n_257_49_95));
   INV_X1 i_257_49_97 (.A(n_255), .ZN(n_257_49_96));
   INV_X1 i_257_49_98 (.A(n_256), .ZN(n_257_49_97));
   INV_X1 i_257_49_99 (.A(n_257), .ZN(n_257_49_98));
   INV_X1 i_257_50_0 (.A(n_254), .ZN(n_257_50_0));
   NAND2_X1 i_257_50_1 (.A1(n_257_50_0), .A2(n_255), .ZN(n_257_50_1));
   INV_X1 i_257_50_2 (.A(n_256), .ZN(n_257_50_2));
   NOR2_X1 i_257_50_3 (.A1(n_257_50_1), .A2(n_257_50_2), .ZN(n_257_50_3));
   NAND2_X1 i_257_50_4 (.A1(n_257_50_3), .A2(n_257), .ZN(n_257_50_4));
   INV_X1 i_257_50_5 (.A(n_258), .ZN(n_257_50_5));
   NOR2_X1 i_257_50_6 (.A1(n_257_50_4), .A2(n_257_50_5), .ZN(n_257_50_6));
   NAND2_X1 i_257_50_7 (.A1(CPU_Bus[31]), .A2(n_257_50_6), .ZN(n_257_50_7));
   INV_X1 i_257_50_8 (.A(n_255), .ZN(n_257_50_8));
   NAND2_X1 i_257_50_9 (.A1(n_257_50_0), .A2(n_257_50_8), .ZN(n_257_50_9));
   NOR2_X1 i_257_50_10 (.A1(n_257_50_9), .A2(n_257_50_2), .ZN(n_257_50_10));
   NAND2_X1 i_257_50_11 (.A1(n_257_50_10), .A2(n_257), .ZN(n_257_50_11));
   NOR2_X1 i_257_50_12 (.A1(n_257_50_11), .A2(n_257_50_5), .ZN(n_257_50_12));
   NAND2_X1 i_257_50_13 (.A1(CPU_Bus[29]), .A2(n_257_50_12), .ZN(n_257_50_13));
   NAND2_X1 i_257_50_14 (.A1(n_257_50_7), .A2(n_257_50_13), .ZN(n_257_50_14));
   NOR2_X1 i_257_50_15 (.A1(n_257_50_1), .A2(n_256), .ZN(n_257_50_15));
   NAND2_X1 i_257_50_16 (.A1(n_257_50_15), .A2(n_257), .ZN(n_257_50_16));
   NOR2_X1 i_257_50_17 (.A1(n_257_50_16), .A2(n_257_50_5), .ZN(n_257_50_17));
   NAND2_X1 i_257_50_18 (.A1(CPU_Bus[27]), .A2(n_257_50_17), .ZN(n_257_50_18));
   NOR2_X1 i_257_50_19 (.A1(n_257_50_9), .A2(n_256), .ZN(n_257_50_19));
   NAND2_X1 i_257_50_20 (.A1(n_257_50_19), .A2(n_257), .ZN(n_257_50_20));
   NOR2_X1 i_257_50_21 (.A1(n_257_50_20), .A2(n_257_50_5), .ZN(n_257_50_21));
   NAND2_X1 i_257_50_22 (.A1(CPU_Bus[25]), .A2(n_257_50_21), .ZN(n_257_50_22));
   NAND2_X1 i_257_50_23 (.A1(n_257_50_18), .A2(n_257_50_22), .ZN(n_257_50_23));
   NOR2_X1 i_257_50_24 (.A1(n_257_50_14), .A2(n_257_50_23), .ZN(n_257_50_24));
   INV_X1 i_257_50_25 (.A(n_257), .ZN(n_257_50_25));
   NAND2_X1 i_257_50_26 (.A1(n_257_50_3), .A2(n_257_50_25), .ZN(n_257_50_26));
   NOR2_X1 i_257_50_27 (.A1(n_257_50_26), .A2(n_257_50_5), .ZN(n_257_50_27));
   NAND2_X1 i_257_50_28 (.A1(CPU_Bus[23]), .A2(n_257_50_27), .ZN(n_257_50_28));
   NAND2_X1 i_257_50_29 (.A1(n_257_50_10), .A2(n_257_50_25), .ZN(n_257_50_29));
   NOR2_X1 i_257_50_30 (.A1(n_257_50_29), .A2(n_257_50_5), .ZN(n_257_50_30));
   NAND2_X1 i_257_50_31 (.A1(CPU_Bus[21]), .A2(n_257_50_30), .ZN(n_257_50_31));
   NAND2_X1 i_257_50_32 (.A1(n_257_50_28), .A2(n_257_50_31), .ZN(n_257_50_32));
   NAND2_X1 i_257_50_33 (.A1(n_257_50_15), .A2(n_257_50_25), .ZN(n_257_50_33));
   NOR2_X1 i_257_50_34 (.A1(n_257_50_33), .A2(n_257_50_5), .ZN(n_257_50_34));
   NAND2_X1 i_257_50_35 (.A1(CPU_Bus[19]), .A2(n_257_50_34), .ZN(n_257_50_35));
   NAND2_X1 i_257_50_36 (.A1(n_257_50_19), .A2(n_257_50_25), .ZN(n_257_50_36));
   NOR2_X1 i_257_50_37 (.A1(n_257_50_36), .A2(n_257_50_5), .ZN(n_257_50_37));
   NAND2_X1 i_257_50_38 (.A1(CPU_Bus[17]), .A2(n_257_50_37), .ZN(n_257_50_38));
   NAND2_X1 i_257_50_39 (.A1(n_257_50_35), .A2(n_257_50_38), .ZN(n_257_50_39));
   NOR2_X1 i_257_50_40 (.A1(n_257_50_32), .A2(n_257_50_39), .ZN(n_257_50_40));
   NAND2_X1 i_257_50_41 (.A1(n_257_50_24), .A2(n_257_50_40), .ZN(n_257_50_41));
   NOR2_X1 i_257_50_42 (.A1(n_257_50_4), .A2(n_258), .ZN(n_257_50_42));
   NAND2_X1 i_257_50_43 (.A1(CPU_Bus[15]), .A2(n_257_50_42), .ZN(n_257_50_43));
   NOR2_X1 i_257_50_44 (.A1(n_257_50_11), .A2(n_258), .ZN(n_257_50_44));
   NAND2_X1 i_257_50_45 (.A1(CPU_Bus[13]), .A2(n_257_50_44), .ZN(n_257_50_45));
   NAND2_X1 i_257_50_46 (.A1(n_257_50_43), .A2(n_257_50_45), .ZN(n_257_50_46));
   NOR2_X1 i_257_50_47 (.A1(n_257_50_16), .A2(n_258), .ZN(n_257_50_47));
   NAND2_X1 i_257_50_48 (.A1(CPU_Bus[11]), .A2(n_257_50_47), .ZN(n_257_50_48));
   NOR2_X1 i_257_50_49 (.A1(n_257_50_20), .A2(n_258), .ZN(n_257_50_49));
   NAND2_X1 i_257_50_50 (.A1(CPU_Bus[9]), .A2(n_257_50_49), .ZN(n_257_50_50));
   NAND2_X1 i_257_50_51 (.A1(n_257_50_48), .A2(n_257_50_50), .ZN(n_257_50_51));
   NOR2_X1 i_257_50_52 (.A1(n_257_50_46), .A2(n_257_50_51), .ZN(n_257_50_52));
   NOR2_X1 i_257_50_53 (.A1(n_257_50_26), .A2(n_258), .ZN(n_257_50_53));
   NAND2_X1 i_257_50_54 (.A1(CPU_Bus[7]), .A2(n_257_50_53), .ZN(n_257_50_54));
   NOR2_X1 i_257_50_55 (.A1(n_257_50_29), .A2(n_258), .ZN(n_257_50_55));
   NAND2_X1 i_257_50_56 (.A1(CPU_Bus[5]), .A2(n_257_50_55), .ZN(n_257_50_56));
   NAND2_X1 i_257_50_57 (.A1(n_257_50_54), .A2(n_257_50_56), .ZN(n_257_50_57));
   NOR2_X1 i_257_50_58 (.A1(n_257_50_33), .A2(n_258), .ZN(n_257_50_58));
   NAND2_X1 i_257_50_59 (.A1(CPU_Bus[3]), .A2(n_257_50_58), .ZN(n_257_50_59));
   NOR2_X1 i_257_50_60 (.A1(n_257_50_36), .A2(n_258), .ZN(n_257_50_60));
   NAND2_X1 i_257_50_61 (.A1(CPU_Bus[1]), .A2(n_257_50_60), .ZN(n_257_50_61));
   NAND2_X1 i_257_50_62 (.A1(n_257_50_59), .A2(n_257_50_61), .ZN(n_257_50_62));
   NOR2_X1 i_257_50_63 (.A1(n_257_50_57), .A2(n_257_50_62), .ZN(n_257_50_63));
   NAND2_X1 i_257_50_64 (.A1(n_257_50_52), .A2(n_257_50_63), .ZN(n_257_50_64));
   NOR2_X1 i_257_50_65 (.A1(n_257_50_41), .A2(n_257_50_64), .ZN(n_257_50_65));
   NAND2_X1 i_257_50_66 (.A1(n_257_50_8), .A2(n_254), .ZN(n_257_50_66));
   NOR2_X1 i_257_50_67 (.A1(n_257_50_66), .A2(n_257_50_2), .ZN(n_257_50_67));
   NAND2_X1 i_257_50_68 (.A1(n_257_50_67), .A2(n_257), .ZN(n_257_50_68));
   NOR2_X1 i_257_50_69 (.A1(n_257_50_68), .A2(n_257_50_5), .ZN(n_257_50_69));
   NAND2_X1 i_257_50_70 (.A1(CPU_Bus[30]), .A2(n_257_50_69), .ZN(n_257_50_70));
   NOR2_X1 i_257_50_71 (.A1(n_257_50_66), .A2(n_256), .ZN(n_257_50_71));
   NAND2_X1 i_257_50_72 (.A1(n_257_50_71), .A2(n_257), .ZN(n_257_50_72));
   NOR2_X1 i_257_50_73 (.A1(n_257_50_72), .A2(n_257_50_5), .ZN(n_257_50_73));
   NAND2_X1 i_257_50_74 (.A1(CPU_Bus[26]), .A2(n_257_50_73), .ZN(n_257_50_74));
   NAND2_X1 i_257_50_75 (.A1(n_257_50_70), .A2(n_257_50_74), .ZN(n_257_50_75));
   NAND2_X1 i_257_50_76 (.A1(n_257_50_67), .A2(n_257_50_25), .ZN(n_257_50_76));
   NOR2_X1 i_257_50_77 (.A1(n_257_50_76), .A2(n_257_50_5), .ZN(n_257_50_77));
   NAND2_X1 i_257_50_78 (.A1(CPU_Bus[22]), .A2(n_257_50_77), .ZN(n_257_50_78));
   NAND2_X1 i_257_50_79 (.A1(n_257_50_71), .A2(n_257_50_25), .ZN(n_257_50_79));
   NOR2_X1 i_257_50_80 (.A1(n_257_50_79), .A2(n_257_50_5), .ZN(n_257_50_80));
   NAND2_X1 i_257_50_81 (.A1(CPU_Bus[18]), .A2(n_257_50_80), .ZN(n_257_50_81));
   NAND2_X1 i_257_50_82 (.A1(n_257_50_78), .A2(n_257_50_81), .ZN(n_257_50_82));
   NOR2_X1 i_257_50_83 (.A1(n_257_50_75), .A2(n_257_50_82), .ZN(n_257_50_83));
   NOR2_X1 i_257_50_84 (.A1(n_257_50_68), .A2(n_258), .ZN(n_257_50_84));
   NAND2_X1 i_257_50_85 (.A1(CPU_Bus[14]), .A2(n_257_50_84), .ZN(n_257_50_85));
   NOR2_X1 i_257_50_86 (.A1(n_257_50_72), .A2(n_258), .ZN(n_257_50_86));
   NAND2_X1 i_257_50_87 (.A1(CPU_Bus[10]), .A2(n_257_50_86), .ZN(n_257_50_87));
   NAND2_X1 i_257_50_88 (.A1(n_257_50_85), .A2(n_257_50_87), .ZN(n_257_50_88));
   NOR2_X1 i_257_50_89 (.A1(n_257_50_76), .A2(n_258), .ZN(n_257_50_89));
   NAND2_X1 i_257_50_90 (.A1(CPU_Bus[6]), .A2(n_257_50_89), .ZN(n_257_50_90));
   NOR2_X1 i_257_50_91 (.A1(n_257_50_79), .A2(n_258), .ZN(n_257_50_91));
   NAND2_X1 i_257_50_92 (.A1(CPU_Bus[2]), .A2(n_257_50_91), .ZN(n_257_50_92));
   NAND2_X1 i_257_50_93 (.A1(n_257_50_90), .A2(n_257_50_92), .ZN(n_257_50_93));
   NOR2_X1 i_257_50_94 (.A1(n_257_50_88), .A2(n_257_50_93), .ZN(n_257_50_94));
   NAND2_X1 i_257_50_95 (.A1(n_257_50_83), .A2(n_257_50_94), .ZN(n_257_50_95));
   NAND2_X1 i_257_50_96 (.A1(n_254), .A2(n_255), .ZN(n_257_50_96));
   NOR2_X1 i_257_50_97 (.A1(n_257_50_96), .A2(n_257_50_2), .ZN(n_257_50_97));
   NAND2_X1 i_257_50_98 (.A1(n_257_50_97), .A2(n_257), .ZN(n_257_50_98));
   NOR2_X1 i_257_50_99 (.A1(n_257_50_98), .A2(n_257_50_5), .ZN(n_257_50_99));
   NAND2_X1 i_257_50_100 (.A1(CPU_Bus[0]), .A2(n_257_50_99), .ZN(n_257_50_100));
   NOR2_X1 i_257_50_101 (.A1(n_257_50_96), .A2(n_256), .ZN(n_257_50_101));
   NAND2_X1 i_257_50_102 (.A1(n_257_50_101), .A2(n_257), .ZN(n_257_50_102));
   NOR2_X1 i_257_50_103 (.A1(n_257_50_102), .A2(n_257_50_5), .ZN(n_257_50_103));
   NAND2_X1 i_257_50_104 (.A1(CPU_Bus[28]), .A2(n_257_50_103), .ZN(n_257_50_104));
   NAND2_X1 i_257_50_105 (.A1(n_257_50_100), .A2(n_257_50_104), .ZN(n_257_50_105));
   NAND2_X1 i_257_50_106 (.A1(n_257_50_97), .A2(n_257_50_25), .ZN(n_257_50_106));
   NOR2_X1 i_257_50_107 (.A1(n_257_50_106), .A2(n_257_50_5), .ZN(n_257_50_107));
   NAND2_X1 i_257_50_108 (.A1(CPU_Bus[24]), .A2(n_257_50_107), .ZN(n_257_50_108));
   NAND2_X1 i_257_50_109 (.A1(n_257_50_101), .A2(n_257_50_25), .ZN(n_257_50_109));
   NOR2_X1 i_257_50_110 (.A1(n_257_50_109), .A2(n_257_50_5), .ZN(n_257_50_110));
   NAND2_X1 i_257_50_111 (.A1(CPU_Bus[20]), .A2(n_257_50_110), .ZN(n_257_50_111));
   NAND2_X1 i_257_50_112 (.A1(n_257_50_108), .A2(n_257_50_111), .ZN(n_257_50_112));
   NOR2_X1 i_257_50_113 (.A1(n_257_50_105), .A2(n_257_50_112), .ZN(n_257_50_113));
   NOR2_X1 i_257_50_114 (.A1(n_257_50_98), .A2(n_258), .ZN(n_257_50_114));
   NAND2_X1 i_257_50_115 (.A1(CPU_Bus[16]), .A2(n_257_50_114), .ZN(n_257_50_115));
   NOR2_X1 i_257_50_116 (.A1(n_257_50_102), .A2(n_258), .ZN(n_257_50_116));
   NAND2_X1 i_257_50_117 (.A1(CPU_Bus[12]), .A2(n_257_50_116), .ZN(n_257_50_117));
   NAND2_X1 i_257_50_118 (.A1(n_257_50_115), .A2(n_257_50_117), .ZN(n_257_50_118));
   NOR2_X1 i_257_50_119 (.A1(n_257_50_106), .A2(n_258), .ZN(n_257_50_119));
   NAND2_X1 i_257_50_120 (.A1(CPU_Bus[8]), .A2(n_257_50_119), .ZN(n_257_50_120));
   NOR2_X1 i_257_50_121 (.A1(n_257_50_109), .A2(n_258), .ZN(n_257_50_121));
   NAND2_X1 i_257_50_122 (.A1(CPU_Bus[4]), .A2(n_257_50_121), .ZN(n_257_50_122));
   NAND2_X1 i_257_50_123 (.A1(n_257_50_120), .A2(n_257_50_122), .ZN(n_257_50_123));
   NOR2_X1 i_257_50_124 (.A1(n_257_50_118), .A2(n_257_50_123), .ZN(n_257_50_124));
   NAND2_X1 i_257_50_125 (.A1(n_257_50_113), .A2(n_257_50_124), .ZN(n_257_50_125));
   NOR2_X1 i_257_50_126 (.A1(n_257_50_95), .A2(n_257_50_125), .ZN(n_257_50_126));
   NAND2_X1 i_257_50_127 (.A1(n_257_50_65), .A2(n_257_50_126), .ZN(n_257_382));
   datapath__1_378 i_257_51 (.PacketSize(PacketSize), .p_0({n_257_387, uc_565, 
      uc_566, uc_567, uc_568, uc_569, uc_570, uc_571, uc_572, uc_573, uc_574, 
      uc_575, uc_576, uc_577, uc_578, uc_579, uc_580, uc_581, uc_582, uc_583, 
      uc_584, uc_585, uc_586, uc_587, uc_588, uc_589, uc_590, n_257_386, 
      n_257_385, n_257_384, n_257_383, uc_591}));
   datapath__1_379 i_257_52 (.p_0({uc_592, uc_593, uc_594, uc_595, uc_596, 
      uc_597, uc_598, uc_599, uc_600, uc_601, uc_602, uc_603, uc_604, uc_605, 
      uc_606, uc_607, uc_608, uc_609, uc_610, uc_611, uc_612, uc_613, uc_614, 
      uc_615, uc_616, n_257_387, 1'b0, n_257_386, n_257_385, n_257_384, 
      n_257_383, n_151}), .p_1({n_257_419, n_257_418, n_257_417, n_257_416, 
      n_257_415, n_257_414, n_257_413, n_257_412, n_257_411, n_257_410, 
      n_257_409, n_257_408, n_257_407, n_257_406, n_257_405, n_257_404, 
      n_257_403, n_257_402, n_257_401, n_257_400, n_257_399, n_257_398, 
      n_257_397, n_257_396, n_257_395, n_257_394, n_257_393, n_257_392, 
      n_257_391, n_257_390, n_257_389, n_257_388}));
   NOR2_X1 i_257_53_0 (.A1(n_36), .A2(n_37), .ZN(n_257_53_0));
   NAND4_X1 i_257_53_1 (.A1(n_32), .A2(n_33), .A3(n_34), .A4(n_35), .ZN(
      n_257_53_1));
   INV_X1 i_257_53_2 (.A(n_151), .ZN(n_257_53_2));
   OAI21_X1 i_257_53_3 (.A(n_257_53_0), .B1(n_257_53_1), .B2(n_257_53_2), 
      .ZN(n_257_420));
   NAND4_X1 i_257_54_0 (.A1(n_32), .A2(n_33), .A3(n_34), .A4(n_35), .ZN(
      n_257_54_0));
   NOR2_X1 i_257_54_1 (.A1(n_36), .A2(n_37), .ZN(n_257_54_1));
   NAND2_X1 i_257_54_2 (.A1(n_257_54_0), .A2(n_257_54_1), .ZN(n_257_421));
   OAI21_X1 i_257_55_0 (.A(n_257_55_0), .B1(n_257_55_2), .B2(n_257_55_1), 
      .ZN(n_257_422));
   NOR2_X1 i_257_55_1 (.A1(n_37), .A2(n_36), .ZN(n_257_55_0));
   NAND3_X1 i_257_55_2 (.A1(n_35), .A2(n_33), .A3(n_34), .ZN(n_257_55_1));
   NOR2_X1 i_257_55_3 (.A1(n_32), .A2(n_151), .ZN(n_257_55_2));
   NAND3_X1 i_257_56_0 (.A1(n_33), .A2(n_34), .A3(n_35), .ZN(n_257_56_0));
   NOR2_X1 i_257_56_1 (.A1(n_36), .A2(n_37), .ZN(n_257_56_1));
   NAND2_X1 i_257_56_2 (.A1(n_257_56_0), .A2(n_257_56_1), .ZN(n_257_423));
   OAI21_X1 i_257_57_0 (.A(n_257_57_0), .B1(n_257_57_2), .B2(n_257_57_1), 
      .ZN(n_257_424));
   NOR2_X1 i_257_57_1 (.A1(n_37), .A2(n_36), .ZN(n_257_57_0));
   NAND2_X1 i_257_57_2 (.A1(n_35), .A2(n_34), .ZN(n_257_57_1));
   AOI21_X1 i_257_57_3 (.A(n_33), .B1(n_32), .B2(n_151), .ZN(n_257_57_2));
   OAI211_X1 i_257_58_0 (.A(n_35), .B(n_34), .C1(n_32), .C2(n_33), .ZN(
      n_257_58_0));
   NOR2_X1 i_257_58_1 (.A1(n_36), .A2(n_37), .ZN(n_257_58_1));
   NAND2_X1 i_257_58_2 (.A1(n_257_58_0), .A2(n_257_58_1), .ZN(n_257_425));
   OR3_X1 i_257_59_0 (.A1(n_151), .A2(n_32), .A3(n_33), .ZN(n_257_59_0));
   NAND3_X1 i_257_59_1 (.A1(n_257_59_0), .A2(n_34), .A3(n_35), .ZN(n_257_59_1));
   NOR2_X1 i_257_59_2 (.A1(n_36), .A2(n_37), .ZN(n_257_59_2));
   NAND2_X1 i_257_59_3 (.A1(n_257_59_1), .A2(n_257_59_2), .ZN(n_257_426));
   INV_X1 i_257_60_0 (.A(n_257_60_0), .ZN(n_257_427));
   AOI211_X1 i_257_60_1 (.A(n_37), .B(n_36), .C1(n_35), .C2(n_34), .ZN(
      n_257_60_0));
   AND3_X1 i_257_61_0 (.A1(n_151), .A2(n_32), .A3(n_33), .ZN(n_257_61_0));
   OAI21_X1 i_257_61_1 (.A(n_35), .B1(n_257_61_0), .B2(n_34), .ZN(n_257_61_1));
   NOR2_X1 i_257_61_2 (.A1(n_36), .A2(n_37), .ZN(n_257_61_2));
   NAND2_X1 i_257_61_3 (.A1(n_257_61_1), .A2(n_257_61_2), .ZN(n_257_428));
   NOR2_X1 i_257_62_0 (.A1(n_36), .A2(n_37), .ZN(n_257_62_0));
   AOI21_X1 i_257_62_1 (.A(n_34), .B1(n_32), .B2(n_33), .ZN(n_257_62_1));
   INV_X1 i_257_62_2 (.A(n_35), .ZN(n_257_62_2));
   OAI21_X1 i_257_62_3 (.A(n_257_62_0), .B1(n_257_62_1), .B2(n_257_62_2), 
      .ZN(n_257_429));
   OAI21_X1 i_257_63_0 (.A(n_33), .B1(n_151), .B2(n_32), .ZN(n_257_63_0));
   INV_X1 i_257_63_1 (.A(n_257_63_0), .ZN(n_257_63_1));
   OAI21_X1 i_257_63_2 (.A(n_35), .B1(n_257_63_1), .B2(n_34), .ZN(n_257_63_2));
   NOR2_X1 i_257_63_3 (.A1(n_36), .A2(n_37), .ZN(n_257_63_3));
   NAND2_X1 i_257_63_4 (.A1(n_257_63_2), .A2(n_257_63_3), .ZN(n_257_430));
   OAI21_X1 i_257_64_0 (.A(n_35), .B1(n_33), .B2(n_34), .ZN(n_257_64_0));
   NOR2_X1 i_257_64_1 (.A1(n_36), .A2(n_37), .ZN(n_257_64_1));
   NAND2_X1 i_257_64_2 (.A1(n_257_64_0), .A2(n_257_64_1), .ZN(n_257_431));
   NAND3_X1 i_257_65_0 (.A1(n_257_65_4), .A2(n_257_65_5), .A3(n_257_65_0), 
      .ZN(n_257_432));
   OAI21_X1 i_257_65_1 (.A(n_35), .B1(n_34), .B2(n_257_65_1), .ZN(n_257_65_0));
   NAND2_X1 i_257_65_2 (.A1(n_257_65_2), .A2(n_257_65_3), .ZN(n_257_65_1));
   NAND2_X1 i_257_65_3 (.A1(n_32), .A2(n_151), .ZN(n_257_65_2));
   INV_X1 i_257_65_4 (.A(n_33), .ZN(n_257_65_3));
   INV_X1 i_257_65_5 (.A(n_36), .ZN(n_257_65_4));
   INV_X1 i_257_65_6 (.A(n_37), .ZN(n_257_65_5));
   NOR2_X1 i_257_66_0 (.A1(n_36), .A2(n_37), .ZN(n_257_66_0));
   NOR3_X1 i_257_66_1 (.A1(n_32), .A2(n_33), .A3(n_34), .ZN(n_257_66_1));
   INV_X1 i_257_66_2 (.A(n_35), .ZN(n_257_66_2));
   OAI21_X1 i_257_66_3 (.A(n_257_66_0), .B1(n_257_66_1), .B2(n_257_66_2), 
      .ZN(n_257_433));
   INV_X1 i_257_67_0 (.A(n_254), .ZN(n_257_67_0));
   NAND2_X1 i_257_67_1 (.A1(n_257_67_0), .A2(n_255), .ZN(n_257_67_1));
   INV_X1 i_257_67_2 (.A(n_256), .ZN(n_257_67_2));
   NOR2_X1 i_257_67_3 (.A1(n_257_67_1), .A2(n_257_67_2), .ZN(n_257_67_3));
   NAND2_X1 i_257_67_4 (.A1(n_257_67_3), .A2(n_257), .ZN(n_257_67_4));
   INV_X1 i_257_67_5 (.A(n_258), .ZN(n_257_67_5));
   NOR2_X1 i_257_67_6 (.A1(n_257_67_4), .A2(n_257_67_5), .ZN(n_257_67_6));
   NAND2_X1 i_257_67_7 (.A1(CPU_Bus[13]), .A2(n_257_67_6), .ZN(n_257_67_7));
   INV_X1 i_257_67_8 (.A(n_255), .ZN(n_257_67_8));
   NAND2_X1 i_257_67_9 (.A1(n_257_67_0), .A2(n_257_67_8), .ZN(n_257_67_9));
   NOR2_X1 i_257_67_10 (.A1(n_257_67_9), .A2(n_257_67_2), .ZN(n_257_67_10));
   NAND2_X1 i_257_67_11 (.A1(n_257_67_10), .A2(n_257), .ZN(n_257_67_11));
   NOR2_X1 i_257_67_12 (.A1(n_257_67_11), .A2(n_257_67_5), .ZN(n_257_67_12));
   NAND2_X1 i_257_67_13 (.A1(CPU_Bus[11]), .A2(n_257_67_12), .ZN(n_257_67_13));
   NAND2_X1 i_257_67_14 (.A1(n_257_67_7), .A2(n_257_67_13), .ZN(n_257_67_14));
   NOR2_X1 i_257_67_15 (.A1(n_257_67_1), .A2(n_256), .ZN(n_257_67_15));
   NAND2_X1 i_257_67_16 (.A1(n_257_67_15), .A2(n_257), .ZN(n_257_67_16));
   NOR2_X1 i_257_67_17 (.A1(n_257_67_16), .A2(n_257_67_5), .ZN(n_257_67_17));
   NAND2_X1 i_257_67_18 (.A1(CPU_Bus[9]), .A2(n_257_67_17), .ZN(n_257_67_18));
   NOR2_X1 i_257_67_19 (.A1(n_257_67_9), .A2(n_256), .ZN(n_257_67_19));
   NAND2_X1 i_257_67_20 (.A1(n_257_67_19), .A2(n_257), .ZN(n_257_67_20));
   NOR2_X1 i_257_67_21 (.A1(n_257_67_20), .A2(n_257_67_5), .ZN(n_257_67_21));
   NAND2_X1 i_257_67_22 (.A1(CPU_Bus[7]), .A2(n_257_67_21), .ZN(n_257_67_22));
   NAND2_X1 i_257_67_23 (.A1(n_257_67_18), .A2(n_257_67_22), .ZN(n_257_67_23));
   NOR2_X1 i_257_67_24 (.A1(n_257_67_14), .A2(n_257_67_23), .ZN(n_257_67_24));
   INV_X1 i_257_67_25 (.A(n_257), .ZN(n_257_67_25));
   NAND2_X1 i_257_67_26 (.A1(n_257_67_3), .A2(n_257_67_25), .ZN(n_257_67_26));
   NOR2_X1 i_257_67_27 (.A1(n_257_67_26), .A2(n_257_67_5), .ZN(n_257_67_27));
   NAND2_X1 i_257_67_28 (.A1(CPU_Bus[5]), .A2(n_257_67_27), .ZN(n_257_67_28));
   NAND2_X1 i_257_67_29 (.A1(n_257_67_10), .A2(n_257_67_25), .ZN(n_257_67_29));
   NOR2_X1 i_257_67_30 (.A1(n_257_67_29), .A2(n_257_67_5), .ZN(n_257_67_30));
   NAND2_X1 i_257_67_31 (.A1(CPU_Bus[3]), .A2(n_257_67_30), .ZN(n_257_67_31));
   NAND2_X1 i_257_67_32 (.A1(n_257_67_28), .A2(n_257_67_31), .ZN(n_257_67_32));
   NAND2_X1 i_257_67_33 (.A1(n_257_67_15), .A2(n_257_67_25), .ZN(n_257_67_33));
   NOR2_X1 i_257_67_34 (.A1(n_257_67_33), .A2(n_257_67_5), .ZN(n_257_67_34));
   NAND2_X1 i_257_67_35 (.A1(CPU_Bus[1]), .A2(n_257_67_34), .ZN(n_257_67_35));
   NAND2_X1 i_257_67_36 (.A1(n_257_67_19), .A2(n_257_67_25), .ZN(n_257_67_36));
   NOR2_X1 i_257_67_37 (.A1(n_257_67_36), .A2(n_257_67_5), .ZN(n_257_67_37));
   NAND2_X1 i_257_67_38 (.A1(CPU_Bus[31]), .A2(n_257_67_37), .ZN(n_257_67_38));
   NAND2_X1 i_257_67_39 (.A1(n_257_67_35), .A2(n_257_67_38), .ZN(n_257_67_39));
   NOR2_X1 i_257_67_40 (.A1(n_257_67_32), .A2(n_257_67_39), .ZN(n_257_67_40));
   NAND2_X1 i_257_67_41 (.A1(n_257_67_24), .A2(n_257_67_40), .ZN(n_257_67_41));
   NOR2_X1 i_257_67_42 (.A1(n_257_67_4), .A2(n_258), .ZN(n_257_67_42));
   NAND2_X1 i_257_67_43 (.A1(CPU_Bus[29]), .A2(n_257_67_42), .ZN(n_257_67_43));
   NOR2_X1 i_257_67_44 (.A1(n_257_67_11), .A2(n_258), .ZN(n_257_67_44));
   NAND2_X1 i_257_67_45 (.A1(CPU_Bus[27]), .A2(n_257_67_44), .ZN(n_257_67_45));
   NAND2_X1 i_257_67_46 (.A1(n_257_67_43), .A2(n_257_67_45), .ZN(n_257_67_46));
   NOR2_X1 i_257_67_47 (.A1(n_257_67_16), .A2(n_258), .ZN(n_257_67_47));
   NAND2_X1 i_257_67_48 (.A1(CPU_Bus[25]), .A2(n_257_67_47), .ZN(n_257_67_48));
   NOR2_X1 i_257_67_49 (.A1(n_257_67_20), .A2(n_258), .ZN(n_257_67_49));
   NAND2_X1 i_257_67_50 (.A1(CPU_Bus[23]), .A2(n_257_67_49), .ZN(n_257_67_50));
   NAND2_X1 i_257_67_51 (.A1(n_257_67_48), .A2(n_257_67_50), .ZN(n_257_67_51));
   NOR2_X1 i_257_67_52 (.A1(n_257_67_46), .A2(n_257_67_51), .ZN(n_257_67_52));
   NOR2_X1 i_257_67_53 (.A1(n_257_67_26), .A2(n_258), .ZN(n_257_67_53));
   NAND2_X1 i_257_67_54 (.A1(CPU_Bus[21]), .A2(n_257_67_53), .ZN(n_257_67_54));
   NOR2_X1 i_257_67_55 (.A1(n_257_67_29), .A2(n_258), .ZN(n_257_67_55));
   NAND2_X1 i_257_67_56 (.A1(CPU_Bus[19]), .A2(n_257_67_55), .ZN(n_257_67_56));
   NAND2_X1 i_257_67_57 (.A1(n_257_67_54), .A2(n_257_67_56), .ZN(n_257_67_57));
   NOR2_X1 i_257_67_58 (.A1(n_257_67_33), .A2(n_258), .ZN(n_257_67_58));
   NAND2_X1 i_257_67_59 (.A1(CPU_Bus[17]), .A2(n_257_67_58), .ZN(n_257_67_59));
   NOR2_X1 i_257_67_60 (.A1(n_257_67_36), .A2(n_258), .ZN(n_257_67_60));
   NAND2_X1 i_257_67_61 (.A1(CPU_Bus[15]), .A2(n_257_67_60), .ZN(n_257_67_61));
   NAND2_X1 i_257_67_62 (.A1(n_257_67_59), .A2(n_257_67_61), .ZN(n_257_67_62));
   NOR2_X1 i_257_67_63 (.A1(n_257_67_57), .A2(n_257_67_62), .ZN(n_257_67_63));
   NAND2_X1 i_257_67_64 (.A1(n_257_67_52), .A2(n_257_67_63), .ZN(n_257_67_64));
   NOR2_X1 i_257_67_65 (.A1(n_257_67_41), .A2(n_257_67_64), .ZN(n_257_67_65));
   NAND2_X1 i_257_67_66 (.A1(n_257_67_8), .A2(n_254), .ZN(n_257_67_66));
   NOR2_X1 i_257_67_67 (.A1(n_257_67_66), .A2(n_257_67_2), .ZN(n_257_67_67));
   NAND2_X1 i_257_67_68 (.A1(n_257_67_67), .A2(n_257), .ZN(n_257_67_68));
   NOR2_X1 i_257_67_69 (.A1(n_257_67_68), .A2(n_257_67_5), .ZN(n_257_67_69));
   NAND2_X1 i_257_67_70 (.A1(CPU_Bus[12]), .A2(n_257_67_69), .ZN(n_257_67_70));
   NOR2_X1 i_257_67_71 (.A1(n_257_67_66), .A2(n_256), .ZN(n_257_67_71));
   NAND2_X1 i_257_67_72 (.A1(n_257_67_71), .A2(n_257), .ZN(n_257_67_72));
   NOR2_X1 i_257_67_73 (.A1(n_257_67_72), .A2(n_257_67_5), .ZN(n_257_67_73));
   NAND2_X1 i_257_67_74 (.A1(CPU_Bus[8]), .A2(n_257_67_73), .ZN(n_257_67_74));
   NAND2_X1 i_257_67_75 (.A1(n_257_67_70), .A2(n_257_67_74), .ZN(n_257_67_75));
   NAND2_X1 i_257_67_76 (.A1(n_257_67_67), .A2(n_257_67_25), .ZN(n_257_67_76));
   NOR2_X1 i_257_67_77 (.A1(n_257_67_76), .A2(n_257_67_5), .ZN(n_257_67_77));
   NAND2_X1 i_257_67_78 (.A1(CPU_Bus[4]), .A2(n_257_67_77), .ZN(n_257_67_78));
   NAND2_X1 i_257_67_79 (.A1(n_257_67_71), .A2(n_257_67_25), .ZN(n_257_67_79));
   NOR2_X1 i_257_67_80 (.A1(n_257_67_79), .A2(n_257_67_5), .ZN(n_257_67_80));
   NAND2_X1 i_257_67_81 (.A1(CPU_Bus[0]), .A2(n_257_67_80), .ZN(n_257_67_81));
   NAND2_X1 i_257_67_82 (.A1(n_257_67_78), .A2(n_257_67_81), .ZN(n_257_67_82));
   NOR2_X1 i_257_67_83 (.A1(n_257_67_75), .A2(n_257_67_82), .ZN(n_257_67_83));
   NOR2_X1 i_257_67_84 (.A1(n_257_67_68), .A2(n_258), .ZN(n_257_67_84));
   NAND2_X1 i_257_67_85 (.A1(CPU_Bus[28]), .A2(n_257_67_84), .ZN(n_257_67_85));
   NOR2_X1 i_257_67_86 (.A1(n_257_67_72), .A2(n_258), .ZN(n_257_67_86));
   NAND2_X1 i_257_67_87 (.A1(CPU_Bus[24]), .A2(n_257_67_86), .ZN(n_257_67_87));
   NAND2_X1 i_257_67_88 (.A1(n_257_67_85), .A2(n_257_67_87), .ZN(n_257_67_88));
   NOR2_X1 i_257_67_89 (.A1(n_257_67_76), .A2(n_258), .ZN(n_257_67_89));
   NAND2_X1 i_257_67_90 (.A1(CPU_Bus[20]), .A2(n_257_67_89), .ZN(n_257_67_90));
   NOR2_X1 i_257_67_91 (.A1(n_257_67_79), .A2(n_258), .ZN(n_257_67_91));
   NAND2_X1 i_257_67_92 (.A1(CPU_Bus[16]), .A2(n_257_67_91), .ZN(n_257_67_92));
   NAND2_X1 i_257_67_93 (.A1(n_257_67_90), .A2(n_257_67_92), .ZN(n_257_67_93));
   NOR2_X1 i_257_67_94 (.A1(n_257_67_88), .A2(n_257_67_93), .ZN(n_257_67_94));
   NAND2_X1 i_257_67_95 (.A1(n_257_67_83), .A2(n_257_67_94), .ZN(n_257_67_95));
   NAND2_X1 i_257_67_96 (.A1(n_254), .A2(n_255), .ZN(n_257_67_96));
   NOR2_X1 i_257_67_97 (.A1(n_257_67_96), .A2(n_257_67_2), .ZN(n_257_67_97));
   NAND2_X1 i_257_67_98 (.A1(n_257_67_97), .A2(n_257), .ZN(n_257_67_98));
   NOR2_X1 i_257_67_99 (.A1(n_257_67_98), .A2(n_257_67_5), .ZN(n_257_67_99));
   NAND2_X1 i_257_67_100 (.A1(CPU_Bus[14]), .A2(n_257_67_99), .ZN(n_257_67_100));
   NOR2_X1 i_257_67_101 (.A1(n_257_67_96), .A2(n_256), .ZN(n_257_67_101));
   NAND2_X1 i_257_67_102 (.A1(n_257_67_101), .A2(n_257), .ZN(n_257_67_102));
   NOR2_X1 i_257_67_103 (.A1(n_257_67_102), .A2(n_257_67_5), .ZN(n_257_67_103));
   NAND2_X1 i_257_67_104 (.A1(CPU_Bus[10]), .A2(n_257_67_103), .ZN(n_257_67_104));
   NAND2_X1 i_257_67_105 (.A1(n_257_67_100), .A2(n_257_67_104), .ZN(n_257_67_105));
   NAND2_X1 i_257_67_106 (.A1(n_257_67_97), .A2(n_257_67_25), .ZN(n_257_67_106));
   NOR2_X1 i_257_67_107 (.A1(n_257_67_106), .A2(n_257_67_5), .ZN(n_257_67_107));
   NAND2_X1 i_257_67_108 (.A1(CPU_Bus[6]), .A2(n_257_67_107), .ZN(n_257_67_108));
   NAND2_X1 i_257_67_109 (.A1(n_257_67_101), .A2(n_257_67_25), .ZN(n_257_67_109));
   NOR2_X1 i_257_67_110 (.A1(n_257_67_109), .A2(n_257_67_5), .ZN(n_257_67_110));
   NAND2_X1 i_257_67_111 (.A1(CPU_Bus[2]), .A2(n_257_67_110), .ZN(n_257_67_111));
   NAND2_X1 i_257_67_112 (.A1(n_257_67_108), .A2(n_257_67_111), .ZN(n_257_67_112));
   NOR2_X1 i_257_67_113 (.A1(n_257_67_105), .A2(n_257_67_112), .ZN(n_257_67_113));
   NOR2_X1 i_257_67_114 (.A1(n_257_67_98), .A2(n_258), .ZN(n_257_67_114));
   NAND2_X1 i_257_67_115 (.A1(CPU_Bus[30]), .A2(n_257_67_114), .ZN(n_257_67_115));
   NOR2_X1 i_257_67_116 (.A1(n_257_67_102), .A2(n_258), .ZN(n_257_67_116));
   NAND2_X1 i_257_67_117 (.A1(CPU_Bus[26]), .A2(n_257_67_116), .ZN(n_257_67_117));
   NAND2_X1 i_257_67_118 (.A1(n_257_67_115), .A2(n_257_67_117), .ZN(n_257_67_118));
   NOR2_X1 i_257_67_119 (.A1(n_257_67_106), .A2(n_258), .ZN(n_257_67_119));
   NAND2_X1 i_257_67_120 (.A1(CPU_Bus[22]), .A2(n_257_67_119), .ZN(n_257_67_120));
   NOR2_X1 i_257_67_121 (.A1(n_257_67_109), .A2(n_258), .ZN(n_257_67_121));
   NAND2_X1 i_257_67_122 (.A1(CPU_Bus[18]), .A2(n_257_67_121), .ZN(n_257_67_122));
   NAND2_X1 i_257_67_123 (.A1(n_257_67_120), .A2(n_257_67_122), .ZN(n_257_67_123));
   NOR2_X1 i_257_67_124 (.A1(n_257_67_118), .A2(n_257_67_123), .ZN(n_257_67_124));
   NAND2_X1 i_257_67_125 (.A1(n_257_67_113), .A2(n_257_67_124), .ZN(n_257_67_125));
   NOR2_X1 i_257_67_126 (.A1(n_257_67_95), .A2(n_257_67_125), .ZN(n_257_67_126));
   NAND2_X1 i_257_67_127 (.A1(n_257_67_65), .A2(n_257_67_126), .ZN(n_257_434));
   OAI211_X1 i_257_68_0 (.A(n_34), .B(n_33), .C1(n_151), .C2(n_32), .ZN(
      n_257_68_0));
   NOR3_X1 i_257_68_1 (.A1(n_35), .A2(n_36), .A3(n_37), .ZN(n_257_68_1));
   NAND2_X1 i_257_68_2 (.A1(n_257_68_0), .A2(n_257_68_1), .ZN(n_257_435));
   NOR3_X1 i_257_69_0 (.A1(n_35), .A2(n_36), .A3(n_37), .ZN(n_257_69_0));
   NAND2_X1 i_257_69_1 (.A1(n_33), .A2(n_34), .ZN(n_257_69_1));
   NAND2_X1 i_257_69_2 (.A1(n_257_69_0), .A2(n_257_69_1), .ZN(n_257_436));
   OAI21_X1 i_257_70_0 (.A(n_34), .B1(n_32), .B2(n_33), .ZN(n_257_70_0));
   NOR3_X1 i_257_70_1 (.A1(n_35), .A2(n_36), .A3(n_37), .ZN(n_257_70_1));
   NAND2_X1 i_257_70_2 (.A1(n_257_70_0), .A2(n_257_70_1), .ZN(n_257_437));
   NAND3_X1 i_257_71_0 (.A1(n_151), .A2(n_32), .A3(n_33), .ZN(n_257_71_0));
   NOR4_X1 i_257_71_1 (.A1(n_34), .A2(n_35), .A3(n_36), .A4(n_37), .ZN(
      n_257_71_1));
   NAND2_X1 i_257_71_2 (.A1(n_257_71_0), .A2(n_257_71_1), .ZN(n_257_438));
   NOR4_X1 i_257_72_0 (.A1(n_34), .A2(n_35), .A3(n_36), .A4(n_37), .ZN(
      n_257_72_0));
   NAND2_X1 i_257_72_1 (.A1(n_32), .A2(n_33), .ZN(n_257_72_1));
   NAND2_X1 i_257_72_2 (.A1(n_257_72_0), .A2(n_257_72_1), .ZN(n_257_439));
   NOR4_X1 i_257_73_0 (.A1(n_34), .A2(n_35), .A3(n_36), .A4(n_37), .ZN(
      n_257_73_0));
   OAI21_X1 i_257_73_1 (.A(n_33), .B1(n_151), .B2(n_32), .ZN(n_257_73_1));
   NAND2_X1 i_257_73_2 (.A1(n_257_73_0), .A2(n_257_73_1), .ZN(n_257_440));
   OR4_X1 i_257_74_0 (.A1(n_34), .A2(n_35), .A3(n_36), .A4(n_37), .ZN(n_257_74_0));
   OR2_X1 i_257_74_1 (.A1(n_257_74_0), .A2(n_33), .ZN(n_257_441));
   HA_X1 i_257_75_0 (.A(PacketSize[2]), .B(n_257_75_256), .CO(n_257_75_1), 
      .S(n_257_75_0));
   HA_X1 i_257_75_1 (.A(PacketSize[2]), .B(PacketSize[1]), .CO(n_257_75_3), 
      .S(n_257_75_2));
   HA_X1 i_257_75_2 (.A(PacketSize[1]), .B(PacketSize[0]), .CO(n_257_75_5), 
      .S(n_257_75_4));
   HA_X1 i_257_75_3 (.A(PacketSize[2]), .B(n_257_75_5), .CO(n_257_75_7), 
      .S(n_257_75_6));
   HA_X1 i_257_75_4 (.A(PacketSize[4]), .B(PacketSize[3]), .CO(n_257_75_9), 
      .S(n_257_75_8));
   HA_X1 i_257_75_5 (.A(PacketSize[3]), .B(n_257_75_254), .CO(n_257_75_11), 
      .S(n_257_75_10));
   HA_X1 i_257_75_6 (.A(PacketSize[3]), .B(n_257_75_307), .CO(n_257_75_13), 
      .S(n_257_75_12));
   HA_X1 i_257_75_7 (.A(PacketSize[3]), .B(n_257_75_127), .CO(n_257_75_15), 
      .S(n_257_75_14));
   HA_X1 i_257_75_8 (.A(PacketSize[4]), .B(n_257_75_19), .CO(n_257_75_17), 
      .S(n_257_75_16));
   HA_X1 i_257_75_9 (.A(PacketSize[3]), .B(PacketSize[2]), .CO(n_257_75_19), 
      .S(n_257_75_18));
   HA_X1 i_257_75_10 (.A(PacketSize[3]), .B(n_257_75_1), .CO(n_257_75_21), 
      .S(n_257_75_20));
   HA_X1 i_257_75_11 (.A(PacketSize[3]), .B(n_257_75_3), .CO(n_257_75_23), 
      .S(n_257_75_22));
   HA_X1 i_257_75_12 (.A(PacketSize[3]), .B(n_257_75_7), .CO(n_257_75_25), 
      .S(n_257_75_24));
   HA_X1 i_257_75_13 (.A(PacketSize[4]), .B(n_257_75_76), .CO(n_257_75_27), 
      .S(n_257_75_26));
   HA_X1 i_257_75_14 (.A(PacketSize[4]), .B(n_257_75_265), .CO(n_257_75_29), 
      .S(n_257_75_28));
   HA_X1 i_257_75_15 (.A(PacketSize[4]), .B(n_257_75_13), .CO(n_257_75_31), 
      .S(n_257_75_30));
   HA_X1 i_257_75_16 (.A(PacketSize[4]), .B(n_257_75_264), .CO(n_257_75_33), 
      .S(n_257_75_32));
   NAND3_X1 i_257_75_17 (.A1(n_257_75_306), .A2(n_257_75_304), .A3(n_257_75_303), 
      .ZN(n_257_444));
   OAI21_X1 i_257_75_18 (.A(n_257_75_304), .B1(n_257_75_294), .B2(n_257_75_34), 
      .ZN(n_257_449));
   NAND2_X1 i_257_75_19 (.A1(n_257_75_304), .A2(n_257_75_34), .ZN(n_257_448));
   NAND3_X1 i_257_75_20 (.A1(n_33), .A2(n_32), .A3(n_34), .ZN(n_257_75_34));
   AOI21_X1 i_257_75_21 (.A(n_257_75_304), .B1(n_257_75_302), .B2(n_257_75_35), 
      .ZN(n_257_451));
   NOR2_X1 i_257_75_22 (.A1(n_34), .A2(n_257_484), .ZN(n_257_75_35));
   INV_X1 i_257_75_23 (.A(n_257_75_304), .ZN(n_257_450));
   NOR2_X1 i_257_75_24 (.A1(n_257_75_246), .A2(n_257_75_36), .ZN(n_257_452));
   NOR2_X1 i_257_75_25 (.A1(n_257_75_247), .A2(n_257_75_36), .ZN(n_257_453));
   NOR2_X1 i_257_75_26 (.A1(n_257_75_248), .A2(n_257_75_36), .ZN(n_257_454));
   NOR2_X1 i_257_75_27 (.A1(n_257_75_249), .A2(n_257_75_36), .ZN(n_257_455));
   NOR2_X1 i_257_75_28 (.A1(n_257_75_250), .A2(n_257_75_36), .ZN(n_257_456));
   NOR2_X1 i_257_75_29 (.A1(n_257_75_252), .A2(n_257_75_36), .ZN(n_257_457));
   NOR2_X1 i_257_75_30 (.A1(n_257_75_254), .A2(n_257_75_36), .ZN(n_257_458));
   NOR2_X1 i_257_75_31 (.A1(n_257_75_258), .A2(n_257_75_36), .ZN(n_257_459));
   OR2_X1 i_257_75_32 (.A1(n_257_1093), .A2(n_257_75_38), .ZN(n_257_75_36));
   NOR2_X1 i_257_75_33 (.A1(n_257_75_246), .A2(n_257_75_37), .ZN(n_257_460));
   NOR2_X1 i_257_75_34 (.A1(n_257_75_247), .A2(n_257_75_37), .ZN(n_257_461));
   NOR2_X1 i_257_75_35 (.A1(n_257_75_248), .A2(n_257_75_37), .ZN(n_257_462));
   NOR2_X1 i_257_75_36 (.A1(n_257_75_249), .A2(n_257_75_37), .ZN(n_257_463));
   NOR2_X1 i_257_75_37 (.A1(n_257_75_250), .A2(n_257_75_37), .ZN(n_257_464));
   NOR2_X1 i_257_75_38 (.A1(n_257_75_252), .A2(n_257_75_37), .ZN(n_257_465));
   NOR2_X1 i_257_75_39 (.A1(n_257_75_254), .A2(n_257_75_37), .ZN(n_257_466));
   NOR2_X1 i_257_75_40 (.A1(n_257_75_258), .A2(n_257_75_37), .ZN(n_257_467));
   OR2_X1 i_257_75_41 (.A1(n_257_75_261), .A2(n_257_75_38), .ZN(n_257_75_37));
   NAND2_X1 i_257_75_42 (.A1(n_257_75_266), .A2(n_257_75_42), .ZN(n_257_75_38));
   NOR2_X1 i_257_75_43 (.A1(n_257_75_246), .A2(n_257_75_39), .ZN(n_257_468));
   NOR2_X1 i_257_75_44 (.A1(n_257_75_247), .A2(n_257_75_39), .ZN(n_257_469));
   NOR2_X1 i_257_75_45 (.A1(n_257_75_248), .A2(n_257_75_39), .ZN(n_257_470));
   NOR2_X1 i_257_75_46 (.A1(n_257_75_249), .A2(n_257_75_39), .ZN(n_257_471));
   NOR2_X1 i_257_75_47 (.A1(n_257_75_250), .A2(n_257_75_39), .ZN(n_257_472));
   NOR2_X1 i_257_75_48 (.A1(n_257_75_252), .A2(n_257_75_39), .ZN(n_257_473));
   NOR2_X1 i_257_75_49 (.A1(n_257_75_254), .A2(n_257_75_39), .ZN(n_257_474));
   NOR2_X1 i_257_75_50 (.A1(n_257_75_258), .A2(n_257_75_39), .ZN(n_257_475));
   OR2_X1 i_257_75_51 (.A1(n_257_1093), .A2(n_257_75_41), .ZN(n_257_75_39));
   NOR2_X1 i_257_75_52 (.A1(n_257_75_246), .A2(n_257_75_40), .ZN(n_257_476));
   NOR2_X1 i_257_75_53 (.A1(n_257_75_247), .A2(n_257_75_40), .ZN(n_257_477));
   NOR2_X1 i_257_75_54 (.A1(n_257_75_248), .A2(n_257_75_40), .ZN(n_257_478));
   NOR2_X1 i_257_75_55 (.A1(n_257_75_249), .A2(n_257_75_40), .ZN(n_257_479));
   NOR2_X1 i_257_75_56 (.A1(n_257_75_250), .A2(n_257_75_40), .ZN(n_257_480));
   NOR2_X1 i_257_75_57 (.A1(n_257_75_252), .A2(n_257_75_40), .ZN(n_257_481));
   NOR2_X1 i_257_75_58 (.A1(n_257_75_254), .A2(n_257_75_40), .ZN(n_257_482));
   NOR2_X1 i_257_75_59 (.A1(n_257_75_258), .A2(n_257_75_40), .ZN(n_257_483));
   OR2_X1 i_257_75_60 (.A1(n_257_75_261), .A2(n_257_75_41), .ZN(n_257_75_40));
   NAND2_X1 i_257_75_61 (.A1(n_257_75_32), .A2(n_257_75_42), .ZN(n_257_75_41));
   XOR2_X1 i_257_75_62 (.A(PacketSize[5]), .B(n_257_75_33), .Z(n_257_75_42));
   NOR2_X1 i_257_75_63 (.A1(n_257_75_254), .A2(n_257_75_43), .ZN(n_257_485));
   NOR2_X1 i_257_75_64 (.A1(n_257_75_258), .A2(n_257_75_43), .ZN(n_257_486));
   NOR2_X1 i_257_75_65 (.A1(n_257_75_246), .A2(n_257_75_43), .ZN(n_257_487));
   NOR2_X1 i_257_75_66 (.A1(n_257_75_247), .A2(n_257_75_43), .ZN(n_257_488));
   NOR2_X1 i_257_75_67 (.A1(n_257_75_248), .A2(n_257_75_43), .ZN(n_257_489));
   NOR2_X1 i_257_75_68 (.A1(n_257_75_249), .A2(n_257_75_43), .ZN(n_257_490));
   NOR2_X1 i_257_75_69 (.A1(n_257_75_250), .A2(n_257_75_43), .ZN(n_257_491));
   NOR2_X1 i_257_75_70 (.A1(n_257_75_252), .A2(n_257_75_43), .ZN(n_257_492));
   NAND3_X1 i_257_75_71 (.A1(PacketSize[5]), .A2(PacketSize[4]), .A3(
      n_257_75_297), .ZN(n_257_75_43));
   NOR2_X1 i_257_75_72 (.A1(n_257_75_254), .A2(n_257_75_44), .ZN(n_257_493));
   NOR2_X1 i_257_75_73 (.A1(n_257_75_258), .A2(n_257_75_44), .ZN(n_257_494));
   NOR2_X1 i_257_75_74 (.A1(n_257_75_246), .A2(n_257_75_44), .ZN(n_257_495));
   NOR2_X1 i_257_75_75 (.A1(n_257_75_247), .A2(n_257_75_44), .ZN(n_257_496));
   NOR2_X1 i_257_75_76 (.A1(n_257_75_248), .A2(n_257_75_44), .ZN(n_257_497));
   NOR2_X1 i_257_75_77 (.A1(n_257_75_249), .A2(n_257_75_44), .ZN(n_257_498));
   NOR2_X1 i_257_75_78 (.A1(n_257_75_250), .A2(n_257_75_44), .ZN(n_257_499));
   NOR2_X1 i_257_75_79 (.A1(n_257_75_252), .A2(n_257_75_44), .ZN(n_257_500));
   NAND3_X1 i_257_75_80 (.A1(PacketSize[5]), .A2(PacketSize[4]), .A3(
      PacketSize[3]), .ZN(n_257_75_44));
   NOR2_X1 i_257_75_81 (.A1(n_257_75_248), .A2(n_257_75_45), .ZN(n_257_501));
   NOR2_X1 i_257_75_82 (.A1(n_257_75_249), .A2(n_257_75_45), .ZN(n_257_502));
   NOR2_X1 i_257_75_83 (.A1(n_257_75_250), .A2(n_257_75_45), .ZN(n_257_503));
   NOR2_X1 i_257_75_84 (.A1(n_257_75_252), .A2(n_257_75_45), .ZN(n_257_504));
   NOR2_X1 i_257_75_85 (.A1(n_257_75_254), .A2(n_257_75_45), .ZN(n_257_505));
   NOR2_X1 i_257_75_86 (.A1(n_257_75_258), .A2(n_257_75_45), .ZN(n_257_506));
   NOR2_X1 i_257_75_87 (.A1(n_257_75_246), .A2(n_257_75_45), .ZN(n_257_507));
   NOR2_X1 i_257_75_88 (.A1(n_257_75_247), .A2(n_257_75_45), .ZN(n_257_508));
   NAND3_X1 i_257_75_89 (.A1(n_257_75_278), .A2(n_257_75_49), .A3(n_257_75_276), 
      .ZN(n_257_75_45));
   NOR2_X1 i_257_75_90 (.A1(n_257_75_248), .A2(n_257_75_46), .ZN(n_257_509));
   NOR2_X1 i_257_75_91 (.A1(n_257_75_249), .A2(n_257_75_46), .ZN(n_257_510));
   NOR2_X1 i_257_75_92 (.A1(n_257_75_250), .A2(n_257_75_46), .ZN(n_257_511));
   NOR2_X1 i_257_75_93 (.A1(n_257_75_252), .A2(n_257_75_46), .ZN(n_257_512));
   NOR2_X1 i_257_75_94 (.A1(n_257_75_254), .A2(n_257_75_46), .ZN(n_257_513));
   NOR2_X1 i_257_75_95 (.A1(n_257_75_258), .A2(n_257_75_46), .ZN(n_257_514));
   NOR2_X1 i_257_75_96 (.A1(n_257_75_246), .A2(n_257_75_46), .ZN(n_257_515));
   NOR2_X1 i_257_75_97 (.A1(n_257_75_247), .A2(n_257_75_46), .ZN(n_257_516));
   NAND3_X1 i_257_75_98 (.A1(n_257_75_278), .A2(n_257_75_49), .A3(n_257_75_18), 
      .ZN(n_257_75_46));
   NOR2_X1 i_257_75_99 (.A1(n_257_75_248), .A2(n_257_75_47), .ZN(n_257_517));
   NOR2_X1 i_257_75_100 (.A1(n_257_75_249), .A2(n_257_75_47), .ZN(n_257_518));
   NOR2_X1 i_257_75_101 (.A1(n_257_75_250), .A2(n_257_75_47), .ZN(n_257_519));
   NOR2_X1 i_257_75_102 (.A1(n_257_75_252), .A2(n_257_75_47), .ZN(n_257_520));
   NOR2_X1 i_257_75_103 (.A1(n_257_75_254), .A2(n_257_75_47), .ZN(n_257_521));
   NOR2_X1 i_257_75_104 (.A1(n_257_75_258), .A2(n_257_75_47), .ZN(n_257_522));
   NOR2_X1 i_257_75_105 (.A1(n_257_75_246), .A2(n_257_75_47), .ZN(n_257_523));
   NOR2_X1 i_257_75_106 (.A1(n_257_75_247), .A2(n_257_75_47), .ZN(n_257_524));
   NAND3_X1 i_257_75_107 (.A1(n_257_75_16), .A2(n_257_75_49), .A3(n_257_75_276), 
      .ZN(n_257_75_47));
   NOR2_X1 i_257_75_108 (.A1(n_257_75_248), .A2(n_257_75_48), .ZN(n_257_525));
   NOR2_X1 i_257_75_109 (.A1(n_257_75_249), .A2(n_257_75_48), .ZN(n_257_526));
   NOR2_X1 i_257_75_110 (.A1(n_257_75_250), .A2(n_257_75_48), .ZN(n_257_527));
   NOR2_X1 i_257_75_111 (.A1(n_257_75_252), .A2(n_257_75_48), .ZN(n_257_528));
   NOR2_X1 i_257_75_112 (.A1(n_257_75_254), .A2(n_257_75_48), .ZN(n_257_529));
   NOR2_X1 i_257_75_113 (.A1(n_257_75_258), .A2(n_257_75_48), .ZN(n_257_530));
   NOR2_X1 i_257_75_114 (.A1(n_257_75_246), .A2(n_257_75_48), .ZN(n_257_531));
   NOR2_X1 i_257_75_115 (.A1(n_257_75_247), .A2(n_257_75_48), .ZN(n_257_532));
   NAND3_X1 i_257_75_116 (.A1(n_257_75_16), .A2(n_257_75_49), .A3(n_257_75_18), 
      .ZN(n_257_75_48));
   XOR2_X1 i_257_75_117 (.A(PacketSize[5]), .B(n_257_75_17), .Z(n_257_75_49));
   NOR2_X1 i_257_75_118 (.A1(n_257_75_246), .A2(n_257_75_50), .ZN(n_257_533));
   NOR2_X1 i_257_75_119 (.A1(n_257_75_247), .A2(n_257_75_50), .ZN(n_257_534));
   NOR2_X1 i_257_75_120 (.A1(n_257_75_248), .A2(n_257_75_50), .ZN(n_257_535));
   NOR2_X1 i_257_75_121 (.A1(n_257_75_249), .A2(n_257_75_50), .ZN(n_257_536));
   NOR2_X1 i_257_75_122 (.A1(n_257_75_250), .A2(n_257_75_50), .ZN(n_257_537));
   NOR2_X1 i_257_75_123 (.A1(n_257_75_252), .A2(n_257_75_50), .ZN(n_257_538));
   NOR2_X1 i_257_75_124 (.A1(n_257_75_254), .A2(n_257_75_50), .ZN(n_257_539));
   NOR2_X1 i_257_75_125 (.A1(n_257_75_258), .A2(n_257_75_50), .ZN(n_257_540));
   NAND3_X1 i_257_75_126 (.A1(n_257_75_267), .A2(n_257_75_54), .A3(n_257_75_282), 
      .ZN(n_257_75_50));
   NOR2_X1 i_257_75_127 (.A1(n_257_75_246), .A2(n_257_75_51), .ZN(n_257_541));
   NOR2_X1 i_257_75_128 (.A1(n_257_75_247), .A2(n_257_75_51), .ZN(n_257_542));
   NOR2_X1 i_257_75_129 (.A1(n_257_75_248), .A2(n_257_75_51), .ZN(n_257_543));
   NOR2_X1 i_257_75_130 (.A1(n_257_75_249), .A2(n_257_75_51), .ZN(n_257_544));
   NOR2_X1 i_257_75_131 (.A1(n_257_75_250), .A2(n_257_75_51), .ZN(n_257_545));
   NOR2_X1 i_257_75_132 (.A1(n_257_75_252), .A2(n_257_75_51), .ZN(n_257_546));
   NOR2_X1 i_257_75_133 (.A1(n_257_75_254), .A2(n_257_75_51), .ZN(n_257_547));
   NOR2_X1 i_257_75_134 (.A1(n_257_75_258), .A2(n_257_75_51), .ZN(n_257_548));
   NAND3_X1 i_257_75_135 (.A1(n_257_75_267), .A2(n_257_75_54), .A3(n_257_75_12), 
      .ZN(n_257_75_51));
   NOR2_X1 i_257_75_136 (.A1(n_257_75_246), .A2(n_257_75_52), .ZN(n_257_549));
   NOR2_X1 i_257_75_137 (.A1(n_257_75_247), .A2(n_257_75_52), .ZN(n_257_550));
   NOR2_X1 i_257_75_138 (.A1(n_257_75_248), .A2(n_257_75_52), .ZN(n_257_551));
   NOR2_X1 i_257_75_139 (.A1(n_257_75_249), .A2(n_257_75_52), .ZN(n_257_552));
   NOR2_X1 i_257_75_140 (.A1(n_257_75_250), .A2(n_257_75_52), .ZN(n_257_553));
   NOR2_X1 i_257_75_141 (.A1(n_257_75_252), .A2(n_257_75_52), .ZN(n_257_554));
   NOR2_X1 i_257_75_142 (.A1(n_257_75_254), .A2(n_257_75_52), .ZN(n_257_555));
   NOR2_X1 i_257_75_143 (.A1(n_257_75_258), .A2(n_257_75_52), .ZN(n_257_556));
   NAND3_X1 i_257_75_144 (.A1(n_257_75_30), .A2(n_257_75_54), .A3(n_257_75_282), 
      .ZN(n_257_75_52));
   NOR2_X1 i_257_75_145 (.A1(n_257_75_246), .A2(n_257_75_53), .ZN(n_257_557));
   NOR2_X1 i_257_75_146 (.A1(n_257_75_247), .A2(n_257_75_53), .ZN(n_257_558));
   NOR2_X1 i_257_75_147 (.A1(n_257_75_248), .A2(n_257_75_53), .ZN(n_257_559));
   NOR2_X1 i_257_75_148 (.A1(n_257_75_249), .A2(n_257_75_53), .ZN(n_257_560));
   NOR2_X1 i_257_75_149 (.A1(n_257_75_250), .A2(n_257_75_53), .ZN(n_257_561));
   NOR2_X1 i_257_75_150 (.A1(n_257_75_252), .A2(n_257_75_53), .ZN(n_257_562));
   NOR2_X1 i_257_75_151 (.A1(n_257_75_254), .A2(n_257_75_53), .ZN(n_257_563));
   NOR2_X1 i_257_75_152 (.A1(n_257_75_258), .A2(n_257_75_53), .ZN(n_257_564));
   NAND3_X1 i_257_75_153 (.A1(n_257_75_30), .A2(n_257_75_54), .A3(n_257_75_12), 
      .ZN(n_257_75_53));
   XOR2_X1 i_257_75_154 (.A(PacketSize[5]), .B(n_257_75_31), .Z(n_257_75_54));
   NOR2_X1 i_257_75_155 (.A1(n_257_75_254), .A2(n_257_75_55), .ZN(n_257_565));
   NOR2_X1 i_257_75_156 (.A1(n_257_75_258), .A2(n_257_75_55), .ZN(n_257_566));
   NOR2_X1 i_257_75_157 (.A1(n_257_75_246), .A2(n_257_75_55), .ZN(n_257_567));
   NOR2_X1 i_257_75_158 (.A1(n_257_75_247), .A2(n_257_75_55), .ZN(n_257_568));
   NOR2_X1 i_257_75_159 (.A1(n_257_75_248), .A2(n_257_75_55), .ZN(n_257_569));
   NOR2_X1 i_257_75_160 (.A1(n_257_75_249), .A2(n_257_75_55), .ZN(n_257_570));
   NOR2_X1 i_257_75_161 (.A1(n_257_75_250), .A2(n_257_75_55), .ZN(n_257_571));
   NOR2_X1 i_257_75_162 (.A1(n_257_75_252), .A2(n_257_75_55), .ZN(n_257_572));
   OR2_X1 i_257_75_163 (.A1(n_257_75_297), .A2(n_257_75_57), .ZN(n_257_75_55));
   NOR2_X1 i_257_75_164 (.A1(n_257_75_254), .A2(n_257_75_56), .ZN(n_257_573));
   NOR2_X1 i_257_75_165 (.A1(n_257_75_258), .A2(n_257_75_56), .ZN(n_257_574));
   NOR2_X1 i_257_75_166 (.A1(n_257_75_246), .A2(n_257_75_56), .ZN(n_257_575));
   NOR2_X1 i_257_75_167 (.A1(n_257_75_247), .A2(n_257_75_56), .ZN(n_257_576));
   NOR2_X1 i_257_75_168 (.A1(n_257_75_248), .A2(n_257_75_56), .ZN(n_257_577));
   NOR2_X1 i_257_75_169 (.A1(n_257_75_249), .A2(n_257_75_56), .ZN(n_257_578));
   NOR2_X1 i_257_75_170 (.A1(n_257_75_250), .A2(n_257_75_56), .ZN(n_257_579));
   NOR2_X1 i_257_75_171 (.A1(n_257_75_252), .A2(n_257_75_56), .ZN(n_257_580));
   OR2_X1 i_257_75_172 (.A1(PacketSize[3]), .A2(n_257_75_57), .ZN(n_257_75_56));
   NAND2_X1 i_257_75_173 (.A1(n_257_75_286), .A2(n_257_75_61), .ZN(n_257_75_57));
   NOR2_X1 i_257_75_174 (.A1(n_257_75_254), .A2(n_257_75_58), .ZN(n_257_581));
   NOR2_X1 i_257_75_175 (.A1(n_257_75_258), .A2(n_257_75_58), .ZN(n_257_582));
   NOR2_X1 i_257_75_176 (.A1(n_257_75_246), .A2(n_257_75_58), .ZN(n_257_583));
   NOR2_X1 i_257_75_177 (.A1(n_257_75_247), .A2(n_257_75_58), .ZN(n_257_584));
   NOR2_X1 i_257_75_178 (.A1(n_257_75_248), .A2(n_257_75_58), .ZN(n_257_585));
   NOR2_X1 i_257_75_179 (.A1(n_257_75_249), .A2(n_257_75_58), .ZN(n_257_586));
   NOR2_X1 i_257_75_180 (.A1(n_257_75_250), .A2(n_257_75_58), .ZN(n_257_587));
   NOR2_X1 i_257_75_181 (.A1(n_257_75_252), .A2(n_257_75_58), .ZN(n_257_588));
   OR2_X1 i_257_75_182 (.A1(n_257_75_297), .A2(n_257_75_60), .ZN(n_257_75_58));
   NOR2_X1 i_257_75_183 (.A1(n_257_75_254), .A2(n_257_75_59), .ZN(n_257_589));
   NOR2_X1 i_257_75_184 (.A1(n_257_75_258), .A2(n_257_75_59), .ZN(n_257_590));
   NOR2_X1 i_257_75_185 (.A1(n_257_75_246), .A2(n_257_75_59), .ZN(n_257_591));
   NOR2_X1 i_257_75_186 (.A1(n_257_75_247), .A2(n_257_75_59), .ZN(n_257_592));
   NOR2_X1 i_257_75_187 (.A1(n_257_75_248), .A2(n_257_75_59), .ZN(n_257_593));
   NOR2_X1 i_257_75_188 (.A1(n_257_75_249), .A2(n_257_75_59), .ZN(n_257_594));
   NOR2_X1 i_257_75_189 (.A1(n_257_75_250), .A2(n_257_75_59), .ZN(n_257_595));
   NOR2_X1 i_257_75_190 (.A1(n_257_75_252), .A2(n_257_75_59), .ZN(n_257_596));
   OR2_X1 i_257_75_191 (.A1(PacketSize[3]), .A2(n_257_75_60), .ZN(n_257_75_59));
   NAND2_X1 i_257_75_192 (.A1(n_257_75_8), .A2(n_257_75_61), .ZN(n_257_75_60));
   XOR2_X1 i_257_75_193 (.A(PacketSize[5]), .B(n_257_75_9), .Z(n_257_75_61));
   NOR2_X1 i_257_75_194 (.A1(n_257_75_248), .A2(n_257_75_62), .ZN(n_257_597));
   NOR2_X1 i_257_75_195 (.A1(n_257_75_249), .A2(n_257_75_62), .ZN(n_257_598));
   NOR2_X1 i_257_75_196 (.A1(n_257_75_250), .A2(n_257_75_62), .ZN(n_257_599));
   NOR2_X1 i_257_75_197 (.A1(n_257_75_252), .A2(n_257_75_62), .ZN(n_257_600));
   NOR2_X1 i_257_75_198 (.A1(n_257_75_254), .A2(n_257_75_62), .ZN(n_257_601));
   NOR2_X1 i_257_75_199 (.A1(n_257_75_258), .A2(n_257_75_62), .ZN(n_257_602));
   NOR2_X1 i_257_75_200 (.A1(n_257_75_246), .A2(n_257_75_62), .ZN(n_257_603));
   NOR2_X1 i_257_75_201 (.A1(n_257_75_247), .A2(n_257_75_62), .ZN(n_257_604));
   NAND3_X1 i_257_75_202 (.A1(n_257_75_268), .A2(n_257_75_66), .A3(n_257_75_67), 
      .ZN(n_257_75_62));
   NOR2_X1 i_257_75_203 (.A1(n_257_75_248), .A2(n_257_75_63), .ZN(n_257_605));
   NOR2_X1 i_257_75_204 (.A1(n_257_75_249), .A2(n_257_75_63), .ZN(n_257_606));
   NOR2_X1 i_257_75_205 (.A1(n_257_75_250), .A2(n_257_75_63), .ZN(n_257_607));
   NOR2_X1 i_257_75_206 (.A1(n_257_75_252), .A2(n_257_75_63), .ZN(n_257_608));
   NOR2_X1 i_257_75_207 (.A1(n_257_75_254), .A2(n_257_75_63), .ZN(n_257_609));
   NOR2_X1 i_257_75_208 (.A1(n_257_75_258), .A2(n_257_75_63), .ZN(n_257_610));
   NOR2_X1 i_257_75_209 (.A1(n_257_75_246), .A2(n_257_75_63), .ZN(n_257_611));
   NOR2_X1 i_257_75_210 (.A1(n_257_75_247), .A2(n_257_75_63), .ZN(n_257_612));
   NAND3_X1 i_257_75_211 (.A1(n_257_75_268), .A2(n_257_75_66), .A3(n_257_75_68), 
      .ZN(n_257_75_63));
   NOR2_X1 i_257_75_212 (.A1(n_257_75_248), .A2(n_257_75_64), .ZN(n_257_613));
   NOR2_X1 i_257_75_213 (.A1(n_257_75_249), .A2(n_257_75_64), .ZN(n_257_614));
   NOR2_X1 i_257_75_214 (.A1(n_257_75_250), .A2(n_257_75_64), .ZN(n_257_615));
   NOR2_X1 i_257_75_215 (.A1(n_257_75_252), .A2(n_257_75_64), .ZN(n_257_616));
   NOR2_X1 i_257_75_216 (.A1(n_257_75_254), .A2(n_257_75_64), .ZN(n_257_617));
   NOR2_X1 i_257_75_217 (.A1(n_257_75_258), .A2(n_257_75_64), .ZN(n_257_618));
   NOR2_X1 i_257_75_218 (.A1(n_257_75_246), .A2(n_257_75_64), .ZN(n_257_619));
   NOR2_X1 i_257_75_219 (.A1(n_257_75_247), .A2(n_257_75_64), .ZN(n_257_620));
   NAND3_X1 i_257_75_220 (.A1(n_257_75_28), .A2(n_257_75_66), .A3(n_257_75_67), 
      .ZN(n_257_75_64));
   NOR2_X1 i_257_75_221 (.A1(n_257_75_248), .A2(n_257_75_65), .ZN(n_257_621));
   NOR2_X1 i_257_75_222 (.A1(n_257_75_249), .A2(n_257_75_65), .ZN(n_257_622));
   NOR2_X1 i_257_75_223 (.A1(n_257_75_250), .A2(n_257_75_65), .ZN(n_257_623));
   NOR2_X1 i_257_75_224 (.A1(n_257_75_252), .A2(n_257_75_65), .ZN(n_257_624));
   NOR2_X1 i_257_75_225 (.A1(n_257_75_254), .A2(n_257_75_65), .ZN(n_257_625));
   NOR2_X1 i_257_75_226 (.A1(n_257_75_258), .A2(n_257_75_65), .ZN(n_257_626));
   NOR2_X1 i_257_75_227 (.A1(n_257_75_246), .A2(n_257_75_65), .ZN(n_257_627));
   NOR2_X1 i_257_75_228 (.A1(n_257_75_247), .A2(n_257_75_65), .ZN(n_257_628));
   NAND3_X1 i_257_75_229 (.A1(n_257_75_28), .A2(n_257_75_66), .A3(n_257_75_68), 
      .ZN(n_257_75_65));
   XOR2_X1 i_257_75_230 (.A(PacketSize[5]), .B(n_257_75_29), .Z(n_257_75_66));
   INV_X1 i_257_75_231 (.A(n_257_75_68), .ZN(n_257_75_67));
   OAI21_X1 i_257_75_232 (.A(n_257_75_265), .B1(n_257_75_297), .B2(n_257_75_296), 
      .ZN(n_257_75_68));
   NOR2_X1 i_257_75_233 (.A1(n_257_75_140), .A2(n_257_75_69), .ZN(n_257_629));
   NOR2_X1 i_257_75_234 (.A1(n_257_75_141), .A2(n_257_75_69), .ZN(n_257_630));
   NOR2_X1 i_257_75_235 (.A1(n_257_75_142), .A2(n_257_75_69), .ZN(n_257_631));
   NOR2_X1 i_257_75_236 (.A1(n_257_75_143), .A2(n_257_75_69), .ZN(n_257_632));
   NOR2_X1 i_257_75_237 (.A1(n_257_75_144), .A2(n_257_75_69), .ZN(n_257_633));
   NOR2_X1 i_257_75_238 (.A1(n_257_75_145), .A2(n_257_75_69), .ZN(n_257_634));
   NOR2_X1 i_257_75_239 (.A1(n_257_75_146), .A2(n_257_75_69), .ZN(n_257_635));
   NOR2_X1 i_257_75_240 (.A1(n_257_75_151), .A2(n_257_75_69), .ZN(n_257_636));
   NAND3_X1 i_257_75_241 (.A1(n_257_75_269), .A2(n_257_75_73), .A3(n_257_75_74), 
      .ZN(n_257_75_69));
   NOR2_X1 i_257_75_242 (.A1(n_257_75_140), .A2(n_257_75_70), .ZN(n_257_637));
   NOR2_X1 i_257_75_243 (.A1(n_257_75_141), .A2(n_257_75_70), .ZN(n_257_638));
   NOR2_X1 i_257_75_244 (.A1(n_257_75_142), .A2(n_257_75_70), .ZN(n_257_639));
   NOR2_X1 i_257_75_245 (.A1(n_257_75_143), .A2(n_257_75_70), .ZN(n_257_640));
   NOR2_X1 i_257_75_246 (.A1(n_257_75_144), .A2(n_257_75_70), .ZN(n_257_641));
   NOR2_X1 i_257_75_247 (.A1(n_257_75_145), .A2(n_257_75_70), .ZN(n_257_642));
   NOR2_X1 i_257_75_248 (.A1(n_257_75_146), .A2(n_257_75_70), .ZN(n_257_643));
   NOR2_X1 i_257_75_249 (.A1(n_257_75_151), .A2(n_257_75_70), .ZN(n_257_644));
   NAND3_X1 i_257_75_250 (.A1(n_257_75_269), .A2(n_257_75_73), .A3(n_257_75_75), 
      .ZN(n_257_75_70));
   NOR2_X1 i_257_75_251 (.A1(n_257_75_140), .A2(n_257_75_71), .ZN(n_257_645));
   NOR2_X1 i_257_75_252 (.A1(n_257_75_141), .A2(n_257_75_71), .ZN(n_257_646));
   NOR2_X1 i_257_75_253 (.A1(n_257_75_142), .A2(n_257_75_71), .ZN(n_257_647));
   NOR2_X1 i_257_75_254 (.A1(n_257_75_143), .A2(n_257_75_71), .ZN(n_257_648));
   NOR2_X1 i_257_75_255 (.A1(n_257_75_144), .A2(n_257_75_71), .ZN(n_257_649));
   NOR2_X1 i_257_75_256 (.A1(n_257_75_145), .A2(n_257_75_71), .ZN(n_257_650));
   NOR2_X1 i_257_75_257 (.A1(n_257_75_146), .A2(n_257_75_71), .ZN(n_257_651));
   NOR2_X1 i_257_75_258 (.A1(n_257_75_151), .A2(n_257_75_71), .ZN(n_257_652));
   NAND3_X1 i_257_75_259 (.A1(n_257_75_26), .A2(n_257_75_73), .A3(n_257_75_74), 
      .ZN(n_257_75_71));
   NOR2_X1 i_257_75_260 (.A1(n_257_75_140), .A2(n_257_75_72), .ZN(n_257_653));
   NOR2_X1 i_257_75_261 (.A1(n_257_75_141), .A2(n_257_75_72), .ZN(n_257_654));
   NOR2_X1 i_257_75_262 (.A1(n_257_75_142), .A2(n_257_75_72), .ZN(n_257_655));
   NOR2_X1 i_257_75_263 (.A1(n_257_75_143), .A2(n_257_75_72), .ZN(n_257_656));
   NOR2_X1 i_257_75_264 (.A1(n_257_75_144), .A2(n_257_75_72), .ZN(n_257_657));
   NOR2_X1 i_257_75_265 (.A1(n_257_75_145), .A2(n_257_75_72), .ZN(n_257_658));
   NOR2_X1 i_257_75_266 (.A1(n_257_75_146), .A2(n_257_75_72), .ZN(n_257_659));
   NOR2_X1 i_257_75_267 (.A1(n_257_75_151), .A2(n_257_75_72), .ZN(n_257_660));
   NAND3_X1 i_257_75_268 (.A1(n_257_75_26), .A2(n_257_75_73), .A3(n_257_75_75), 
      .ZN(n_257_75_72));
   XOR2_X1 i_257_75_269 (.A(PacketSize[5]), .B(n_257_75_27), .Z(n_257_75_73));
   INV_X1 i_257_75_270 (.A(n_257_75_75), .ZN(n_257_75_74));
   OAI21_X1 i_257_75_271 (.A(n_257_75_76), .B1(n_257_75_297), .B2(n_257_75_255), 
      .ZN(n_257_75_75));
   NAND2_X1 i_257_75_272 (.A1(n_257_75_297), .A2(n_257_75_255), .ZN(n_257_75_76));
   NOR2_X1 i_257_75_273 (.A1(n_257_75_254), .A2(n_257_75_77), .ZN(n_257_661));
   NOR2_X1 i_257_75_274 (.A1(n_257_75_258), .A2(n_257_75_77), .ZN(n_257_662));
   NOR2_X1 i_257_75_275 (.A1(n_257_75_246), .A2(n_257_75_77), .ZN(n_257_663));
   NOR2_X1 i_257_75_276 (.A1(n_257_75_247), .A2(n_257_75_77), .ZN(n_257_664));
   NOR2_X1 i_257_75_277 (.A1(n_257_75_248), .A2(n_257_75_77), .ZN(n_257_665));
   NOR2_X1 i_257_75_278 (.A1(n_257_75_249), .A2(n_257_75_77), .ZN(n_257_666));
   NOR2_X1 i_257_75_279 (.A1(n_257_75_250), .A2(n_257_75_77), .ZN(n_257_667));
   NOR2_X1 i_257_75_280 (.A1(n_257_75_252), .A2(n_257_75_77), .ZN(n_257_668));
   NAND3_X1 i_257_75_281 (.A1(PacketSize[5]), .A2(n_257_75_322), .A3(
      PacketSize[3]), .ZN(n_257_75_77));
   NOR2_X1 i_257_75_282 (.A1(n_257_75_157), .A2(n_257_75_78), .ZN(n_257_669));
   NOR2_X1 i_257_75_283 (.A1(n_257_75_158), .A2(n_257_75_78), .ZN(n_257_670));
   NOR2_X1 i_257_75_284 (.A1(n_257_75_159), .A2(n_257_75_78), .ZN(n_257_671));
   NOR2_X1 i_257_75_285 (.A1(n_257_75_160), .A2(n_257_75_78), .ZN(n_257_672));
   NOR2_X1 i_257_75_286 (.A1(n_257_75_161), .A2(n_257_75_78), .ZN(n_257_673));
   NOR2_X1 i_257_75_287 (.A1(n_257_75_162), .A2(n_257_75_78), .ZN(n_257_674));
   NOR2_X1 i_257_75_288 (.A1(n_257_75_163), .A2(n_257_75_78), .ZN(n_257_675));
   NOR2_X1 i_257_75_289 (.A1(n_257_75_172), .A2(n_257_75_78), .ZN(n_257_676));
   OR2_X1 i_257_75_290 (.A1(n_257_75_24), .A2(n_257_75_80), .ZN(n_257_75_78));
   NOR2_X1 i_257_75_291 (.A1(n_257_75_157), .A2(n_257_75_79), .ZN(n_257_677));
   NOR2_X1 i_257_75_292 (.A1(n_257_75_158), .A2(n_257_75_79), .ZN(n_257_678));
   NOR2_X1 i_257_75_293 (.A1(n_257_75_159), .A2(n_257_75_79), .ZN(n_257_679));
   NOR2_X1 i_257_75_294 (.A1(n_257_75_160), .A2(n_257_75_79), .ZN(n_257_680));
   NOR2_X1 i_257_75_295 (.A1(n_257_75_161), .A2(n_257_75_79), .ZN(n_257_681));
   NOR2_X1 i_257_75_296 (.A1(n_257_75_162), .A2(n_257_75_79), .ZN(n_257_682));
   NOR2_X1 i_257_75_297 (.A1(n_257_75_163), .A2(n_257_75_79), .ZN(n_257_683));
   NOR2_X1 i_257_75_298 (.A1(n_257_75_172), .A2(n_257_75_79), .ZN(n_257_684));
   OR2_X1 i_257_75_299 (.A1(n_257_75_270), .A2(n_257_75_80), .ZN(n_257_75_79));
   OR2_X1 i_257_75_300 (.A1(n_257_75_85), .A2(n_257_75_84), .ZN(n_257_75_80));
   NOR2_X1 i_257_75_301 (.A1(n_257_75_157), .A2(n_257_75_81), .ZN(n_257_685));
   NOR2_X1 i_257_75_302 (.A1(n_257_75_158), .A2(n_257_75_81), .ZN(n_257_686));
   NOR2_X1 i_257_75_303 (.A1(n_257_75_159), .A2(n_257_75_81), .ZN(n_257_687));
   NOR2_X1 i_257_75_304 (.A1(n_257_75_160), .A2(n_257_75_81), .ZN(n_257_688));
   NOR2_X1 i_257_75_305 (.A1(n_257_75_161), .A2(n_257_75_81), .ZN(n_257_689));
   NOR2_X1 i_257_75_306 (.A1(n_257_75_162), .A2(n_257_75_81), .ZN(n_257_690));
   NOR2_X1 i_257_75_307 (.A1(n_257_75_163), .A2(n_257_75_81), .ZN(n_257_691));
   NOR2_X1 i_257_75_308 (.A1(n_257_75_172), .A2(n_257_75_81), .ZN(n_257_692));
   OR2_X1 i_257_75_309 (.A1(n_257_75_24), .A2(n_257_75_83), .ZN(n_257_75_81));
   NOR2_X1 i_257_75_310 (.A1(n_257_75_82), .A2(n_257_75_157), .ZN(n_257_693));
   NOR2_X1 i_257_75_311 (.A1(n_257_75_82), .A2(n_257_75_158), .ZN(n_257_694));
   NOR2_X1 i_257_75_312 (.A1(n_257_75_82), .A2(n_257_75_159), .ZN(n_257_695));
   NOR2_X1 i_257_75_313 (.A1(n_257_75_82), .A2(n_257_75_160), .ZN(n_257_696));
   NOR2_X1 i_257_75_314 (.A1(n_257_75_82), .A2(n_257_75_161), .ZN(n_257_697));
   NOR2_X1 i_257_75_315 (.A1(n_257_75_82), .A2(n_257_75_162), .ZN(n_257_698));
   NOR2_X1 i_257_75_316 (.A1(n_257_75_82), .A2(n_257_75_163), .ZN(n_257_699));
   NOR2_X1 i_257_75_317 (.A1(n_257_75_172), .A2(n_257_75_82), .ZN(n_257_700));
   OR2_X1 i_257_75_318 (.A1(n_257_75_270), .A2(n_257_75_83), .ZN(n_257_75_82));
   OAI21_X1 i_257_75_319 (.A(n_257_75_84), .B1(n_257_75_298), .B2(n_257_75_85), 
      .ZN(n_257_75_83));
   OAI21_X1 i_257_75_320 (.A(n_257_75_298), .B1(n_257_75_322), .B2(n_257_75_271), 
      .ZN(n_257_75_84));
   NOR2_X1 i_257_75_321 (.A1(PacketSize[4]), .A2(n_257_75_25), .ZN(n_257_75_85));
   NOR2_X1 i_257_75_322 (.A1(n_257_75_176), .A2(n_257_75_86), .ZN(n_257_701));
   NOR2_X1 i_257_75_323 (.A1(n_257_75_177), .A2(n_257_75_86), .ZN(n_257_702));
   NOR2_X1 i_257_75_324 (.A1(n_257_75_178), .A2(n_257_75_86), .ZN(n_257_703));
   NOR2_X1 i_257_75_325 (.A1(n_257_75_179), .A2(n_257_75_86), .ZN(n_257_704));
   NOR2_X1 i_257_75_326 (.A1(n_257_75_180), .A2(n_257_75_86), .ZN(n_257_705));
   NOR2_X1 i_257_75_327 (.A1(n_257_75_181), .A2(n_257_75_86), .ZN(n_257_706));
   NOR2_X1 i_257_75_328 (.A1(n_257_75_182), .A2(n_257_75_86), .ZN(n_257_707));
   NOR2_X1 i_257_75_329 (.A1(n_257_75_191), .A2(n_257_75_86), .ZN(n_257_708));
   OR2_X1 i_257_75_330 (.A1(n_257_75_22), .A2(n_257_75_88), .ZN(n_257_75_86));
   NOR2_X1 i_257_75_331 (.A1(n_257_75_176), .A2(n_257_75_87), .ZN(n_257_709));
   NOR2_X1 i_257_75_332 (.A1(n_257_75_177), .A2(n_257_75_87), .ZN(n_257_710));
   NOR2_X1 i_257_75_333 (.A1(n_257_75_178), .A2(n_257_75_87), .ZN(n_257_711));
   NOR2_X1 i_257_75_334 (.A1(n_257_75_179), .A2(n_257_75_87), .ZN(n_257_712));
   NOR2_X1 i_257_75_335 (.A1(n_257_75_180), .A2(n_257_75_87), .ZN(n_257_713));
   NOR2_X1 i_257_75_336 (.A1(n_257_75_181), .A2(n_257_75_87), .ZN(n_257_714));
   NOR2_X1 i_257_75_337 (.A1(n_257_75_182), .A2(n_257_75_87), .ZN(n_257_715));
   NOR2_X1 i_257_75_338 (.A1(n_257_75_191), .A2(n_257_75_87), .ZN(n_257_716));
   OR2_X1 i_257_75_339 (.A1(n_257_75_272), .A2(n_257_75_88), .ZN(n_257_75_87));
   OR2_X1 i_257_75_340 (.A1(n_257_75_93), .A2(n_257_75_92), .ZN(n_257_75_88));
   NOR2_X1 i_257_75_341 (.A1(n_257_75_176), .A2(n_257_75_89), .ZN(n_257_717));
   NOR2_X1 i_257_75_342 (.A1(n_257_75_177), .A2(n_257_75_89), .ZN(n_257_718));
   NOR2_X1 i_257_75_343 (.A1(n_257_75_178), .A2(n_257_75_89), .ZN(n_257_719));
   NOR2_X1 i_257_75_344 (.A1(n_257_75_179), .A2(n_257_75_89), .ZN(n_257_720));
   NOR2_X1 i_257_75_345 (.A1(n_257_75_180), .A2(n_257_75_89), .ZN(n_257_721));
   NOR2_X1 i_257_75_346 (.A1(n_257_75_181), .A2(n_257_75_89), .ZN(n_257_722));
   NOR2_X1 i_257_75_347 (.A1(n_257_75_182), .A2(n_257_75_89), .ZN(n_257_723));
   NOR2_X1 i_257_75_348 (.A1(n_257_75_191), .A2(n_257_75_89), .ZN(n_257_724));
   OR2_X1 i_257_75_349 (.A1(n_257_75_22), .A2(n_257_75_91), .ZN(n_257_75_89));
   NOR2_X1 i_257_75_350 (.A1(n_257_75_90), .A2(n_257_75_176), .ZN(n_257_725));
   NOR2_X1 i_257_75_351 (.A1(n_257_75_90), .A2(n_257_75_177), .ZN(n_257_726));
   NOR2_X1 i_257_75_352 (.A1(n_257_75_90), .A2(n_257_75_178), .ZN(n_257_727));
   NOR2_X1 i_257_75_353 (.A1(n_257_75_90), .A2(n_257_75_179), .ZN(n_257_728));
   NOR2_X1 i_257_75_354 (.A1(n_257_75_90), .A2(n_257_75_180), .ZN(n_257_729));
   NOR2_X1 i_257_75_355 (.A1(n_257_75_90), .A2(n_257_75_181), .ZN(n_257_730));
   NOR2_X1 i_257_75_356 (.A1(n_257_75_90), .A2(n_257_75_182), .ZN(n_257_731));
   NOR2_X1 i_257_75_357 (.A1(n_257_75_191), .A2(n_257_75_90), .ZN(n_257_732));
   OR2_X1 i_257_75_358 (.A1(n_257_75_272), .A2(n_257_75_91), .ZN(n_257_75_90));
   OAI21_X1 i_257_75_359 (.A(n_257_75_92), .B1(n_257_75_298), .B2(n_257_75_93), 
      .ZN(n_257_75_91));
   OAI21_X1 i_257_75_360 (.A(n_257_75_298), .B1(n_257_75_322), .B2(n_257_75_273), 
      .ZN(n_257_75_92));
   NOR2_X1 i_257_75_361 (.A1(PacketSize[4]), .A2(n_257_75_23), .ZN(n_257_75_93));
   NOR2_X1 i_257_75_362 (.A1(n_257_75_195), .A2(n_257_75_94), .ZN(n_257_733));
   NOR2_X1 i_257_75_363 (.A1(n_257_75_196), .A2(n_257_75_94), .ZN(n_257_734));
   NOR2_X1 i_257_75_364 (.A1(n_257_75_197), .A2(n_257_75_94), .ZN(n_257_735));
   NOR2_X1 i_257_75_365 (.A1(n_257_75_198), .A2(n_257_75_94), .ZN(n_257_736));
   NOR2_X1 i_257_75_366 (.A1(n_257_75_199), .A2(n_257_75_94), .ZN(n_257_737));
   NOR2_X1 i_257_75_367 (.A1(n_257_75_201), .A2(n_257_75_94), .ZN(n_257_738));
   NOR2_X1 i_257_75_368 (.A1(n_257_75_203), .A2(n_257_75_94), .ZN(n_257_739));
   NOR2_X1 i_257_75_369 (.A1(n_257_75_213), .A2(n_257_75_94), .ZN(n_257_740));
   OR2_X1 i_257_75_370 (.A1(n_257_75_20), .A2(n_257_75_96), .ZN(n_257_75_94));
   NOR2_X1 i_257_75_371 (.A1(n_257_75_195), .A2(n_257_75_95), .ZN(n_257_741));
   NOR2_X1 i_257_75_372 (.A1(n_257_75_196), .A2(n_257_75_95), .ZN(n_257_742));
   NOR2_X1 i_257_75_373 (.A1(n_257_75_197), .A2(n_257_75_95), .ZN(n_257_743));
   NOR2_X1 i_257_75_374 (.A1(n_257_75_198), .A2(n_257_75_95), .ZN(n_257_744));
   NOR2_X1 i_257_75_375 (.A1(n_257_75_199), .A2(n_257_75_95), .ZN(n_257_745));
   NOR2_X1 i_257_75_376 (.A1(n_257_75_201), .A2(n_257_75_95), .ZN(n_257_746));
   NOR2_X1 i_257_75_377 (.A1(n_257_75_203), .A2(n_257_75_95), .ZN(n_257_747));
   NOR2_X1 i_257_75_378 (.A1(n_257_75_213), .A2(n_257_75_95), .ZN(n_257_748));
   OR2_X1 i_257_75_379 (.A1(n_257_75_274), .A2(n_257_75_96), .ZN(n_257_75_95));
   OR2_X1 i_257_75_380 (.A1(n_257_75_101), .A2(n_257_75_100), .ZN(n_257_75_96));
   NOR2_X1 i_257_75_381 (.A1(n_257_75_195), .A2(n_257_75_97), .ZN(n_257_749));
   NOR2_X1 i_257_75_382 (.A1(n_257_75_196), .A2(n_257_75_97), .ZN(n_257_750));
   NOR2_X1 i_257_75_383 (.A1(n_257_75_197), .A2(n_257_75_97), .ZN(n_257_751));
   NOR2_X1 i_257_75_384 (.A1(n_257_75_198), .A2(n_257_75_97), .ZN(n_257_752));
   NOR2_X1 i_257_75_385 (.A1(n_257_75_199), .A2(n_257_75_97), .ZN(n_257_753));
   NOR2_X1 i_257_75_386 (.A1(n_257_75_201), .A2(n_257_75_97), .ZN(n_257_754));
   NOR2_X1 i_257_75_387 (.A1(n_257_75_203), .A2(n_257_75_97), .ZN(n_257_755));
   NOR2_X1 i_257_75_388 (.A1(n_257_75_213), .A2(n_257_75_97), .ZN(n_257_756));
   OR2_X1 i_257_75_389 (.A1(n_257_75_20), .A2(n_257_75_99), .ZN(n_257_75_97));
   NOR2_X1 i_257_75_390 (.A1(n_257_75_98), .A2(n_257_75_195), .ZN(n_257_757));
   NOR2_X1 i_257_75_391 (.A1(n_257_75_98), .A2(n_257_75_196), .ZN(n_257_758));
   NOR2_X1 i_257_75_392 (.A1(n_257_75_98), .A2(n_257_75_197), .ZN(n_257_759));
   NOR2_X1 i_257_75_393 (.A1(n_257_75_98), .A2(n_257_75_198), .ZN(n_257_760));
   NOR2_X1 i_257_75_394 (.A1(n_257_75_98), .A2(n_257_75_199), .ZN(n_257_761));
   NOR2_X1 i_257_75_395 (.A1(n_257_75_98), .A2(n_257_75_201), .ZN(n_257_762));
   NOR2_X1 i_257_75_396 (.A1(n_257_75_98), .A2(n_257_75_203), .ZN(n_257_763));
   NOR2_X1 i_257_75_397 (.A1(n_257_75_213), .A2(n_257_75_98), .ZN(n_257_764));
   OR2_X1 i_257_75_398 (.A1(n_257_75_274), .A2(n_257_75_99), .ZN(n_257_75_98));
   OAI21_X1 i_257_75_399 (.A(n_257_75_100), .B1(n_257_75_298), .B2(n_257_75_101), 
      .ZN(n_257_75_99));
   OAI21_X1 i_257_75_400 (.A(n_257_75_298), .B1(n_257_75_322), .B2(n_257_75_275), 
      .ZN(n_257_75_100));
   NOR2_X1 i_257_75_401 (.A1(PacketSize[4]), .A2(n_257_75_21), .ZN(n_257_75_101));
   NOR2_X1 i_257_75_402 (.A1(n_257_75_248), .A2(n_257_75_102), .ZN(n_257_765));
   NOR2_X1 i_257_75_403 (.A1(n_257_75_249), .A2(n_257_75_102), .ZN(n_257_766));
   NOR2_X1 i_257_75_404 (.A1(n_257_75_250), .A2(n_257_75_102), .ZN(n_257_767));
   NOR2_X1 i_257_75_405 (.A1(n_257_75_252), .A2(n_257_75_102), .ZN(n_257_768));
   NOR2_X1 i_257_75_406 (.A1(n_257_75_254), .A2(n_257_75_102), .ZN(n_257_769));
   NOR2_X1 i_257_75_407 (.A1(n_257_75_258), .A2(n_257_75_102), .ZN(n_257_770));
   NOR2_X1 i_257_75_408 (.A1(n_257_75_246), .A2(n_257_75_102), .ZN(n_257_771));
   NOR2_X1 i_257_75_409 (.A1(n_257_75_247), .A2(n_257_75_102), .ZN(n_257_772));
   OR2_X1 i_257_75_410 (.A1(n_257_75_18), .A2(n_257_75_104), .ZN(n_257_75_102));
   NOR2_X1 i_257_75_411 (.A1(n_257_75_248), .A2(n_257_75_103), .ZN(n_257_773));
   NOR2_X1 i_257_75_412 (.A1(n_257_75_249), .A2(n_257_75_103), .ZN(n_257_774));
   NOR2_X1 i_257_75_413 (.A1(n_257_75_250), .A2(n_257_75_103), .ZN(n_257_775));
   NOR2_X1 i_257_75_414 (.A1(n_257_75_252), .A2(n_257_75_103), .ZN(n_257_776));
   NOR2_X1 i_257_75_415 (.A1(n_257_75_254), .A2(n_257_75_103), .ZN(n_257_777));
   NOR2_X1 i_257_75_416 (.A1(n_257_75_258), .A2(n_257_75_103), .ZN(n_257_778));
   NOR2_X1 i_257_75_417 (.A1(n_257_75_246), .A2(n_257_75_103), .ZN(n_257_779));
   NOR2_X1 i_257_75_418 (.A1(n_257_75_247), .A2(n_257_75_103), .ZN(n_257_780));
   OR2_X1 i_257_75_419 (.A1(n_257_75_276), .A2(n_257_75_104), .ZN(n_257_75_103));
   OR2_X1 i_257_75_420 (.A1(n_257_75_109), .A2(n_257_75_108), .ZN(n_257_75_104));
   NOR2_X1 i_257_75_421 (.A1(n_257_75_248), .A2(n_257_75_105), .ZN(n_257_781));
   NOR2_X1 i_257_75_422 (.A1(n_257_75_249), .A2(n_257_75_105), .ZN(n_257_782));
   NOR2_X1 i_257_75_423 (.A1(n_257_75_250), .A2(n_257_75_105), .ZN(n_257_783));
   NOR2_X1 i_257_75_424 (.A1(n_257_75_252), .A2(n_257_75_105), .ZN(n_257_784));
   NOR2_X1 i_257_75_425 (.A1(n_257_75_254), .A2(n_257_75_105), .ZN(n_257_785));
   NOR2_X1 i_257_75_426 (.A1(n_257_75_258), .A2(n_257_75_105), .ZN(n_257_786));
   NOR2_X1 i_257_75_427 (.A1(n_257_75_246), .A2(n_257_75_105), .ZN(n_257_787));
   NOR2_X1 i_257_75_428 (.A1(n_257_75_247), .A2(n_257_75_105), .ZN(n_257_788));
   OR2_X1 i_257_75_429 (.A1(n_257_75_18), .A2(n_257_75_107), .ZN(n_257_75_105));
   NOR2_X1 i_257_75_430 (.A1(n_257_75_248), .A2(n_257_75_106), .ZN(n_257_789));
   NOR2_X1 i_257_75_431 (.A1(n_257_75_249), .A2(n_257_75_106), .ZN(n_257_790));
   NOR2_X1 i_257_75_432 (.A1(n_257_75_250), .A2(n_257_75_106), .ZN(n_257_791));
   NOR2_X1 i_257_75_433 (.A1(n_257_75_252), .A2(n_257_75_106), .ZN(n_257_792));
   NOR2_X1 i_257_75_434 (.A1(n_257_75_254), .A2(n_257_75_106), .ZN(n_257_793));
   NOR2_X1 i_257_75_435 (.A1(n_257_75_258), .A2(n_257_75_106), .ZN(n_257_794));
   NOR2_X1 i_257_75_436 (.A1(n_257_75_246), .A2(n_257_75_106), .ZN(n_257_795));
   NOR2_X1 i_257_75_437 (.A1(n_257_75_247), .A2(n_257_75_106), .ZN(n_257_796));
   OR2_X1 i_257_75_438 (.A1(n_257_75_276), .A2(n_257_75_107), .ZN(n_257_75_106));
   OAI21_X1 i_257_75_439 (.A(n_257_75_108), .B1(n_257_75_298), .B2(n_257_75_109), 
      .ZN(n_257_75_107));
   OAI21_X1 i_257_75_440 (.A(n_257_75_298), .B1(n_257_75_322), .B2(n_257_75_277), 
      .ZN(n_257_75_108));
   NOR2_X1 i_257_75_441 (.A1(PacketSize[4]), .A2(n_257_75_19), .ZN(n_257_75_109));
   NOR2_X1 i_257_75_442 (.A1(n_257_75_114), .A2(n_257_75_110), .ZN(n_257_797));
   NOR2_X1 i_257_75_443 (.A1(n_257_75_115), .A2(n_257_75_110), .ZN(n_257_798));
   NOR2_X1 i_257_75_444 (.A1(n_257_75_116), .A2(n_257_75_110), .ZN(n_257_799));
   NOR2_X1 i_257_75_445 (.A1(n_257_75_117), .A2(n_257_75_110), .ZN(n_257_800));
   NOR2_X1 i_257_75_446 (.A1(n_257_75_118), .A2(n_257_75_110), .ZN(n_257_801));
   NOR2_X1 i_257_75_447 (.A1(n_257_75_119), .A2(n_257_75_110), .ZN(n_257_802));
   NOR2_X1 i_257_75_448 (.A1(n_257_75_120), .A2(n_257_75_110), .ZN(n_257_803));
   NOR2_X1 i_257_75_449 (.A1(n_257_75_125), .A2(n_257_75_110), .ZN(n_257_804));
   OR2_X1 i_257_75_450 (.A1(n_257_75_14), .A2(n_257_75_112), .ZN(n_257_75_110));
   NOR2_X1 i_257_75_451 (.A1(n_257_75_114), .A2(n_257_75_111), .ZN(n_257_805));
   NOR2_X1 i_257_75_452 (.A1(n_257_75_115), .A2(n_257_75_111), .ZN(n_257_806));
   NOR2_X1 i_257_75_453 (.A1(n_257_75_116), .A2(n_257_75_111), .ZN(n_257_807));
   NOR2_X1 i_257_75_454 (.A1(n_257_75_117), .A2(n_257_75_111), .ZN(n_257_808));
   NOR2_X1 i_257_75_455 (.A1(n_257_75_118), .A2(n_257_75_111), .ZN(n_257_809));
   NOR2_X1 i_257_75_456 (.A1(n_257_75_119), .A2(n_257_75_111), .ZN(n_257_810));
   NOR2_X1 i_257_75_457 (.A1(n_257_75_120), .A2(n_257_75_111), .ZN(n_257_811));
   NOR2_X1 i_257_75_458 (.A1(n_257_75_125), .A2(n_257_75_111), .ZN(n_257_812));
   OR2_X1 i_257_75_459 (.A1(n_257_75_279), .A2(n_257_75_112), .ZN(n_257_75_111));
   OR2_X1 i_257_75_460 (.A1(n_257_75_124), .A2(n_257_75_123), .ZN(n_257_75_112));
   NOR2_X1 i_257_75_461 (.A1(n_257_75_114), .A2(n_257_75_113), .ZN(n_257_813));
   NOR2_X1 i_257_75_462 (.A1(n_257_75_115), .A2(n_257_75_113), .ZN(n_257_814));
   NOR2_X1 i_257_75_463 (.A1(n_257_75_116), .A2(n_257_75_113), .ZN(n_257_815));
   NOR2_X1 i_257_75_464 (.A1(n_257_75_117), .A2(n_257_75_113), .ZN(n_257_816));
   NOR2_X1 i_257_75_465 (.A1(n_257_75_118), .A2(n_257_75_113), .ZN(n_257_817));
   NOR2_X1 i_257_75_466 (.A1(n_257_75_119), .A2(n_257_75_113), .ZN(n_257_818));
   NOR2_X1 i_257_75_467 (.A1(n_257_75_120), .A2(n_257_75_113), .ZN(n_257_819));
   NOR2_X1 i_257_75_468 (.A1(n_257_75_125), .A2(n_257_75_113), .ZN(n_257_820));
   OR2_X1 i_257_75_469 (.A1(n_257_75_14), .A2(n_257_75_122), .ZN(n_257_75_113));
   NOR2_X1 i_257_75_470 (.A1(n_257_75_121), .A2(n_257_75_114), .ZN(n_257_821));
   OR3_X1 i_257_75_471 (.A1(n_151), .A2(n_257_75_4), .A3(n_257_75_126), .ZN(
      n_257_75_114));
   NOR2_X1 i_257_75_472 (.A1(n_257_75_121), .A2(n_257_75_115), .ZN(n_257_822));
   OR3_X1 i_257_75_473 (.A1(n_257_75_294), .A2(n_257_75_4), .A3(n_257_75_126), 
      .ZN(n_257_75_115));
   NOR2_X1 i_257_75_474 (.A1(n_257_75_121), .A2(n_257_75_116), .ZN(n_257_823));
   OR3_X1 i_257_75_475 (.A1(n_151), .A2(n_257_75_287), .A3(n_257_75_126), 
      .ZN(n_257_75_116));
   NOR2_X1 i_257_75_476 (.A1(n_257_75_121), .A2(n_257_75_117), .ZN(n_257_824));
   OR3_X1 i_257_75_477 (.A1(n_257_75_294), .A2(n_257_75_287), .A3(n_257_75_126), 
      .ZN(n_257_75_117));
   NOR2_X1 i_257_75_478 (.A1(n_257_75_121), .A2(n_257_75_118), .ZN(n_257_825));
   NAND3_X1 i_257_75_479 (.A1(n_257_75_294), .A2(n_257_75_287), .A3(n_257_75_126), 
      .ZN(n_257_75_118));
   NOR2_X1 i_257_75_480 (.A1(n_257_75_121), .A2(n_257_75_119), .ZN(n_257_826));
   NAND3_X1 i_257_75_481 (.A1(n_151), .A2(n_257_75_287), .A3(n_257_75_126), 
      .ZN(n_257_75_119));
   NOR2_X1 i_257_75_482 (.A1(n_257_75_121), .A2(n_257_75_120), .ZN(n_257_827));
   NAND3_X1 i_257_75_483 (.A1(n_257_75_294), .A2(n_257_75_4), .A3(n_257_75_126), 
      .ZN(n_257_75_120));
   NOR2_X1 i_257_75_484 (.A1(n_257_75_125), .A2(n_257_75_121), .ZN(n_257_828));
   OR2_X1 i_257_75_485 (.A1(n_257_75_279), .A2(n_257_75_122), .ZN(n_257_75_121));
   OAI21_X1 i_257_75_486 (.A(n_257_75_123), .B1(n_257_75_298), .B2(n_257_75_124), 
      .ZN(n_257_75_122));
   OAI21_X1 i_257_75_487 (.A(n_257_75_298), .B1(n_257_75_322), .B2(n_257_75_280), 
      .ZN(n_257_75_123));
   NOR2_X1 i_257_75_488 (.A1(PacketSize[4]), .A2(n_257_75_15), .ZN(n_257_75_124));
   NAND3_X1 i_257_75_489 (.A1(n_151), .A2(n_257_75_4), .A3(n_257_75_126), 
      .ZN(n_257_75_125));
   OAI21_X1 i_257_75_490 (.A(n_257_75_127), .B1(n_257_75_296), .B2(n_257_75_281), 
      .ZN(n_257_75_126));
   NAND2_X1 i_257_75_491 (.A1(n_257_75_296), .A2(n_257_75_281), .ZN(n_257_75_127));
   NOR2_X1 i_257_75_492 (.A1(n_257_75_246), .A2(n_257_75_128), .ZN(n_257_829));
   NOR2_X1 i_257_75_493 (.A1(n_257_75_247), .A2(n_257_75_128), .ZN(n_257_830));
   NOR2_X1 i_257_75_494 (.A1(n_257_75_248), .A2(n_257_75_128), .ZN(n_257_831));
   NOR2_X1 i_257_75_495 (.A1(n_257_75_249), .A2(n_257_75_128), .ZN(n_257_832));
   NOR2_X1 i_257_75_496 (.A1(n_257_75_250), .A2(n_257_75_128), .ZN(n_257_833));
   NOR2_X1 i_257_75_497 (.A1(n_257_75_252), .A2(n_257_75_128), .ZN(n_257_834));
   NOR2_X1 i_257_75_498 (.A1(n_257_75_254), .A2(n_257_75_128), .ZN(n_257_835));
   NOR2_X1 i_257_75_499 (.A1(n_257_75_258), .A2(n_257_75_128), .ZN(n_257_836));
   OR2_X1 i_257_75_500 (.A1(n_257_75_12), .A2(n_257_75_130), .ZN(n_257_75_128));
   NOR2_X1 i_257_75_501 (.A1(n_257_75_246), .A2(n_257_75_129), .ZN(n_257_837));
   NOR2_X1 i_257_75_502 (.A1(n_257_75_247), .A2(n_257_75_129), .ZN(n_257_838));
   NOR2_X1 i_257_75_503 (.A1(n_257_75_248), .A2(n_257_75_129), .ZN(n_257_839));
   NOR2_X1 i_257_75_504 (.A1(n_257_75_249), .A2(n_257_75_129), .ZN(n_257_840));
   NOR2_X1 i_257_75_505 (.A1(n_257_75_250), .A2(n_257_75_129), .ZN(n_257_841));
   NOR2_X1 i_257_75_506 (.A1(n_257_75_252), .A2(n_257_75_129), .ZN(n_257_842));
   NOR2_X1 i_257_75_507 (.A1(n_257_75_254), .A2(n_257_75_129), .ZN(n_257_843));
   NOR2_X1 i_257_75_508 (.A1(n_257_75_258), .A2(n_257_75_129), .ZN(n_257_844));
   OR2_X1 i_257_75_509 (.A1(n_257_75_282), .A2(n_257_75_130), .ZN(n_257_75_129));
   OR2_X1 i_257_75_510 (.A1(n_257_75_135), .A2(n_257_75_134), .ZN(n_257_75_130));
   NOR2_X1 i_257_75_511 (.A1(n_257_75_246), .A2(n_257_75_131), .ZN(n_257_845));
   NOR2_X1 i_257_75_512 (.A1(n_257_75_247), .A2(n_257_75_131), .ZN(n_257_846));
   NOR2_X1 i_257_75_513 (.A1(n_257_75_248), .A2(n_257_75_131), .ZN(n_257_847));
   NOR2_X1 i_257_75_514 (.A1(n_257_75_249), .A2(n_257_75_131), .ZN(n_257_848));
   NOR2_X1 i_257_75_515 (.A1(n_257_75_250), .A2(n_257_75_131), .ZN(n_257_849));
   NOR2_X1 i_257_75_516 (.A1(n_257_75_252), .A2(n_257_75_131), .ZN(n_257_850));
   NOR2_X1 i_257_75_517 (.A1(n_257_75_254), .A2(n_257_75_131), .ZN(n_257_851));
   NOR2_X1 i_257_75_518 (.A1(n_257_75_258), .A2(n_257_75_131), .ZN(n_257_852));
   OR2_X1 i_257_75_519 (.A1(n_257_75_12), .A2(n_257_75_133), .ZN(n_257_75_131));
   NOR2_X1 i_257_75_520 (.A1(n_257_75_246), .A2(n_257_75_132), .ZN(n_257_853));
   NOR2_X1 i_257_75_521 (.A1(n_257_75_247), .A2(n_257_75_132), .ZN(n_257_854));
   NOR2_X1 i_257_75_522 (.A1(n_257_75_248), .A2(n_257_75_132), .ZN(n_257_855));
   NOR2_X1 i_257_75_523 (.A1(n_257_75_249), .A2(n_257_75_132), .ZN(n_257_856));
   NOR2_X1 i_257_75_524 (.A1(n_257_75_250), .A2(n_257_75_132), .ZN(n_257_857));
   NOR2_X1 i_257_75_525 (.A1(n_257_75_252), .A2(n_257_75_132), .ZN(n_257_858));
   NOR2_X1 i_257_75_526 (.A1(n_257_75_254), .A2(n_257_75_132), .ZN(n_257_859));
   NOR2_X1 i_257_75_527 (.A1(n_257_75_258), .A2(n_257_75_132), .ZN(n_257_860));
   OR2_X1 i_257_75_528 (.A1(n_257_75_282), .A2(n_257_75_133), .ZN(n_257_75_132));
   OAI21_X1 i_257_75_529 (.A(n_257_75_134), .B1(n_257_75_298), .B2(n_257_75_135), 
      .ZN(n_257_75_133));
   OAI21_X1 i_257_75_530 (.A(n_257_75_298), .B1(n_257_75_322), .B2(n_257_75_283), 
      .ZN(n_257_75_134));
   NOR2_X1 i_257_75_531 (.A1(PacketSize[4]), .A2(n_257_75_13), .ZN(n_257_75_135));
   NOR2_X1 i_257_75_532 (.A1(n_257_75_140), .A2(n_257_75_136), .ZN(n_257_861));
   NOR2_X1 i_257_75_533 (.A1(n_257_75_141), .A2(n_257_75_136), .ZN(n_257_862));
   NOR2_X1 i_257_75_534 (.A1(n_257_75_142), .A2(n_257_75_136), .ZN(n_257_863));
   NOR2_X1 i_257_75_535 (.A1(n_257_75_143), .A2(n_257_75_136), .ZN(n_257_864));
   NOR2_X1 i_257_75_536 (.A1(n_257_75_144), .A2(n_257_75_136), .ZN(n_257_865));
   NOR2_X1 i_257_75_537 (.A1(n_257_75_145), .A2(n_257_75_136), .ZN(n_257_866));
   NOR2_X1 i_257_75_538 (.A1(n_257_75_146), .A2(n_257_75_136), .ZN(n_257_867));
   NOR2_X1 i_257_75_539 (.A1(n_257_75_151), .A2(n_257_75_136), .ZN(n_257_868));
   OR2_X1 i_257_75_540 (.A1(n_257_75_10), .A2(n_257_75_138), .ZN(n_257_75_136));
   NOR2_X1 i_257_75_541 (.A1(n_257_75_140), .A2(n_257_75_137), .ZN(n_257_869));
   NOR2_X1 i_257_75_542 (.A1(n_257_75_141), .A2(n_257_75_137), .ZN(n_257_870));
   NOR2_X1 i_257_75_543 (.A1(n_257_75_142), .A2(n_257_75_137), .ZN(n_257_871));
   NOR2_X1 i_257_75_544 (.A1(n_257_75_143), .A2(n_257_75_137), .ZN(n_257_872));
   NOR2_X1 i_257_75_545 (.A1(n_257_75_144), .A2(n_257_75_137), .ZN(n_257_873));
   NOR2_X1 i_257_75_546 (.A1(n_257_75_145), .A2(n_257_75_137), .ZN(n_257_874));
   NOR2_X1 i_257_75_547 (.A1(n_257_75_146), .A2(n_257_75_137), .ZN(n_257_875));
   NOR2_X1 i_257_75_548 (.A1(n_257_75_151), .A2(n_257_75_137), .ZN(n_257_876));
   OR2_X1 i_257_75_549 (.A1(n_257_75_284), .A2(n_257_75_138), .ZN(n_257_75_137));
   OR2_X1 i_257_75_550 (.A1(n_257_75_150), .A2(n_257_75_149), .ZN(n_257_75_138));
   NOR2_X1 i_257_75_551 (.A1(n_257_75_140), .A2(n_257_75_139), .ZN(n_257_877));
   NOR2_X1 i_257_75_552 (.A1(n_257_75_141), .A2(n_257_75_139), .ZN(n_257_878));
   NOR2_X1 i_257_75_553 (.A1(n_257_75_142), .A2(n_257_75_139), .ZN(n_257_879));
   NOR2_X1 i_257_75_554 (.A1(n_257_75_143), .A2(n_257_75_139), .ZN(n_257_880));
   NOR2_X1 i_257_75_555 (.A1(n_257_75_144), .A2(n_257_75_139), .ZN(n_257_881));
   NOR2_X1 i_257_75_556 (.A1(n_257_75_145), .A2(n_257_75_139), .ZN(n_257_882));
   NOR2_X1 i_257_75_557 (.A1(n_257_75_146), .A2(n_257_75_139), .ZN(n_257_883));
   NOR2_X1 i_257_75_558 (.A1(n_257_75_151), .A2(n_257_75_139), .ZN(n_257_884));
   OR2_X1 i_257_75_559 (.A1(n_257_75_10), .A2(n_257_75_148), .ZN(n_257_75_139));
   NOR2_X1 i_257_75_560 (.A1(n_257_75_147), .A2(n_257_75_140), .ZN(n_257_885));
   NAND3_X1 i_257_75_561 (.A1(n_257_75_294), .A2(n_257_75_216), .A3(n_257_75_296), 
      .ZN(n_257_75_140));
   NOR2_X1 i_257_75_562 (.A1(n_257_75_147), .A2(n_257_75_141), .ZN(n_257_886));
   NAND3_X1 i_257_75_563 (.A1(n_151), .A2(n_257_75_216), .A3(n_257_75_296), 
      .ZN(n_257_75_141));
   NOR2_X1 i_257_75_564 (.A1(n_257_75_147), .A2(n_257_75_142), .ZN(n_257_887));
   OR2_X1 i_257_75_565 (.A1(n_257_75_204), .A2(n_257_75_152), .ZN(n_257_75_142));
   NOR2_X1 i_257_75_566 (.A1(n_257_75_147), .A2(n_257_75_143), .ZN(n_257_888));
   OR2_X1 i_257_75_567 (.A1(n_257_75_214), .A2(n_257_75_152), .ZN(n_257_75_143));
   NOR2_X1 i_257_75_568 (.A1(n_257_75_147), .A2(n_257_75_144), .ZN(n_257_889));
   NAND3_X1 i_257_75_569 (.A1(n_257_75_294), .A2(n_257_75_216), .A3(
      PacketSize[2]), .ZN(n_257_75_144));
   NOR2_X1 i_257_75_570 (.A1(n_257_75_147), .A2(n_257_75_145), .ZN(n_257_890));
   NAND3_X1 i_257_75_571 (.A1(n_151), .A2(n_257_75_216), .A3(PacketSize[2]), 
      .ZN(n_257_75_145));
   NOR2_X1 i_257_75_572 (.A1(n_257_75_147), .A2(n_257_75_146), .ZN(n_257_891));
   NAND3_X1 i_257_75_573 (.A1(n_257_75_294), .A2(n_257_75_215), .A3(n_257_75_152), 
      .ZN(n_257_75_146));
   NOR2_X1 i_257_75_574 (.A1(n_257_75_151), .A2(n_257_75_147), .ZN(n_257_892));
   OR2_X1 i_257_75_575 (.A1(n_257_75_284), .A2(n_257_75_148), .ZN(n_257_75_147));
   OAI21_X1 i_257_75_576 (.A(n_257_75_149), .B1(n_257_75_298), .B2(n_257_75_150), 
      .ZN(n_257_75_148));
   OAI21_X1 i_257_75_577 (.A(n_257_75_298), .B1(n_257_75_322), .B2(n_257_75_285), 
      .ZN(n_257_75_149));
   NOR2_X1 i_257_75_578 (.A1(PacketSize[4]), .A2(n_257_75_11), .ZN(n_257_75_150));
   NAND3_X1 i_257_75_579 (.A1(n_151), .A2(n_257_75_215), .A3(n_257_75_152), 
      .ZN(n_257_75_151));
   OAI21_X1 i_257_75_580 (.A(n_257_75_254), .B1(n_257_75_296), .B2(n_257_75_257), 
      .ZN(n_257_75_152));
   NOR2_X1 i_257_75_581 (.A1(n_257_75_246), .A2(n_257_75_153), .ZN(n_257_893));
   NOR2_X1 i_257_75_582 (.A1(n_257_75_247), .A2(n_257_75_153), .ZN(n_257_894));
   NOR2_X1 i_257_75_583 (.A1(n_257_75_248), .A2(n_257_75_153), .ZN(n_257_895));
   NOR2_X1 i_257_75_584 (.A1(n_257_75_249), .A2(n_257_75_153), .ZN(n_257_896));
   NOR2_X1 i_257_75_585 (.A1(n_257_75_250), .A2(n_257_75_153), .ZN(n_257_897));
   NOR2_X1 i_257_75_586 (.A1(n_257_75_252), .A2(n_257_75_153), .ZN(n_257_898));
   NAND3_X1 i_257_75_587 (.A1(n_257_75_322), .A2(n_257_75_297), .A3(
      PacketSize[5]), .ZN(n_257_75_153));
   NOR2_X1 i_257_75_588 (.A1(n_257_75_157), .A2(n_257_75_154), .ZN(n_257_899));
   NOR2_X1 i_257_75_589 (.A1(n_257_75_158), .A2(n_257_75_154), .ZN(n_257_900));
   NOR2_X1 i_257_75_590 (.A1(n_257_75_159), .A2(n_257_75_154), .ZN(n_257_901));
   NOR2_X1 i_257_75_591 (.A1(n_257_75_160), .A2(n_257_75_154), .ZN(n_257_902));
   NOR2_X1 i_257_75_592 (.A1(n_257_75_161), .A2(n_257_75_154), .ZN(n_257_903));
   NOR2_X1 i_257_75_593 (.A1(n_257_75_162), .A2(n_257_75_154), .ZN(n_257_904));
   NOR2_X1 i_257_75_594 (.A1(n_257_75_163), .A2(n_257_75_154), .ZN(n_257_905));
   NOR2_X1 i_257_75_595 (.A1(n_257_75_172), .A2(n_257_75_154), .ZN(n_257_906));
   NAND3_X1 i_257_75_596 (.A1(n_257_75_298), .A2(n_257_75_322), .A3(n_257_75_170), 
      .ZN(n_257_75_154));
   NOR2_X1 i_257_75_597 (.A1(n_257_75_157), .A2(n_257_75_155), .ZN(n_257_907));
   NOR2_X1 i_257_75_598 (.A1(n_257_75_158), .A2(n_257_75_155), .ZN(n_257_908));
   NOR2_X1 i_257_75_599 (.A1(n_257_75_159), .A2(n_257_75_155), .ZN(n_257_909));
   NOR2_X1 i_257_75_600 (.A1(n_257_75_160), .A2(n_257_75_155), .ZN(n_257_910));
   NOR2_X1 i_257_75_601 (.A1(n_257_75_161), .A2(n_257_75_155), .ZN(n_257_911));
   NOR2_X1 i_257_75_602 (.A1(n_257_75_162), .A2(n_257_75_155), .ZN(n_257_912));
   NOR2_X1 i_257_75_603 (.A1(n_257_75_163), .A2(n_257_75_155), .ZN(n_257_913));
   NOR2_X1 i_257_75_604 (.A1(n_257_75_172), .A2(n_257_75_155), .ZN(n_257_914));
   OR3_X1 i_257_75_605 (.A1(PacketSize[5]), .A2(n_257_75_170), .A3(n_257_75_167), 
      .ZN(n_257_75_155));
   NOR2_X1 i_257_75_606 (.A1(n_257_75_157), .A2(n_257_75_156), .ZN(n_257_915));
   NOR2_X1 i_257_75_607 (.A1(n_257_75_158), .A2(n_257_75_156), .ZN(n_257_916));
   NOR2_X1 i_257_75_608 (.A1(n_257_75_159), .A2(n_257_75_156), .ZN(n_257_917));
   NOR2_X1 i_257_75_609 (.A1(n_257_75_160), .A2(n_257_75_156), .ZN(n_257_918));
   NOR2_X1 i_257_75_610 (.A1(n_257_75_161), .A2(n_257_75_156), .ZN(n_257_919));
   NOR2_X1 i_257_75_611 (.A1(n_257_75_162), .A2(n_257_75_156), .ZN(n_257_920));
   NOR2_X1 i_257_75_612 (.A1(n_257_75_163), .A2(n_257_75_156), .ZN(n_257_921));
   NOR2_X1 i_257_75_613 (.A1(n_257_75_172), .A2(n_257_75_156), .ZN(n_257_922));
   NAND2_X1 i_257_75_614 (.A1(n_257_75_170), .A2(n_257_75_165), .ZN(n_257_75_156));
   NOR2_X1 i_257_75_615 (.A1(n_257_75_164), .A2(n_257_75_157), .ZN(n_257_923));
   OR3_X1 i_257_75_616 (.A1(n_151), .A2(n_257_75_4), .A3(n_257_75_6), .ZN(
      n_257_75_157));
   NOR2_X1 i_257_75_617 (.A1(n_257_75_164), .A2(n_257_75_158), .ZN(n_257_924));
   OR3_X1 i_257_75_618 (.A1(n_257_75_294), .A2(n_257_75_4), .A3(n_257_75_6), 
      .ZN(n_257_75_158));
   NOR2_X1 i_257_75_619 (.A1(n_257_75_164), .A2(n_257_75_159), .ZN(n_257_925));
   OR3_X1 i_257_75_620 (.A1(n_151), .A2(n_257_75_287), .A3(n_257_75_6), .ZN(
      n_257_75_159));
   NOR2_X1 i_257_75_621 (.A1(n_257_75_164), .A2(n_257_75_160), .ZN(n_257_926));
   OR3_X1 i_257_75_622 (.A1(n_257_75_294), .A2(n_257_75_287), .A3(n_257_75_6), 
      .ZN(n_257_75_160));
   NOR2_X1 i_257_75_623 (.A1(n_257_75_164), .A2(n_257_75_161), .ZN(n_257_927));
   NAND3_X1 i_257_75_624 (.A1(n_257_75_294), .A2(n_257_75_287), .A3(n_257_75_6), 
      .ZN(n_257_75_161));
   NOR2_X1 i_257_75_625 (.A1(n_257_75_164), .A2(n_257_75_162), .ZN(n_257_928));
   NAND3_X1 i_257_75_626 (.A1(n_151), .A2(n_257_75_287), .A3(n_257_75_6), 
      .ZN(n_257_75_162));
   NOR2_X1 i_257_75_627 (.A1(n_257_75_164), .A2(n_257_75_163), .ZN(n_257_929));
   NAND3_X1 i_257_75_628 (.A1(n_257_75_294), .A2(n_257_75_4), .A3(n_257_75_6), 
      .ZN(n_257_75_163));
   NOR2_X1 i_257_75_629 (.A1(n_257_75_172), .A2(n_257_75_164), .ZN(n_257_930));
   OR2_X1 i_257_75_630 (.A1(n_257_75_170), .A2(n_257_75_166), .ZN(n_257_75_164));
   INV_X1 i_257_75_631 (.A(n_257_75_166), .ZN(n_257_75_165));
   OAI221_X1 i_257_75_632 (.A(n_257_75_167), .B1(n_257_75_7), .B2(n_257_75_263), 
      .C1(n_257_75_298), .C2(n_257_75_168), .ZN(n_257_75_166));
   OAI21_X1 i_257_75_633 (.A(n_257_75_169), .B1(n_257_75_322), .B2(n_257_75_171), 
      .ZN(n_257_75_167));
   INV_X1 i_257_75_634 (.A(n_257_75_169), .ZN(n_257_75_168));
   NAND2_X1 i_257_75_635 (.A1(n_257_75_322), .A2(n_257_75_171), .ZN(n_257_75_169));
   AOI21_X1 i_257_75_636 (.A(n_257_75_171), .B1(PacketSize[3]), .B2(n_257_75_7), 
      .ZN(n_257_75_170));
   NOR2_X1 i_257_75_637 (.A1(PacketSize[3]), .A2(n_257_75_7), .ZN(n_257_75_171));
   NAND3_X1 i_257_75_638 (.A1(n_151), .A2(n_257_75_4), .A3(n_257_75_6), .ZN(
      n_257_75_172));
   NOR2_X1 i_257_75_639 (.A1(n_257_75_176), .A2(n_257_75_173), .ZN(n_257_931));
   NOR2_X1 i_257_75_640 (.A1(n_257_75_177), .A2(n_257_75_173), .ZN(n_257_932));
   NOR2_X1 i_257_75_641 (.A1(n_257_75_178), .A2(n_257_75_173), .ZN(n_257_933));
   NOR2_X1 i_257_75_642 (.A1(n_257_75_179), .A2(n_257_75_173), .ZN(n_257_934));
   NOR2_X1 i_257_75_643 (.A1(n_257_75_180), .A2(n_257_75_173), .ZN(n_257_935));
   NOR2_X1 i_257_75_644 (.A1(n_257_75_181), .A2(n_257_75_173), .ZN(n_257_936));
   NOR2_X1 i_257_75_645 (.A1(n_257_75_182), .A2(n_257_75_173), .ZN(n_257_937));
   NOR2_X1 i_257_75_646 (.A1(n_257_75_191), .A2(n_257_75_173), .ZN(n_257_938));
   NAND3_X1 i_257_75_647 (.A1(n_257_75_298), .A2(n_257_75_322), .A3(n_257_75_189), 
      .ZN(n_257_75_173));
   NOR2_X1 i_257_75_648 (.A1(n_257_75_176), .A2(n_257_75_174), .ZN(n_257_939));
   NOR2_X1 i_257_75_649 (.A1(n_257_75_177), .A2(n_257_75_174), .ZN(n_257_940));
   NOR2_X1 i_257_75_650 (.A1(n_257_75_178), .A2(n_257_75_174), .ZN(n_257_941));
   NOR2_X1 i_257_75_651 (.A1(n_257_75_179), .A2(n_257_75_174), .ZN(n_257_942));
   NOR2_X1 i_257_75_652 (.A1(n_257_75_180), .A2(n_257_75_174), .ZN(n_257_943));
   NOR2_X1 i_257_75_653 (.A1(n_257_75_181), .A2(n_257_75_174), .ZN(n_257_944));
   NOR2_X1 i_257_75_654 (.A1(n_257_75_182), .A2(n_257_75_174), .ZN(n_257_945));
   NOR2_X1 i_257_75_655 (.A1(n_257_75_191), .A2(n_257_75_174), .ZN(n_257_946));
   OR3_X1 i_257_75_656 (.A1(PacketSize[5]), .A2(n_257_75_189), .A3(n_257_75_186), 
      .ZN(n_257_75_174));
   NOR2_X1 i_257_75_657 (.A1(n_257_75_176), .A2(n_257_75_175), .ZN(n_257_947));
   NOR2_X1 i_257_75_658 (.A1(n_257_75_177), .A2(n_257_75_175), .ZN(n_257_948));
   NOR2_X1 i_257_75_659 (.A1(n_257_75_178), .A2(n_257_75_175), .ZN(n_257_949));
   NOR2_X1 i_257_75_660 (.A1(n_257_75_179), .A2(n_257_75_175), .ZN(n_257_950));
   NOR2_X1 i_257_75_661 (.A1(n_257_75_180), .A2(n_257_75_175), .ZN(n_257_951));
   NOR2_X1 i_257_75_662 (.A1(n_257_75_181), .A2(n_257_75_175), .ZN(n_257_952));
   NOR2_X1 i_257_75_663 (.A1(n_257_75_182), .A2(n_257_75_175), .ZN(n_257_953));
   NOR2_X1 i_257_75_664 (.A1(n_257_75_191), .A2(n_257_75_175), .ZN(n_257_954));
   NAND2_X1 i_257_75_665 (.A1(n_257_75_189), .A2(n_257_75_184), .ZN(n_257_75_175));
   NOR2_X1 i_257_75_666 (.A1(n_257_75_183), .A2(n_257_75_176), .ZN(n_257_955));
   OR2_X1 i_257_75_667 (.A1(n_257_75_2), .A2(n_257_75_251), .ZN(n_257_75_176));
   NOR2_X1 i_257_75_668 (.A1(n_257_75_183), .A2(n_257_75_177), .ZN(n_257_956));
   NAND2_X1 i_257_75_669 (.A1(n_257_75_288), .A2(n_257_75_253), .ZN(n_257_75_177));
   NOR2_X1 i_257_75_670 (.A1(n_257_75_183), .A2(n_257_75_178), .ZN(n_257_957));
   NAND2_X1 i_257_75_671 (.A1(n_257_75_288), .A2(n_257_75_257), .ZN(n_257_75_178));
   NOR2_X1 i_257_75_672 (.A1(n_257_75_183), .A2(n_257_75_179), .ZN(n_257_958));
   NAND3_X1 i_257_75_673 (.A1(n_257_1091), .A2(PacketSize[0]), .A3(n_257_75_288), 
      .ZN(n_257_75_179));
   NOR2_X1 i_257_75_674 (.A1(n_257_75_183), .A2(n_257_75_180), .ZN(n_257_959));
   OR2_X1 i_257_75_675 (.A1(n_257_75_288), .A2(n_257_75_251), .ZN(n_257_75_180));
   NOR2_X1 i_257_75_676 (.A1(n_257_75_183), .A2(n_257_75_181), .ZN(n_257_960));
   NAND2_X1 i_257_75_677 (.A1(n_257_75_2), .A2(n_257_75_253), .ZN(n_257_75_181));
   NOR2_X1 i_257_75_678 (.A1(n_257_75_183), .A2(n_257_75_182), .ZN(n_257_961));
   NAND2_X1 i_257_75_679 (.A1(n_257_75_2), .A2(n_257_75_257), .ZN(n_257_75_182));
   NOR2_X1 i_257_75_680 (.A1(n_257_75_191), .A2(n_257_75_183), .ZN(n_257_962));
   OR2_X1 i_257_75_681 (.A1(n_257_75_189), .A2(n_257_75_185), .ZN(n_257_75_183));
   INV_X1 i_257_75_682 (.A(n_257_75_185), .ZN(n_257_75_184));
   OAI221_X1 i_257_75_683 (.A(n_257_75_186), .B1(n_257_75_3), .B2(n_257_75_263), 
      .C1(n_257_75_298), .C2(n_257_75_187), .ZN(n_257_75_185));
   OAI21_X1 i_257_75_684 (.A(n_257_75_188), .B1(n_257_75_322), .B2(n_257_75_190), 
      .ZN(n_257_75_186));
   INV_X1 i_257_75_685 (.A(n_257_75_188), .ZN(n_257_75_187));
   NAND2_X1 i_257_75_686 (.A1(n_257_75_322), .A2(n_257_75_190), .ZN(n_257_75_188));
   AOI21_X1 i_257_75_687 (.A(n_257_75_190), .B1(PacketSize[3]), .B2(n_257_75_3), 
      .ZN(n_257_75_189));
   NOR2_X1 i_257_75_688 (.A1(PacketSize[3]), .A2(n_257_75_3), .ZN(n_257_75_190));
   NAND3_X1 i_257_75_689 (.A1(n_257_1091), .A2(PacketSize[0]), .A3(n_257_75_2), 
      .ZN(n_257_75_191));
   NOR2_X1 i_257_75_690 (.A1(n_257_75_195), .A2(n_257_75_192), .ZN(n_257_963));
   NOR2_X1 i_257_75_691 (.A1(n_257_75_196), .A2(n_257_75_192), .ZN(n_257_964));
   NOR2_X1 i_257_75_692 (.A1(n_257_75_197), .A2(n_257_75_192), .ZN(n_257_965));
   NOR2_X1 i_257_75_693 (.A1(n_257_75_198), .A2(n_257_75_192), .ZN(n_257_966));
   NOR2_X1 i_257_75_694 (.A1(n_257_75_199), .A2(n_257_75_192), .ZN(n_257_967));
   NOR2_X1 i_257_75_695 (.A1(n_257_75_201), .A2(n_257_75_192), .ZN(n_257_968));
   NOR2_X1 i_257_75_696 (.A1(n_257_75_203), .A2(n_257_75_192), .ZN(n_257_969));
   NOR2_X1 i_257_75_697 (.A1(n_257_75_213), .A2(n_257_75_192), .ZN(n_257_970));
   NAND3_X1 i_257_75_698 (.A1(n_257_75_298), .A2(n_257_75_322), .A3(n_257_75_211), 
      .ZN(n_257_75_192));
   NOR2_X1 i_257_75_699 (.A1(n_257_75_195), .A2(n_257_75_193), .ZN(n_257_971));
   NOR2_X1 i_257_75_700 (.A1(n_257_75_196), .A2(n_257_75_193), .ZN(n_257_972));
   NOR2_X1 i_257_75_701 (.A1(n_257_75_197), .A2(n_257_75_193), .ZN(n_257_973));
   NOR2_X1 i_257_75_702 (.A1(n_257_75_198), .A2(n_257_75_193), .ZN(n_257_974));
   NOR2_X1 i_257_75_703 (.A1(n_257_75_199), .A2(n_257_75_193), .ZN(n_257_975));
   NOR2_X1 i_257_75_704 (.A1(n_257_75_201), .A2(n_257_75_193), .ZN(n_257_976));
   NOR2_X1 i_257_75_705 (.A1(n_257_75_203), .A2(n_257_75_193), .ZN(n_257_977));
   NOR2_X1 i_257_75_706 (.A1(n_257_75_213), .A2(n_257_75_193), .ZN(n_257_978));
   OR3_X1 i_257_75_707 (.A1(PacketSize[5]), .A2(n_257_75_211), .A3(n_257_75_208), 
      .ZN(n_257_75_193));
   NOR2_X1 i_257_75_708 (.A1(n_257_75_195), .A2(n_257_75_194), .ZN(n_257_979));
   NOR2_X1 i_257_75_709 (.A1(n_257_75_196), .A2(n_257_75_194), .ZN(n_257_980));
   NOR2_X1 i_257_75_710 (.A1(n_257_75_197), .A2(n_257_75_194), .ZN(n_257_981));
   NOR2_X1 i_257_75_711 (.A1(n_257_75_198), .A2(n_257_75_194), .ZN(n_257_982));
   NOR2_X1 i_257_75_712 (.A1(n_257_75_199), .A2(n_257_75_194), .ZN(n_257_983));
   NOR2_X1 i_257_75_713 (.A1(n_257_75_201), .A2(n_257_75_194), .ZN(n_257_984));
   NOR2_X1 i_257_75_714 (.A1(n_257_75_203), .A2(n_257_75_194), .ZN(n_257_985));
   NOR2_X1 i_257_75_715 (.A1(n_257_75_213), .A2(n_257_75_194), .ZN(n_257_986));
   NAND2_X1 i_257_75_716 (.A1(n_257_75_211), .A2(n_257_75_206), .ZN(n_257_75_194));
   NOR2_X1 i_257_75_717 (.A1(n_257_75_205), .A2(n_257_75_195), .ZN(n_257_987));
   OR2_X1 i_257_75_718 (.A1(n_257_75_0), .A2(n_257_75_200), .ZN(n_257_75_195));
   NOR2_X1 i_257_75_719 (.A1(n_257_75_205), .A2(n_257_75_196), .ZN(n_257_988));
   OR2_X1 i_257_75_720 (.A1(n_257_75_0), .A2(n_257_75_202), .ZN(n_257_75_196));
   NOR2_X1 i_257_75_721 (.A1(n_257_75_205), .A2(n_257_75_197), .ZN(n_257_989));
   OR2_X1 i_257_75_722 (.A1(n_257_75_0), .A2(n_257_75_204), .ZN(n_257_75_197));
   NOR2_X1 i_257_75_723 (.A1(n_257_75_205), .A2(n_257_75_198), .ZN(n_257_990));
   OR2_X1 i_257_75_724 (.A1(n_257_75_0), .A2(n_257_75_214), .ZN(n_257_75_198));
   NOR2_X1 i_257_75_725 (.A1(n_257_75_205), .A2(n_257_75_199), .ZN(n_257_991));
   NAND3_X1 i_257_75_726 (.A1(n_257_75_294), .A2(n_257_75_216), .A3(n_257_75_0), 
      .ZN(n_257_75_199));
   NAND2_X1 i_257_75_727 (.A1(n_257_75_294), .A2(n_257_75_216), .ZN(n_257_75_200));
   NOR2_X1 i_257_75_728 (.A1(n_257_75_205), .A2(n_257_75_201), .ZN(n_257_992));
   NAND3_X1 i_257_75_729 (.A1(n_151), .A2(n_257_75_216), .A3(n_257_75_0), 
      .ZN(n_257_75_201));
   NAND2_X1 i_257_75_730 (.A1(n_151), .A2(n_257_75_216), .ZN(n_257_75_202));
   NOR2_X1 i_257_75_731 (.A1(n_257_75_205), .A2(n_257_75_203), .ZN(n_257_993));
   NAND3_X1 i_257_75_732 (.A1(n_257_75_294), .A2(n_257_75_215), .A3(n_257_75_0), 
      .ZN(n_257_75_203));
   NAND2_X1 i_257_75_733 (.A1(n_257_75_294), .A2(n_257_75_215), .ZN(n_257_75_204));
   NOR2_X1 i_257_75_734 (.A1(n_257_75_213), .A2(n_257_75_205), .ZN(n_257_994));
   OR2_X1 i_257_75_735 (.A1(n_257_75_211), .A2(n_257_75_207), .ZN(n_257_75_205));
   INV_X1 i_257_75_736 (.A(n_257_75_207), .ZN(n_257_75_206));
   OAI221_X1 i_257_75_737 (.A(n_257_75_208), .B1(n_257_75_1), .B2(n_257_75_263), 
      .C1(n_257_75_298), .C2(n_257_75_209), .ZN(n_257_75_207));
   OAI21_X1 i_257_75_738 (.A(n_257_75_210), .B1(n_257_75_322), .B2(n_257_75_212), 
      .ZN(n_257_75_208));
   INV_X1 i_257_75_739 (.A(n_257_75_210), .ZN(n_257_75_209));
   NAND2_X1 i_257_75_740 (.A1(n_257_75_322), .A2(n_257_75_212), .ZN(n_257_75_210));
   AOI21_X1 i_257_75_741 (.A(n_257_75_212), .B1(PacketSize[3]), .B2(n_257_75_1), 
      .ZN(n_257_75_211));
   NOR2_X1 i_257_75_742 (.A1(PacketSize[3]), .A2(n_257_75_1), .ZN(n_257_75_212));
   NAND3_X1 i_257_75_743 (.A1(n_151), .A2(n_257_75_215), .A3(n_257_75_0), 
      .ZN(n_257_75_213));
   NAND2_X1 i_257_75_744 (.A1(n_151), .A2(n_257_75_215), .ZN(n_257_75_214));
   INV_X1 i_257_75_745 (.A(n_257_75_216), .ZN(n_257_75_215));
   NOR2_X1 i_257_75_746 (.A1(n_257_75_257), .A2(n_257_75_253), .ZN(n_257_75_216));
   NOR2_X1 i_257_75_747 (.A1(n_257_75_220), .A2(n_257_75_217), .ZN(n_257_995));
   NOR2_X1 i_257_75_748 (.A1(n_257_75_221), .A2(n_257_75_217), .ZN(n_257_996));
   NOR2_X1 i_257_75_749 (.A1(n_257_75_222), .A2(n_257_75_217), .ZN(n_257_997));
   NOR2_X1 i_257_75_750 (.A1(n_257_75_223), .A2(n_257_75_217), .ZN(n_257_998));
   NOR2_X1 i_257_75_751 (.A1(n_257_75_224), .A2(n_257_75_217), .ZN(n_257_999));
   NOR2_X1 i_257_75_752 (.A1(n_257_75_225), .A2(n_257_75_217), .ZN(n_257_1000));
   NOR2_X1 i_257_75_753 (.A1(n_257_75_226), .A2(n_257_75_217), .ZN(n_257_1001));
   NOR2_X1 i_257_75_754 (.A1(n_257_75_229), .A2(n_257_75_217), .ZN(n_257_1002));
   NAND3_X1 i_257_75_755 (.A1(n_257_75_291), .A2(n_257_75_228), .A3(n_257_75_290), 
      .ZN(n_257_75_217));
   NOR2_X1 i_257_75_756 (.A1(n_257_75_220), .A2(n_257_75_218), .ZN(n_257_1003));
   NOR2_X1 i_257_75_757 (.A1(n_257_75_221), .A2(n_257_75_218), .ZN(n_257_1004));
   NOR2_X1 i_257_75_758 (.A1(n_257_75_222), .A2(n_257_75_218), .ZN(n_257_1005));
   NOR2_X1 i_257_75_759 (.A1(n_257_75_223), .A2(n_257_75_218), .ZN(n_257_1006));
   NOR2_X1 i_257_75_760 (.A1(n_257_75_224), .A2(n_257_75_218), .ZN(n_257_1007));
   NOR2_X1 i_257_75_761 (.A1(n_257_75_225), .A2(n_257_75_218), .ZN(n_257_1008));
   NOR2_X1 i_257_75_762 (.A1(n_257_75_226), .A2(n_257_75_218), .ZN(n_257_1009));
   NOR2_X1 i_257_75_763 (.A1(n_257_75_229), .A2(n_257_75_218), .ZN(n_257_1010));
   NAND3_X1 i_257_75_764 (.A1(n_257_75_291), .A2(n_257_75_228), .A3(n_257_7), 
      .ZN(n_257_75_218));
   NOR2_X1 i_257_75_765 (.A1(n_257_75_220), .A2(n_257_75_219), .ZN(n_257_1011));
   NOR2_X1 i_257_75_766 (.A1(n_257_75_221), .A2(n_257_75_219), .ZN(n_257_1012));
   NOR2_X1 i_257_75_767 (.A1(n_257_75_222), .A2(n_257_75_219), .ZN(n_257_1013));
   NOR2_X1 i_257_75_768 (.A1(n_257_75_223), .A2(n_257_75_219), .ZN(n_257_1014));
   NOR2_X1 i_257_75_769 (.A1(n_257_75_224), .A2(n_257_75_219), .ZN(n_257_1015));
   NOR2_X1 i_257_75_770 (.A1(n_257_75_225), .A2(n_257_75_219), .ZN(n_257_1016));
   NOR2_X1 i_257_75_771 (.A1(n_257_75_226), .A2(n_257_75_219), .ZN(n_257_1017));
   NOR2_X1 i_257_75_772 (.A1(n_257_75_229), .A2(n_257_75_219), .ZN(n_257_1018));
   NAND3_X1 i_257_75_773 (.A1(n_257_8), .A2(n_257_75_228), .A3(n_257_75_290), 
      .ZN(n_257_75_219));
   NOR2_X1 i_257_75_774 (.A1(n_257_75_227), .A2(n_257_75_220), .ZN(n_257_1019));
   NAND2_X1 i_257_75_775 (.A1(n_257_75_289), .A2(n_257_75_257), .ZN(n_257_75_220));
   NOR2_X1 i_257_75_776 (.A1(n_257_75_227), .A2(n_257_75_221), .ZN(n_257_1020));
   NAND3_X1 i_257_75_777 (.A1(n_257_1091), .A2(PacketSize[0]), .A3(n_257_75_289), 
      .ZN(n_257_75_221));
   NOR2_X1 i_257_75_778 (.A1(n_257_75_227), .A2(n_257_75_222), .ZN(n_257_1021));
   OR2_X1 i_257_75_779 (.A1(n_257_6), .A2(n_257_75_251), .ZN(n_257_75_222));
   NOR2_X1 i_257_75_780 (.A1(n_257_75_227), .A2(n_257_75_223), .ZN(n_257_1022));
   NAND2_X1 i_257_75_781 (.A1(n_257_75_289), .A2(n_257_75_253), .ZN(n_257_75_223));
   NOR2_X1 i_257_75_782 (.A1(n_257_75_227), .A2(n_257_75_224), .ZN(n_257_1023));
   NAND2_X1 i_257_75_783 (.A1(n_257_6), .A2(n_257_75_257), .ZN(n_257_75_224));
   NOR2_X1 i_257_75_784 (.A1(n_257_75_227), .A2(n_257_75_225), .ZN(n_257_1024));
   NAND3_X1 i_257_75_785 (.A1(n_257_1091), .A2(PacketSize[0]), .A3(n_257_6), 
      .ZN(n_257_75_225));
   NOR2_X1 i_257_75_786 (.A1(n_257_75_227), .A2(n_257_75_226), .ZN(n_257_1025));
   OR2_X1 i_257_75_787 (.A1(n_257_75_289), .A2(n_257_75_251), .ZN(n_257_75_226));
   NOR2_X1 i_257_75_788 (.A1(n_257_75_229), .A2(n_257_75_227), .ZN(n_257_1026));
   NAND3_X1 i_257_75_789 (.A1(n_257_8), .A2(n_257_75_228), .A3(n_257_7), 
      .ZN(n_257_75_227));
   NOR3_X1 i_257_75_790 (.A1(n_257_11), .A2(n_257_9), .A3(n_257_10), .ZN(
      n_257_75_228));
   NAND2_X1 i_257_75_791 (.A1(n_257_6), .A2(n_257_75_253), .ZN(n_257_75_229));
   NOR2_X1 i_257_75_792 (.A1(n_257_75_233), .A2(n_257_75_230), .ZN(n_257_1027));
   NOR2_X1 i_257_75_793 (.A1(n_257_75_234), .A2(n_257_75_230), .ZN(n_257_1028));
   NOR2_X1 i_257_75_794 (.A1(n_257_75_235), .A2(n_257_75_230), .ZN(n_257_1029));
   NOR2_X1 i_257_75_795 (.A1(n_257_75_236), .A2(n_257_75_230), .ZN(n_257_1030));
   NOR2_X1 i_257_75_796 (.A1(n_257_75_237), .A2(n_257_75_230), .ZN(n_257_1031));
   NOR2_X1 i_257_75_797 (.A1(n_257_75_238), .A2(n_257_75_230), .ZN(n_257_1032));
   NOR2_X1 i_257_75_798 (.A1(n_257_75_239), .A2(n_257_75_230), .ZN(n_257_1033));
   NOR2_X1 i_257_75_799 (.A1(n_257_75_242), .A2(n_257_75_230), .ZN(n_257_1034));
   NAND3_X1 i_257_75_800 (.A1(n_257_75_293), .A2(n_257_75_241), .A3(n_257_75_292), 
      .ZN(n_257_75_230));
   NOR2_X1 i_257_75_801 (.A1(n_257_75_233), .A2(n_257_75_231), .ZN(n_257_1035));
   NOR2_X1 i_257_75_802 (.A1(n_257_75_234), .A2(n_257_75_231), .ZN(n_257_1036));
   NOR2_X1 i_257_75_803 (.A1(n_257_75_235), .A2(n_257_75_231), .ZN(n_257_1037));
   NOR2_X1 i_257_75_804 (.A1(n_257_75_236), .A2(n_257_75_231), .ZN(n_257_1038));
   NOR2_X1 i_257_75_805 (.A1(n_257_75_237), .A2(n_257_75_231), .ZN(n_257_1039));
   NOR2_X1 i_257_75_806 (.A1(n_257_75_238), .A2(n_257_75_231), .ZN(n_257_1040));
   NOR2_X1 i_257_75_807 (.A1(n_257_75_239), .A2(n_257_75_231), .ZN(n_257_1041));
   NOR2_X1 i_257_75_808 (.A1(n_257_75_242), .A2(n_257_75_231), .ZN(n_257_1042));
   NAND3_X1 i_257_75_809 (.A1(n_257_75_293), .A2(n_257_75_241), .A3(n_257_1), 
      .ZN(n_257_75_231));
   NOR2_X1 i_257_75_810 (.A1(n_257_75_233), .A2(n_257_75_232), .ZN(n_257_1043));
   NOR2_X1 i_257_75_811 (.A1(n_257_75_234), .A2(n_257_75_232), .ZN(n_257_1044));
   NOR2_X1 i_257_75_812 (.A1(n_257_75_235), .A2(n_257_75_232), .ZN(n_257_1045));
   NOR2_X1 i_257_75_813 (.A1(n_257_75_236), .A2(n_257_75_232), .ZN(n_257_1046));
   NOR2_X1 i_257_75_814 (.A1(n_257_75_237), .A2(n_257_75_232), .ZN(n_257_1047));
   NOR2_X1 i_257_75_815 (.A1(n_257_75_238), .A2(n_257_75_232), .ZN(n_257_1048));
   NOR2_X1 i_257_75_816 (.A1(n_257_75_239), .A2(n_257_75_232), .ZN(n_257_1049));
   NOR2_X1 i_257_75_817 (.A1(n_257_75_242), .A2(n_257_75_232), .ZN(n_257_1050));
   NAND3_X1 i_257_75_818 (.A1(n_257_2), .A2(n_257_75_241), .A3(n_257_75_292), 
      .ZN(n_257_75_232));
   NOR2_X1 i_257_75_819 (.A1(n_257_75_240), .A2(n_257_75_233), .ZN(n_257_1051));
   OR3_X1 i_257_75_820 (.A1(n_257_75_295), .A2(n_151), .A3(n_257_0), .ZN(
      n_257_75_233));
   NOR2_X1 i_257_75_821 (.A1(n_257_75_240), .A2(n_257_75_234), .ZN(n_257_1052));
   OR3_X1 i_257_75_822 (.A1(n_257_75_295), .A2(n_257_75_294), .A3(n_257_0), 
      .ZN(n_257_75_234));
   NOR2_X1 i_257_75_823 (.A1(n_257_75_240), .A2(n_257_75_235), .ZN(n_257_1053));
   OR3_X1 i_257_75_824 (.A1(n_32), .A2(n_151), .A3(n_257_0), .ZN(n_257_75_235));
   NOR2_X1 i_257_75_825 (.A1(n_257_75_240), .A2(n_257_75_236), .ZN(n_257_1054));
   OR3_X1 i_257_75_826 (.A1(n_32), .A2(n_257_75_294), .A3(n_257_0), .ZN(
      n_257_75_236));
   NOR2_X1 i_257_75_827 (.A1(n_257_75_240), .A2(n_257_75_237), .ZN(n_257_1055));
   NAND3_X1 i_257_75_828 (.A1(n_32), .A2(n_257_75_294), .A3(n_257_0), .ZN(
      n_257_75_237));
   NOR2_X1 i_257_75_829 (.A1(n_257_75_240), .A2(n_257_75_238), .ZN(n_257_1056));
   NAND3_X1 i_257_75_830 (.A1(n_32), .A2(n_151), .A3(n_257_0), .ZN(n_257_75_238));
   NOR2_X1 i_257_75_831 (.A1(n_257_75_240), .A2(n_257_75_239), .ZN(n_257_1057));
   NAND3_X1 i_257_75_832 (.A1(n_257_75_295), .A2(n_257_75_294), .A3(n_257_0), 
      .ZN(n_257_75_239));
   NOR2_X1 i_257_75_833 (.A1(n_257_75_242), .A2(n_257_75_240), .ZN(n_257_1058));
   NAND3_X1 i_257_75_834 (.A1(n_257_2), .A2(n_257_75_241), .A3(n_257_1), 
      .ZN(n_257_75_240));
   NOR3_X1 i_257_75_835 (.A1(n_257_5), .A2(n_257_3), .A3(n_257_4), .ZN(
      n_257_75_241));
   NAND3_X1 i_257_75_836 (.A1(n_257_75_295), .A2(n_151), .A3(n_257_0), .ZN(
      n_257_75_242));
   NOR2_X1 i_257_75_837 (.A1(n_257_75_246), .A2(n_257_75_243), .ZN(n_257_1059));
   NOR2_X1 i_257_75_838 (.A1(n_257_75_247), .A2(n_257_75_243), .ZN(n_257_1060));
   NOR2_X1 i_257_75_839 (.A1(n_257_75_248), .A2(n_257_75_243), .ZN(n_257_1061));
   NOR2_X1 i_257_75_840 (.A1(n_257_75_249), .A2(n_257_75_243), .ZN(n_257_1062));
   NOR2_X1 i_257_75_841 (.A1(n_257_75_250), .A2(n_257_75_243), .ZN(n_257_1063));
   NOR2_X1 i_257_75_842 (.A1(n_257_75_252), .A2(n_257_75_243), .ZN(n_257_1064));
   NOR2_X1 i_257_75_843 (.A1(n_257_75_254), .A2(n_257_75_243), .ZN(n_257_1065));
   NOR2_X1 i_257_75_844 (.A1(n_257_75_258), .A2(n_257_75_243), .ZN(n_257_1066));
   NAND3_X1 i_257_75_845 (.A1(n_257_75_298), .A2(n_257_75_322), .A3(n_257_75_261), 
      .ZN(n_257_75_243));
   NOR2_X1 i_257_75_846 (.A1(n_257_75_246), .A2(n_257_75_244), .ZN(n_257_1067));
   NOR2_X1 i_257_75_847 (.A1(n_257_75_247), .A2(n_257_75_244), .ZN(n_257_1068));
   NOR2_X1 i_257_75_848 (.A1(n_257_75_248), .A2(n_257_75_244), .ZN(n_257_1069));
   NOR2_X1 i_257_75_849 (.A1(n_257_75_249), .A2(n_257_75_244), .ZN(n_257_1070));
   NOR2_X1 i_257_75_850 (.A1(n_257_75_250), .A2(n_257_75_244), .ZN(n_257_1071));
   NOR2_X1 i_257_75_851 (.A1(n_257_75_252), .A2(n_257_75_244), .ZN(n_257_1072));
   NOR2_X1 i_257_75_852 (.A1(n_257_75_254), .A2(n_257_75_244), .ZN(n_257_1073));
   NOR2_X1 i_257_75_853 (.A1(n_257_75_258), .A2(n_257_75_244), .ZN(n_257_1074));
   OR3_X1 i_257_75_854 (.A1(PacketSize[5]), .A2(n_257_75_261), .A3(n_257_1094), 
      .ZN(n_257_75_244));
   NOR2_X1 i_257_75_855 (.A1(n_257_75_246), .A2(n_257_75_245), .ZN(n_257_1075));
   NOR2_X1 i_257_75_856 (.A1(n_257_75_247), .A2(n_257_75_245), .ZN(n_257_1076));
   NOR2_X1 i_257_75_857 (.A1(n_257_75_248), .A2(n_257_75_245), .ZN(n_257_1077));
   NOR2_X1 i_257_75_858 (.A1(n_257_75_249), .A2(n_257_75_245), .ZN(n_257_1078));
   NOR2_X1 i_257_75_859 (.A1(n_257_75_250), .A2(n_257_75_245), .ZN(n_257_1079));
   NOR2_X1 i_257_75_860 (.A1(n_257_75_252), .A2(n_257_75_245), .ZN(n_257_1080));
   NOR2_X1 i_257_75_861 (.A1(n_257_75_254), .A2(n_257_75_245), .ZN(n_257_1081));
   NOR2_X1 i_257_75_862 (.A1(n_257_75_258), .A2(n_257_75_245), .ZN(n_257_1082));
   OR2_X1 i_257_75_863 (.A1(n_257_1093), .A2(n_257_75_260), .ZN(n_257_75_245));
   NOR2_X1 i_257_75_864 (.A1(n_257_75_259), .A2(n_257_75_246), .ZN(n_257_1083));
   OR2_X1 i_257_75_865 (.A1(PacketSize[2]), .A2(n_257_75_251), .ZN(n_257_75_246));
   NOR2_X1 i_257_75_866 (.A1(n_257_75_259), .A2(n_257_75_247), .ZN(n_257_1084));
   NAND2_X1 i_257_75_867 (.A1(n_257_75_296), .A2(n_257_75_253), .ZN(n_257_75_247));
   NOR2_X1 i_257_75_868 (.A1(n_257_75_259), .A2(n_257_75_248), .ZN(n_257_1085));
   NAND2_X1 i_257_75_869 (.A1(PacketSize[2]), .A2(n_257_75_257), .ZN(
      n_257_75_248));
   NOR2_X1 i_257_75_870 (.A1(n_257_75_259), .A2(n_257_75_249), .ZN(n_257_1086));
   NAND3_X1 i_257_75_871 (.A1(n_257_1091), .A2(PacketSize[0]), .A3(PacketSize[2]), 
      .ZN(n_257_75_249));
   NOR2_X1 i_257_75_872 (.A1(n_257_75_259), .A2(n_257_75_250), .ZN(n_257_1087));
   OR2_X1 i_257_75_873 (.A1(n_257_75_296), .A2(n_257_75_251), .ZN(n_257_75_250));
   OR2_X1 i_257_75_874 (.A1(n_257_1091), .A2(PacketSize[0]), .ZN(n_257_75_251));
   NOR2_X1 i_257_75_875 (.A1(n_257_75_259), .A2(n_257_75_252), .ZN(n_257_1088));
   NAND2_X1 i_257_75_876 (.A1(PacketSize[2]), .A2(n_257_75_253), .ZN(
      n_257_75_252));
   AND2_X1 i_257_75_877 (.A1(PacketSize[1]), .A2(PacketSize[0]), .ZN(
      n_257_75_253));
   NOR2_X1 i_257_75_878 (.A1(n_257_75_259), .A2(n_257_75_254), .ZN(n_257_1089));
   INV_X1 i_257_75_879 (.A(n_257_75_255), .ZN(n_257_75_254));
   NOR2_X1 i_257_75_880 (.A1(PacketSize[2]), .A2(n_257_75_256), .ZN(n_257_75_255));
   INV_X1 i_257_75_881 (.A(n_257_75_257), .ZN(n_257_75_256));
   NOR2_X1 i_257_75_882 (.A1(PacketSize[1]), .A2(PacketSize[0]), .ZN(
      n_257_75_257));
   NOR2_X1 i_257_75_883 (.A1(n_257_75_259), .A2(n_257_75_258), .ZN(n_257_1090));
   NAND2_X1 i_257_75_884 (.A1(PacketSize[0]), .A2(n_257_75_320), .ZN(
      n_257_75_258));
   OR2_X1 i_257_75_885 (.A1(n_257_75_261), .A2(n_257_75_260), .ZN(n_257_75_259));
   NAND2_X1 i_257_75_886 (.A1(n_257_75_262), .A2(n_257_1094), .ZN(n_257_75_260));
   OAI21_X1 i_257_75_887 (.A(n_257_75_307), .B1(n_257_75_296), .B2(n_257_1091), 
      .ZN(n_257_1092));
   INV_X1 i_257_75_888 (.A(n_257_1093), .ZN(n_257_75_261));
   OAI21_X1 i_257_75_889 (.A(n_257_75_264), .B1(n_257_75_297), .B2(n_257_75_320), 
      .ZN(n_257_1093));
   OAI21_X1 i_257_75_890 (.A(n_257_75_319), .B1(n_257_75_322), .B2(n_257_75_300), 
      .ZN(n_257_1094));
   INV_X1 i_257_75_891 (.A(n_257_75_262), .ZN(n_257_1095));
   AOI21_X1 i_257_75_892 (.A(n_257_1096), .B1(PacketSize[5]), .B2(n_257_75_319), 
      .ZN(n_257_75_262));
   NAND3_X1 i_257_75_893 (.A1(n_257_75_322), .A2(n_257_75_297), .A3(n_257_75_298), 
      .ZN(n_257_75_263));
   INV_X1 i_257_75_894 (.A(n_257_75_300), .ZN(n_257_75_264));
   NAND2_X1 i_257_75_895 (.A1(n_257_75_297), .A2(n_257_75_296), .ZN(n_257_75_265));
   INV_X1 i_257_75_896 (.A(n_257_75_32), .ZN(n_257_75_266));
   INV_X1 i_257_75_897 (.A(n_257_75_30), .ZN(n_257_75_267));
   INV_X1 i_257_75_898 (.A(n_257_75_28), .ZN(n_257_75_268));
   INV_X1 i_257_75_899 (.A(n_257_75_26), .ZN(n_257_75_269));
   INV_X1 i_257_75_900 (.A(n_257_75_24), .ZN(n_257_75_270));
   INV_X1 i_257_75_901 (.A(n_257_75_25), .ZN(n_257_75_271));
   INV_X1 i_257_75_902 (.A(n_257_75_22), .ZN(n_257_75_272));
   INV_X1 i_257_75_903 (.A(n_257_75_23), .ZN(n_257_75_273));
   INV_X1 i_257_75_904 (.A(n_257_75_20), .ZN(n_257_75_274));
   INV_X1 i_257_75_905 (.A(n_257_75_21), .ZN(n_257_75_275));
   INV_X1 i_257_75_906 (.A(n_257_75_18), .ZN(n_257_75_276));
   INV_X1 i_257_75_907 (.A(n_257_75_19), .ZN(n_257_75_277));
   INV_X1 i_257_75_908 (.A(n_257_75_16), .ZN(n_257_75_278));
   INV_X1 i_257_75_909 (.A(n_257_75_14), .ZN(n_257_75_279));
   INV_X1 i_257_75_910 (.A(n_257_75_15), .ZN(n_257_75_280));
   INV_X1 i_257_75_911 (.A(n_257_75_5), .ZN(n_257_75_281));
   INV_X1 i_257_75_912 (.A(n_257_75_12), .ZN(n_257_75_282));
   INV_X1 i_257_75_913 (.A(n_257_75_13), .ZN(n_257_75_283));
   INV_X1 i_257_75_914 (.A(n_257_75_10), .ZN(n_257_75_284));
   INV_X1 i_257_75_915 (.A(n_257_75_11), .ZN(n_257_75_285));
   INV_X1 i_257_75_916 (.A(n_257_75_8), .ZN(n_257_75_286));
   INV_X1 i_257_75_917 (.A(n_257_75_4), .ZN(n_257_75_287));
   INV_X1 i_257_75_918 (.A(n_257_75_2), .ZN(n_257_75_288));
   INV_X1 i_257_75_919 (.A(n_257_6), .ZN(n_257_75_289));
   INV_X1 i_257_75_920 (.A(n_257_7), .ZN(n_257_75_290));
   INV_X1 i_257_75_921 (.A(n_257_8), .ZN(n_257_75_291));
   INV_X1 i_257_75_922 (.A(n_257_1), .ZN(n_257_75_292));
   INV_X1 i_257_75_923 (.A(n_257_2), .ZN(n_257_75_293));
   INV_X1 i_257_75_924 (.A(n_151), .ZN(n_257_75_294));
   INV_X1 i_257_75_925 (.A(n_32), .ZN(n_257_75_295));
   INV_X1 i_257_75_926 (.A(PacketSize[1]), .ZN(n_257_1091));
   INV_X1 i_257_75_927 (.A(PacketSize[2]), .ZN(n_257_75_296));
   INV_X1 i_257_75_928 (.A(PacketSize[3]), .ZN(n_257_75_297));
   INV_X1 i_257_75_929 (.A(PacketSize[5]), .ZN(n_257_75_298));
   NAND4_X1 i_257_75_930 (.A1(n_257_75_315), .A2(n_257_75_316), .A3(n_257_75_306), 
      .A4(n_257_75_299), .ZN(n_257_443));
   NOR2_X1 i_257_75_931 (.A1(n_33), .A2(n_32), .ZN(n_257_75_299));
   NAND3_X1 i_257_75_932 (.A1(n_257_75_315), .A2(n_257_75_316), .A3(n_257_75_306), 
      .ZN(n_257_445));
   INV_X1 i_257_75_933 (.A(n_257_75_315), .ZN(n_257_484));
   INV_X1 i_257_75_934 (.A(n_257_75_301), .ZN(n_257_75_300));
   NAND2_X1 i_257_75_935 (.A1(n_257_75_320), .A2(n_257_75_321), .ZN(n_257_75_301));
   INV_X1 i_257_75_936 (.A(n_257_75_309), .ZN(n_257_75_302));
   INV_X1 i_257_75_937 (.A(n_257_75_311), .ZN(n_257_75_303));
   INV_X1 i_257_75_938 (.A(n_257_75_305), .ZN(n_257_75_304));
   NAND2_X1 i_257_75_939 (.A1(n_257_75_315), .A2(n_257_75_316), .ZN(n_257_75_305));
   INV_X1 i_257_75_940 (.A(n_34), .ZN(n_257_75_306));
   INV_X1 i_257_75_941 (.A(n_257_75_320), .ZN(n_257_75_307));
   NAND3_X1 i_257_75_942 (.A1(n_257_75_318), .A2(n_257_75_323), .A3(
      PacketSize[0]), .ZN(n_257_442));
   NAND3_X1 i_257_75_943 (.A1(n_257_75_315), .A2(n_257_75_316), .A3(n_257_75_308), 
      .ZN(n_257_446));
   NAND2_X1 i_257_75_944 (.A1(n_34), .A2(n_257_75_309), .ZN(n_257_75_308));
   NAND3_X1 i_257_75_945 (.A1(n_257_75_314), .A2(n_257_75_313), .A3(n_257_75_312), 
      .ZN(n_257_75_309));
   NAND3_X1 i_257_75_946 (.A1(n_257_75_315), .A2(n_257_75_316), .A3(n_257_75_310), 
      .ZN(n_257_447));
   NAND2_X1 i_257_75_947 (.A1(n_34), .A2(n_257_75_311), .ZN(n_257_75_310));
   OAI21_X1 i_257_75_948 (.A(n_257_75_314), .B1(n_257_75_313), .B2(n_257_75_312), 
      .ZN(n_257_75_311));
   INV_X1 i_257_75_949 (.A(n_151), .ZN(n_257_75_312));
   INV_X1 i_257_75_950 (.A(n_32), .ZN(n_257_75_313));
   INV_X1 i_257_75_951 (.A(n_33), .ZN(n_257_75_314));
   NOR2_X1 i_257_75_952 (.A1(n_36), .A2(n_37), .ZN(n_257_75_315));
   INV_X1 i_257_75_953 (.A(n_35), .ZN(n_257_75_316));
   INV_X1 i_257_75_954 (.A(n_257_75_317), .ZN(n_257_1096));
   NAND2_X1 i_257_75_955 (.A1(n_257_75_318), .A2(n_257_75_323), .ZN(n_257_75_317));
   INV_X1 i_257_75_956 (.A(n_257_75_319), .ZN(n_257_75_318));
   NAND3_X1 i_257_75_957 (.A1(n_257_75_320), .A2(n_257_75_322), .A3(n_257_75_321), 
      .ZN(n_257_75_319));
   NOR2_X1 i_257_75_958 (.A1(PacketSize[2]), .A2(PacketSize[1]), .ZN(
      n_257_75_320));
   INV_X1 i_257_75_959 (.A(PacketSize[3]), .ZN(n_257_75_321));
   INV_X1 i_257_75_960 (.A(PacketSize[4]), .ZN(n_257_75_322));
   INV_X1 i_257_75_961 (.A(PacketSize[5]), .ZN(n_257_75_323));
   NAND2_X1 i_257_76_0 (.A1(n_257_995), .A2(n_257_444), .ZN(n_257_76_0));
   NAND2_X1 i_257_76_1 (.A1(n_257_441), .A2(n_257_963), .ZN(n_257_76_1));
   NOR2_X1 i_257_76_2 (.A1(n_257_1059), .A2(n_257_76_17412), .ZN(n_257_76_2));
   INV_X1 i_257_76_3 (.A(n_257_76_2), .ZN(n_257_76_3));
   INV_X1 i_257_76_4 (.A(n_257_931), .ZN(n_257_76_4));
   NOR2_X1 i_257_76_5 (.A1(n_257_76_3), .A2(n_257_76_4), .ZN(n_257_76_5));
   NAND2_X1 i_257_76_6 (.A1(n_257_440), .A2(n_257_76_5), .ZN(n_257_76_6));
   INV_X1 i_257_76_7 (.A(n_257_76_6), .ZN(n_257_76_7));
   NAND2_X1 i_257_76_8 (.A1(n_257_76_1), .A2(n_257_76_7), .ZN(n_257_76_8));
   INV_X1 i_257_76_9 (.A(n_257_76_8), .ZN(n_257_76_9));
   NAND2_X1 i_257_76_10 (.A1(n_257_76_0), .A2(n_257_76_9), .ZN(n_257_76_10));
   INV_X1 i_257_76_11 (.A(n_257_76_10), .ZN(n_257_76_11));
   NAND2_X1 i_257_76_12 (.A1(n_257_1027), .A2(n_257_443), .ZN(n_257_76_12));
   NAND2_X1 i_257_76_13 (.A1(n_257_76_11), .A2(n_257_76_12), .ZN(n_257_76_13));
   INV_X1 i_257_76_14 (.A(n_257_76_13), .ZN(n_257_76_14));
   NAND2_X1 i_257_76_15 (.A1(n_257_17), .A2(n_257_76_14), .ZN(n_257_76_15));
   NAND2_X1 i_257_76_16 (.A1(n_257_451), .A2(n_257_452), .ZN(n_257_76_16));
   NAND2_X1 i_257_76_17 (.A1(n_257_861), .A2(n_257_445), .ZN(n_257_76_17));
   NAND2_X1 i_257_76_18 (.A1(n_257_76_16), .A2(n_257_76_17), .ZN(n_257_76_18));
   NAND2_X1 i_257_76_19 (.A1(n_257_733), .A2(n_257_436), .ZN(n_257_76_19));
   NAND2_X1 i_257_76_20 (.A1(n_257_797), .A2(n_257_437), .ZN(n_257_76_20));
   NAND3_X1 i_257_76_21 (.A1(n_257_76_19), .A2(n_257_76_20), .A3(n_257_76_1), 
      .ZN(n_257_76_21));
   NOR2_X1 i_257_76_22 (.A1(n_257_76_18), .A2(n_257_76_21), .ZN(n_257_76_22));
   NAND2_X1 i_257_76_23 (.A1(n_257_669), .A2(n_257_448), .ZN(n_257_76_23));
   NAND2_X1 i_257_76_24 (.A1(n_257_629), .A2(n_257_450), .ZN(n_257_76_24));
   NAND2_X1 i_257_76_25 (.A1(n_257_440), .A2(n_257_931), .ZN(n_257_76_25));
   NAND2_X1 i_257_76_26 (.A1(n_257_438), .A2(n_257_1065), .ZN(n_257_76_26));
   NAND3_X1 i_257_76_27 (.A1(n_257_76_24), .A2(n_257_76_25), .A3(n_257_76_26), 
      .ZN(n_257_76_27));
   INV_X1 i_257_76_28 (.A(n_257_76_27), .ZN(n_257_76_28));
   NAND2_X1 i_257_76_29 (.A1(n_257_447), .A2(n_257_765), .ZN(n_257_76_29));
   NAND2_X1 i_257_76_30 (.A1(n_257_439), .A2(n_257_899), .ZN(n_257_76_30));
   NAND2_X1 i_257_76_31 (.A1(n_257_701), .A2(n_257_435), .ZN(n_257_76_31));
   NAND2_X1 i_257_76_32 (.A1(n_257_597), .A2(n_257_442), .ZN(n_257_76_32));
   NOR2_X1 i_257_76_33 (.A1(n_257_76_32), .A2(n_257_1059), .ZN(n_257_76_33));
   NAND2_X1 i_257_76_34 (.A1(n_257_432), .A2(n_257_76_33), .ZN(n_257_76_34));
   INV_X1 i_257_76_35 (.A(n_257_76_34), .ZN(n_257_76_35));
   NAND3_X1 i_257_76_36 (.A1(n_257_76_30), .A2(n_257_76_31), .A3(n_257_76_35), 
      .ZN(n_257_76_36));
   INV_X1 i_257_76_37 (.A(n_257_76_36), .ZN(n_257_76_37));
   NAND3_X1 i_257_76_38 (.A1(n_257_76_28), .A2(n_257_76_29), .A3(n_257_76_37), 
      .ZN(n_257_76_38));
   NAND2_X1 i_257_76_39 (.A1(n_257_35), .A2(n_257_433), .ZN(n_257_76_39));
   NAND2_X1 i_257_76_40 (.A1(n_257_446), .A2(n_257_829), .ZN(n_257_76_40));
   NAND2_X1 i_257_76_41 (.A1(n_257_449), .A2(n_257_1073), .ZN(n_257_76_41));
   NAND3_X1 i_257_76_42 (.A1(n_257_76_39), .A2(n_257_76_40), .A3(n_257_76_41), 
      .ZN(n_257_76_42));
   NOR2_X1 i_257_76_43 (.A1(n_257_76_38), .A2(n_257_76_42), .ZN(n_257_76_43));
   NAND3_X1 i_257_76_44 (.A1(n_257_76_22), .A2(n_257_76_23), .A3(n_257_76_43), 
      .ZN(n_257_76_44));
   INV_X1 i_257_76_45 (.A(n_257_76_44), .ZN(n_257_76_45));
   NAND2_X1 i_257_76_46 (.A1(n_257_76_45), .A2(n_257_76_0), .ZN(n_257_76_46));
   INV_X1 i_257_76_47 (.A(n_257_76_12), .ZN(n_257_76_47));
   NOR2_X1 i_257_76_48 (.A1(n_257_76_46), .A2(n_257_76_47), .ZN(n_257_76_48));
   NAND2_X1 i_257_76_49 (.A1(n_257_68), .A2(n_257_76_48), .ZN(n_257_76_49));
   NAND4_X1 i_257_76_50 (.A1(n_257_76_17), .A2(n_257_76_19), .A3(n_257_76_20), 
      .A4(n_257_76_1), .ZN(n_257_76_50));
   INV_X1 i_257_76_51 (.A(n_257_76_50), .ZN(n_257_76_51));
   NAND2_X1 i_257_76_52 (.A1(n_257_76_40), .A2(n_257_76_41), .ZN(n_257_76_52));
   INV_X1 i_257_76_53 (.A(n_257_76_52), .ZN(n_257_76_53));
   NAND2_X1 i_257_76_54 (.A1(n_257_76_29), .A2(n_257_76_25), .ZN(n_257_76_54));
   INV_X1 i_257_76_55 (.A(n_257_76_54), .ZN(n_257_76_55));
   NAND2_X1 i_257_76_56 (.A1(n_257_76_26), .A2(n_257_76_30), .ZN(n_257_76_56));
   NAND2_X1 i_257_76_57 (.A1(n_257_450), .A2(n_257_76_2), .ZN(n_257_76_57));
   INV_X1 i_257_76_58 (.A(n_257_76_57), .ZN(n_257_76_58));
   NAND3_X1 i_257_76_59 (.A1(n_257_76_31), .A2(n_257_629), .A3(n_257_76_58), 
      .ZN(n_257_76_59));
   NOR2_X1 i_257_76_60 (.A1(n_257_76_56), .A2(n_257_76_59), .ZN(n_257_76_60));
   NAND3_X1 i_257_76_61 (.A1(n_257_76_53), .A2(n_257_76_55), .A3(n_257_76_60), 
      .ZN(n_257_76_61));
   INV_X1 i_257_76_62 (.A(n_257_76_61), .ZN(n_257_76_62));
   NAND2_X1 i_257_76_63 (.A1(n_257_76_51), .A2(n_257_76_62), .ZN(n_257_76_63));
   INV_X1 i_257_76_64 (.A(n_257_76_23), .ZN(n_257_76_64));
   NOR2_X1 i_257_76_65 (.A1(n_257_76_63), .A2(n_257_76_64), .ZN(n_257_76_65));
   NAND2_X1 i_257_76_66 (.A1(n_257_76_0), .A2(n_257_76_65), .ZN(n_257_76_66));
   NOR2_X1 i_257_76_67 (.A1(n_257_76_66), .A2(n_257_76_47), .ZN(n_257_76_67));
   NAND2_X1 i_257_76_68 (.A1(n_257_28), .A2(n_257_76_67), .ZN(n_257_76_68));
   NAND3_X1 i_257_76_69 (.A1(n_257_76_15), .A2(n_257_76_49), .A3(n_257_76_68), 
      .ZN(n_257_76_69));
   INV_X1 i_257_76_70 (.A(n_257_76_25), .ZN(n_257_76_70));
   NAND3_X1 i_257_76_71 (.A1(n_257_439), .A2(n_257_899), .A3(n_257_76_2), 
      .ZN(n_257_76_71));
   NOR2_X1 i_257_76_72 (.A1(n_257_76_70), .A2(n_257_76_71), .ZN(n_257_76_72));
   NAND2_X1 i_257_76_73 (.A1(n_257_76_1), .A2(n_257_76_72), .ZN(n_257_76_73));
   INV_X1 i_257_76_74 (.A(n_257_76_73), .ZN(n_257_76_74));
   NAND2_X1 i_257_76_75 (.A1(n_257_76_0), .A2(n_257_76_74), .ZN(n_257_76_75));
   INV_X1 i_257_76_76 (.A(n_257_76_75), .ZN(n_257_76_76));
   NAND2_X1 i_257_76_77 (.A1(n_257_76_76), .A2(n_257_76_12), .ZN(n_257_76_77));
   INV_X1 i_257_76_78 (.A(n_257_76_77), .ZN(n_257_76_78));
   NAND2_X1 i_257_76_79 (.A1(n_257_18), .A2(n_257_76_78), .ZN(n_257_76_79));
   NAND2_X1 i_257_76_80 (.A1(n_257_829), .A2(n_257_76_2), .ZN(n_257_76_80));
   INV_X1 i_257_76_81 (.A(n_257_76_80), .ZN(n_257_76_81));
   NAND3_X1 i_257_76_82 (.A1(n_257_76_26), .A2(n_257_76_30), .A3(n_257_76_81), 
      .ZN(n_257_76_82));
   NAND2_X1 i_257_76_83 (.A1(n_257_446), .A2(n_257_76_25), .ZN(n_257_76_83));
   NOR2_X1 i_257_76_84 (.A1(n_257_76_82), .A2(n_257_76_83), .ZN(n_257_76_84));
   NAND3_X1 i_257_76_85 (.A1(n_257_76_84), .A2(n_257_76_17), .A3(n_257_76_1), 
      .ZN(n_257_76_85));
   INV_X1 i_257_76_86 (.A(n_257_76_85), .ZN(n_257_76_86));
   NAND2_X1 i_257_76_87 (.A1(n_257_76_0), .A2(n_257_76_86), .ZN(n_257_76_87));
   INV_X1 i_257_76_88 (.A(n_257_76_87), .ZN(n_257_76_88));
   NAND2_X1 i_257_76_89 (.A1(n_257_76_88), .A2(n_257_76_12), .ZN(n_257_76_89));
   INV_X1 i_257_76_90 (.A(n_257_76_89), .ZN(n_257_76_90));
   NAND2_X1 i_257_76_91 (.A1(n_257_21), .A2(n_257_76_90), .ZN(n_257_76_91));
   NAND2_X1 i_257_76_92 (.A1(n_257_113), .A2(n_257_430), .ZN(n_257_76_92));
   NAND3_X1 i_257_76_93 (.A1(n_257_76_16), .A2(n_257_76_17), .A3(n_257_76_92), 
      .ZN(n_257_76_93));
   NAND4_X1 i_257_76_94 (.A1(n_257_76_1), .A2(n_257_76_40), .A3(n_257_76_41), 
      .A4(n_257_76_29), .ZN(n_257_76_94));
   NOR2_X1 i_257_76_95 (.A1(n_257_76_93), .A2(n_257_76_94), .ZN(n_257_76_95));
   NAND2_X1 i_257_76_96 (.A1(n_257_152), .A2(n_257_429), .ZN(n_257_76_96));
   NAND2_X1 i_257_76_97 (.A1(n_257_75), .A2(n_257_431), .ZN(n_257_76_97));
   NAND3_X1 i_257_76_98 (.A1(n_257_76_95), .A2(n_257_76_96), .A3(n_257_76_97), 
      .ZN(n_257_76_98));
   NAND2_X1 i_257_76_99 (.A1(n_257_192), .A2(n_257_427), .ZN(n_257_76_99));
   NAND4_X1 i_257_76_100 (.A1(n_257_76_99), .A2(n_257_76_24), .A3(n_257_76_25), 
      .A4(n_257_76_26), .ZN(n_257_76_100));
   NAND2_X1 i_257_76_101 (.A1(n_257_423), .A2(n_257_76_2), .ZN(n_257_76_101));
   INV_X1 i_257_76_102 (.A(n_257_76_101), .ZN(n_257_76_102));
   NAND2_X1 i_257_76_103 (.A1(n_257_432), .A2(n_257_597), .ZN(n_257_76_103));
   NAND2_X1 i_257_76_104 (.A1(n_257_428), .A2(n_257_565), .ZN(n_257_76_104));
   NAND3_X1 i_257_76_105 (.A1(n_257_76_102), .A2(n_257_76_103), .A3(n_257_76_104), 
      .ZN(n_257_76_105));
   INV_X1 i_257_76_106 (.A(n_257_76_105), .ZN(n_257_76_106));
   NAND2_X1 i_257_76_107 (.A1(n_257_501), .A2(n_257_424), .ZN(n_257_76_107));
   NAND4_X1 i_257_76_108 (.A1(n_257_76_30), .A2(n_257_76_106), .A3(n_257_76_107), 
      .A4(n_257_76_31), .ZN(n_257_76_108));
   NOR2_X1 i_257_76_109 (.A1(n_257_76_100), .A2(n_257_76_108), .ZN(n_257_76_109));
   NAND2_X1 i_257_76_110 (.A1(n_257_76_19), .A2(n_257_76_20), .ZN(n_257_76_110));
   INV_X1 i_257_76_111 (.A(n_257_76_110), .ZN(n_257_76_111));
   NAND2_X1 i_257_76_112 (.A1(n_257_533), .A2(n_257_426), .ZN(n_257_76_112));
   NAND3_X1 i_257_76_113 (.A1(n_257_76_39), .A2(n_257_76_112), .A3(n_257_272), 
      .ZN(n_257_76_113));
   INV_X1 i_257_76_114 (.A(n_257_76_113), .ZN(n_257_76_114));
   NAND3_X1 i_257_76_115 (.A1(n_257_76_109), .A2(n_257_76_111), .A3(n_257_76_114), 
      .ZN(n_257_76_115));
   INV_X1 i_257_76_116 (.A(n_257_76_115), .ZN(n_257_76_116));
   NAND2_X1 i_257_76_117 (.A1(n_257_76_116), .A2(n_257_76_23), .ZN(n_257_76_117));
   NOR2_X1 i_257_76_118 (.A1(n_257_76_98), .A2(n_257_76_117), .ZN(n_257_76_118));
   NAND2_X1 i_257_76_119 (.A1(n_257_232), .A2(n_257_425), .ZN(n_257_76_119));
   NAND2_X1 i_257_76_120 (.A1(n_257_76_119), .A2(n_257_76_0), .ZN(n_257_76_120));
   INV_X1 i_257_76_121 (.A(n_257_76_120), .ZN(n_257_76_121));
   NAND3_X1 i_257_76_122 (.A1(n_257_76_118), .A2(n_257_76_121), .A3(n_257_76_12), 
      .ZN(n_257_76_122));
   INV_X1 i_257_76_123 (.A(n_257_76_122), .ZN(n_257_76_123));
   NAND2_X1 i_257_76_124 (.A1(n_257_304), .A2(n_257_76_123), .ZN(n_257_76_124));
   NAND3_X1 i_257_76_125 (.A1(n_257_76_79), .A2(n_257_76_91), .A3(n_257_76_124), 
      .ZN(n_257_76_125));
   NOR2_X1 i_257_76_126 (.A1(n_257_76_69), .A2(n_257_76_125), .ZN(n_257_76_126));
   NAND2_X1 i_257_76_127 (.A1(n_257_963), .A2(n_257_76_2), .ZN(n_257_76_127));
   INV_X1 i_257_76_128 (.A(n_257_76_127), .ZN(n_257_76_128));
   NAND2_X1 i_257_76_129 (.A1(n_257_441), .A2(n_257_76_128), .ZN(n_257_76_129));
   INV_X1 i_257_76_130 (.A(n_257_76_129), .ZN(n_257_76_130));
   NAND2_X1 i_257_76_131 (.A1(n_257_76_0), .A2(n_257_76_130), .ZN(n_257_76_131));
   INV_X1 i_257_76_132 (.A(n_257_76_131), .ZN(n_257_76_132));
   NAND2_X1 i_257_76_133 (.A1(n_257_76_132), .A2(n_257_76_12), .ZN(n_257_76_133));
   INV_X1 i_257_76_134 (.A(n_257_76_133), .ZN(n_257_76_134));
   NAND2_X1 i_257_76_135 (.A1(n_257_16), .A2(n_257_76_134), .ZN(n_257_76_135));
   NAND3_X1 i_257_76_136 (.A1(n_257_76_17), .A2(n_257_76_19), .A3(n_257_76_20), 
      .ZN(n_257_76_136));
   NAND2_X1 i_257_76_137 (.A1(n_257_76_40), .A2(n_257_76_29), .ZN(n_257_76_137));
   INV_X1 i_257_76_138 (.A(n_257_76_137), .ZN(n_257_76_138));
   NAND2_X1 i_257_76_139 (.A1(n_257_435), .A2(n_257_76_2), .ZN(n_257_76_139));
   INV_X1 i_257_76_140 (.A(n_257_76_139), .ZN(n_257_76_140));
   NAND2_X1 i_257_76_141 (.A1(n_257_701), .A2(n_257_76_140), .ZN(n_257_76_141));
   INV_X1 i_257_76_142 (.A(n_257_76_141), .ZN(n_257_76_142));
   NAND4_X1 i_257_76_143 (.A1(n_257_76_25), .A2(n_257_76_26), .A3(n_257_76_30), 
      .A4(n_257_76_142), .ZN(n_257_76_143));
   INV_X1 i_257_76_144 (.A(n_257_76_143), .ZN(n_257_76_144));
   NAND3_X1 i_257_76_145 (.A1(n_257_76_138), .A2(n_257_76_1), .A3(n_257_76_144), 
      .ZN(n_257_76_145));
   NOR2_X1 i_257_76_146 (.A1(n_257_76_136), .A2(n_257_76_145), .ZN(n_257_76_146));
   NAND2_X1 i_257_76_147 (.A1(n_257_76_0), .A2(n_257_76_146), .ZN(n_257_76_147));
   INV_X1 i_257_76_148 (.A(n_257_76_147), .ZN(n_257_76_148));
   NAND2_X1 i_257_76_149 (.A1(n_257_76_148), .A2(n_257_76_12), .ZN(n_257_76_149));
   INV_X1 i_257_76_150 (.A(n_257_76_149), .ZN(n_257_76_150));
   NAND2_X1 i_257_76_151 (.A1(n_257_25), .A2(n_257_76_150), .ZN(n_257_76_151));
   NAND2_X1 i_257_76_152 (.A1(n_257_442), .A2(n_257_565), .ZN(n_257_76_152));
   NOR2_X1 i_257_76_153 (.A1(n_257_76_152), .A2(n_257_1059), .ZN(n_257_76_153));
   NAND2_X1 i_257_76_154 (.A1(n_257_428), .A2(n_257_76_153), .ZN(n_257_76_154));
   INV_X1 i_257_76_155 (.A(n_257_76_154), .ZN(n_257_76_155));
   NAND2_X1 i_257_76_156 (.A1(n_257_76_155), .A2(n_257_76_103), .ZN(n_257_76_156));
   INV_X1 i_257_76_157 (.A(n_257_76_156), .ZN(n_257_76_157));
   NAND3_X1 i_257_76_158 (.A1(n_257_76_30), .A2(n_257_76_31), .A3(n_257_76_157), 
      .ZN(n_257_76_158));
   INV_X1 i_257_76_159 (.A(n_257_76_158), .ZN(n_257_76_159));
   NAND3_X1 i_257_76_160 (.A1(n_257_76_28), .A2(n_257_76_29), .A3(n_257_76_159), 
      .ZN(n_257_76_160));
   NOR2_X1 i_257_76_161 (.A1(n_257_76_160), .A2(n_257_76_42), .ZN(n_257_76_161));
   INV_X1 i_257_76_162 (.A(n_257_76_93), .ZN(n_257_76_162));
   INV_X1 i_257_76_163 (.A(n_257_76_21), .ZN(n_257_76_163));
   NAND4_X1 i_257_76_164 (.A1(n_257_76_161), .A2(n_257_76_162), .A3(n_257_76_97), 
      .A4(n_257_76_163), .ZN(n_257_76_164));
   NAND2_X1 i_257_76_165 (.A1(n_257_76_23), .A2(n_257_76_96), .ZN(n_257_76_165));
   NOR2_X1 i_257_76_166 (.A1(n_257_76_164), .A2(n_257_76_165), .ZN(n_257_76_166));
   NAND3_X1 i_257_76_167 (.A1(n_257_76_166), .A2(n_257_76_12), .A3(n_257_76_0), 
      .ZN(n_257_76_167));
   INV_X1 i_257_76_168 (.A(n_257_76_167), .ZN(n_257_76_168));
   NAND2_X1 i_257_76_169 (.A1(n_257_185), .A2(n_257_76_168), .ZN(n_257_76_169));
   NAND3_X1 i_257_76_170 (.A1(n_257_76_135), .A2(n_257_76_151), .A3(n_257_76_169), 
      .ZN(n_257_76_170));
   NAND2_X1 i_257_76_171 (.A1(n_257_1059), .A2(n_257_442), .ZN(n_257_76_171));
   INV_X1 i_257_76_172 (.A(n_257_76_171), .ZN(n_257_76_172));
   NAND2_X1 i_257_76_173 (.A1(n_257_13), .A2(n_257_76_172), .ZN(n_257_76_173));
   NAND2_X1 i_257_76_174 (.A1(n_257_445), .A2(n_257_76_2), .ZN(n_257_76_174));
   INV_X1 i_257_76_175 (.A(n_257_76_174), .ZN(n_257_76_175));
   NAND4_X1 i_257_76_176 (.A1(n_257_76_25), .A2(n_257_76_26), .A3(n_257_76_30), 
      .A4(n_257_76_175), .ZN(n_257_76_176));
   INV_X1 i_257_76_177 (.A(n_257_76_176), .ZN(n_257_76_177));
   NAND3_X1 i_257_76_178 (.A1(n_257_76_177), .A2(n_257_76_1), .A3(n_257_861), 
      .ZN(n_257_76_178));
   INV_X1 i_257_76_179 (.A(n_257_76_178), .ZN(n_257_76_179));
   NAND2_X1 i_257_76_180 (.A1(n_257_76_0), .A2(n_257_76_179), .ZN(n_257_76_180));
   INV_X1 i_257_76_181 (.A(n_257_76_180), .ZN(n_257_76_181));
   NAND2_X1 i_257_76_182 (.A1(n_257_76_181), .A2(n_257_76_12), .ZN(n_257_76_182));
   INV_X1 i_257_76_183 (.A(n_257_76_182), .ZN(n_257_76_183));
   NAND2_X1 i_257_76_184 (.A1(n_257_20), .A2(n_257_76_183), .ZN(n_257_76_184));
   NAND2_X1 i_257_76_185 (.A1(n_257_76_173), .A2(n_257_76_184), .ZN(n_257_76_185));
   NOR2_X1 i_257_76_186 (.A1(n_257_76_170), .A2(n_257_76_185), .ZN(n_257_76_186));
   NAND2_X1 i_257_76_187 (.A1(n_257_436), .A2(n_257_76_2), .ZN(n_257_76_187));
   INV_X1 i_257_76_188 (.A(n_257_76_187), .ZN(n_257_76_188));
   NAND4_X1 i_257_76_189 (.A1(n_257_76_25), .A2(n_257_76_26), .A3(n_257_76_30), 
      .A4(n_257_76_188), .ZN(n_257_76_189));
   INV_X1 i_257_76_190 (.A(n_257_76_189), .ZN(n_257_76_190));
   NAND4_X1 i_257_76_191 (.A1(n_257_76_190), .A2(n_257_733), .A3(n_257_76_40), 
      .A4(n_257_76_29), .ZN(n_257_76_191));
   NAND3_X1 i_257_76_192 (.A1(n_257_76_17), .A2(n_257_76_20), .A3(n_257_76_1), 
      .ZN(n_257_76_192));
   NOR2_X1 i_257_76_193 (.A1(n_257_76_191), .A2(n_257_76_192), .ZN(n_257_76_193));
   NAND2_X1 i_257_76_194 (.A1(n_257_76_0), .A2(n_257_76_193), .ZN(n_257_76_194));
   INV_X1 i_257_76_195 (.A(n_257_76_194), .ZN(n_257_76_195));
   NAND2_X1 i_257_76_196 (.A1(n_257_76_195), .A2(n_257_76_12), .ZN(n_257_76_196));
   INV_X1 i_257_76_197 (.A(n_257_76_196), .ZN(n_257_76_197));
   NAND2_X1 i_257_76_198 (.A1(n_257_24), .A2(n_257_76_197), .ZN(n_257_76_198));
   INV_X1 i_257_76_199 (.A(n_257_76_39), .ZN(n_257_76_199));
   NAND2_X1 i_257_76_200 (.A1(n_257_76_99), .A2(n_257_533), .ZN(n_257_76_200));
   NOR2_X1 i_257_76_201 (.A1(n_257_76_199), .A2(n_257_76_200), .ZN(n_257_76_201));
   NAND2_X1 i_257_76_202 (.A1(n_257_426), .A2(n_257_76_2), .ZN(n_257_76_202));
   INV_X1 i_257_76_203 (.A(n_257_76_202), .ZN(n_257_76_203));
   NAND3_X1 i_257_76_204 (.A1(n_257_76_103), .A2(n_257_76_203), .A3(n_257_76_104), 
      .ZN(n_257_76_204));
   INV_X1 i_257_76_205 (.A(n_257_76_204), .ZN(n_257_76_205));
   NAND3_X1 i_257_76_206 (.A1(n_257_76_30), .A2(n_257_76_31), .A3(n_257_76_205), 
      .ZN(n_257_76_206));
   NOR2_X1 i_257_76_207 (.A1(n_257_76_27), .A2(n_257_76_206), .ZN(n_257_76_207));
   NAND4_X1 i_257_76_208 (.A1(n_257_76_201), .A2(n_257_76_207), .A3(n_257_76_19), 
      .A4(n_257_76_20), .ZN(n_257_76_208));
   INV_X1 i_257_76_209 (.A(n_257_76_208), .ZN(n_257_76_209));
   NAND2_X1 i_257_76_210 (.A1(n_257_76_23), .A2(n_257_76_209), .ZN(n_257_76_210));
   NOR2_X1 i_257_76_211 (.A1(n_257_76_98), .A2(n_257_76_210), .ZN(n_257_76_211));
   NAND3_X1 i_257_76_212 (.A1(n_257_76_211), .A2(n_257_76_12), .A3(n_257_76_0), 
      .ZN(n_257_76_212));
   INV_X1 i_257_76_213 (.A(n_257_76_212), .ZN(n_257_76_213));
   NAND2_X1 i_257_76_214 (.A1(n_257_225), .A2(n_257_76_213), .ZN(n_257_76_214));
   NAND2_X1 i_257_76_215 (.A1(n_257_443), .A2(n_257_76_2), .ZN(n_257_76_215));
   INV_X1 i_257_76_216 (.A(n_257_76_215), .ZN(n_257_76_216));
   NAND2_X1 i_257_76_217 (.A1(n_257_1027), .A2(n_257_76_216), .ZN(n_257_76_217));
   INV_X1 i_257_76_218 (.A(n_257_76_217), .ZN(n_257_76_218));
   NAND2_X1 i_257_76_219 (.A1(n_257_14), .A2(n_257_76_218), .ZN(n_257_76_219));
   NAND3_X1 i_257_76_220 (.A1(n_257_76_198), .A2(n_257_76_214), .A3(n_257_76_219), 
      .ZN(n_257_76_220));
   NAND2_X1 i_257_76_221 (.A1(n_257_76_40), .A2(n_257_797), .ZN(n_257_76_221));
   INV_X1 i_257_76_222 (.A(n_257_76_221), .ZN(n_257_76_222));
   NAND2_X1 i_257_76_223 (.A1(n_257_437), .A2(n_257_76_2), .ZN(n_257_76_223));
   INV_X1 i_257_76_224 (.A(n_257_76_223), .ZN(n_257_76_224));
   NAND4_X1 i_257_76_225 (.A1(n_257_76_25), .A2(n_257_76_26), .A3(n_257_76_30), 
      .A4(n_257_76_224), .ZN(n_257_76_225));
   INV_X1 i_257_76_226 (.A(n_257_76_225), .ZN(n_257_76_226));
   NAND4_X1 i_257_76_227 (.A1(n_257_76_222), .A2(n_257_76_17), .A3(n_257_76_1), 
      .A4(n_257_76_226), .ZN(n_257_76_227));
   INV_X1 i_257_76_228 (.A(n_257_76_227), .ZN(n_257_76_228));
   NAND2_X1 i_257_76_229 (.A1(n_257_76_0), .A2(n_257_76_228), .ZN(n_257_76_229));
   INV_X1 i_257_76_230 (.A(n_257_76_229), .ZN(n_257_76_230));
   NAND2_X1 i_257_76_231 (.A1(n_257_76_230), .A2(n_257_76_12), .ZN(n_257_76_231));
   INV_X1 i_257_76_232 (.A(n_257_76_231), .ZN(n_257_76_232));
   NAND2_X1 i_257_76_233 (.A1(n_257_22), .A2(n_257_76_232), .ZN(n_257_76_233));
   NAND2_X1 i_257_76_234 (.A1(n_257_444), .A2(n_257_76_2), .ZN(n_257_76_234));
   INV_X1 i_257_76_235 (.A(n_257_76_234), .ZN(n_257_76_235));
   NAND2_X1 i_257_76_236 (.A1(n_257_995), .A2(n_257_76_235), .ZN(n_257_76_236));
   INV_X1 i_257_76_237 (.A(n_257_76_236), .ZN(n_257_76_237));
   NAND2_X1 i_257_76_238 (.A1(n_257_76_12), .A2(n_257_76_237), .ZN(n_257_76_238));
   INV_X1 i_257_76_239 (.A(n_257_76_238), .ZN(n_257_76_239));
   NAND2_X1 i_257_76_240 (.A1(n_257_15), .A2(n_257_76_239), .ZN(n_257_76_240));
   NAND2_X1 i_257_76_241 (.A1(n_257_76_233), .A2(n_257_76_240), .ZN(n_257_76_241));
   NOR2_X1 i_257_76_242 (.A1(n_257_76_220), .A2(n_257_76_241), .ZN(n_257_76_242));
   NAND3_X1 i_257_76_243 (.A1(n_257_76_126), .A2(n_257_76_186), .A3(n_257_76_242), 
      .ZN(n_257_76_243));
   INV_X1 i_257_76_244 (.A(n_257_76_243), .ZN(n_257_76_244));
   NAND2_X1 i_257_76_245 (.A1(n_257_433), .A2(n_257_76_2), .ZN(n_257_76_245));
   INV_X1 i_257_76_246 (.A(n_257_76_245), .ZN(n_257_76_246));
   NAND3_X1 i_257_76_247 (.A1(n_257_76_30), .A2(n_257_76_31), .A3(n_257_76_246), 
      .ZN(n_257_76_247));
   INV_X1 i_257_76_248 (.A(n_257_76_247), .ZN(n_257_76_248));
   NAND3_X1 i_257_76_249 (.A1(n_257_76_28), .A2(n_257_35), .A3(n_257_76_248), 
      .ZN(n_257_76_249));
   NAND3_X1 i_257_76_250 (.A1(n_257_76_40), .A2(n_257_76_41), .A3(n_257_76_29), 
      .ZN(n_257_76_250));
   NOR2_X1 i_257_76_251 (.A1(n_257_76_249), .A2(n_257_76_250), .ZN(n_257_76_251));
   NAND3_X1 i_257_76_252 (.A1(n_257_76_22), .A2(n_257_76_23), .A3(n_257_76_251), 
      .ZN(n_257_76_252));
   INV_X1 i_257_76_253 (.A(n_257_76_252), .ZN(n_257_76_253));
   NAND2_X1 i_257_76_254 (.A1(n_257_76_253), .A2(n_257_76_0), .ZN(n_257_76_254));
   NOR2_X1 i_257_76_255 (.A1(n_257_76_254), .A2(n_257_76_47), .ZN(n_257_76_255));
   NAND2_X1 i_257_76_256 (.A1(n_257_67), .A2(n_257_76_255), .ZN(n_257_76_256));
   NAND2_X1 i_257_76_257 (.A1(n_257_76_20), .A2(n_257_76_1), .ZN(n_257_76_257));
   INV_X1 i_257_76_258 (.A(n_257_76_257), .ZN(n_257_76_258));
   NAND2_X1 i_257_76_259 (.A1(n_257_431), .A2(n_257_76_2), .ZN(n_257_76_259));
   INV_X1 i_257_76_260 (.A(n_257_76_259), .ZN(n_257_76_260));
   NAND2_X1 i_257_76_261 (.A1(n_257_76_103), .A2(n_257_76_260), .ZN(n_257_76_261));
   INV_X1 i_257_76_262 (.A(n_257_76_261), .ZN(n_257_76_262));
   NAND3_X1 i_257_76_263 (.A1(n_257_76_30), .A2(n_257_76_31), .A3(n_257_76_262), 
      .ZN(n_257_76_263));
   INV_X1 i_257_76_264 (.A(n_257_76_263), .ZN(n_257_76_264));
   NAND3_X1 i_257_76_265 (.A1(n_257_76_28), .A2(n_257_76_29), .A3(n_257_76_264), 
      .ZN(n_257_76_265));
   INV_X1 i_257_76_266 (.A(n_257_76_265), .ZN(n_257_76_266));
   INV_X1 i_257_76_267 (.A(n_257_76_42), .ZN(n_257_76_267));
   NAND3_X1 i_257_76_268 (.A1(n_257_76_258), .A2(n_257_76_266), .A3(n_257_76_267), 
      .ZN(n_257_76_268));
   NAND4_X1 i_257_76_269 (.A1(n_257_75), .A2(n_257_76_16), .A3(n_257_76_17), 
      .A4(n_257_76_19), .ZN(n_257_76_269));
   NOR2_X1 i_257_76_270 (.A1(n_257_76_268), .A2(n_257_76_269), .ZN(n_257_76_270));
   NAND3_X1 i_257_76_271 (.A1(n_257_76_270), .A2(n_257_76_0), .A3(n_257_76_23), 
      .ZN(n_257_76_271));
   NOR2_X1 i_257_76_272 (.A1(n_257_76_47), .A2(n_257_76_271), .ZN(n_257_76_272));
   NAND2_X1 i_257_76_273 (.A1(n_257_107), .A2(n_257_76_272), .ZN(n_257_76_273));
   NAND2_X1 i_257_76_274 (.A1(n_257_76_97), .A2(n_257_152), .ZN(n_257_76_274));
   INV_X1 i_257_76_275 (.A(n_257_76_274), .ZN(n_257_76_275));
   NAND3_X1 i_257_76_276 (.A1(n_257_76_92), .A2(n_257_76_19), .A3(n_257_76_20), 
      .ZN(n_257_76_276));
   NOR2_X1 i_257_76_277 (.A1(n_257_76_276), .A2(n_257_76_18), .ZN(n_257_76_277));
   NAND2_X1 i_257_76_278 (.A1(n_257_429), .A2(n_257_76_2), .ZN(n_257_76_278));
   INV_X1 i_257_76_279 (.A(n_257_76_278), .ZN(n_257_76_279));
   NAND2_X1 i_257_76_280 (.A1(n_257_76_279), .A2(n_257_76_103), .ZN(n_257_76_280));
   INV_X1 i_257_76_281 (.A(n_257_76_280), .ZN(n_257_76_281));
   NAND3_X1 i_257_76_282 (.A1(n_257_76_30), .A2(n_257_76_31), .A3(n_257_76_281), 
      .ZN(n_257_76_282));
   INV_X1 i_257_76_283 (.A(n_257_76_282), .ZN(n_257_76_283));
   NAND4_X1 i_257_76_284 (.A1(n_257_76_28), .A2(n_257_76_283), .A3(n_257_76_41), 
      .A4(n_257_76_29), .ZN(n_257_76_284));
   NAND3_X1 i_257_76_285 (.A1(n_257_76_1), .A2(n_257_76_39), .A3(n_257_76_40), 
      .ZN(n_257_76_285));
   NOR2_X1 i_257_76_286 (.A1(n_257_76_284), .A2(n_257_76_285), .ZN(n_257_76_286));
   NAND4_X1 i_257_76_287 (.A1(n_257_76_275), .A2(n_257_76_277), .A3(n_257_76_286), 
      .A4(n_257_76_23), .ZN(n_257_76_287));
   INV_X1 i_257_76_288 (.A(n_257_76_287), .ZN(n_257_76_288));
   NAND3_X1 i_257_76_289 (.A1(n_257_76_288), .A2(n_257_76_12), .A3(n_257_76_0), 
      .ZN(n_257_76_289));
   INV_X1 i_257_76_290 (.A(n_257_76_289), .ZN(n_257_76_290));
   NAND2_X1 i_257_76_291 (.A1(n_257_184), .A2(n_257_76_290), .ZN(n_257_76_291));
   NAND3_X1 i_257_76_292 (.A1(n_257_76_256), .A2(n_257_76_273), .A3(n_257_76_291), 
      .ZN(n_257_76_292));
   INV_X1 i_257_76_293 (.A(n_257_76_292), .ZN(n_257_76_293));
   NOR2_X1 i_257_76_294 (.A1(n_257_76_3), .A2(n_257_76_3603), .ZN(n_257_76_294));
   NAND2_X1 i_257_76_295 (.A1(n_257_438), .A2(n_257_76_294), .ZN(n_257_76_295));
   INV_X1 i_257_76_296 (.A(n_257_76_295), .ZN(n_257_76_296));
   NAND3_X1 i_257_76_297 (.A1(n_257_76_296), .A2(n_257_76_25), .A3(n_257_76_30), 
      .ZN(n_257_76_297));
   INV_X1 i_257_76_298 (.A(n_257_76_297), .ZN(n_257_76_298));
   NAND2_X1 i_257_76_299 (.A1(n_257_76_1), .A2(n_257_76_298), .ZN(n_257_76_299));
   INV_X1 i_257_76_300 (.A(n_257_76_299), .ZN(n_257_76_300));
   NAND2_X1 i_257_76_301 (.A1(n_257_76_0), .A2(n_257_76_300), .ZN(n_257_76_301));
   INV_X1 i_257_76_302 (.A(n_257_76_301), .ZN(n_257_76_302));
   NAND2_X1 i_257_76_303 (.A1(n_257_76_302), .A2(n_257_76_12), .ZN(n_257_76_303));
   INV_X1 i_257_76_304 (.A(n_257_76_303), .ZN(n_257_76_304));
   NAND2_X1 i_257_76_305 (.A1(n_257_19), .A2(n_257_76_304), .ZN(n_257_76_305));
   NAND4_X1 i_257_76_306 (.A1(n_257_76_16), .A2(n_257_76_17), .A3(n_257_76_92), 
      .A4(n_257_76_19), .ZN(n_257_76_306));
   INV_X1 i_257_76_307 (.A(n_257_76_306), .ZN(n_257_76_307));
   NAND2_X1 i_257_76_308 (.A1(n_257_310), .A2(n_257_422), .ZN(n_257_76_308));
   NAND2_X1 i_257_76_309 (.A1(n_257_76_308), .A2(n_257_76_24), .ZN(n_257_76_309));
   INV_X1 i_257_76_310 (.A(n_257_76_309), .ZN(n_257_76_310));
   INV_X1 i_257_76_311 (.A(n_257_1059), .ZN(n_257_76_311));
   INV_X1 i_257_76_312 (.A(n_257_565), .ZN(n_257_76_312));
   NAND3_X1 i_257_76_313 (.A1(n_257_76_311), .A2(n_257_76_312), .A3(n_257_442), 
      .ZN(n_257_76_313));
   OAI21_X1 i_257_76_314 (.A(n_257_76_313), .B1(n_257_428), .B2(n_257_76_3), 
      .ZN(n_257_76_314));
   NAND3_X1 i_257_76_315 (.A1(n_257_76_314), .A2(n_257_420), .A3(n_257_76_103), 
      .ZN(n_257_76_315));
   INV_X1 i_257_76_316 (.A(n_257_76_315), .ZN(n_257_76_316));
   NAND3_X1 i_257_76_317 (.A1(n_257_76_25), .A2(n_257_76_26), .A3(n_257_76_316), 
      .ZN(n_257_76_317));
   INV_X1 i_257_76_318 (.A(n_257_76_317), .ZN(n_257_76_318));
   NAND4_X1 i_257_76_319 (.A1(n_257_76_30), .A2(n_257_76_107), .A3(n_257_76_31), 
      .A4(n_257_1089), .ZN(n_257_76_319));
   INV_X1 i_257_76_320 (.A(n_257_76_319), .ZN(n_257_76_320));
   NAND3_X1 i_257_76_321 (.A1(n_257_76_310), .A2(n_257_76_318), .A3(n_257_76_320), 
      .ZN(n_257_76_321));
   NAND4_X1 i_257_76_322 (.A1(n_257_76_40), .A2(n_257_76_41), .A3(n_257_76_29), 
      .A4(n_257_76_99), .ZN(n_257_76_322));
   NOR2_X1 i_257_76_323 (.A1(n_257_76_321), .A2(n_257_76_322), .ZN(n_257_76_323));
   NAND3_X1 i_257_76_324 (.A1(n_257_76_1), .A2(n_257_76_39), .A3(n_257_76_112), 
      .ZN(n_257_76_324));
   NAND2_X1 i_257_76_325 (.A1(n_257_272), .A2(n_257_423), .ZN(n_257_76_325));
   NAND2_X1 i_257_76_326 (.A1(n_257_76_325), .A2(n_257_76_20), .ZN(n_257_76_326));
   NOR2_X1 i_257_76_327 (.A1(n_257_76_324), .A2(n_257_76_326), .ZN(n_257_76_327));
   NAND4_X1 i_257_76_328 (.A1(n_257_76_307), .A2(n_257_76_323), .A3(n_257_76_327), 
      .A4(n_257_76_97), .ZN(n_257_76_328));
   NAND2_X1 i_257_76_329 (.A1(n_257_349), .A2(n_257_421), .ZN(n_257_76_329));
   NAND3_X1 i_257_76_330 (.A1(n_257_76_23), .A2(n_257_76_96), .A3(n_257_76_329), 
      .ZN(n_257_76_330));
   NOR2_X1 i_257_76_331 (.A1(n_257_76_328), .A2(n_257_76_330), .ZN(n_257_76_331));
   NAND3_X1 i_257_76_332 (.A1(n_257_76_331), .A2(n_257_76_121), .A3(n_257_76_12), 
      .ZN(n_257_76_332));
   INV_X1 i_257_76_333 (.A(n_257_76_332), .ZN(n_257_76_333));
   NAND2_X1 i_257_76_334 (.A1(n_257_382), .A2(n_257_76_333), .ZN(n_257_76_334));
   NAND3_X1 i_257_76_335 (.A1(n_257_76_16), .A2(n_257_76_17), .A3(n_257_76_19), 
      .ZN(n_257_76_335));
   INV_X1 i_257_76_336 (.A(n_257_76_335), .ZN(n_257_76_336));
   NAND4_X1 i_257_76_337 (.A1(n_257_76_20), .A2(n_257_76_1), .A3(n_257_76_39), 
      .A4(n_257_113), .ZN(n_257_76_337));
   INV_X1 i_257_76_338 (.A(n_257_76_337), .ZN(n_257_76_338));
   NAND2_X1 i_257_76_339 (.A1(n_257_76_24), .A2(n_257_76_25), .ZN(n_257_76_339));
   INV_X1 i_257_76_340 (.A(n_257_76_339), .ZN(n_257_76_340));
   INV_X1 i_257_76_341 (.A(n_257_76_56), .ZN(n_257_76_341));
   NAND2_X1 i_257_76_342 (.A1(n_257_430), .A2(n_257_76_2), .ZN(n_257_76_342));
   INV_X1 i_257_76_343 (.A(n_257_76_342), .ZN(n_257_76_343));
   NAND2_X1 i_257_76_344 (.A1(n_257_76_103), .A2(n_257_76_343), .ZN(n_257_76_344));
   INV_X1 i_257_76_345 (.A(n_257_76_344), .ZN(n_257_76_345));
   NAND2_X1 i_257_76_346 (.A1(n_257_76_31), .A2(n_257_76_345), .ZN(n_257_76_346));
   INV_X1 i_257_76_347 (.A(n_257_76_346), .ZN(n_257_76_347));
   NAND3_X1 i_257_76_348 (.A1(n_257_76_340), .A2(n_257_76_341), .A3(n_257_76_347), 
      .ZN(n_257_76_348));
   NOR2_X1 i_257_76_349 (.A1(n_257_76_348), .A2(n_257_76_250), .ZN(n_257_76_349));
   NAND4_X1 i_257_76_350 (.A1(n_257_76_336), .A2(n_257_76_97), .A3(n_257_76_338), 
      .A4(n_257_76_349), .ZN(n_257_76_350));
   INV_X1 i_257_76_351 (.A(n_257_76_350), .ZN(n_257_76_351));
   NAND3_X1 i_257_76_352 (.A1(n_257_76_351), .A2(n_257_76_0), .A3(n_257_76_23), 
      .ZN(n_257_76_352));
   NOR2_X1 i_257_76_353 (.A1(n_257_76_352), .A2(n_257_76_47), .ZN(n_257_76_353));
   NAND2_X1 i_257_76_354 (.A1(n_257_145), .A2(n_257_76_353), .ZN(n_257_76_354));
   NAND3_X1 i_257_76_355 (.A1(n_257_76_305), .A2(n_257_76_334), .A3(n_257_76_354), 
      .ZN(n_257_76_355));
   INV_X1 i_257_76_356 (.A(n_257_76_355), .ZN(n_257_76_356));
   NAND3_X1 i_257_76_357 (.A1(n_257_447), .A2(n_257_76_25), .A3(n_257_76_26), 
      .ZN(n_257_76_357));
   INV_X1 i_257_76_358 (.A(n_257_76_357), .ZN(n_257_76_358));
   INV_X1 i_257_76_359 (.A(n_257_765), .ZN(n_257_76_359));
   NOR2_X1 i_257_76_360 (.A1(n_257_76_3), .A2(n_257_76_359), .ZN(n_257_76_360));
   NAND2_X1 i_257_76_361 (.A1(n_257_76_30), .A2(n_257_76_360), .ZN(n_257_76_361));
   INV_X1 i_257_76_362 (.A(n_257_76_361), .ZN(n_257_76_362));
   NAND4_X1 i_257_76_363 (.A1(n_257_76_1), .A2(n_257_76_358), .A3(n_257_76_40), 
      .A4(n_257_76_362), .ZN(n_257_76_363));
   NAND2_X1 i_257_76_364 (.A1(n_257_76_17), .A2(n_257_76_20), .ZN(n_257_76_364));
   NOR2_X1 i_257_76_365 (.A1(n_257_76_363), .A2(n_257_76_364), .ZN(n_257_76_365));
   NAND2_X1 i_257_76_366 (.A1(n_257_76_0), .A2(n_257_76_365), .ZN(n_257_76_366));
   INV_X1 i_257_76_367 (.A(n_257_76_366), .ZN(n_257_76_367));
   NAND2_X1 i_257_76_368 (.A1(n_257_76_367), .A2(n_257_76_12), .ZN(n_257_76_368));
   INV_X1 i_257_76_369 (.A(n_257_76_368), .ZN(n_257_76_369));
   NAND3_X1 i_257_76_370 (.A1(n_257_449), .A2(n_257_76_25), .A3(n_257_76_26), 
      .ZN(n_257_76_370));
   NAND2_X1 i_257_76_371 (.A1(n_257_1073), .A2(n_257_76_2), .ZN(n_257_76_371));
   INV_X1 i_257_76_372 (.A(n_257_76_371), .ZN(n_257_76_372));
   NAND3_X1 i_257_76_373 (.A1(n_257_76_30), .A2(n_257_76_372), .A3(n_257_76_31), 
      .ZN(n_257_76_373));
   NOR2_X1 i_257_76_374 (.A1(n_257_76_370), .A2(n_257_76_373), .ZN(n_257_76_374));
   NAND3_X1 i_257_76_375 (.A1(n_257_76_374), .A2(n_257_76_138), .A3(n_257_76_1), 
      .ZN(n_257_76_375));
   INV_X1 i_257_76_376 (.A(n_257_76_375), .ZN(n_257_76_376));
   INV_X1 i_257_76_377 (.A(n_257_76_136), .ZN(n_257_76_377));
   NAND2_X1 i_257_76_378 (.A1(n_257_76_376), .A2(n_257_76_377), .ZN(n_257_76_378));
   NOR2_X1 i_257_76_379 (.A1(n_257_76_378), .A2(n_257_76_64), .ZN(n_257_76_379));
   NAND2_X1 i_257_76_380 (.A1(n_257_76_0), .A2(n_257_76_379), .ZN(n_257_76_380));
   NOR2_X1 i_257_76_381 (.A1(n_257_76_380), .A2(n_257_76_47), .ZN(n_257_76_381));
   AOI22_X1 i_257_76_382 (.A1(n_257_23), .A2(n_257_76_369), .B1(n_257_27), 
      .B2(n_257_76_381), .ZN(n_257_76_382));
   NAND3_X1 i_257_76_383 (.A1(n_257_76_293), .A2(n_257_76_356), .A3(n_257_76_382), 
      .ZN(n_257_76_383));
   NAND3_X1 i_257_76_384 (.A1(n_257_76_26), .A2(n_257_448), .A3(n_257_76_30), 
      .ZN(n_257_76_384));
   NAND2_X1 i_257_76_385 (.A1(n_257_76_17760), .A2(n_257_76_2), .ZN(n_257_76_385));
   OAI21_X1 i_257_76_386 (.A(n_257_76_385), .B1(n_257_701), .B2(n_257_76_3), 
      .ZN(n_257_76_386));
   NAND2_X1 i_257_76_387 (.A1(n_257_76_25), .A2(n_257_76_386), .ZN(n_257_76_387));
   NOR2_X1 i_257_76_388 (.A1(n_257_76_384), .A2(n_257_76_387), .ZN(n_257_76_388));
   NAND3_X1 i_257_76_389 (.A1(n_257_76_388), .A2(n_257_76_138), .A3(n_257_76_1), 
      .ZN(n_257_76_389));
   INV_X1 i_257_76_390 (.A(n_257_76_389), .ZN(n_257_76_390));
   NAND3_X1 i_257_76_391 (.A1(n_257_76_390), .A2(n_257_669), .A3(n_257_76_377), 
      .ZN(n_257_76_391));
   INV_X1 i_257_76_392 (.A(n_257_76_391), .ZN(n_257_76_392));
   NAND2_X1 i_257_76_393 (.A1(n_257_76_0), .A2(n_257_76_392), .ZN(n_257_76_393));
   NOR2_X1 i_257_76_394 (.A1(n_257_76_47), .A2(n_257_76_393), .ZN(n_257_76_394));
   NAND2_X1 i_257_76_395 (.A1(n_257_26), .A2(n_257_76_394), .ZN(n_257_76_395));
   NAND2_X1 i_257_76_396 (.A1(n_257_425), .A2(n_257_76_2), .ZN(n_257_76_396));
   INV_X1 i_257_76_397 (.A(n_257_76_396), .ZN(n_257_76_397));
   NAND3_X1 i_257_76_398 (.A1(n_257_76_397), .A2(n_257_76_103), .A3(n_257_76_104), 
      .ZN(n_257_76_398));
   INV_X1 i_257_76_399 (.A(n_257_76_398), .ZN(n_257_76_399));
   NAND3_X1 i_257_76_400 (.A1(n_257_76_30), .A2(n_257_76_31), .A3(n_257_76_399), 
      .ZN(n_257_76_400));
   INV_X1 i_257_76_401 (.A(n_257_76_400), .ZN(n_257_76_401));
   NAND4_X1 i_257_76_402 (.A1(n_257_76_28), .A2(n_257_76_401), .A3(n_257_76_29), 
      .A4(n_257_76_99), .ZN(n_257_76_402));
   NAND4_X1 i_257_76_403 (.A1(n_257_76_39), .A2(n_257_76_112), .A3(n_257_76_40), 
      .A4(n_257_76_41), .ZN(n_257_76_403));
   NOR2_X1 i_257_76_404 (.A1(n_257_76_402), .A2(n_257_76_403), .ZN(n_257_76_404));
   NAND4_X1 i_257_76_405 (.A1(n_257_76_404), .A2(n_257_76_162), .A3(n_257_76_97), 
      .A4(n_257_76_163), .ZN(n_257_76_405));
   INV_X1 i_257_76_406 (.A(n_257_76_405), .ZN(n_257_76_406));
   INV_X1 i_257_76_407 (.A(n_257_76_165), .ZN(n_257_76_407));
   NAND3_X1 i_257_76_408 (.A1(n_257_76_406), .A2(n_257_76_407), .A3(n_257_232), 
      .ZN(n_257_76_408));
   NAND2_X1 i_257_76_409 (.A1(n_257_76_12), .A2(n_257_76_0), .ZN(n_257_76_409));
   NOR2_X1 i_257_76_410 (.A1(n_257_76_408), .A2(n_257_76_409), .ZN(n_257_76_410));
   NAND2_X1 i_257_76_411 (.A1(n_257_264), .A2(n_257_76_410), .ZN(n_257_76_411));
   NAND4_X1 i_257_76_412 (.A1(n_257_76_308), .A2(n_257_76_24), .A3(n_257_76_25), 
      .A4(n_257_76_26), .ZN(n_257_76_412));
   NAND2_X1 i_257_76_413 (.A1(n_257_421), .A2(n_257_76_2), .ZN(n_257_76_413));
   INV_X1 i_257_76_414 (.A(n_257_76_413), .ZN(n_257_76_414));
   NAND3_X1 i_257_76_415 (.A1(n_257_76_414), .A2(n_257_76_103), .A3(n_257_76_104), 
      .ZN(n_257_76_415));
   INV_X1 i_257_76_416 (.A(n_257_76_415), .ZN(n_257_76_416));
   NAND4_X1 i_257_76_417 (.A1(n_257_76_30), .A2(n_257_76_416), .A3(n_257_76_107), 
      .A4(n_257_76_31), .ZN(n_257_76_417));
   NOR2_X1 i_257_76_418 (.A1(n_257_76_412), .A2(n_257_76_417), .ZN(n_257_76_418));
   NAND3_X1 i_257_76_419 (.A1(n_257_76_39), .A2(n_257_76_112), .A3(n_257_76_40), 
      .ZN(n_257_76_419));
   INV_X1 i_257_76_420 (.A(n_257_76_419), .ZN(n_257_76_420));
   NAND3_X1 i_257_76_421 (.A1(n_257_76_41), .A2(n_257_76_29), .A3(n_257_76_99), 
      .ZN(n_257_76_421));
   INV_X1 i_257_76_422 (.A(n_257_76_421), .ZN(n_257_76_422));
   NAND3_X1 i_257_76_423 (.A1(n_257_76_418), .A2(n_257_76_420), .A3(n_257_76_422), 
      .ZN(n_257_76_423));
   NAND4_X1 i_257_76_424 (.A1(n_257_76_19), .A2(n_257_76_325), .A3(n_257_76_20), 
      .A4(n_257_76_1), .ZN(n_257_76_424));
   NOR2_X1 i_257_76_425 (.A1(n_257_76_423), .A2(n_257_76_424), .ZN(n_257_76_425));
   NAND3_X1 i_257_76_426 (.A1(n_257_76_162), .A2(n_257_76_97), .A3(n_257_349), 
      .ZN(n_257_76_426));
   INV_X1 i_257_76_427 (.A(n_257_76_426), .ZN(n_257_76_427));
   NAND4_X1 i_257_76_428 (.A1(n_257_76_425), .A2(n_257_76_427), .A3(n_257_76_23), 
      .A4(n_257_76_96), .ZN(n_257_76_428));
   INV_X1 i_257_76_429 (.A(n_257_76_428), .ZN(n_257_76_429));
   NAND3_X1 i_257_76_430 (.A1(n_257_76_429), .A2(n_257_76_121), .A3(n_257_76_12), 
      .ZN(n_257_76_430));
   INV_X1 i_257_76_431 (.A(n_257_76_430), .ZN(n_257_76_431));
   NAND2_X1 i_257_76_432 (.A1(n_257_381), .A2(n_257_76_431), .ZN(n_257_76_432));
   NAND3_X1 i_257_76_433 (.A1(n_257_76_395), .A2(n_257_76_411), .A3(n_257_76_432), 
      .ZN(n_257_76_433));
   INV_X1 i_257_76_434 (.A(n_257_76_433), .ZN(n_257_76_434));
   NAND4_X1 i_257_76_435 (.A1(n_257_76_39), .A2(n_257_76_40), .A3(n_257_76_41), 
      .A4(n_257_76_29), .ZN(n_257_76_435));
   NAND2_X1 i_257_76_436 (.A1(n_257_76_314), .A2(n_257_76_103), .ZN(n_257_76_436));
   INV_X1 i_257_76_437 (.A(n_257_76_436), .ZN(n_257_76_437));
   NAND3_X1 i_257_76_438 (.A1(n_257_76_26), .A2(n_257_76_30), .A3(n_257_76_437), 
      .ZN(n_257_76_438));
   INV_X1 i_257_76_439 (.A(n_257_76_438), .ZN(n_257_76_439));
   NAND3_X1 i_257_76_440 (.A1(n_257_192), .A2(n_257_76_31), .A3(n_257_427), 
      .ZN(n_257_76_440));
   INV_X1 i_257_76_441 (.A(n_257_76_440), .ZN(n_257_76_441));
   NAND3_X1 i_257_76_442 (.A1(n_257_76_439), .A2(n_257_76_340), .A3(n_257_76_441), 
      .ZN(n_257_76_442));
   NOR2_X1 i_257_76_443 (.A1(n_257_76_435), .A2(n_257_76_442), .ZN(n_257_76_443));
   NAND4_X1 i_257_76_444 (.A1(n_257_76_443), .A2(n_257_76_162), .A3(n_257_76_97), 
      .A4(n_257_76_163), .ZN(n_257_76_444));
   NOR2_X1 i_257_76_445 (.A1(n_257_76_444), .A2(n_257_76_165), .ZN(n_257_76_445));
   NAND3_X1 i_257_76_446 (.A1(n_257_76_445), .A2(n_257_76_12), .A3(n_257_76_0), 
      .ZN(n_257_76_446));
   INV_X1 i_257_76_447 (.A(n_257_76_446), .ZN(n_257_76_447));
   NAND2_X1 i_257_76_448 (.A1(n_257_224), .A2(n_257_76_447), .ZN(n_257_76_448));
   NAND2_X1 i_257_76_449 (.A1(n_257_452), .A2(n_257_76_2), .ZN(n_257_76_449));
   INV_X1 i_257_76_450 (.A(n_257_76_449), .ZN(n_257_76_450));
   NAND2_X1 i_257_76_451 (.A1(n_257_76_450), .A2(n_257_76_31), .ZN(n_257_76_451));
   INV_X1 i_257_76_452 (.A(n_257_76_451), .ZN(n_257_76_452));
   NAND3_X1 i_257_76_453 (.A1(n_257_76_340), .A2(n_257_76_341), .A3(n_257_76_452), 
      .ZN(n_257_76_453));
   NOR2_X1 i_257_76_454 (.A1(n_257_76_453), .A2(n_257_76_250), .ZN(n_257_76_454));
   NAND2_X1 i_257_76_455 (.A1(n_257_76_17), .A2(n_257_76_19), .ZN(n_257_76_455));
   INV_X1 i_257_76_456 (.A(n_257_76_455), .ZN(n_257_76_456));
   NAND3_X1 i_257_76_457 (.A1(n_257_76_20), .A2(n_257_76_1), .A3(n_257_451), 
      .ZN(n_257_76_457));
   INV_X1 i_257_76_458 (.A(n_257_76_457), .ZN(n_257_76_458));
   NAND3_X1 i_257_76_459 (.A1(n_257_76_454), .A2(n_257_76_456), .A3(n_257_76_458), 
      .ZN(n_257_76_459));
   NOR2_X1 i_257_76_460 (.A1(n_257_76_459), .A2(n_257_76_64), .ZN(n_257_76_460));
   NAND2_X1 i_257_76_461 (.A1(n_257_76_460), .A2(n_257_76_0), .ZN(n_257_76_461));
   NOR2_X1 i_257_76_462 (.A1(n_257_76_461), .A2(n_257_76_47), .ZN(n_257_76_462));
   NAND2_X1 i_257_76_463 (.A1(n_257_434), .A2(n_257_76_462), .ZN(n_257_76_463));
   NOR2_X1 i_257_76_464 (.A1(n_257_76_324), .A2(n_257_76_110), .ZN(n_257_76_464));
   NAND3_X1 i_257_76_465 (.A1(n_257_76_314), .A2(n_257_76_103), .A3(n_257_424), 
      .ZN(n_257_76_465));
   INV_X1 i_257_76_466 (.A(n_257_76_465), .ZN(n_257_76_466));
   NAND2_X1 i_257_76_467 (.A1(n_257_76_24), .A2(n_257_76_466), .ZN(n_257_76_467));
   INV_X1 i_257_76_468 (.A(n_257_76_467), .ZN(n_257_76_468));
   NAND2_X1 i_257_76_469 (.A1(n_257_76_25), .A2(n_257_76_26), .ZN(n_257_76_469));
   INV_X1 i_257_76_470 (.A(n_257_76_469), .ZN(n_257_76_470));
   NAND3_X1 i_257_76_471 (.A1(n_257_76_30), .A2(n_257_76_31), .A3(n_257_501), 
      .ZN(n_257_76_471));
   INV_X1 i_257_76_472 (.A(n_257_76_471), .ZN(n_257_76_472));
   NAND3_X1 i_257_76_473 (.A1(n_257_76_468), .A2(n_257_76_470), .A3(n_257_76_472), 
      .ZN(n_257_76_473));
   NOR2_X1 i_257_76_474 (.A1(n_257_76_322), .A2(n_257_76_473), .ZN(n_257_76_474));
   NAND4_X1 i_257_76_475 (.A1(n_257_76_464), .A2(n_257_76_474), .A3(n_257_76_162), 
      .A4(n_257_76_97), .ZN(n_257_76_475));
   NOR2_X1 i_257_76_476 (.A1(n_257_76_475), .A2(n_257_76_165), .ZN(n_257_76_476));
   NAND4_X1 i_257_76_477 (.A1(n_257_76_476), .A2(n_257_76_12), .A3(n_257_76_119), 
      .A4(n_257_76_0), .ZN(n_257_76_477));
   INV_X1 i_257_76_478 (.A(n_257_76_477), .ZN(n_257_76_478));
   NAND2_X1 i_257_76_479 (.A1(n_257_265), .A2(n_257_76_478), .ZN(n_257_76_479));
   NAND3_X1 i_257_76_480 (.A1(n_257_76_448), .A2(n_257_76_463), .A3(n_257_76_479), 
      .ZN(n_257_76_480));
   INV_X1 i_257_76_481 (.A(n_257_76_480), .ZN(n_257_76_481));
   NAND3_X1 i_257_76_482 (.A1(n_257_76_314), .A2(n_257_76_103), .A3(n_257_422), 
      .ZN(n_257_76_482));
   INV_X1 i_257_76_483 (.A(n_257_76_482), .ZN(n_257_76_483));
   NAND4_X1 i_257_76_484 (.A1(n_257_76_483), .A2(n_257_76_107), .A3(n_257_76_31), 
      .A4(n_257_310), .ZN(n_257_76_484));
   INV_X1 i_257_76_485 (.A(n_257_76_484), .ZN(n_257_76_485));
   NAND2_X1 i_257_76_486 (.A1(n_257_76_99), .A2(n_257_76_24), .ZN(n_257_76_486));
   INV_X1 i_257_76_487 (.A(n_257_76_486), .ZN(n_257_76_487));
   NAND3_X1 i_257_76_488 (.A1(n_257_76_25), .A2(n_257_76_26), .A3(n_257_76_30), 
      .ZN(n_257_76_488));
   INV_X1 i_257_76_489 (.A(n_257_76_488), .ZN(n_257_76_489));
   NAND3_X1 i_257_76_490 (.A1(n_257_76_485), .A2(n_257_76_487), .A3(n_257_76_489), 
      .ZN(n_257_76_490));
   NAND4_X1 i_257_76_491 (.A1(n_257_76_112), .A2(n_257_76_40), .A3(n_257_76_41), 
      .A4(n_257_76_29), .ZN(n_257_76_491));
   NOR2_X1 i_257_76_492 (.A1(n_257_76_490), .A2(n_257_76_491), .ZN(n_257_76_492));
   NAND3_X1 i_257_76_493 (.A1(n_257_76_20), .A2(n_257_76_1), .A3(n_257_76_39), 
      .ZN(n_257_76_493));
   NAND2_X1 i_257_76_494 (.A1(n_257_76_19), .A2(n_257_76_325), .ZN(n_257_76_494));
   NOR2_X1 i_257_76_495 (.A1(n_257_76_493), .A2(n_257_76_494), .ZN(n_257_76_495));
   NAND4_X1 i_257_76_496 (.A1(n_257_76_492), .A2(n_257_76_495), .A3(n_257_76_162), 
      .A4(n_257_76_97), .ZN(n_257_76_496));
   NOR2_X1 i_257_76_497 (.A1(n_257_76_496), .A2(n_257_76_165), .ZN(n_257_76_497));
   NAND4_X1 i_257_76_498 (.A1(n_257_76_497), .A2(n_257_76_12), .A3(n_257_76_119), 
      .A4(n_257_76_0), .ZN(n_257_76_498));
   INV_X1 i_257_76_499 (.A(n_257_76_498), .ZN(n_257_76_499));
   NAND2_X1 i_257_76_500 (.A1(n_257_342), .A2(n_257_76_499), .ZN(n_257_76_500));
   NAND2_X1 i_257_76_501 (.A1(n_257_452), .A2(n_257_442), .ZN(n_257_76_501));
   INV_X1 i_257_76_502 (.A(n_257_76_501), .ZN(n_257_76_502));
   AOI22_X1 i_257_76_503 (.A1(n_257_451), .A2(n_257_76_502), .B1(n_257_861), 
      .B2(n_257_76_17903), .ZN(n_257_76_503));
   AOI22_X1 i_257_76_504 (.A1(n_257_113), .A2(n_257_76_17925), .B1(n_257_733), 
      .B2(n_257_76_17935), .ZN(n_257_76_504));
   NAND2_X1 i_257_76_505 (.A1(n_257_76_503), .A2(n_257_76_504), .ZN(n_257_76_505));
   NAND2_X1 i_257_76_506 (.A1(n_257_75), .A2(n_257_76_17932), .ZN(n_257_76_506));
   INV_X1 i_257_76_507 (.A(n_257_76_506), .ZN(n_257_76_507));
   NOR2_X1 i_257_76_508 (.A1(n_257_76_505), .A2(n_257_76_507), .ZN(n_257_76_508));
   NAND2_X1 i_257_76_509 (.A1(n_257_629), .A2(n_257_76_17928), .ZN(n_257_76_509));
   NAND3_X1 i_257_76_510 (.A1(n_257_439), .A2(n_257_899), .A3(n_257_442), 
      .ZN(n_257_76_510));
   NAND2_X1 i_257_76_511 (.A1(n_257_76_509), .A2(n_257_76_510), .ZN(n_257_76_511));
   NAND2_X1 i_257_76_512 (.A1(n_257_422), .A2(n_257_442), .ZN(n_257_76_512));
   INV_X1 i_257_76_513 (.A(n_257_76_512), .ZN(n_257_76_513));
   NAND2_X1 i_257_76_514 (.A1(n_257_310), .A2(n_257_76_513), .ZN(n_257_76_514));
   INV_X1 i_257_76_515 (.A(n_257_76_514), .ZN(n_257_76_515));
   NOR2_X1 i_257_76_516 (.A1(n_257_76_511), .A2(n_257_76_515), .ZN(n_257_76_516));
   INV_X1 i_257_76_517 (.A(n_257_76_32), .ZN(n_257_76_517));
   NAND2_X1 i_257_76_518 (.A1(n_257_432), .A2(n_257_76_517), .ZN(n_257_76_518));
   NAND2_X1 i_257_76_519 (.A1(n_257_76_518), .A2(n_257_76_154), .ZN(n_257_76_519));
   NAND3_X1 i_257_76_520 (.A1(n_257_388), .A2(n_257_76_2), .A3(n_257_484), 
      .ZN(n_257_76_520));
   INV_X1 i_257_76_521 (.A(Small_Packet_Data_Size[0]), .ZN(n_257_76_521));
   NAND2_X1 i_257_76_522 (.A1(n_257_76_520), .A2(n_257_76_18059), .ZN(
      n_257_76_522));
   NOR2_X1 i_257_76_523 (.A1(n_257_76_519), .A2(n_257_76_522), .ZN(n_257_76_523));
   NAND2_X1 i_257_76_524 (.A1(n_257_701), .A2(n_257_76_15655), .ZN(n_257_76_524));
   NAND2_X1 i_257_76_525 (.A1(n_257_76_523), .A2(n_257_76_524), .ZN(n_257_76_525));
   NAND2_X1 i_257_76_526 (.A1(n_257_442), .A2(n_257_931), .ZN(n_257_76_526));
   INV_X1 i_257_76_527 (.A(n_257_76_526), .ZN(n_257_76_527));
   NAND2_X1 i_257_76_528 (.A1(n_257_440), .A2(n_257_76_527), .ZN(n_257_76_528));
   NAND2_X1 i_257_76_529 (.A1(n_257_438), .A2(n_257_76_3760), .ZN(n_257_76_529));
   NAND2_X1 i_257_76_530 (.A1(n_257_76_528), .A2(n_257_76_529), .ZN(n_257_76_530));
   NOR2_X1 i_257_76_531 (.A1(n_257_76_525), .A2(n_257_76_530), .ZN(n_257_76_531));
   NAND2_X1 i_257_76_532 (.A1(n_257_76_516), .A2(n_257_76_531), .ZN(n_257_76_532));
   INV_X1 i_257_76_533 (.A(n_257_76_532), .ZN(n_257_76_533));
   NAND3_X1 i_257_76_534 (.A1(n_257_192), .A2(n_257_76_437), .A3(n_257_427), 
      .ZN(n_257_76_534));
   NAND2_X1 i_257_76_535 (.A1(n_257_765), .A2(n_257_442), .ZN(n_257_76_535));
   INV_X1 i_257_76_536 (.A(n_257_76_535), .ZN(n_257_76_536));
   NAND2_X1 i_257_76_537 (.A1(n_257_447), .A2(n_257_76_536), .ZN(n_257_76_537));
   NAND2_X1 i_257_76_538 (.A1(n_257_76_534), .A2(n_257_76_537), .ZN(n_257_76_538));
   INV_X1 i_257_76_539 (.A(n_257_501), .ZN(n_257_76_539));
   OAI22_X1 i_257_76_540 (.A1(n_257_76_315), .A2(n_257_76_16925), .B1(
      n_257_76_465), .B2(n_257_76_539), .ZN(n_257_76_540));
   NOR2_X1 i_257_76_541 (.A1(n_257_76_538), .A2(n_257_76_540), .ZN(n_257_76_541));
   NAND2_X1 i_257_76_542 (.A1(n_257_76_533), .A2(n_257_76_541), .ZN(n_257_76_542));
   NAND2_X1 i_257_76_543 (.A1(n_257_829), .A2(n_257_442), .ZN(n_257_76_543));
   INV_X1 i_257_76_544 (.A(n_257_76_543), .ZN(n_257_76_544));
   NAND2_X1 i_257_76_545 (.A1(n_257_446), .A2(n_257_76_544), .ZN(n_257_76_545));
   NAND2_X1 i_257_76_546 (.A1(n_257_449), .A2(n_257_76_8280), .ZN(n_257_76_546));
   NAND2_X1 i_257_76_547 (.A1(n_257_76_545), .A2(n_257_76_546), .ZN(n_257_76_547));
   NAND2_X1 i_257_76_548 (.A1(n_257_35), .A2(n_257_76_17918), .ZN(n_257_76_548));
   INV_X1 i_257_76_549 (.A(n_257_76_548), .ZN(n_257_76_549));
   NOR2_X1 i_257_76_550 (.A1(n_257_76_547), .A2(n_257_76_549), .ZN(n_257_76_550));
   NAND2_X1 i_257_76_551 (.A1(n_257_963), .A2(n_257_442), .ZN(n_257_76_551));
   INV_X1 i_257_76_552 (.A(n_257_76_551), .ZN(n_257_76_552));
   AOI22_X1 i_257_76_553 (.A1(n_257_797), .A2(n_257_76_17952), .B1(n_257_441), 
      .B2(n_257_76_552), .ZN(n_257_76_553));
   NAND2_X1 i_257_76_554 (.A1(n_257_76_550), .A2(n_257_76_553), .ZN(n_257_76_554));
   NOR2_X1 i_257_76_555 (.A1(n_257_76_542), .A2(n_257_76_554), .ZN(n_257_76_555));
   NAND2_X1 i_257_76_556 (.A1(n_257_76_508), .A2(n_257_76_555), .ZN(n_257_76_556));
   INV_X1 i_257_76_557 (.A(n_257_152), .ZN(n_257_76_557));
   OAI21_X1 i_257_76_558 (.A(n_257_76_208), .B1(n_257_76_557), .B2(
      n_257_76_17660), .ZN(n_257_76_558));
   INV_X1 i_257_76_559 (.A(n_257_76_558), .ZN(n_257_76_559));
   NAND2_X1 i_257_76_560 (.A1(n_257_669), .A2(n_257_76_17958), .ZN(n_257_76_560));
   NAND2_X1 i_257_76_561 (.A1(n_257_76_115), .A2(n_257_76_560), .ZN(n_257_76_561));
   INV_X1 i_257_76_562 (.A(n_257_76_561), .ZN(n_257_76_562));
   NAND2_X1 i_257_76_563 (.A1(n_257_76_559), .A2(n_257_76_562), .ZN(n_257_76_563));
   NOR2_X1 i_257_76_564 (.A1(n_257_76_556), .A2(n_257_76_563), .ZN(n_257_76_564));
   AOI22_X1 i_257_76_565 (.A1(n_257_1027), .A2(n_257_76_17969), .B1(n_257_995), 
      .B2(n_257_76_17964), .ZN(n_257_76_565));
   NAND2_X1 i_257_76_566 (.A1(n_257_76_564), .A2(n_257_76_565), .ZN(n_257_76_566));
   NAND2_X1 i_257_76_567 (.A1(n_257_76_408), .A2(n_257_76_428), .ZN(n_257_76_567));
   NOR2_X1 i_257_76_568 (.A1(n_257_76_566), .A2(n_257_76_567), .ZN(n_257_76_568));
   NAND2_X1 i_257_76_569 (.A1(n_257_76_0), .A2(n_257_76_407), .ZN(n_257_76_569));
   INV_X1 i_257_76_570 (.A(n_257_76_569), .ZN(n_257_76_570));
   NAND2_X1 i_257_76_571 (.A1(n_257_76_41), .A2(n_257_76_29), .ZN(n_257_76_571));
   INV_X1 i_257_76_572 (.A(n_257_76_571), .ZN(n_257_76_572));
   NAND2_X1 i_257_76_573 (.A1(n_257_76_572), .A2(n_257_76_40), .ZN(n_257_76_573));
   NAND2_X1 i_257_76_574 (.A1(n_257_76_39), .A2(n_257_76_112), .ZN(n_257_76_574));
   NOR2_X1 i_257_76_575 (.A1(n_257_76_573), .A2(n_257_76_574), .ZN(n_257_76_575));
   INV_X1 i_257_76_576 (.A(n_257_76_520), .ZN(n_257_76_576));
   NAND2_X1 i_257_76_577 (.A1(n_257_76_104), .A2(n_257_76_576), .ZN(n_257_76_577));
   INV_X1 i_257_76_578 (.A(n_257_76_103), .ZN(n_257_76_578));
   NOR2_X1 i_257_76_579 (.A1(n_257_76_577), .A2(n_257_76_578), .ZN(n_257_76_579));
   NAND2_X1 i_257_76_580 (.A1(n_257_1089), .A2(n_257_420), .ZN(n_257_76_580));
   NAND2_X1 i_257_76_581 (.A1(n_257_76_579), .A2(n_257_76_580), .ZN(n_257_76_581));
   NAND2_X1 i_257_76_582 (.A1(n_257_76_107), .A2(n_257_76_31), .ZN(n_257_76_582));
   NOR2_X1 i_257_76_583 (.A1(n_257_76_581), .A2(n_257_76_582), .ZN(n_257_76_583));
   NAND2_X1 i_257_76_584 (.A1(n_257_76_583), .A2(n_257_76_341), .ZN(n_257_76_584));
   NAND2_X1 i_257_76_585 (.A1(n_257_76_99), .A2(n_257_76_308), .ZN(n_257_76_585));
   INV_X1 i_257_76_586 (.A(n_257_76_585), .ZN(n_257_76_586));
   NAND2_X1 i_257_76_587 (.A1(n_257_76_586), .A2(n_257_76_340), .ZN(n_257_76_587));
   NOR2_X1 i_257_76_588 (.A1(n_257_76_584), .A2(n_257_76_587), .ZN(n_257_76_588));
   NAND2_X1 i_257_76_589 (.A1(n_257_76_575), .A2(n_257_76_588), .ZN(n_257_76_589));
   INV_X1 i_257_76_590 (.A(n_257_76_325), .ZN(n_257_76_590));
   NOR2_X1 i_257_76_591 (.A1(n_257_76_257), .A2(n_257_76_590), .ZN(n_257_76_591));
   NAND2_X1 i_257_76_592 (.A1(n_257_76_92), .A2(n_257_76_19), .ZN(n_257_76_592));
   INV_X1 i_257_76_593 (.A(n_257_76_592), .ZN(n_257_76_593));
   NAND2_X1 i_257_76_594 (.A1(n_257_76_591), .A2(n_257_76_593), .ZN(n_257_76_594));
   NOR2_X1 i_257_76_595 (.A1(n_257_76_589), .A2(n_257_76_594), .ZN(n_257_76_595));
   INV_X1 i_257_76_596 (.A(n_257_76_18), .ZN(n_257_76_596));
   NAND2_X1 i_257_76_597 (.A1(n_257_76_97), .A2(n_257_76_596), .ZN(n_257_76_597));
   INV_X1 i_257_76_598 (.A(n_257_76_329), .ZN(n_257_76_598));
   NOR2_X1 i_257_76_599 (.A1(n_257_76_597), .A2(n_257_76_598), .ZN(n_257_76_599));
   NAND2_X1 i_257_76_600 (.A1(n_257_76_595), .A2(n_257_76_599), .ZN(n_257_76_600));
   INV_X1 i_257_76_601 (.A(n_257_76_600), .ZN(n_257_76_601));
   NAND2_X1 i_257_76_602 (.A1(n_257_76_570), .A2(n_257_76_601), .ZN(n_257_76_602));
   NAND2_X1 i_257_76_603 (.A1(n_257_76_12), .A2(n_257_76_119), .ZN(n_257_76_603));
   NOR2_X1 i_257_76_604 (.A1(n_257_76_602), .A2(n_257_76_603), .ZN(n_257_76_604));
   AOI21_X1 i_257_76_605 (.A(n_257_76_568), .B1(n_257_12), .B2(n_257_76_604), 
      .ZN(n_257_76_605));
   NAND2_X1 i_257_76_606 (.A1(n_257_76_500), .A2(n_257_76_605), .ZN(n_257_76_606));
   INV_X1 i_257_76_607 (.A(n_257_76_606), .ZN(n_257_76_607));
   NAND3_X1 i_257_76_608 (.A1(n_257_76_434), .A2(n_257_76_481), .A3(n_257_76_607), 
      .ZN(n_257_76_608));
   NOR2_X1 i_257_76_609 (.A1(n_257_76_383), .A2(n_257_76_608), .ZN(n_257_76_609));
   NAND2_X1 i_257_76_610 (.A1(n_257_76_244), .A2(n_257_76_609), .ZN(n_0));
   NAND2_X1 i_257_76_611 (.A1(n_257_996), .A2(n_257_444), .ZN(n_257_76_610));
   NAND2_X1 i_257_76_612 (.A1(n_257_441), .A2(n_257_964), .ZN(n_257_76_611));
   NOR2_X1 i_257_76_613 (.A1(n_257_1060), .A2(n_257_76_17412), .ZN(n_257_76_612));
   INV_X1 i_257_76_614 (.A(n_257_76_612), .ZN(n_257_76_613));
   INV_X1 i_257_76_615 (.A(n_257_932), .ZN(n_257_76_614));
   NOR2_X1 i_257_76_616 (.A1(n_257_76_613), .A2(n_257_76_614), .ZN(n_257_76_615));
   NAND2_X1 i_257_76_617 (.A1(n_257_440), .A2(n_257_76_615), .ZN(n_257_76_616));
   INV_X1 i_257_76_618 (.A(n_257_76_616), .ZN(n_257_76_617));
   NAND2_X1 i_257_76_619 (.A1(n_257_76_611), .A2(n_257_76_617), .ZN(n_257_76_618));
   INV_X1 i_257_76_620 (.A(n_257_76_618), .ZN(n_257_76_619));
   NAND2_X1 i_257_76_621 (.A1(n_257_76_610), .A2(n_257_76_619), .ZN(n_257_76_620));
   INV_X1 i_257_76_622 (.A(n_257_76_620), .ZN(n_257_76_621));
   NAND2_X1 i_257_76_623 (.A1(n_257_1028), .A2(n_257_443), .ZN(n_257_76_622));
   NAND2_X1 i_257_76_624 (.A1(n_257_76_621), .A2(n_257_76_622), .ZN(n_257_76_623));
   INV_X1 i_257_76_625 (.A(n_257_76_623), .ZN(n_257_76_624));
   NAND2_X1 i_257_76_626 (.A1(n_257_17), .A2(n_257_76_624), .ZN(n_257_76_625));
   INV_X1 i_257_76_627 (.A(n_257_76_622), .ZN(n_257_76_626));
   NAND2_X1 i_257_76_628 (.A1(n_257_862), .A2(n_257_445), .ZN(n_257_76_627));
   NAND2_X1 i_257_76_629 (.A1(n_257_798), .A2(n_257_437), .ZN(n_257_76_628));
   NAND3_X1 i_257_76_630 (.A1(n_257_76_627), .A2(n_257_76_611), .A3(n_257_76_628), 
      .ZN(n_257_76_629));
   NAND2_X1 i_257_76_631 (.A1(n_257_451), .A2(n_257_453), .ZN(n_257_76_630));
   NAND2_X1 i_257_76_632 (.A1(n_257_734), .A2(n_257_436), .ZN(n_257_76_631));
   NAND2_X1 i_257_76_633 (.A1(n_257_76_630), .A2(n_257_76_631), .ZN(n_257_76_632));
   NOR2_X1 i_257_76_634 (.A1(n_257_76_629), .A2(n_257_76_632), .ZN(n_257_76_633));
   NAND2_X1 i_257_76_635 (.A1(n_257_670), .A2(n_257_448), .ZN(n_257_76_634));
   NAND2_X1 i_257_76_636 (.A1(n_257_36), .A2(n_257_433), .ZN(n_257_76_635));
   NAND2_X1 i_257_76_637 (.A1(n_257_446), .A2(n_257_830), .ZN(n_257_76_636));
   NAND2_X1 i_257_76_638 (.A1(n_257_449), .A2(n_257_1074), .ZN(n_257_76_637));
   NAND2_X1 i_257_76_639 (.A1(n_257_447), .A2(n_257_766), .ZN(n_257_76_638));
   NAND4_X1 i_257_76_640 (.A1(n_257_76_635), .A2(n_257_76_636), .A3(n_257_76_637), 
      .A4(n_257_76_638), .ZN(n_257_76_639));
   NAND2_X1 i_257_76_641 (.A1(n_257_438), .A2(n_257_1066), .ZN(n_257_76_640));
   NAND2_X1 i_257_76_642 (.A1(n_257_439), .A2(n_257_900), .ZN(n_257_76_641));
   INV_X1 i_257_76_643 (.A(n_257_598), .ZN(n_257_76_642));
   NOR2_X1 i_257_76_644 (.A1(n_257_76_613), .A2(n_257_76_642), .ZN(n_257_76_643));
   NAND2_X1 i_257_76_645 (.A1(n_257_432), .A2(n_257_76_643), .ZN(n_257_76_644));
   INV_X1 i_257_76_646 (.A(n_257_76_644), .ZN(n_257_76_645));
   NAND3_X1 i_257_76_647 (.A1(n_257_76_640), .A2(n_257_76_641), .A3(n_257_76_645), 
      .ZN(n_257_76_646));
   INV_X1 i_257_76_648 (.A(n_257_76_646), .ZN(n_257_76_647));
   NAND2_X1 i_257_76_649 (.A1(n_257_440), .A2(n_257_932), .ZN(n_257_76_648));
   NAND2_X1 i_257_76_650 (.A1(n_257_702), .A2(n_257_435), .ZN(n_257_76_649));
   NAND2_X1 i_257_76_651 (.A1(n_257_76_648), .A2(n_257_76_649), .ZN(n_257_76_650));
   INV_X1 i_257_76_652 (.A(n_257_76_650), .ZN(n_257_76_651));
   NAND2_X1 i_257_76_653 (.A1(n_257_630), .A2(n_257_450), .ZN(n_257_76_652));
   NAND3_X1 i_257_76_654 (.A1(n_257_76_647), .A2(n_257_76_651), .A3(n_257_76_652), 
      .ZN(n_257_76_653));
   NOR2_X1 i_257_76_655 (.A1(n_257_76_639), .A2(n_257_76_653), .ZN(n_257_76_654));
   NAND3_X1 i_257_76_656 (.A1(n_257_76_633), .A2(n_257_76_634), .A3(n_257_76_654), 
      .ZN(n_257_76_655));
   INV_X1 i_257_76_657 (.A(n_257_76_655), .ZN(n_257_76_656));
   NAND2_X1 i_257_76_658 (.A1(n_257_76_656), .A2(n_257_76_610), .ZN(n_257_76_657));
   NOR2_X1 i_257_76_659 (.A1(n_257_76_626), .A2(n_257_76_657), .ZN(n_257_76_658));
   NAND2_X1 i_257_76_660 (.A1(n_257_68), .A2(n_257_76_658), .ZN(n_257_76_659));
   NAND2_X1 i_257_76_661 (.A1(n_257_450), .A2(n_257_76_612), .ZN(n_257_76_660));
   INV_X1 i_257_76_662 (.A(n_257_76_660), .ZN(n_257_76_661));
   NAND3_X1 i_257_76_663 (.A1(n_257_76_641), .A2(n_257_630), .A3(n_257_76_661), 
      .ZN(n_257_76_662));
   NAND2_X1 i_257_76_664 (.A1(n_257_76_649), .A2(n_257_76_640), .ZN(n_257_76_663));
   NOR2_X1 i_257_76_665 (.A1(n_257_76_662), .A2(n_257_76_663), .ZN(n_257_76_664));
   NAND2_X1 i_257_76_666 (.A1(n_257_76_636), .A2(n_257_76_637), .ZN(n_257_76_665));
   INV_X1 i_257_76_667 (.A(n_257_76_665), .ZN(n_257_76_666));
   NAND2_X1 i_257_76_668 (.A1(n_257_76_638), .A2(n_257_76_648), .ZN(n_257_76_667));
   INV_X1 i_257_76_669 (.A(n_257_76_667), .ZN(n_257_76_668));
   NAND3_X1 i_257_76_670 (.A1(n_257_76_664), .A2(n_257_76_666), .A3(n_257_76_668), 
      .ZN(n_257_76_669));
   INV_X1 i_257_76_671 (.A(n_257_76_669), .ZN(n_257_76_670));
   NAND4_X1 i_257_76_672 (.A1(n_257_76_631), .A2(n_257_76_627), .A3(n_257_76_611), 
      .A4(n_257_76_628), .ZN(n_257_76_671));
   INV_X1 i_257_76_673 (.A(n_257_76_671), .ZN(n_257_76_672));
   NAND2_X1 i_257_76_674 (.A1(n_257_76_670), .A2(n_257_76_672), .ZN(n_257_76_673));
   INV_X1 i_257_76_675 (.A(n_257_76_634), .ZN(n_257_76_674));
   NOR2_X1 i_257_76_676 (.A1(n_257_76_673), .A2(n_257_76_674), .ZN(n_257_76_675));
   NAND2_X1 i_257_76_677 (.A1(n_257_76_610), .A2(n_257_76_675), .ZN(n_257_76_676));
   NOR2_X1 i_257_76_678 (.A1(n_257_76_676), .A2(n_257_76_626), .ZN(n_257_76_677));
   NAND2_X1 i_257_76_679 (.A1(n_257_28), .A2(n_257_76_677), .ZN(n_257_76_678));
   NAND3_X1 i_257_76_680 (.A1(n_257_76_625), .A2(n_257_76_659), .A3(n_257_76_678), 
      .ZN(n_257_76_679));
   INV_X1 i_257_76_681 (.A(n_257_76_648), .ZN(n_257_76_680));
   NAND3_X1 i_257_76_682 (.A1(n_257_439), .A2(n_257_900), .A3(n_257_76_612), 
      .ZN(n_257_76_681));
   NOR2_X1 i_257_76_683 (.A1(n_257_76_680), .A2(n_257_76_681), .ZN(n_257_76_682));
   NAND2_X1 i_257_76_684 (.A1(n_257_76_611), .A2(n_257_76_682), .ZN(n_257_76_683));
   INV_X1 i_257_76_685 (.A(n_257_76_683), .ZN(n_257_76_684));
   NAND2_X1 i_257_76_686 (.A1(n_257_76_610), .A2(n_257_76_684), .ZN(n_257_76_685));
   INV_X1 i_257_76_687 (.A(n_257_76_685), .ZN(n_257_76_686));
   NAND2_X1 i_257_76_688 (.A1(n_257_76_686), .A2(n_257_76_622), .ZN(n_257_76_687));
   INV_X1 i_257_76_689 (.A(n_257_76_687), .ZN(n_257_76_688));
   NAND2_X1 i_257_76_690 (.A1(n_257_18), .A2(n_257_76_688), .ZN(n_257_76_689));
   NAND2_X1 i_257_76_691 (.A1(n_257_830), .A2(n_257_76_612), .ZN(n_257_76_690));
   INV_X1 i_257_76_692 (.A(n_257_76_690), .ZN(n_257_76_691));
   NAND3_X1 i_257_76_693 (.A1(n_257_76_640), .A2(n_257_76_641), .A3(n_257_76_691), 
      .ZN(n_257_76_692));
   NAND2_X1 i_257_76_694 (.A1(n_257_446), .A2(n_257_76_648), .ZN(n_257_76_693));
   NOR2_X1 i_257_76_695 (.A1(n_257_76_692), .A2(n_257_76_693), .ZN(n_257_76_694));
   NAND3_X1 i_257_76_696 (.A1(n_257_76_694), .A2(n_257_76_627), .A3(n_257_76_611), 
      .ZN(n_257_76_695));
   INV_X1 i_257_76_697 (.A(n_257_76_695), .ZN(n_257_76_696));
   NAND2_X1 i_257_76_698 (.A1(n_257_76_610), .A2(n_257_76_696), .ZN(n_257_76_697));
   INV_X1 i_257_76_699 (.A(n_257_76_697), .ZN(n_257_76_698));
   NAND2_X1 i_257_76_700 (.A1(n_257_76_698), .A2(n_257_76_622), .ZN(n_257_76_699));
   INV_X1 i_257_76_701 (.A(n_257_76_699), .ZN(n_257_76_700));
   NAND2_X1 i_257_76_702 (.A1(n_257_21), .A2(n_257_76_700), .ZN(n_257_76_701));
   NAND2_X1 i_257_76_703 (.A1(n_257_193), .A2(n_257_427), .ZN(n_257_76_702));
   NAND4_X1 i_257_76_704 (.A1(n_257_76_652), .A2(n_257_76_702), .A3(n_257_76_648), 
      .A4(n_257_76_649), .ZN(n_257_76_703));
   INV_X1 i_257_76_705 (.A(n_257_76_703), .ZN(n_257_76_704));
   NAND2_X1 i_257_76_706 (.A1(n_257_423), .A2(n_257_76_612), .ZN(n_257_76_705));
   INV_X1 i_257_76_707 (.A(n_257_76_705), .ZN(n_257_76_706));
   NAND2_X1 i_257_76_708 (.A1(n_257_432), .A2(n_257_598), .ZN(n_257_76_707));
   NAND2_X1 i_257_76_709 (.A1(n_257_428), .A2(n_257_566), .ZN(n_257_76_708));
   NAND3_X1 i_257_76_710 (.A1(n_257_76_706), .A2(n_257_76_707), .A3(n_257_76_708), 
      .ZN(n_257_76_709));
   INV_X1 i_257_76_711 (.A(n_257_76_709), .ZN(n_257_76_710));
   NAND2_X1 i_257_76_712 (.A1(n_257_502), .A2(n_257_424), .ZN(n_257_76_711));
   NAND4_X1 i_257_76_713 (.A1(n_257_76_640), .A2(n_257_76_641), .A3(n_257_76_710), 
      .A4(n_257_76_711), .ZN(n_257_76_712));
   INV_X1 i_257_76_714 (.A(n_257_76_712), .ZN(n_257_76_713));
   NAND3_X1 i_257_76_715 (.A1(n_257_76_704), .A2(n_257_273), .A3(n_257_76_713), 
      .ZN(n_257_76_714));
   NAND2_X1 i_257_76_716 (.A1(n_257_534), .A2(n_257_426), .ZN(n_257_76_715));
   NAND3_X1 i_257_76_717 (.A1(n_257_76_628), .A2(n_257_76_635), .A3(n_257_76_715), 
      .ZN(n_257_76_716));
   NAND2_X1 i_257_76_718 (.A1(n_257_76_631), .A2(n_257_76_627), .ZN(n_257_76_717));
   NOR3_X1 i_257_76_719 (.A1(n_257_76_714), .A2(n_257_76_716), .A3(n_257_76_717), 
      .ZN(n_257_76_718));
   NAND2_X1 i_257_76_720 (.A1(n_257_76_610), .A2(n_257_76_718), .ZN(n_257_76_719));
   INV_X1 i_257_76_721 (.A(n_257_76_719), .ZN(n_257_76_720));
   NAND3_X1 i_257_76_722 (.A1(n_257_76_636), .A2(n_257_76_637), .A3(n_257_76_638), 
      .ZN(n_257_76_721));
   INV_X1 i_257_76_723 (.A(n_257_76_611), .ZN(n_257_76_722));
   NOR2_X1 i_257_76_724 (.A1(n_257_76_721), .A2(n_257_76_722), .ZN(n_257_76_723));
   NAND2_X1 i_257_76_725 (.A1(n_257_76), .A2(n_257_431), .ZN(n_257_76_724));
   NAND2_X1 i_257_76_726 (.A1(n_257_114), .A2(n_257_430), .ZN(n_257_76_725));
   NAND2_X1 i_257_76_727 (.A1(n_257_76_630), .A2(n_257_76_725), .ZN(n_257_76_726));
   INV_X1 i_257_76_728 (.A(n_257_76_726), .ZN(n_257_76_727));
   NAND3_X1 i_257_76_729 (.A1(n_257_76_723), .A2(n_257_76_724), .A3(n_257_76_727), 
      .ZN(n_257_76_728));
   INV_X1 i_257_76_730 (.A(n_257_76_728), .ZN(n_257_76_729));
   NAND2_X1 i_257_76_731 (.A1(n_257_233), .A2(n_257_425), .ZN(n_257_76_730));
   NAND2_X1 i_257_76_732 (.A1(n_257_153), .A2(n_257_429), .ZN(n_257_76_731));
   NAND4_X1 i_257_76_733 (.A1(n_257_76_729), .A2(n_257_76_730), .A3(n_257_76_731), 
      .A4(n_257_76_634), .ZN(n_257_76_732));
   INV_X1 i_257_76_734 (.A(n_257_76_732), .ZN(n_257_76_733));
   NAND3_X1 i_257_76_735 (.A1(n_257_76_720), .A2(n_257_76_622), .A3(n_257_76_733), 
      .ZN(n_257_76_734));
   INV_X1 i_257_76_736 (.A(n_257_76_734), .ZN(n_257_76_735));
   NAND2_X1 i_257_76_737 (.A1(n_257_304), .A2(n_257_76_735), .ZN(n_257_76_736));
   NAND3_X1 i_257_76_738 (.A1(n_257_76_689), .A2(n_257_76_701), .A3(n_257_76_736), 
      .ZN(n_257_76_737));
   NOR2_X1 i_257_76_739 (.A1(n_257_76_679), .A2(n_257_76_737), .ZN(n_257_76_738));
   NAND2_X1 i_257_76_740 (.A1(n_257_964), .A2(n_257_76_612), .ZN(n_257_76_739));
   INV_X1 i_257_76_741 (.A(n_257_76_739), .ZN(n_257_76_740));
   NAND2_X1 i_257_76_742 (.A1(n_257_441), .A2(n_257_76_740), .ZN(n_257_76_741));
   INV_X1 i_257_76_743 (.A(n_257_76_741), .ZN(n_257_76_742));
   NAND2_X1 i_257_76_744 (.A1(n_257_76_610), .A2(n_257_76_742), .ZN(n_257_76_743));
   INV_X1 i_257_76_745 (.A(n_257_76_743), .ZN(n_257_76_744));
   NAND2_X1 i_257_76_746 (.A1(n_257_76_744), .A2(n_257_76_622), .ZN(n_257_76_745));
   INV_X1 i_257_76_747 (.A(n_257_76_745), .ZN(n_257_76_746));
   NAND2_X1 i_257_76_748 (.A1(n_257_16), .A2(n_257_76_746), .ZN(n_257_76_747));
   NAND2_X1 i_257_76_749 (.A1(n_257_76_636), .A2(n_257_76_638), .ZN(n_257_76_748));
   INV_X1 i_257_76_750 (.A(n_257_76_748), .ZN(n_257_76_749));
   NAND2_X1 i_257_76_751 (.A1(n_257_435), .A2(n_257_76_612), .ZN(n_257_76_750));
   INV_X1 i_257_76_752 (.A(n_257_76_750), .ZN(n_257_76_751));
   NAND2_X1 i_257_76_753 (.A1(n_257_702), .A2(n_257_76_751), .ZN(n_257_76_752));
   INV_X1 i_257_76_754 (.A(n_257_76_752), .ZN(n_257_76_753));
   NAND4_X1 i_257_76_755 (.A1(n_257_76_753), .A2(n_257_76_648), .A3(n_257_76_640), 
      .A4(n_257_76_641), .ZN(n_257_76_754));
   INV_X1 i_257_76_756 (.A(n_257_76_754), .ZN(n_257_76_755));
   NAND3_X1 i_257_76_757 (.A1(n_257_76_749), .A2(n_257_76_755), .A3(n_257_76_628), 
      .ZN(n_257_76_756));
   NAND3_X1 i_257_76_758 (.A1(n_257_76_631), .A2(n_257_76_627), .A3(n_257_76_611), 
      .ZN(n_257_76_757));
   NOR2_X1 i_257_76_759 (.A1(n_257_76_756), .A2(n_257_76_757), .ZN(n_257_76_758));
   NAND2_X1 i_257_76_760 (.A1(n_257_76_610), .A2(n_257_76_758), .ZN(n_257_76_759));
   INV_X1 i_257_76_761 (.A(n_257_76_759), .ZN(n_257_76_760));
   NAND2_X1 i_257_76_762 (.A1(n_257_76_760), .A2(n_257_76_622), .ZN(n_257_76_761));
   INV_X1 i_257_76_763 (.A(n_257_76_761), .ZN(n_257_76_762));
   NAND2_X1 i_257_76_764 (.A1(n_257_25), .A2(n_257_76_762), .ZN(n_257_76_763));
   NAND2_X1 i_257_76_765 (.A1(n_257_442), .A2(n_257_566), .ZN(n_257_76_764));
   NOR2_X1 i_257_76_766 (.A1(n_257_76_764), .A2(n_257_1060), .ZN(n_257_76_765));
   NAND2_X1 i_257_76_767 (.A1(n_257_428), .A2(n_257_76_765), .ZN(n_257_76_766));
   INV_X1 i_257_76_768 (.A(n_257_76_766), .ZN(n_257_76_767));
   NAND2_X1 i_257_76_769 (.A1(n_257_76_707), .A2(n_257_76_767), .ZN(n_257_76_768));
   INV_X1 i_257_76_770 (.A(n_257_76_768), .ZN(n_257_76_769));
   NAND3_X1 i_257_76_771 (.A1(n_257_76_640), .A2(n_257_76_641), .A3(n_257_76_769), 
      .ZN(n_257_76_770));
   INV_X1 i_257_76_772 (.A(n_257_76_770), .ZN(n_257_76_771));
   NAND3_X1 i_257_76_773 (.A1(n_257_76_771), .A2(n_257_76_651), .A3(n_257_76_652), 
      .ZN(n_257_76_772));
   NOR2_X1 i_257_76_774 (.A1(n_257_76_772), .A2(n_257_76_721), .ZN(n_257_76_773));
   NAND4_X1 i_257_76_775 (.A1(n_257_76_627), .A2(n_257_76_611), .A3(n_257_76_628), 
      .A4(n_257_76_635), .ZN(n_257_76_774));
   INV_X1 i_257_76_776 (.A(n_257_76_774), .ZN(n_257_76_775));
   NAND3_X1 i_257_76_777 (.A1(n_257_76_630), .A2(n_257_76_725), .A3(n_257_76_631), 
      .ZN(n_257_76_776));
   INV_X1 i_257_76_778 (.A(n_257_76_776), .ZN(n_257_76_777));
   NAND4_X1 i_257_76_779 (.A1(n_257_76_773), .A2(n_257_76_775), .A3(n_257_76_777), 
      .A4(n_257_76_724), .ZN(n_257_76_778));
   NAND2_X1 i_257_76_780 (.A1(n_257_76_731), .A2(n_257_76_634), .ZN(n_257_76_779));
   NOR2_X1 i_257_76_781 (.A1(n_257_76_778), .A2(n_257_76_779), .ZN(n_257_76_780));
   NAND3_X1 i_257_76_782 (.A1(n_257_76_780), .A2(n_257_76_622), .A3(n_257_76_610), 
      .ZN(n_257_76_781));
   INV_X1 i_257_76_783 (.A(n_257_76_781), .ZN(n_257_76_782));
   NAND2_X1 i_257_76_784 (.A1(n_257_185), .A2(n_257_76_782), .ZN(n_257_76_783));
   NAND3_X1 i_257_76_785 (.A1(n_257_76_747), .A2(n_257_76_763), .A3(n_257_76_783), 
      .ZN(n_257_76_784));
   NAND2_X1 i_257_76_786 (.A1(n_257_1060), .A2(n_257_442), .ZN(n_257_76_785));
   INV_X1 i_257_76_787 (.A(n_257_76_785), .ZN(n_257_76_786));
   NAND2_X1 i_257_76_788 (.A1(n_257_13), .A2(n_257_76_786), .ZN(n_257_76_787));
   NAND2_X1 i_257_76_789 (.A1(n_257_76_648), .A2(n_257_76_640), .ZN(n_257_76_788));
   INV_X1 i_257_76_790 (.A(n_257_76_788), .ZN(n_257_76_789));
   NAND2_X1 i_257_76_791 (.A1(n_257_445), .A2(n_257_76_612), .ZN(n_257_76_790));
   INV_X1 i_257_76_792 (.A(n_257_76_790), .ZN(n_257_76_791));
   NAND2_X1 i_257_76_793 (.A1(n_257_76_641), .A2(n_257_76_791), .ZN(n_257_76_792));
   INV_X1 i_257_76_794 (.A(n_257_76_792), .ZN(n_257_76_793));
   NAND3_X1 i_257_76_795 (.A1(n_257_76_789), .A2(n_257_862), .A3(n_257_76_793), 
      .ZN(n_257_76_794));
   NOR2_X1 i_257_76_796 (.A1(n_257_76_794), .A2(n_257_76_722), .ZN(n_257_76_795));
   NAND2_X1 i_257_76_797 (.A1(n_257_76_610), .A2(n_257_76_795), .ZN(n_257_76_796));
   INV_X1 i_257_76_798 (.A(n_257_76_796), .ZN(n_257_76_797));
   NAND2_X1 i_257_76_799 (.A1(n_257_76_797), .A2(n_257_76_622), .ZN(n_257_76_798));
   INV_X1 i_257_76_800 (.A(n_257_76_798), .ZN(n_257_76_799));
   NAND2_X1 i_257_76_801 (.A1(n_257_20), .A2(n_257_76_799), .ZN(n_257_76_800));
   NAND2_X1 i_257_76_802 (.A1(n_257_76_787), .A2(n_257_76_800), .ZN(n_257_76_801));
   NOR2_X1 i_257_76_803 (.A1(n_257_76_784), .A2(n_257_76_801), .ZN(n_257_76_802));
   NAND2_X1 i_257_76_804 (.A1(n_257_436), .A2(n_257_76_612), .ZN(n_257_76_803));
   INV_X1 i_257_76_805 (.A(n_257_76_803), .ZN(n_257_76_804));
   NAND4_X1 i_257_76_806 (.A1(n_257_76_648), .A2(n_257_76_640), .A3(n_257_76_641), 
      .A4(n_257_76_804), .ZN(n_257_76_805));
   INV_X1 i_257_76_807 (.A(n_257_76_805), .ZN(n_257_76_806));
   NAND4_X1 i_257_76_808 (.A1(n_257_76_806), .A2(n_257_734), .A3(n_257_76_636), 
      .A4(n_257_76_638), .ZN(n_257_76_807));
   NOR2_X1 i_257_76_809 (.A1(n_257_76_807), .A2(n_257_76_629), .ZN(n_257_76_808));
   NAND2_X1 i_257_76_810 (.A1(n_257_76_610), .A2(n_257_76_808), .ZN(n_257_76_809));
   INV_X1 i_257_76_811 (.A(n_257_76_809), .ZN(n_257_76_810));
   NAND2_X1 i_257_76_812 (.A1(n_257_76_810), .A2(n_257_76_622), .ZN(n_257_76_811));
   INV_X1 i_257_76_813 (.A(n_257_76_811), .ZN(n_257_76_812));
   NAND2_X1 i_257_76_814 (.A1(n_257_24), .A2(n_257_76_812), .ZN(n_257_76_813));
   NAND4_X1 i_257_76_815 (.A1(n_257_534), .A2(n_257_76_652), .A3(n_257_76_702), 
      .A4(n_257_76_648), .ZN(n_257_76_814));
   NAND2_X1 i_257_76_816 (.A1(n_257_426), .A2(n_257_76_612), .ZN(n_257_76_815));
   INV_X1 i_257_76_817 (.A(n_257_76_815), .ZN(n_257_76_816));
   NAND3_X1 i_257_76_818 (.A1(n_257_76_707), .A2(n_257_76_816), .A3(n_257_76_708), 
      .ZN(n_257_76_817));
   INV_X1 i_257_76_819 (.A(n_257_76_817), .ZN(n_257_76_818));
   NAND4_X1 i_257_76_820 (.A1(n_257_76_649), .A2(n_257_76_640), .A3(n_257_76_641), 
      .A4(n_257_76_818), .ZN(n_257_76_819));
   NOR2_X1 i_257_76_821 (.A1(n_257_76_814), .A2(n_257_76_819), .ZN(n_257_76_820));
   INV_X1 i_257_76_822 (.A(n_257_76_717), .ZN(n_257_76_821));
   NAND2_X1 i_257_76_823 (.A1(n_257_76_628), .A2(n_257_76_635), .ZN(n_257_76_822));
   INV_X1 i_257_76_824 (.A(n_257_76_822), .ZN(n_257_76_823));
   NAND3_X1 i_257_76_825 (.A1(n_257_76_820), .A2(n_257_76_821), .A3(n_257_76_823), 
      .ZN(n_257_76_824));
   INV_X1 i_257_76_826 (.A(n_257_76_824), .ZN(n_257_76_825));
   NAND2_X1 i_257_76_827 (.A1(n_257_76_610), .A2(n_257_76_825), .ZN(n_257_76_826));
   INV_X1 i_257_76_828 (.A(n_257_76_826), .ZN(n_257_76_827));
   INV_X1 i_257_76_829 (.A(n_257_76_721), .ZN(n_257_76_828));
   NAND4_X1 i_257_76_830 (.A1(n_257_76_828), .A2(n_257_76_630), .A3(n_257_76_725), 
      .A4(n_257_76_611), .ZN(n_257_76_829));
   INV_X1 i_257_76_831 (.A(n_257_76_829), .ZN(n_257_76_830));
   NAND4_X1 i_257_76_832 (.A1(n_257_76_731), .A2(n_257_76_634), .A3(n_257_76_830), 
      .A4(n_257_76_724), .ZN(n_257_76_831));
   INV_X1 i_257_76_833 (.A(n_257_76_831), .ZN(n_257_76_832));
   NAND3_X1 i_257_76_834 (.A1(n_257_76_827), .A2(n_257_76_622), .A3(n_257_76_832), 
      .ZN(n_257_76_833));
   INV_X1 i_257_76_835 (.A(n_257_76_833), .ZN(n_257_76_834));
   NAND2_X1 i_257_76_836 (.A1(n_257_225), .A2(n_257_76_834), .ZN(n_257_76_835));
   NAND2_X1 i_257_76_837 (.A1(n_257_443), .A2(n_257_76_612), .ZN(n_257_76_836));
   INV_X1 i_257_76_838 (.A(n_257_76_836), .ZN(n_257_76_837));
   NAND2_X1 i_257_76_839 (.A1(n_257_1028), .A2(n_257_76_837), .ZN(n_257_76_838));
   INV_X1 i_257_76_840 (.A(n_257_76_838), .ZN(n_257_76_839));
   NAND2_X1 i_257_76_841 (.A1(n_257_14), .A2(n_257_76_839), .ZN(n_257_76_840));
   NAND3_X1 i_257_76_842 (.A1(n_257_76_813), .A2(n_257_76_835), .A3(n_257_76_840), 
      .ZN(n_257_76_841));
   NAND2_X1 i_257_76_843 (.A1(n_257_76_636), .A2(n_257_798), .ZN(n_257_76_842));
   INV_X1 i_257_76_844 (.A(n_257_76_842), .ZN(n_257_76_843));
   NAND2_X1 i_257_76_845 (.A1(n_257_437), .A2(n_257_76_612), .ZN(n_257_76_844));
   INV_X1 i_257_76_846 (.A(n_257_76_844), .ZN(n_257_76_845));
   NAND4_X1 i_257_76_847 (.A1(n_257_76_648), .A2(n_257_76_640), .A3(n_257_76_641), 
      .A4(n_257_76_845), .ZN(n_257_76_846));
   INV_X1 i_257_76_848 (.A(n_257_76_846), .ZN(n_257_76_847));
   NAND4_X1 i_257_76_849 (.A1(n_257_76_843), .A2(n_257_76_847), .A3(n_257_76_627), 
      .A4(n_257_76_611), .ZN(n_257_76_848));
   INV_X1 i_257_76_850 (.A(n_257_76_848), .ZN(n_257_76_849));
   NAND2_X1 i_257_76_851 (.A1(n_257_76_610), .A2(n_257_76_849), .ZN(n_257_76_850));
   INV_X1 i_257_76_852 (.A(n_257_76_850), .ZN(n_257_76_851));
   NAND2_X1 i_257_76_853 (.A1(n_257_76_851), .A2(n_257_76_622), .ZN(n_257_76_852));
   INV_X1 i_257_76_854 (.A(n_257_76_852), .ZN(n_257_76_853));
   NAND2_X1 i_257_76_855 (.A1(n_257_22), .A2(n_257_76_853), .ZN(n_257_76_854));
   NAND2_X1 i_257_76_856 (.A1(n_257_444), .A2(n_257_76_612), .ZN(n_257_76_855));
   INV_X1 i_257_76_857 (.A(n_257_76_855), .ZN(n_257_76_856));
   NAND2_X1 i_257_76_858 (.A1(n_257_996), .A2(n_257_76_856), .ZN(n_257_76_857));
   INV_X1 i_257_76_859 (.A(n_257_76_857), .ZN(n_257_76_858));
   NAND2_X1 i_257_76_860 (.A1(n_257_76_622), .A2(n_257_76_858), .ZN(n_257_76_859));
   INV_X1 i_257_76_861 (.A(n_257_76_859), .ZN(n_257_76_860));
   NAND2_X1 i_257_76_862 (.A1(n_257_15), .A2(n_257_76_860), .ZN(n_257_76_861));
   NAND2_X1 i_257_76_863 (.A1(n_257_76_854), .A2(n_257_76_861), .ZN(n_257_76_862));
   NOR2_X1 i_257_76_864 (.A1(n_257_76_841), .A2(n_257_76_862), .ZN(n_257_76_863));
   NAND3_X1 i_257_76_865 (.A1(n_257_76_738), .A2(n_257_76_802), .A3(n_257_76_863), 
      .ZN(n_257_76_864));
   INV_X1 i_257_76_866 (.A(n_257_76_864), .ZN(n_257_76_865));
   NAND4_X1 i_257_76_867 (.A1(n_257_76_636), .A2(n_257_76_637), .A3(n_257_76_638), 
      .A4(n_257_36), .ZN(n_257_76_866));
   NAND2_X1 i_257_76_868 (.A1(n_257_433), .A2(n_257_76_612), .ZN(n_257_76_867));
   INV_X1 i_257_76_869 (.A(n_257_76_867), .ZN(n_257_76_868));
   NAND3_X1 i_257_76_870 (.A1(n_257_76_640), .A2(n_257_76_641), .A3(n_257_76_868), 
      .ZN(n_257_76_869));
   INV_X1 i_257_76_871 (.A(n_257_76_869), .ZN(n_257_76_870));
   NAND3_X1 i_257_76_872 (.A1(n_257_76_870), .A2(n_257_76_651), .A3(n_257_76_652), 
      .ZN(n_257_76_871));
   NOR2_X1 i_257_76_873 (.A1(n_257_76_866), .A2(n_257_76_871), .ZN(n_257_76_872));
   NAND3_X1 i_257_76_874 (.A1(n_257_76_633), .A2(n_257_76_634), .A3(n_257_76_872), 
      .ZN(n_257_76_873));
   INV_X1 i_257_76_875 (.A(n_257_76_873), .ZN(n_257_76_874));
   NAND2_X1 i_257_76_876 (.A1(n_257_76_874), .A2(n_257_76_610), .ZN(n_257_76_875));
   NOR2_X1 i_257_76_877 (.A1(n_257_76_626), .A2(n_257_76_875), .ZN(n_257_76_876));
   NAND2_X1 i_257_76_878 (.A1(n_257_67), .A2(n_257_76_876), .ZN(n_257_76_877));
   INV_X1 i_257_76_879 (.A(n_257_76_639), .ZN(n_257_76_878));
   NAND2_X1 i_257_76_880 (.A1(n_257_76_611), .A2(n_257_76_628), .ZN(n_257_76_879));
   INV_X1 i_257_76_881 (.A(n_257_76_879), .ZN(n_257_76_880));
   NAND3_X1 i_257_76_882 (.A1(n_257_76_652), .A2(n_257_76_648), .A3(n_257_76_649), 
      .ZN(n_257_76_881));
   NAND2_X1 i_257_76_883 (.A1(n_257_431), .A2(n_257_76_612), .ZN(n_257_76_882));
   INV_X1 i_257_76_884 (.A(n_257_76_882), .ZN(n_257_76_883));
   NAND2_X1 i_257_76_885 (.A1(n_257_76_707), .A2(n_257_76_883), .ZN(n_257_76_884));
   INV_X1 i_257_76_886 (.A(n_257_76_884), .ZN(n_257_76_885));
   NAND3_X1 i_257_76_887 (.A1(n_257_76_640), .A2(n_257_76_641), .A3(n_257_76_885), 
      .ZN(n_257_76_886));
   NOR2_X1 i_257_76_888 (.A1(n_257_76_881), .A2(n_257_76_886), .ZN(n_257_76_887));
   NAND3_X1 i_257_76_889 (.A1(n_257_76_878), .A2(n_257_76_880), .A3(n_257_76_887), 
      .ZN(n_257_76_888));
   NAND4_X1 i_257_76_890 (.A1(n_257_76), .A2(n_257_76_630), .A3(n_257_76_631), 
      .A4(n_257_76_627), .ZN(n_257_76_889));
   NOR2_X1 i_257_76_891 (.A1(n_257_76_888), .A2(n_257_76_889), .ZN(n_257_76_890));
   NAND3_X1 i_257_76_892 (.A1(n_257_76_890), .A2(n_257_76_610), .A3(n_257_76_634), 
      .ZN(n_257_76_891));
   NOR2_X1 i_257_76_893 (.A1(n_257_76_626), .A2(n_257_76_891), .ZN(n_257_76_892));
   NAND2_X1 i_257_76_894 (.A1(n_257_107), .A2(n_257_76_892), .ZN(n_257_76_893));
   NAND2_X1 i_257_76_895 (.A1(n_257_429), .A2(n_257_76_612), .ZN(n_257_76_894));
   INV_X1 i_257_76_896 (.A(n_257_76_894), .ZN(n_257_76_895));
   NAND2_X1 i_257_76_897 (.A1(n_257_76_895), .A2(n_257_76_707), .ZN(n_257_76_896));
   INV_X1 i_257_76_898 (.A(n_257_76_896), .ZN(n_257_76_897));
   NAND3_X1 i_257_76_899 (.A1(n_257_76_640), .A2(n_257_76_641), .A3(n_257_76_897), 
      .ZN(n_257_76_898));
   INV_X1 i_257_76_900 (.A(n_257_76_898), .ZN(n_257_76_899));
   NAND3_X1 i_257_76_901 (.A1(n_257_76_899), .A2(n_257_76_651), .A3(n_257_76_652), 
      .ZN(n_257_76_900));
   NOR2_X1 i_257_76_902 (.A1(n_257_76_900), .A2(n_257_76_721), .ZN(n_257_76_901));
   NAND4_X1 i_257_76_903 (.A1(n_257_76_901), .A2(n_257_76_775), .A3(n_257_76_777), 
      .A4(n_257_76_724), .ZN(n_257_76_902));
   NAND2_X1 i_257_76_904 (.A1(n_257_76_634), .A2(n_257_153), .ZN(n_257_76_903));
   NOR2_X1 i_257_76_905 (.A1(n_257_76_902), .A2(n_257_76_903), .ZN(n_257_76_904));
   NAND3_X1 i_257_76_906 (.A1(n_257_76_904), .A2(n_257_76_622), .A3(n_257_76_610), 
      .ZN(n_257_76_905));
   INV_X1 i_257_76_907 (.A(n_257_76_905), .ZN(n_257_76_906));
   NAND2_X1 i_257_76_908 (.A1(n_257_184), .A2(n_257_76_906), .ZN(n_257_76_907));
   NAND3_X1 i_257_76_909 (.A1(n_257_76_877), .A2(n_257_76_893), .A3(n_257_76_907), 
      .ZN(n_257_76_908));
   INV_X1 i_257_76_910 (.A(n_257_76_908), .ZN(n_257_76_909));
   NOR2_X1 i_257_76_911 (.A1(n_257_76_613), .A2(n_257_76_4200), .ZN(n_257_76_910));
   NAND2_X1 i_257_76_912 (.A1(n_257_438), .A2(n_257_76_910), .ZN(n_257_76_911));
   INV_X1 i_257_76_913 (.A(n_257_76_911), .ZN(n_257_76_912));
   NAND3_X1 i_257_76_914 (.A1(n_257_76_912), .A2(n_257_76_648), .A3(n_257_76_641), 
      .ZN(n_257_76_913));
   INV_X1 i_257_76_915 (.A(n_257_76_913), .ZN(n_257_76_914));
   NAND2_X1 i_257_76_916 (.A1(n_257_76_611), .A2(n_257_76_914), .ZN(n_257_76_915));
   INV_X1 i_257_76_917 (.A(n_257_76_915), .ZN(n_257_76_916));
   NAND2_X1 i_257_76_918 (.A1(n_257_76_610), .A2(n_257_76_916), .ZN(n_257_76_917));
   INV_X1 i_257_76_919 (.A(n_257_76_917), .ZN(n_257_76_918));
   NAND2_X1 i_257_76_920 (.A1(n_257_76_918), .A2(n_257_76_622), .ZN(n_257_76_919));
   INV_X1 i_257_76_921 (.A(n_257_76_919), .ZN(n_257_76_920));
   NAND2_X1 i_257_76_922 (.A1(n_257_19), .A2(n_257_76_920), .ZN(n_257_76_921));
   NAND2_X1 i_257_76_923 (.A1(n_257_273), .A2(n_257_423), .ZN(n_257_76_922));
   NAND3_X1 i_257_76_924 (.A1(n_257_76_628), .A2(n_257_76_922), .A3(n_257_76_635), 
      .ZN(n_257_76_923));
   NOR2_X1 i_257_76_925 (.A1(n_257_76_757), .A2(n_257_76_923), .ZN(n_257_76_924));
   NAND4_X1 i_257_76_926 (.A1(n_257_76_715), .A2(n_257_76_636), .A3(n_257_76_637), 
      .A4(n_257_76_638), .ZN(n_257_76_925));
   NAND2_X1 i_257_76_927 (.A1(n_257_76_652), .A2(n_257_76_702), .ZN(n_257_76_926));
   INV_X1 i_257_76_928 (.A(n_257_76_926), .ZN(n_257_76_927));
   NAND2_X1 i_257_76_929 (.A1(n_257_76_640), .A2(n_257_76_641), .ZN(n_257_76_928));
   INV_X1 i_257_76_930 (.A(n_257_76_928), .ZN(n_257_76_929));
   NAND3_X1 i_257_76_931 (.A1(n_257_76_927), .A2(n_257_76_651), .A3(n_257_76_929), 
      .ZN(n_257_76_930));
   NOR2_X1 i_257_76_932 (.A1(n_257_76_925), .A2(n_257_76_930), .ZN(n_257_76_931));
   NAND2_X1 i_257_76_933 (.A1(n_257_76_711), .A2(n_257_1090), .ZN(n_257_76_932));
   INV_X1 i_257_76_934 (.A(n_257_76_932), .ZN(n_257_76_933));
   NAND2_X1 i_257_76_935 (.A1(n_257_311), .A2(n_257_422), .ZN(n_257_76_934));
   INV_X1 i_257_76_936 (.A(n_257_1060), .ZN(n_257_76_935));
   INV_X1 i_257_76_937 (.A(n_257_566), .ZN(n_257_76_936));
   NAND3_X1 i_257_76_938 (.A1(n_257_76_935), .A2(n_257_76_936), .A3(n_257_442), 
      .ZN(n_257_76_937));
   OAI21_X1 i_257_76_939 (.A(n_257_76_937), .B1(n_257_428), .B2(n_257_76_613), 
      .ZN(n_257_76_938));
   NAND3_X1 i_257_76_940 (.A1(n_257_76_938), .A2(n_257_420), .A3(n_257_76_707), 
      .ZN(n_257_76_939));
   INV_X1 i_257_76_941 (.A(n_257_76_939), .ZN(n_257_76_940));
   NAND3_X1 i_257_76_942 (.A1(n_257_76_933), .A2(n_257_76_934), .A3(n_257_76_940), 
      .ZN(n_257_76_941));
   INV_X1 i_257_76_943 (.A(n_257_76_941), .ZN(n_257_76_942));
   NAND3_X1 i_257_76_944 (.A1(n_257_76_630), .A2(n_257_76_725), .A3(n_257_76_942), 
      .ZN(n_257_76_943));
   INV_X1 i_257_76_945 (.A(n_257_76_943), .ZN(n_257_76_944));
   NAND4_X1 i_257_76_946 (.A1(n_257_76_924), .A2(n_257_76_931), .A3(n_257_76_944), 
      .A4(n_257_76_724), .ZN(n_257_76_945));
   NAND2_X1 i_257_76_947 (.A1(n_257_350), .A2(n_257_421), .ZN(n_257_76_946));
   NAND3_X1 i_257_76_948 (.A1(n_257_76_731), .A2(n_257_76_634), .A3(n_257_76_946), 
      .ZN(n_257_76_947));
   NOR2_X1 i_257_76_949 (.A1(n_257_76_945), .A2(n_257_76_947), .ZN(n_257_76_948));
   NAND2_X1 i_257_76_950 (.A1(n_257_76_610), .A2(n_257_76_730), .ZN(n_257_76_949));
   INV_X1 i_257_76_951 (.A(n_257_76_949), .ZN(n_257_76_950));
   NAND3_X1 i_257_76_952 (.A1(n_257_76_948), .A2(n_257_76_950), .A3(n_257_76_622), 
      .ZN(n_257_76_951));
   INV_X1 i_257_76_953 (.A(n_257_76_951), .ZN(n_257_76_952));
   NAND2_X1 i_257_76_954 (.A1(n_257_382), .A2(n_257_76_952), .ZN(n_257_76_953));
   NAND4_X1 i_257_76_955 (.A1(n_257_114), .A2(n_257_76_635), .A3(n_257_76_636), 
      .A4(n_257_76_637), .ZN(n_257_76_954));
   INV_X1 i_257_76_956 (.A(n_257_76_954), .ZN(n_257_76_955));
   NAND2_X1 i_257_76_957 (.A1(n_257_430), .A2(n_257_76_612), .ZN(n_257_76_956));
   INV_X1 i_257_76_958 (.A(n_257_76_956), .ZN(n_257_76_957));
   NAND2_X1 i_257_76_959 (.A1(n_257_76_707), .A2(n_257_76_957), .ZN(n_257_76_958));
   INV_X1 i_257_76_960 (.A(n_257_76_958), .ZN(n_257_76_959));
   NAND3_X1 i_257_76_961 (.A1(n_257_76_640), .A2(n_257_76_641), .A3(n_257_76_959), 
      .ZN(n_257_76_960));
   INV_X1 i_257_76_962 (.A(n_257_76_960), .ZN(n_257_76_961));
   NAND4_X1 i_257_76_963 (.A1(n_257_76_961), .A2(n_257_76_651), .A3(n_257_76_638), 
      .A4(n_257_76_652), .ZN(n_257_76_962));
   INV_X1 i_257_76_964 (.A(n_257_76_962), .ZN(n_257_76_963));
   NAND3_X1 i_257_76_965 (.A1(n_257_76_955), .A2(n_257_76_880), .A3(n_257_76_963), 
      .ZN(n_257_76_964));
   NAND3_X1 i_257_76_966 (.A1(n_257_76_630), .A2(n_257_76_631), .A3(n_257_76_627), 
      .ZN(n_257_76_965));
   INV_X1 i_257_76_967 (.A(n_257_76_965), .ZN(n_257_76_966));
   NAND2_X1 i_257_76_968 (.A1(n_257_76_966), .A2(n_257_76_724), .ZN(n_257_76_967));
   NOR2_X1 i_257_76_969 (.A1(n_257_76_964), .A2(n_257_76_967), .ZN(n_257_76_968));
   NAND3_X1 i_257_76_970 (.A1(n_257_76_968), .A2(n_257_76_610), .A3(n_257_76_634), 
      .ZN(n_257_76_969));
   NOR2_X1 i_257_76_971 (.A1(n_257_76_969), .A2(n_257_76_626), .ZN(n_257_76_970));
   NAND2_X1 i_257_76_972 (.A1(n_257_145), .A2(n_257_76_970), .ZN(n_257_76_971));
   NAND3_X1 i_257_76_973 (.A1(n_257_76_921), .A2(n_257_76_953), .A3(n_257_76_971), 
      .ZN(n_257_76_972));
   INV_X1 i_257_76_974 (.A(n_257_76_972), .ZN(n_257_76_973));
   INV_X1 i_257_76_975 (.A(n_257_766), .ZN(n_257_76_974));
   NOR2_X1 i_257_76_976 (.A1(n_257_76_613), .A2(n_257_76_974), .ZN(n_257_76_975));
   NAND3_X1 i_257_76_977 (.A1(n_257_76_640), .A2(n_257_76_641), .A3(n_257_76_975), 
      .ZN(n_257_76_976));
   INV_X1 i_257_76_978 (.A(n_257_76_976), .ZN(n_257_76_977));
   NAND2_X1 i_257_76_979 (.A1(n_257_447), .A2(n_257_76_648), .ZN(n_257_76_978));
   INV_X1 i_257_76_980 (.A(n_257_76_978), .ZN(n_257_76_979));
   NAND3_X1 i_257_76_981 (.A1(n_257_76_977), .A2(n_257_76_979), .A3(n_257_76_636), 
      .ZN(n_257_76_980));
   NOR2_X1 i_257_76_982 (.A1(n_257_76_629), .A2(n_257_76_980), .ZN(n_257_76_981));
   NAND2_X1 i_257_76_983 (.A1(n_257_76_610), .A2(n_257_76_981), .ZN(n_257_76_982));
   INV_X1 i_257_76_984 (.A(n_257_76_982), .ZN(n_257_76_983));
   NAND2_X1 i_257_76_985 (.A1(n_257_76_983), .A2(n_257_76_622), .ZN(n_257_76_984));
   INV_X1 i_257_76_986 (.A(n_257_76_984), .ZN(n_257_76_985));
   NAND3_X1 i_257_76_987 (.A1(n_257_449), .A2(n_257_76_648), .A3(n_257_76_649), 
      .ZN(n_257_76_986));
   NAND2_X1 i_257_76_988 (.A1(n_257_1074), .A2(n_257_76_612), .ZN(n_257_76_987));
   INV_X1 i_257_76_989 (.A(n_257_76_987), .ZN(n_257_76_988));
   NAND3_X1 i_257_76_990 (.A1(n_257_76_640), .A2(n_257_76_641), .A3(n_257_76_988), 
      .ZN(n_257_76_989));
   NOR2_X1 i_257_76_991 (.A1(n_257_76_986), .A2(n_257_76_989), .ZN(n_257_76_990));
   NAND3_X1 i_257_76_992 (.A1(n_257_76_990), .A2(n_257_76_749), .A3(n_257_76_628), 
      .ZN(n_257_76_991));
   INV_X1 i_257_76_993 (.A(n_257_76_991), .ZN(n_257_76_992));
   INV_X1 i_257_76_994 (.A(n_257_76_757), .ZN(n_257_76_993));
   NAND2_X1 i_257_76_995 (.A1(n_257_76_992), .A2(n_257_76_993), .ZN(n_257_76_994));
   NOR2_X1 i_257_76_996 (.A1(n_257_76_994), .A2(n_257_76_674), .ZN(n_257_76_995));
   NAND2_X1 i_257_76_997 (.A1(n_257_76_995), .A2(n_257_76_610), .ZN(n_257_76_996));
   NOR2_X1 i_257_76_998 (.A1(n_257_76_996), .A2(n_257_76_626), .ZN(n_257_76_997));
   AOI22_X1 i_257_76_999 (.A1(n_257_23), .A2(n_257_76_985), .B1(n_257_27), 
      .B2(n_257_76_997), .ZN(n_257_76_998));
   NAND3_X1 i_257_76_1000 (.A1(n_257_76_909), .A2(n_257_76_973), .A3(
      n_257_76_998), .ZN(n_257_76_999));
   NAND2_X1 i_257_76_1001 (.A1(n_257_76_17760), .A2(n_257_76_612), .ZN(
      n_257_76_1000));
   OAI21_X1 i_257_76_1002 (.A(n_257_76_1000), .B1(n_257_702), .B2(n_257_76_613), 
      .ZN(n_257_76_1001));
   NAND2_X1 i_257_76_1003 (.A1(n_257_76_638), .A2(n_257_76_1001), .ZN(
      n_257_76_1002));
   INV_X1 i_257_76_1004 (.A(n_257_76_1002), .ZN(n_257_76_1003));
   NAND4_X1 i_257_76_1005 (.A1(n_257_76_648), .A2(n_257_76_640), .A3(n_257_448), 
      .A4(n_257_76_641), .ZN(n_257_76_1004));
   INV_X1 i_257_76_1006 (.A(n_257_76_1004), .ZN(n_257_76_1005));
   NAND4_X1 i_257_76_1007 (.A1(n_257_76_1003), .A2(n_257_76_1005), .A3(
      n_257_76_628), .A4(n_257_76_636), .ZN(n_257_76_1006));
   INV_X1 i_257_76_1008 (.A(n_257_76_1006), .ZN(n_257_76_1007));
   NAND3_X1 i_257_76_1009 (.A1(n_257_76_1007), .A2(n_257_670), .A3(n_257_76_993), 
      .ZN(n_257_76_1008));
   INV_X1 i_257_76_1010 (.A(n_257_76_1008), .ZN(n_257_76_1009));
   NAND2_X1 i_257_76_1011 (.A1(n_257_76_610), .A2(n_257_76_1009), .ZN(
      n_257_76_1010));
   INV_X1 i_257_76_1012 (.A(n_257_76_1010), .ZN(n_257_76_1011));
   NAND2_X1 i_257_76_1013 (.A1(n_257_76_1011), .A2(n_257_76_622), .ZN(
      n_257_76_1012));
   INV_X1 i_257_76_1014 (.A(n_257_76_1012), .ZN(n_257_76_1013));
   NAND2_X1 i_257_76_1015 (.A1(n_257_26), .A2(n_257_76_1013), .ZN(n_257_76_1014));
   NAND2_X1 i_257_76_1016 (.A1(n_257_76_622), .A2(n_257_76_610), .ZN(
      n_257_76_1015));
   NAND2_X1 i_257_76_1017 (.A1(n_257_425), .A2(n_257_76_612), .ZN(n_257_76_1016));
   INV_X1 i_257_76_1018 (.A(n_257_76_1016), .ZN(n_257_76_1017));
   NAND3_X1 i_257_76_1019 (.A1(n_257_76_1017), .A2(n_257_76_707), .A3(
      n_257_76_708), .ZN(n_257_76_1018));
   INV_X1 i_257_76_1020 (.A(n_257_76_1018), .ZN(n_257_76_1019));
   NAND4_X1 i_257_76_1021 (.A1(n_257_76_649), .A2(n_257_76_640), .A3(
      n_257_76_641), .A4(n_257_76_1019), .ZN(n_257_76_1020));
   NAND3_X1 i_257_76_1022 (.A1(n_257_76_652), .A2(n_257_76_702), .A3(
      n_257_76_648), .ZN(n_257_76_1021));
   NOR2_X1 i_257_76_1023 (.A1(n_257_76_1020), .A2(n_257_76_1021), .ZN(
      n_257_76_1022));
   NAND2_X1 i_257_76_1024 (.A1(n_257_76_635), .A2(n_257_76_715), .ZN(
      n_257_76_1023));
   INV_X1 i_257_76_1025 (.A(n_257_76_1023), .ZN(n_257_76_1024));
   NAND3_X1 i_257_76_1026 (.A1(n_257_76_1022), .A2(n_257_76_828), .A3(
      n_257_76_1024), .ZN(n_257_76_1025));
   NOR2_X1 i_257_76_1027 (.A1(n_257_76_1025), .A2(n_257_76_671), .ZN(
      n_257_76_1026));
   NAND3_X1 i_257_76_1028 (.A1(n_257_233), .A2(n_257_76_724), .A3(n_257_76_727), 
      .ZN(n_257_76_1027));
   INV_X1 i_257_76_1029 (.A(n_257_76_1027), .ZN(n_257_76_1028));
   NAND4_X1 i_257_76_1030 (.A1(n_257_76_1026), .A2(n_257_76_1028), .A3(
      n_257_76_731), .A4(n_257_76_634), .ZN(n_257_76_1029));
   NOR2_X1 i_257_76_1031 (.A1(n_257_76_1015), .A2(n_257_76_1029), .ZN(
      n_257_76_1030));
   NAND2_X1 i_257_76_1032 (.A1(n_257_264), .A2(n_257_76_1030), .ZN(n_257_76_1031));
   NAND3_X1 i_257_76_1033 (.A1(n_257_76_934), .A2(n_257_76_652), .A3(
      n_257_76_702), .ZN(n_257_76_1032));
   NAND3_X1 i_257_76_1034 (.A1(n_257_76_648), .A2(n_257_76_649), .A3(
      n_257_76_640), .ZN(n_257_76_1033));
   NAND2_X1 i_257_76_1035 (.A1(n_257_421), .A2(n_257_76_612), .ZN(n_257_76_1034));
   INV_X1 i_257_76_1036 (.A(n_257_76_1034), .ZN(n_257_76_1035));
   NAND3_X1 i_257_76_1037 (.A1(n_257_76_1035), .A2(n_257_76_707), .A3(
      n_257_76_708), .ZN(n_257_76_1036));
   INV_X1 i_257_76_1038 (.A(n_257_76_1036), .ZN(n_257_76_1037));
   NAND3_X1 i_257_76_1039 (.A1(n_257_76_641), .A2(n_257_76_1037), .A3(
      n_257_76_711), .ZN(n_257_76_1038));
   NOR3_X1 i_257_76_1040 (.A1(n_257_76_1032), .A2(n_257_76_1033), .A3(
      n_257_76_1038), .ZN(n_257_76_1039));
   INV_X1 i_257_76_1041 (.A(n_257_76_923), .ZN(n_257_76_1040));
   INV_X1 i_257_76_1042 (.A(n_257_76_925), .ZN(n_257_76_1041));
   NAND3_X1 i_257_76_1043 (.A1(n_257_76_1039), .A2(n_257_76_1040), .A3(
      n_257_76_1041), .ZN(n_257_76_1042));
   NAND3_X1 i_257_76_1044 (.A1(n_257_76_993), .A2(n_257_76_727), .A3(n_257_350), 
      .ZN(n_257_76_1043));
   NOR2_X1 i_257_76_1045 (.A1(n_257_76_1042), .A2(n_257_76_1043), .ZN(
      n_257_76_1044));
   NAND2_X1 i_257_76_1046 (.A1(n_257_76_730), .A2(n_257_76_731), .ZN(
      n_257_76_1045));
   INV_X1 i_257_76_1047 (.A(n_257_76_1045), .ZN(n_257_76_1046));
   NAND2_X1 i_257_76_1048 (.A1(n_257_76_634), .A2(n_257_76_724), .ZN(
      n_257_76_1047));
   INV_X1 i_257_76_1049 (.A(n_257_76_1047), .ZN(n_257_76_1048));
   NAND3_X1 i_257_76_1050 (.A1(n_257_76_1044), .A2(n_257_76_1046), .A3(
      n_257_76_1048), .ZN(n_257_76_1049));
   NOR2_X1 i_257_76_1051 (.A1(n_257_76_1049), .A2(n_257_76_1015), .ZN(
      n_257_76_1050));
   NAND2_X1 i_257_76_1052 (.A1(n_257_381), .A2(n_257_76_1050), .ZN(n_257_76_1051));
   NAND3_X1 i_257_76_1053 (.A1(n_257_76_1014), .A2(n_257_76_1031), .A3(
      n_257_76_1051), .ZN(n_257_76_1052));
   INV_X1 i_257_76_1054 (.A(n_257_76_1052), .ZN(n_257_76_1053));
   NAND4_X1 i_257_76_1055 (.A1(n_257_193), .A2(n_257_76_938), .A3(n_257_427), 
      .A4(n_257_76_707), .ZN(n_257_76_1054));
   INV_X1 i_257_76_1056 (.A(n_257_76_1054), .ZN(n_257_76_1055));
   NAND4_X1 i_257_76_1057 (.A1(n_257_76_635), .A2(n_257_76_1055), .A3(
      n_257_76_636), .A4(n_257_76_637), .ZN(n_257_76_1056));
   NAND4_X1 i_257_76_1058 (.A1(n_257_76_651), .A2(n_257_76_929), .A3(
      n_257_76_638), .A4(n_257_76_652), .ZN(n_257_76_1057));
   NOR2_X1 i_257_76_1059 (.A1(n_257_76_1056), .A2(n_257_76_1057), .ZN(
      n_257_76_1058));
   INV_X1 i_257_76_1060 (.A(n_257_76_629), .ZN(n_257_76_1059));
   NAND4_X1 i_257_76_1061 (.A1(n_257_76_1058), .A2(n_257_76_777), .A3(
      n_257_76_724), .A4(n_257_76_1059), .ZN(n_257_76_1060));
   NOR2_X1 i_257_76_1062 (.A1(n_257_76_1060), .A2(n_257_76_779), .ZN(
      n_257_76_1061));
   NAND3_X1 i_257_76_1063 (.A1(n_257_76_1061), .A2(n_257_76_622), .A3(
      n_257_76_610), .ZN(n_257_76_1062));
   INV_X1 i_257_76_1064 (.A(n_257_76_1062), .ZN(n_257_76_1063));
   NAND2_X1 i_257_76_1065 (.A1(n_257_224), .A2(n_257_76_1063), .ZN(n_257_76_1064));
   NAND2_X1 i_257_76_1066 (.A1(n_257_453), .A2(n_257_76_612), .ZN(n_257_76_1065));
   INV_X1 i_257_76_1067 (.A(n_257_76_1065), .ZN(n_257_76_1066));
   NAND3_X1 i_257_76_1068 (.A1(n_257_76_640), .A2(n_257_76_641), .A3(
      n_257_76_1066), .ZN(n_257_76_1067));
   INV_X1 i_257_76_1069 (.A(n_257_76_1067), .ZN(n_257_76_1068));
   NAND3_X1 i_257_76_1070 (.A1(n_257_76_1068), .A2(n_257_76_651), .A3(
      n_257_76_652), .ZN(n_257_76_1069));
   NOR2_X1 i_257_76_1071 (.A1(n_257_76_1069), .A2(n_257_76_721), .ZN(
      n_257_76_1070));
   NAND3_X1 i_257_76_1072 (.A1(n_257_76_611), .A2(n_257_76_628), .A3(n_257_451), 
      .ZN(n_257_76_1071));
   INV_X1 i_257_76_1073 (.A(n_257_76_1071), .ZN(n_257_76_1072));
   NAND3_X1 i_257_76_1074 (.A1(n_257_76_1070), .A2(n_257_76_1072), .A3(
      n_257_76_821), .ZN(n_257_76_1073));
   NOR2_X1 i_257_76_1075 (.A1(n_257_76_1073), .A2(n_257_76_674), .ZN(
      n_257_76_1074));
   NAND2_X1 i_257_76_1076 (.A1(n_257_76_610), .A2(n_257_76_1074), .ZN(
      n_257_76_1075));
   NOR2_X1 i_257_76_1077 (.A1(n_257_76_1075), .A2(n_257_76_626), .ZN(
      n_257_76_1076));
   NAND2_X1 i_257_76_1078 (.A1(n_257_434), .A2(n_257_76_1076), .ZN(n_257_76_1077));
   NAND2_X1 i_257_76_1079 (.A1(n_257_76_627), .A2(n_257_76_611), .ZN(
      n_257_76_1078));
   NOR2_X1 i_257_76_1080 (.A1(n_257_76_716), .A2(n_257_76_1078), .ZN(
      n_257_76_1079));
   NAND4_X1 i_257_76_1081 (.A1(n_257_502), .A2(n_257_76_938), .A3(n_257_76_707), 
      .A4(n_257_424), .ZN(n_257_76_1080));
   INV_X1 i_257_76_1082 (.A(n_257_76_1080), .ZN(n_257_76_1081));
   NAND2_X1 i_257_76_1083 (.A1(n_257_76_652), .A2(n_257_76_1081), .ZN(
      n_257_76_1082));
   INV_X1 i_257_76_1084 (.A(n_257_76_1082), .ZN(n_257_76_1083));
   NAND3_X1 i_257_76_1085 (.A1(n_257_76_649), .A2(n_257_76_640), .A3(
      n_257_76_641), .ZN(n_257_76_1084));
   INV_X1 i_257_76_1086 (.A(n_257_76_1084), .ZN(n_257_76_1085));
   NAND2_X1 i_257_76_1087 (.A1(n_257_76_702), .A2(n_257_76_648), .ZN(
      n_257_76_1086));
   INV_X1 i_257_76_1088 (.A(n_257_76_1086), .ZN(n_257_76_1087));
   NAND3_X1 i_257_76_1089 (.A1(n_257_76_1083), .A2(n_257_76_1085), .A3(
      n_257_76_1087), .ZN(n_257_76_1088));
   NOR2_X1 i_257_76_1090 (.A1(n_257_76_1088), .A2(n_257_76_721), .ZN(
      n_257_76_1089));
   NAND4_X1 i_257_76_1091 (.A1(n_257_76_1079), .A2(n_257_76_1089), .A3(
      n_257_76_777), .A4(n_257_76_724), .ZN(n_257_76_1090));
   NOR2_X1 i_257_76_1092 (.A1(n_257_76_1090), .A2(n_257_76_779), .ZN(
      n_257_76_1091));
   NAND3_X1 i_257_76_1093 (.A1(n_257_76_1091), .A2(n_257_76_950), .A3(
      n_257_76_622), .ZN(n_257_76_1092));
   INV_X1 i_257_76_1094 (.A(n_257_76_1092), .ZN(n_257_76_1093));
   NAND2_X1 i_257_76_1095 (.A1(n_257_265), .A2(n_257_76_1093), .ZN(n_257_76_1094));
   NAND3_X1 i_257_76_1096 (.A1(n_257_76_1064), .A2(n_257_76_1077), .A3(
      n_257_76_1094), .ZN(n_257_76_1095));
   INV_X1 i_257_76_1097 (.A(n_257_76_1095), .ZN(n_257_76_1096));
   INV_X1 i_257_76_1098 (.A(n_257_76_724), .ZN(n_257_76_1097));
   NAND4_X1 i_257_76_1099 (.A1(n_257_76_630), .A2(n_257_76_725), .A3(
      n_257_76_631), .A4(n_257_76_627), .ZN(n_257_76_1098));
   NOR2_X1 i_257_76_1100 (.A1(n_257_76_1097), .A2(n_257_76_1098), .ZN(
      n_257_76_1099));
   NOR2_X1 i_257_76_1101 (.A1(n_257_76_1021), .A2(n_257_76_1084), .ZN(
      n_257_76_1100));
   NAND3_X1 i_257_76_1102 (.A1(n_257_76_1100), .A2(n_257_76_828), .A3(
      n_257_76_1024), .ZN(n_257_76_1101));
   NAND3_X1 i_257_76_1103 (.A1(n_257_76_938), .A2(n_257_76_707), .A3(n_257_422), 
      .ZN(n_257_76_1102));
   INV_X1 i_257_76_1104 (.A(n_257_76_1102), .ZN(n_257_76_1103));
   NAND3_X1 i_257_76_1105 (.A1(n_257_76_1103), .A2(n_257_311), .A3(n_257_76_711), 
      .ZN(n_257_76_1104));
   INV_X1 i_257_76_1106 (.A(n_257_76_1104), .ZN(n_257_76_1105));
   NAND4_X1 i_257_76_1107 (.A1(n_257_76_611), .A2(n_257_76_628), .A3(
      n_257_76_922), .A4(n_257_76_1105), .ZN(n_257_76_1106));
   NOR2_X1 i_257_76_1108 (.A1(n_257_76_1101), .A2(n_257_76_1106), .ZN(
      n_257_76_1107));
   NAND4_X1 i_257_76_1109 (.A1(n_257_76_1099), .A2(n_257_76_1107), .A3(
      n_257_76_731), .A4(n_257_76_634), .ZN(n_257_76_1108));
   INV_X1 i_257_76_1110 (.A(n_257_76_1108), .ZN(n_257_76_1109));
   NAND3_X1 i_257_76_1111 (.A1(n_257_76_1109), .A2(n_257_76_950), .A3(
      n_257_76_622), .ZN(n_257_76_1110));
   INV_X1 i_257_76_1112 (.A(n_257_76_1110), .ZN(n_257_76_1111));
   NAND2_X1 i_257_76_1113 (.A1(n_257_342), .A2(n_257_76_1111), .ZN(n_257_76_1112));
   AOI21_X1 i_257_76_1114 (.A(n_257_76_718), .B1(n_257_996), .B2(n_257_76_17964), 
      .ZN(n_257_76_1113));
   NAND2_X1 i_257_76_1115 (.A1(n_257_1028), .A2(n_257_76_17969), .ZN(
      n_257_76_1114));
   NAND2_X1 i_257_76_1116 (.A1(n_257_76_1113), .A2(n_257_76_1114), .ZN(
      n_257_76_1115));
   INV_X1 i_257_76_1117 (.A(n_257_76_1115), .ZN(n_257_76_1116));
   NAND2_X1 i_257_76_1118 (.A1(n_257_453), .A2(n_257_442), .ZN(n_257_76_1117));
   INV_X1 i_257_76_1119 (.A(n_257_76_1117), .ZN(n_257_76_1118));
   NAND2_X1 i_257_76_1120 (.A1(n_257_451), .A2(n_257_76_1118), .ZN(n_257_76_1119));
   NAND2_X1 i_257_76_1121 (.A1(n_257_114), .A2(n_257_76_17925), .ZN(
      n_257_76_1120));
   NAND2_X1 i_257_76_1122 (.A1(n_257_76_1119), .A2(n_257_76_1120), .ZN(
      n_257_76_1121));
   NAND2_X1 i_257_76_1123 (.A1(n_257_734), .A2(n_257_76_17935), .ZN(
      n_257_76_1122));
   NAND2_X1 i_257_76_1124 (.A1(n_257_862), .A2(n_257_76_17903), .ZN(
      n_257_76_1123));
   NAND2_X1 i_257_76_1125 (.A1(n_257_76_1122), .A2(n_257_76_1123), .ZN(
      n_257_76_1124));
   NOR2_X1 i_257_76_1126 (.A1(n_257_76_1121), .A2(n_257_76_1124), .ZN(
      n_257_76_1125));
   NAND2_X1 i_257_76_1127 (.A1(n_257_76), .A2(n_257_76_17932), .ZN(n_257_76_1126));
   NAND2_X1 i_257_76_1128 (.A1(n_257_76_1125), .A2(n_257_76_1126), .ZN(
      n_257_76_1127));
   INV_X1 i_257_76_1129 (.A(n_257_76_1127), .ZN(n_257_76_1128));
   NAND2_X1 i_257_76_1130 (.A1(n_257_964), .A2(n_257_442), .ZN(n_257_76_1129));
   INV_X1 i_257_76_1131 (.A(n_257_76_1129), .ZN(n_257_76_1130));
   NAND2_X1 i_257_76_1132 (.A1(n_257_441), .A2(n_257_76_1130), .ZN(n_257_76_1131));
   NAND2_X1 i_257_76_1133 (.A1(n_257_76_1131), .A2(n_257_76_941), .ZN(
      n_257_76_1132));
   INV_X1 i_257_76_1134 (.A(n_257_76_1132), .ZN(n_257_76_1133));
   NAND2_X1 i_257_76_1135 (.A1(n_257_36), .A2(n_257_76_17918), .ZN(n_257_76_1134));
   NAND2_X1 i_257_76_1136 (.A1(n_257_76_1134), .A2(n_257_76_1104), .ZN(
      n_257_76_1135));
   NAND2_X1 i_257_76_1137 (.A1(n_257_798), .A2(n_257_76_17952), .ZN(
      n_257_76_1136));
   INV_X1 i_257_76_1138 (.A(n_257_76_1136), .ZN(n_257_76_1137));
   NOR2_X1 i_257_76_1139 (.A1(n_257_76_1135), .A2(n_257_76_1137), .ZN(
      n_257_76_1138));
   NAND2_X1 i_257_76_1140 (.A1(n_257_76_1133), .A2(n_257_76_1138), .ZN(
      n_257_76_1139));
   NAND3_X1 i_257_76_1141 (.A1(n_257_439), .A2(n_257_900), .A3(n_257_442), 
      .ZN(n_257_76_1140));
   NAND2_X1 i_257_76_1142 (.A1(n_257_76_1080), .A2(n_257_76_1140), .ZN(
      n_257_76_1141));
   NAND2_X1 i_257_76_1143 (.A1(n_257_630), .A2(n_257_76_17928), .ZN(
      n_257_76_1142));
   INV_X1 i_257_76_1144 (.A(n_257_76_1142), .ZN(n_257_76_1143));
   NOR2_X1 i_257_76_1145 (.A1(n_257_76_1141), .A2(n_257_76_1143), .ZN(
      n_257_76_1144));
   NAND2_X1 i_257_76_1146 (.A1(n_257_438), .A2(n_257_76_4359), .ZN(n_257_76_1145));
   NAND2_X1 i_257_76_1147 (.A1(n_257_598), .A2(n_257_442), .ZN(n_257_76_1146));
   INV_X1 i_257_76_1148 (.A(n_257_76_1146), .ZN(n_257_76_1147));
   NAND2_X1 i_257_76_1149 (.A1(n_257_432), .A2(n_257_76_1147), .ZN(n_257_76_1148));
   NAND2_X1 i_257_76_1150 (.A1(n_257_76_1148), .A2(n_257_76_766), .ZN(
      n_257_76_1149));
   NAND3_X1 i_257_76_1151 (.A1(n_257_76_612), .A2(n_257_389), .A3(n_257_484), 
      .ZN(n_257_76_1150));
   INV_X1 i_257_76_1152 (.A(Small_Packet_Data_Size[1]), .ZN(n_257_76_1151));
   NAND2_X1 i_257_76_1153 (.A1(n_257_76_1150), .A2(n_257_76_18058), .ZN(
      n_257_76_1152));
   NOR2_X1 i_257_76_1154 (.A1(n_257_76_1149), .A2(n_257_76_1152), .ZN(
      n_257_76_1153));
   NAND2_X1 i_257_76_1155 (.A1(n_257_76_1145), .A2(n_257_76_1153), .ZN(
      n_257_76_1154));
   NAND2_X1 i_257_76_1156 (.A1(n_257_442), .A2(n_257_932), .ZN(n_257_76_1155));
   INV_X1 i_257_76_1157 (.A(n_257_76_1155), .ZN(n_257_76_1156));
   NAND2_X1 i_257_76_1158 (.A1(n_257_440), .A2(n_257_76_1156), .ZN(n_257_76_1157));
   NAND2_X1 i_257_76_1159 (.A1(n_257_702), .A2(n_257_76_15655), .ZN(
      n_257_76_1158));
   NAND2_X1 i_257_76_1160 (.A1(n_257_76_1157), .A2(n_257_76_1158), .ZN(
      n_257_76_1159));
   NOR2_X1 i_257_76_1161 (.A1(n_257_76_1154), .A2(n_257_76_1159), .ZN(
      n_257_76_1160));
   NAND2_X1 i_257_76_1162 (.A1(n_257_76_1144), .A2(n_257_76_1160), .ZN(
      n_257_76_1161));
   INV_X1 i_257_76_1163 (.A(n_257_76_1161), .ZN(n_257_76_1162));
   NAND2_X1 i_257_76_1164 (.A1(n_257_830), .A2(n_257_442), .ZN(n_257_76_1163));
   INV_X1 i_257_76_1165 (.A(n_257_76_1163), .ZN(n_257_76_1164));
   NAND2_X1 i_257_76_1166 (.A1(n_257_446), .A2(n_257_76_1164), .ZN(n_257_76_1165));
   NAND2_X1 i_257_76_1167 (.A1(n_257_449), .A2(n_257_76_8828), .ZN(n_257_76_1166));
   NAND2_X1 i_257_76_1168 (.A1(n_257_76_1165), .A2(n_257_76_1166), .ZN(
      n_257_76_1167));
   NAND2_X1 i_257_76_1169 (.A1(n_257_766), .A2(n_257_442), .ZN(n_257_76_1168));
   INV_X1 i_257_76_1170 (.A(n_257_76_1168), .ZN(n_257_76_1169));
   NAND2_X1 i_257_76_1171 (.A1(n_257_447), .A2(n_257_76_1169), .ZN(n_257_76_1170));
   NAND2_X1 i_257_76_1172 (.A1(n_257_76_1170), .A2(n_257_76_1054), .ZN(
      n_257_76_1171));
   NOR2_X1 i_257_76_1173 (.A1(n_257_76_1167), .A2(n_257_76_1171), .ZN(
      n_257_76_1172));
   NAND2_X1 i_257_76_1174 (.A1(n_257_76_1162), .A2(n_257_76_1172), .ZN(
      n_257_76_1173));
   NOR2_X1 i_257_76_1175 (.A1(n_257_76_1139), .A2(n_257_76_1173), .ZN(
      n_257_76_1174));
   NAND2_X1 i_257_76_1176 (.A1(n_257_76_1128), .A2(n_257_76_1174), .ZN(
      n_257_76_1175));
   AOI22_X1 i_257_76_1177 (.A1(n_257_153), .A2(n_257_76_17331), .B1(n_257_670), 
      .B2(n_257_76_17958), .ZN(n_257_76_1176));
   NAND2_X1 i_257_76_1178 (.A1(n_257_76_1176), .A2(n_257_76_824), .ZN(
      n_257_76_1177));
   NOR2_X1 i_257_76_1179 (.A1(n_257_76_1175), .A2(n_257_76_1177), .ZN(
      n_257_76_1178));
   NAND2_X1 i_257_76_1180 (.A1(n_257_76_1116), .A2(n_257_76_1178), .ZN(
      n_257_76_1179));
   NAND2_X1 i_257_76_1181 (.A1(n_257_76_1049), .A2(n_257_76_1029), .ZN(
      n_257_76_1180));
   NOR2_X1 i_257_76_1182 (.A1(n_257_76_1179), .A2(n_257_76_1180), .ZN(
      n_257_76_1181));
   NAND2_X1 i_257_76_1183 (.A1(n_257_76_634), .A2(n_257_76_946), .ZN(
      n_257_76_1182));
   NOR2_X1 i_257_76_1184 (.A1(n_257_76_1045), .A2(n_257_76_1182), .ZN(
      n_257_76_1183));
   NAND2_X1 i_257_76_1185 (.A1(n_257_76_1024), .A2(n_257_76_922), .ZN(
      n_257_76_1184));
   NOR2_X1 i_257_76_1186 (.A1(n_257_76_1184), .A2(n_257_76_879), .ZN(
      n_257_76_1185));
   NAND2_X1 i_257_76_1187 (.A1(n_257_76_934), .A2(n_257_76_652), .ZN(
      n_257_76_1186));
   INV_X1 i_257_76_1188 (.A(n_257_76_638), .ZN(n_257_76_1187));
   NOR2_X1 i_257_76_1189 (.A1(n_257_76_1186), .A2(n_257_76_1187), .ZN(
      n_257_76_1188));
   NAND2_X1 i_257_76_1190 (.A1(n_257_76_666), .A2(n_257_76_1188), .ZN(
      n_257_76_1189));
   NOR2_X1 i_257_76_1191 (.A1(n_257_76_1086), .A2(n_257_76_663), .ZN(
      n_257_76_1190));
   INV_X1 i_257_76_1192 (.A(n_257_76_1150), .ZN(n_257_76_1191));
   NAND2_X1 i_257_76_1193 (.A1(n_257_76_708), .A2(n_257_76_1191), .ZN(
      n_257_76_1192));
   INV_X1 i_257_76_1194 (.A(n_257_76_707), .ZN(n_257_76_1193));
   NOR2_X1 i_257_76_1195 (.A1(n_257_76_1192), .A2(n_257_76_1193), .ZN(
      n_257_76_1194));
   NAND2_X1 i_257_76_1196 (.A1(n_257_76_711), .A2(n_257_76_1194), .ZN(
      n_257_76_1195));
   NAND2_X1 i_257_76_1197 (.A1(n_257_1090), .A2(n_257_420), .ZN(n_257_76_1196));
   NAND2_X1 i_257_76_1198 (.A1(n_257_76_1196), .A2(n_257_76_641), .ZN(
      n_257_76_1197));
   NOR2_X1 i_257_76_1199 (.A1(n_257_76_1195), .A2(n_257_76_1197), .ZN(
      n_257_76_1198));
   NAND2_X1 i_257_76_1200 (.A1(n_257_76_1190), .A2(n_257_76_1198), .ZN(
      n_257_76_1199));
   NOR2_X1 i_257_76_1201 (.A1(n_257_76_1189), .A2(n_257_76_1199), .ZN(
      n_257_76_1200));
   NAND2_X1 i_257_76_1202 (.A1(n_257_76_1185), .A2(n_257_76_1200), .ZN(
      n_257_76_1201));
   NOR2_X1 i_257_76_1203 (.A1(n_257_76_726), .A2(n_257_76_717), .ZN(
      n_257_76_1202));
   NAND2_X1 i_257_76_1204 (.A1(n_257_76_1202), .A2(n_257_76_724), .ZN(
      n_257_76_1203));
   NOR2_X1 i_257_76_1205 (.A1(n_257_76_1201), .A2(n_257_76_1203), .ZN(
      n_257_76_1204));
   NAND2_X1 i_257_76_1206 (.A1(n_257_76_1183), .A2(n_257_76_1204), .ZN(
      n_257_76_1205));
   NOR2_X1 i_257_76_1207 (.A1(n_257_76_1205), .A2(n_257_76_1015), .ZN(
      n_257_76_1206));
   AOI21_X1 i_257_76_1208 (.A(n_257_76_1181), .B1(n_257_12), .B2(n_257_76_1206), 
      .ZN(n_257_76_1207));
   NAND2_X1 i_257_76_1209 (.A1(n_257_76_1112), .A2(n_257_76_1207), .ZN(
      n_257_76_1208));
   INV_X1 i_257_76_1210 (.A(n_257_76_1208), .ZN(n_257_76_1209));
   NAND3_X1 i_257_76_1211 (.A1(n_257_76_1053), .A2(n_257_76_1096), .A3(
      n_257_76_1209), .ZN(n_257_76_1210));
   NOR2_X1 i_257_76_1212 (.A1(n_257_76_999), .A2(n_257_76_1210), .ZN(
      n_257_76_1211));
   NAND2_X1 i_257_76_1213 (.A1(n_257_76_865), .A2(n_257_76_1211), .ZN(n_1));
   NAND2_X1 i_257_76_1214 (.A1(n_257_1029), .A2(n_257_443), .ZN(n_257_76_1212));
   NAND2_X1 i_257_76_1215 (.A1(n_257_997), .A2(n_257_444), .ZN(n_257_76_1213));
   NAND2_X1 i_257_76_1216 (.A1(n_257_441), .A2(n_257_965), .ZN(n_257_76_1214));
   INV_X1 i_257_76_1217 (.A(n_257_1061), .ZN(n_257_76_1215));
   NAND2_X1 i_257_76_1218 (.A1(n_257_442), .A2(n_257_76_1215), .ZN(n_257_76_1216));
   INV_X1 i_257_76_1219 (.A(n_257_933), .ZN(n_257_76_1217));
   NOR2_X1 i_257_76_1220 (.A1(n_257_76_1216), .A2(n_257_76_1217), .ZN(
      n_257_76_1218));
   NAND2_X1 i_257_76_1221 (.A1(n_257_440), .A2(n_257_76_1218), .ZN(n_257_76_1219));
   INV_X1 i_257_76_1222 (.A(n_257_76_1219), .ZN(n_257_76_1220));
   NAND2_X1 i_257_76_1223 (.A1(n_257_76_1214), .A2(n_257_76_1220), .ZN(
      n_257_76_1221));
   INV_X1 i_257_76_1224 (.A(n_257_76_1221), .ZN(n_257_76_1222));
   NAND3_X1 i_257_76_1225 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1222), .ZN(n_257_76_1223));
   INV_X1 i_257_76_1226 (.A(n_257_76_1223), .ZN(n_257_76_1224));
   NAND2_X1 i_257_76_1227 (.A1(n_257_17), .A2(n_257_76_1224), .ZN(n_257_76_1225));
   INV_X1 i_257_76_1228 (.A(n_257_76_1216), .ZN(n_257_76_1226));
   NAND2_X1 i_257_76_1229 (.A1(n_257_443), .A2(n_257_76_1226), .ZN(n_257_76_1227));
   INV_X1 i_257_76_1230 (.A(n_257_76_1227), .ZN(n_257_76_1228));
   NAND2_X1 i_257_76_1231 (.A1(n_257_1029), .A2(n_257_76_1228), .ZN(
      n_257_76_1229));
   INV_X1 i_257_76_1232 (.A(n_257_76_1229), .ZN(n_257_76_1230));
   NAND2_X1 i_257_76_1233 (.A1(n_257_14), .A2(n_257_76_1230), .ZN(n_257_76_1231));
   NAND2_X1 i_257_76_1234 (.A1(n_257_671), .A2(n_257_448), .ZN(n_257_76_1232));
   NAND2_X1 i_257_76_1235 (.A1(n_257_735), .A2(n_257_436), .ZN(n_257_76_1233));
   NAND2_X1 i_257_76_1236 (.A1(n_257_863), .A2(n_257_445), .ZN(n_257_76_1234));
   NAND2_X1 i_257_76_1237 (.A1(n_257_446), .A2(n_257_831), .ZN(n_257_76_1235));
   NAND3_X1 i_257_76_1238 (.A1(n_257_76_1233), .A2(n_257_76_1234), .A3(
      n_257_76_1235), .ZN(n_257_76_1236));
   INV_X1 i_257_76_1239 (.A(n_257_76_1214), .ZN(n_257_76_1237));
   NOR2_X1 i_257_76_1240 (.A1(n_257_76_1236), .A2(n_257_76_1237), .ZN(
      n_257_76_1238));
   NAND2_X1 i_257_76_1241 (.A1(n_257_449), .A2(n_257_1075), .ZN(n_257_76_1239));
   NAND2_X1 i_257_76_1242 (.A1(n_257_447), .A2(n_257_767), .ZN(n_257_76_1240));
   NAND2_X1 i_257_76_1243 (.A1(n_257_799), .A2(n_257_437), .ZN(n_257_76_1241));
   NAND3_X1 i_257_76_1244 (.A1(n_257_76_1239), .A2(n_257_76_1240), .A3(
      n_257_76_1241), .ZN(n_257_76_1242));
   NAND2_X1 i_257_76_1245 (.A1(n_257_703), .A2(n_257_435), .ZN(n_257_76_1243));
   NAND2_X1 i_257_76_1246 (.A1(n_257_450), .A2(n_257_76_1226), .ZN(n_257_76_1244));
   INV_X1 i_257_76_1247 (.A(n_257_76_1244), .ZN(n_257_76_1245));
   NAND3_X1 i_257_76_1248 (.A1(n_257_631), .A2(n_257_76_1243), .A3(n_257_76_1245), 
      .ZN(n_257_76_1246));
   INV_X1 i_257_76_1249 (.A(n_257_76_1246), .ZN(n_257_76_1247));
   NAND2_X1 i_257_76_1250 (.A1(n_257_440), .A2(n_257_933), .ZN(n_257_76_1248));
   NAND2_X1 i_257_76_1251 (.A1(n_257_438), .A2(n_257_1067), .ZN(n_257_76_1249));
   NAND2_X1 i_257_76_1252 (.A1(n_257_439), .A2(n_257_901), .ZN(n_257_76_1250));
   NAND4_X1 i_257_76_1253 (.A1(n_257_76_1247), .A2(n_257_76_1248), .A3(
      n_257_76_1249), .A4(n_257_76_1250), .ZN(n_257_76_1251));
   NOR2_X1 i_257_76_1254 (.A1(n_257_76_1242), .A2(n_257_76_1251), .ZN(
      n_257_76_1252));
   NAND3_X1 i_257_76_1255 (.A1(n_257_76_1232), .A2(n_257_76_1238), .A3(
      n_257_76_1252), .ZN(n_257_76_1253));
   INV_X1 i_257_76_1256 (.A(n_257_76_1253), .ZN(n_257_76_1254));
   NAND3_X1 i_257_76_1257 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1254), .ZN(n_257_76_1255));
   INV_X1 i_257_76_1258 (.A(n_257_76_1255), .ZN(n_257_76_1256));
   NAND2_X1 i_257_76_1259 (.A1(n_257_28), .A2(n_257_76_1256), .ZN(n_257_76_1257));
   NAND3_X1 i_257_76_1260 (.A1(n_257_76_1225), .A2(n_257_76_1231), .A3(
      n_257_76_1257), .ZN(n_257_76_1258));
   NAND3_X1 i_257_76_1261 (.A1(n_257_446), .A2(n_257_76_1248), .A3(n_257_76_1249), 
      .ZN(n_257_76_1259));
   INV_X1 i_257_76_1262 (.A(n_257_76_1259), .ZN(n_257_76_1260));
   NAND2_X1 i_257_76_1263 (.A1(n_257_831), .A2(n_257_76_1226), .ZN(n_257_76_1261));
   INV_X1 i_257_76_1264 (.A(n_257_76_1261), .ZN(n_257_76_1262));
   NAND2_X1 i_257_76_1265 (.A1(n_257_76_1250), .A2(n_257_76_1262), .ZN(
      n_257_76_1263));
   INV_X1 i_257_76_1266 (.A(n_257_76_1263), .ZN(n_257_76_1264));
   NAND4_X1 i_257_76_1267 (.A1(n_257_76_1214), .A2(n_257_76_1260), .A3(
      n_257_76_1234), .A4(n_257_76_1264), .ZN(n_257_76_1265));
   INV_X1 i_257_76_1268 (.A(n_257_76_1265), .ZN(n_257_76_1266));
   NAND3_X1 i_257_76_1269 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1266), .ZN(n_257_76_1267));
   INV_X1 i_257_76_1270 (.A(n_257_76_1267), .ZN(n_257_76_1268));
   NAND2_X1 i_257_76_1271 (.A1(n_257_21), .A2(n_257_76_1268), .ZN(n_257_76_1269));
   INV_X1 i_257_76_1272 (.A(n_257_76_1248), .ZN(n_257_76_1270));
   NAND3_X1 i_257_76_1273 (.A1(n_257_439), .A2(n_257_901), .A3(n_257_76_1226), 
      .ZN(n_257_76_1271));
   NOR2_X1 i_257_76_1274 (.A1(n_257_76_1270), .A2(n_257_76_1271), .ZN(
      n_257_76_1272));
   NAND2_X1 i_257_76_1275 (.A1(n_257_76_1214), .A2(n_257_76_1272), .ZN(
      n_257_76_1273));
   INV_X1 i_257_76_1276 (.A(n_257_76_1273), .ZN(n_257_76_1274));
   NAND3_X1 i_257_76_1277 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1274), .ZN(n_257_76_1275));
   INV_X1 i_257_76_1278 (.A(n_257_76_1275), .ZN(n_257_76_1276));
   NAND2_X1 i_257_76_1279 (.A1(n_257_18), .A2(n_257_76_1276), .ZN(n_257_76_1277));
   NAND2_X1 i_257_76_1280 (.A1(n_257_234), .A2(n_257_425), .ZN(n_257_76_1278));
   NAND2_X1 i_257_76_1281 (.A1(n_257_76_1232), .A2(n_257_76_1278), .ZN(
      n_257_76_1279));
   NAND2_X1 i_257_76_1282 (.A1(n_257_428), .A2(n_257_567), .ZN(n_257_76_1280));
   INV_X1 i_257_76_1283 (.A(n_257_76_1280), .ZN(n_257_76_1281));
   NAND2_X1 i_257_76_1284 (.A1(n_257_423), .A2(n_257_76_1226), .ZN(n_257_76_1282));
   NOR2_X1 i_257_76_1285 (.A1(n_257_76_1281), .A2(n_257_76_1282), .ZN(
      n_257_76_1283));
   NAND2_X1 i_257_76_1286 (.A1(n_257_432), .A2(n_257_599), .ZN(n_257_76_1284));
   NAND3_X1 i_257_76_1287 (.A1(n_257_76_1243), .A2(n_257_76_1283), .A3(
      n_257_76_1284), .ZN(n_257_76_1285));
   INV_X1 i_257_76_1288 (.A(n_257_76_1285), .ZN(n_257_76_1286));
   NAND2_X1 i_257_76_1289 (.A1(n_257_194), .A2(n_257_427), .ZN(n_257_76_1287));
   NAND2_X1 i_257_76_1290 (.A1(n_257_503), .A2(n_257_424), .ZN(n_257_76_1288));
   NAND4_X1 i_257_76_1291 (.A1(n_257_76_1286), .A2(n_257_76_1250), .A3(
      n_257_76_1287), .A4(n_257_76_1288), .ZN(n_257_76_1289));
   NAND2_X1 i_257_76_1292 (.A1(n_257_631), .A2(n_257_450), .ZN(n_257_76_1290));
   NAND3_X1 i_257_76_1293 (.A1(n_257_274), .A2(n_257_76_1249), .A3(n_257_76_1290), 
      .ZN(n_257_76_1291));
   NOR2_X1 i_257_76_1294 (.A1(n_257_76_1289), .A2(n_257_76_1291), .ZN(
      n_257_76_1292));
   NAND2_X1 i_257_76_1295 (.A1(n_257_115), .A2(n_257_430), .ZN(n_257_76_1293));
   NAND3_X1 i_257_76_1296 (.A1(n_257_76_1293), .A2(n_257_76_1233), .A3(
      n_257_76_1234), .ZN(n_257_76_1294));
   INV_X1 i_257_76_1297 (.A(n_257_76_1294), .ZN(n_257_76_1295));
   NAND2_X1 i_257_76_1298 (.A1(n_257_535), .A2(n_257_426), .ZN(n_257_76_1296));
   NAND2_X1 i_257_76_1299 (.A1(n_257_37), .A2(n_257_433), .ZN(n_257_76_1297));
   NAND4_X1 i_257_76_1300 (.A1(n_257_76_1241), .A2(n_257_76_1296), .A3(
      n_257_76_1297), .A4(n_257_76_1248), .ZN(n_257_76_1298));
   INV_X1 i_257_76_1301 (.A(n_257_76_1298), .ZN(n_257_76_1299));
   NAND3_X1 i_257_76_1302 (.A1(n_257_76_1292), .A2(n_257_76_1295), .A3(
      n_257_76_1299), .ZN(n_257_76_1300));
   NOR2_X1 i_257_76_1303 (.A1(n_257_76_1279), .A2(n_257_76_1300), .ZN(
      n_257_76_1301));
   NAND2_X1 i_257_76_1304 (.A1(n_257_451), .A2(n_257_454), .ZN(n_257_76_1302));
   NAND2_X1 i_257_76_1305 (.A1(n_257_76_1214), .A2(n_257_76_1302), .ZN(
      n_257_76_1303));
   NAND3_X1 i_257_76_1306 (.A1(n_257_76_1235), .A2(n_257_76_1239), .A3(
      n_257_76_1240), .ZN(n_257_76_1304));
   NOR2_X1 i_257_76_1307 (.A1(n_257_76_1303), .A2(n_257_76_1304), .ZN(
      n_257_76_1305));
   NAND2_X1 i_257_76_1308 (.A1(n_257_154), .A2(n_257_429), .ZN(n_257_76_1306));
   NAND2_X1 i_257_76_1309 (.A1(n_257_77), .A2(n_257_431), .ZN(n_257_76_1307));
   NAND3_X1 i_257_76_1310 (.A1(n_257_76_1305), .A2(n_257_76_1306), .A3(
      n_257_76_1307), .ZN(n_257_76_1308));
   INV_X1 i_257_76_1311 (.A(n_257_76_1308), .ZN(n_257_76_1309));
   NAND4_X1 i_257_76_1312 (.A1(n_257_76_1212), .A2(n_257_76_1301), .A3(
      n_257_76_1213), .A4(n_257_76_1309), .ZN(n_257_76_1310));
   INV_X1 i_257_76_1313 (.A(n_257_76_1310), .ZN(n_257_76_1311));
   NAND2_X1 i_257_76_1314 (.A1(n_257_304), .A2(n_257_76_1311), .ZN(n_257_76_1312));
   NAND3_X1 i_257_76_1315 (.A1(n_257_76_1269), .A2(n_257_76_1277), .A3(
      n_257_76_1312), .ZN(n_257_76_1313));
   NOR2_X1 i_257_76_1316 (.A1(n_257_76_1258), .A2(n_257_76_1313), .ZN(
      n_257_76_1314));
   NAND2_X1 i_257_76_1317 (.A1(n_257_965), .A2(n_257_76_1226), .ZN(n_257_76_1315));
   INV_X1 i_257_76_1318 (.A(n_257_76_1315), .ZN(n_257_76_1316));
   NAND2_X1 i_257_76_1319 (.A1(n_257_441), .A2(n_257_76_1316), .ZN(n_257_76_1317));
   INV_X1 i_257_76_1320 (.A(n_257_76_1317), .ZN(n_257_76_1318));
   NAND3_X1 i_257_76_1321 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1318), .ZN(n_257_76_1319));
   INV_X1 i_257_76_1322 (.A(n_257_76_1319), .ZN(n_257_76_1320));
   NAND2_X1 i_257_76_1323 (.A1(n_257_16), .A2(n_257_76_1320), .ZN(n_257_76_1321));
   NAND2_X1 i_257_76_1324 (.A1(n_257_76_1248), .A2(n_257_76_1249), .ZN(
      n_257_76_1322));
   INV_X1 i_257_76_1325 (.A(n_257_76_1322), .ZN(n_257_76_1323));
   NAND3_X1 i_257_76_1326 (.A1(n_257_703), .A2(n_257_435), .A3(n_257_76_1226), 
      .ZN(n_257_76_1324));
   INV_X1 i_257_76_1327 (.A(n_257_76_1324), .ZN(n_257_76_1325));
   NAND2_X1 i_257_76_1328 (.A1(n_257_76_1250), .A2(n_257_76_1325), .ZN(
      n_257_76_1326));
   INV_X1 i_257_76_1329 (.A(n_257_76_1326), .ZN(n_257_76_1327));
   NAND4_X1 i_257_76_1330 (.A1(n_257_76_1323), .A2(n_257_76_1240), .A3(
      n_257_76_1241), .A4(n_257_76_1327), .ZN(n_257_76_1328));
   NOR3_X1 i_257_76_1331 (.A1(n_257_76_1328), .A2(n_257_76_1236), .A3(
      n_257_76_1237), .ZN(n_257_76_1329));
   NAND3_X1 i_257_76_1332 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1329), .ZN(n_257_76_1330));
   INV_X1 i_257_76_1333 (.A(n_257_76_1330), .ZN(n_257_76_1331));
   NAND2_X1 i_257_76_1334 (.A1(n_257_25), .A2(n_257_76_1331), .ZN(n_257_76_1332));
   NAND3_X1 i_257_76_1335 (.A1(n_257_76_1232), .A2(n_257_76_1306), .A3(
      n_257_76_1307), .ZN(n_257_76_1333));
   NAND2_X1 i_257_76_1336 (.A1(n_257_76_1233), .A2(n_257_76_1234), .ZN(
      n_257_76_1334));
   NOR2_X1 i_257_76_1337 (.A1(n_257_76_1304), .A2(n_257_76_1334), .ZN(
      n_257_76_1335));
   NAND3_X1 i_257_76_1338 (.A1(n_257_76_1214), .A2(n_257_76_1302), .A3(
      n_257_76_1293), .ZN(n_257_76_1336));
   INV_X1 i_257_76_1339 (.A(n_257_76_1336), .ZN(n_257_76_1337));
   NAND3_X1 i_257_76_1340 (.A1(n_257_76_1297), .A2(n_257_76_1248), .A3(
      n_257_76_1249), .ZN(n_257_76_1338));
   INV_X1 i_257_76_1341 (.A(n_257_76_1338), .ZN(n_257_76_1339));
   NAND3_X1 i_257_76_1342 (.A1(n_257_442), .A2(n_257_567), .A3(n_257_76_1215), 
      .ZN(n_257_76_1340));
   INV_X1 i_257_76_1343 (.A(n_257_76_1340), .ZN(n_257_76_1341));
   NAND2_X1 i_257_76_1344 (.A1(n_257_428), .A2(n_257_76_1341), .ZN(n_257_76_1342));
   INV_X1 i_257_76_1345 (.A(n_257_76_1342), .ZN(n_257_76_1343));
   NAND3_X1 i_257_76_1346 (.A1(n_257_76_1243), .A2(n_257_76_1284), .A3(
      n_257_76_1343), .ZN(n_257_76_1344));
   INV_X1 i_257_76_1347 (.A(n_257_76_1344), .ZN(n_257_76_1345));
   NAND3_X1 i_257_76_1348 (.A1(n_257_76_1345), .A2(n_257_76_1290), .A3(
      n_257_76_1250), .ZN(n_257_76_1346));
   INV_X1 i_257_76_1349 (.A(n_257_76_1346), .ZN(n_257_76_1347));
   NAND3_X1 i_257_76_1350 (.A1(n_257_76_1339), .A2(n_257_76_1347), .A3(
      n_257_76_1241), .ZN(n_257_76_1348));
   INV_X1 i_257_76_1351 (.A(n_257_76_1348), .ZN(n_257_76_1349));
   NAND3_X1 i_257_76_1352 (.A1(n_257_76_1335), .A2(n_257_76_1337), .A3(
      n_257_76_1349), .ZN(n_257_76_1350));
   NOR2_X1 i_257_76_1353 (.A1(n_257_76_1333), .A2(n_257_76_1350), .ZN(
      n_257_76_1351));
   NAND3_X1 i_257_76_1354 (.A1(n_257_76_1351), .A2(n_257_76_1212), .A3(
      n_257_76_1213), .ZN(n_257_76_1352));
   INV_X1 i_257_76_1355 (.A(n_257_76_1352), .ZN(n_257_76_1353));
   NAND2_X1 i_257_76_1356 (.A1(n_257_185), .A2(n_257_76_1353), .ZN(n_257_76_1354));
   NAND3_X1 i_257_76_1357 (.A1(n_257_76_1321), .A2(n_257_76_1332), .A3(
      n_257_76_1354), .ZN(n_257_76_1355));
   NAND2_X1 i_257_76_1358 (.A1(n_257_442), .A2(n_257_1061), .ZN(n_257_76_1356));
   INV_X1 i_257_76_1359 (.A(n_257_76_1356), .ZN(n_257_76_1357));
   NAND2_X1 i_257_76_1360 (.A1(n_257_13), .A2(n_257_76_1357), .ZN(n_257_76_1358));
   NAND3_X1 i_257_76_1361 (.A1(n_257_863), .A2(n_257_76_1248), .A3(n_257_76_1249), 
      .ZN(n_257_76_1359));
   INV_X1 i_257_76_1362 (.A(n_257_76_1359), .ZN(n_257_76_1360));
   NAND2_X1 i_257_76_1363 (.A1(n_257_445), .A2(n_257_76_1226), .ZN(n_257_76_1361));
   INV_X1 i_257_76_1364 (.A(n_257_76_1361), .ZN(n_257_76_1362));
   NAND2_X1 i_257_76_1365 (.A1(n_257_76_1250), .A2(n_257_76_1362), .ZN(
      n_257_76_1363));
   INV_X1 i_257_76_1366 (.A(n_257_76_1363), .ZN(n_257_76_1364));
   NAND3_X1 i_257_76_1367 (.A1(n_257_76_1214), .A2(n_257_76_1360), .A3(
      n_257_76_1364), .ZN(n_257_76_1365));
   INV_X1 i_257_76_1368 (.A(n_257_76_1365), .ZN(n_257_76_1366));
   NAND3_X1 i_257_76_1369 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1366), .ZN(n_257_76_1367));
   INV_X1 i_257_76_1370 (.A(n_257_76_1367), .ZN(n_257_76_1368));
   NAND2_X1 i_257_76_1371 (.A1(n_257_20), .A2(n_257_76_1368), .ZN(n_257_76_1369));
   NAND2_X1 i_257_76_1372 (.A1(n_257_76_1358), .A2(n_257_76_1369), .ZN(
      n_257_76_1370));
   NOR2_X1 i_257_76_1373 (.A1(n_257_76_1355), .A2(n_257_76_1370), .ZN(
      n_257_76_1371));
   NAND2_X1 i_257_76_1374 (.A1(n_257_76_1232), .A2(n_257_76_1306), .ZN(
      n_257_76_1372));
   NAND2_X1 i_257_76_1375 (.A1(n_257_426), .A2(n_257_76_1226), .ZN(n_257_76_1373));
   NOR2_X1 i_257_76_1376 (.A1(n_257_76_1281), .A2(n_257_76_1373), .ZN(
      n_257_76_1374));
   NAND3_X1 i_257_76_1377 (.A1(n_257_76_1243), .A2(n_257_76_1374), .A3(
      n_257_76_1284), .ZN(n_257_76_1375));
   INV_X1 i_257_76_1378 (.A(n_257_76_1375), .ZN(n_257_76_1376));
   NAND4_X1 i_257_76_1379 (.A1(n_257_76_1376), .A2(n_257_76_1290), .A3(
      n_257_76_1250), .A4(n_257_76_1287), .ZN(n_257_76_1377));
   NAND3_X1 i_257_76_1380 (.A1(n_257_76_1248), .A2(n_257_76_1249), .A3(n_257_535), 
      .ZN(n_257_76_1378));
   NOR2_X1 i_257_76_1381 (.A1(n_257_76_1377), .A2(n_257_76_1378), .ZN(
      n_257_76_1379));
   NAND2_X1 i_257_76_1382 (.A1(n_257_76_1293), .A2(n_257_76_1233), .ZN(
      n_257_76_1380));
   INV_X1 i_257_76_1383 (.A(n_257_76_1380), .ZN(n_257_76_1381));
   NAND3_X1 i_257_76_1384 (.A1(n_257_76_1234), .A2(n_257_76_1241), .A3(
      n_257_76_1297), .ZN(n_257_76_1382));
   INV_X1 i_257_76_1385 (.A(n_257_76_1382), .ZN(n_257_76_1383));
   NAND3_X1 i_257_76_1386 (.A1(n_257_76_1379), .A2(n_257_76_1381), .A3(
      n_257_76_1383), .ZN(n_257_76_1384));
   INV_X1 i_257_76_1387 (.A(n_257_76_1303), .ZN(n_257_76_1385));
   INV_X1 i_257_76_1388 (.A(n_257_76_1304), .ZN(n_257_76_1386));
   NAND3_X1 i_257_76_1389 (.A1(n_257_76_1385), .A2(n_257_76_1307), .A3(
      n_257_76_1386), .ZN(n_257_76_1387));
   NOR3_X1 i_257_76_1390 (.A1(n_257_76_1372), .A2(n_257_76_1384), .A3(
      n_257_76_1387), .ZN(n_257_76_1388));
   NAND3_X1 i_257_76_1391 (.A1(n_257_76_1388), .A2(n_257_76_1212), .A3(
      n_257_76_1213), .ZN(n_257_76_1389));
   INV_X1 i_257_76_1392 (.A(n_257_76_1389), .ZN(n_257_76_1390));
   NAND2_X1 i_257_76_1393 (.A1(n_257_225), .A2(n_257_76_1390), .ZN(n_257_76_1391));
   NAND2_X1 i_257_76_1394 (.A1(n_257_735), .A2(n_257_76_1248), .ZN(n_257_76_1392));
   INV_X1 i_257_76_1395 (.A(n_257_76_1392), .ZN(n_257_76_1393));
   NAND2_X1 i_257_76_1396 (.A1(n_257_436), .A2(n_257_76_1226), .ZN(n_257_76_1394));
   INV_X1 i_257_76_1397 (.A(n_257_76_1394), .ZN(n_257_76_1395));
   NAND3_X1 i_257_76_1398 (.A1(n_257_76_1249), .A2(n_257_76_1250), .A3(
      n_257_76_1395), .ZN(n_257_76_1396));
   INV_X1 i_257_76_1399 (.A(n_257_76_1396), .ZN(n_257_76_1397));
   NAND4_X1 i_257_76_1400 (.A1(n_257_76_1393), .A2(n_257_76_1397), .A3(
      n_257_76_1240), .A4(n_257_76_1241), .ZN(n_257_76_1398));
   NAND3_X1 i_257_76_1401 (.A1(n_257_76_1214), .A2(n_257_76_1234), .A3(
      n_257_76_1235), .ZN(n_257_76_1399));
   NOR2_X1 i_257_76_1402 (.A1(n_257_76_1398), .A2(n_257_76_1399), .ZN(
      n_257_76_1400));
   NAND3_X1 i_257_76_1403 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1400), .ZN(n_257_76_1401));
   INV_X1 i_257_76_1404 (.A(n_257_76_1401), .ZN(n_257_76_1402));
   NAND2_X1 i_257_76_1405 (.A1(n_257_24), .A2(n_257_76_1402), .ZN(n_257_76_1403));
   NOR2_X1 i_257_76_1406 (.A1(n_257_76_1303), .A2(n_257_76_1236), .ZN(
      n_257_76_1404));
   NAND2_X1 i_257_76_1407 (.A1(n_257_76_1297), .A2(n_257_76_1248), .ZN(
      n_257_76_1405));
   INV_X1 i_257_76_1408 (.A(n_257_76_1405), .ZN(n_257_76_1406));
   NAND2_X1 i_257_76_1409 (.A1(n_257_76_1249), .A2(n_257_76_1290), .ZN(
      n_257_76_1407));
   INV_X1 i_257_76_1410 (.A(n_257_76_1407), .ZN(n_257_76_1408));
   INV_X1 i_257_76_1411 (.A(n_257_599), .ZN(n_257_76_1409));
   NOR2_X1 i_257_76_1412 (.A1(n_257_76_1216), .A2(n_257_76_1409), .ZN(
      n_257_76_1410));
   NAND2_X1 i_257_76_1413 (.A1(n_257_432), .A2(n_257_76_1410), .ZN(n_257_76_1411));
   INV_X1 i_257_76_1414 (.A(n_257_76_1411), .ZN(n_257_76_1412));
   NAND2_X1 i_257_76_1415 (.A1(n_257_76_1243), .A2(n_257_76_1412), .ZN(
      n_257_76_1413));
   INV_X1 i_257_76_1416 (.A(n_257_76_1413), .ZN(n_257_76_1414));
   NAND2_X1 i_257_76_1417 (.A1(n_257_76_1250), .A2(n_257_76_1414), .ZN(
      n_257_76_1415));
   INV_X1 i_257_76_1418 (.A(n_257_76_1415), .ZN(n_257_76_1416));
   NAND3_X1 i_257_76_1419 (.A1(n_257_76_1406), .A2(n_257_76_1408), .A3(
      n_257_76_1416), .ZN(n_257_76_1417));
   NOR2_X1 i_257_76_1420 (.A1(n_257_76_1417), .A2(n_257_76_1242), .ZN(
      n_257_76_1418));
   NAND3_X1 i_257_76_1421 (.A1(n_257_76_1232), .A2(n_257_76_1404), .A3(
      n_257_76_1418), .ZN(n_257_76_1419));
   INV_X1 i_257_76_1422 (.A(n_257_76_1419), .ZN(n_257_76_1420));
   NAND3_X1 i_257_76_1423 (.A1(n_257_76_1212), .A2(n_257_76_1420), .A3(
      n_257_76_1213), .ZN(n_257_76_1421));
   INV_X1 i_257_76_1424 (.A(n_257_76_1421), .ZN(n_257_76_1422));
   NAND2_X1 i_257_76_1425 (.A1(n_257_68), .A2(n_257_76_1422), .ZN(n_257_76_1423));
   NAND3_X1 i_257_76_1426 (.A1(n_257_76_1391), .A2(n_257_76_1403), .A3(
      n_257_76_1423), .ZN(n_257_76_1424));
   NAND2_X1 i_257_76_1427 (.A1(n_257_437), .A2(n_257_76_1226), .ZN(n_257_76_1425));
   INV_X1 i_257_76_1428 (.A(n_257_76_1425), .ZN(n_257_76_1426));
   NAND3_X1 i_257_76_1429 (.A1(n_257_76_1249), .A2(n_257_76_1250), .A3(
      n_257_76_1426), .ZN(n_257_76_1427));
   NAND2_X1 i_257_76_1430 (.A1(n_257_799), .A2(n_257_76_1248), .ZN(n_257_76_1428));
   NOR2_X1 i_257_76_1431 (.A1(n_257_76_1427), .A2(n_257_76_1428), .ZN(
      n_257_76_1429));
   NAND2_X1 i_257_76_1432 (.A1(n_257_76_1234), .A2(n_257_76_1235), .ZN(
      n_257_76_1430));
   INV_X1 i_257_76_1433 (.A(n_257_76_1430), .ZN(n_257_76_1431));
   NAND3_X1 i_257_76_1434 (.A1(n_257_76_1429), .A2(n_257_76_1431), .A3(
      n_257_76_1214), .ZN(n_257_76_1432));
   INV_X1 i_257_76_1435 (.A(n_257_76_1432), .ZN(n_257_76_1433));
   NAND3_X1 i_257_76_1436 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1433), .ZN(n_257_76_1434));
   INV_X1 i_257_76_1437 (.A(n_257_76_1434), .ZN(n_257_76_1435));
   NAND2_X1 i_257_76_1438 (.A1(n_257_22), .A2(n_257_76_1435), .ZN(n_257_76_1436));
   NAND2_X1 i_257_76_1439 (.A1(n_257_444), .A2(n_257_76_1226), .ZN(n_257_76_1437));
   INV_X1 i_257_76_1440 (.A(n_257_76_1437), .ZN(n_257_76_1438));
   NAND2_X1 i_257_76_1441 (.A1(n_257_997), .A2(n_257_76_1438), .ZN(n_257_76_1439));
   INV_X1 i_257_76_1442 (.A(n_257_76_1439), .ZN(n_257_76_1440));
   NAND2_X1 i_257_76_1443 (.A1(n_257_76_1212), .A2(n_257_76_1440), .ZN(
      n_257_76_1441));
   INV_X1 i_257_76_1444 (.A(n_257_76_1441), .ZN(n_257_76_1442));
   NAND2_X1 i_257_76_1445 (.A1(n_257_15), .A2(n_257_76_1442), .ZN(n_257_76_1443));
   NAND2_X1 i_257_76_1446 (.A1(n_257_76_1436), .A2(n_257_76_1443), .ZN(
      n_257_76_1444));
   NOR2_X1 i_257_76_1447 (.A1(n_257_76_1424), .A2(n_257_76_1444), .ZN(
      n_257_76_1445));
   NAND3_X1 i_257_76_1448 (.A1(n_257_76_1314), .A2(n_257_76_1371), .A3(
      n_257_76_1445), .ZN(n_257_76_1446));
   INV_X1 i_257_76_1449 (.A(n_257_76_1446), .ZN(n_257_76_1447));
   NAND3_X1 i_257_76_1450 (.A1(n_257_76_1248), .A2(n_257_76_1249), .A3(
      n_257_76_1290), .ZN(n_257_76_1448));
   INV_X1 i_257_76_1451 (.A(n_257_76_1448), .ZN(n_257_76_1449));
   NAND2_X1 i_257_76_1452 (.A1(n_257_433), .A2(n_257_76_1226), .ZN(n_257_76_1450));
   INV_X1 i_257_76_1453 (.A(n_257_76_1450), .ZN(n_257_76_1451));
   NAND2_X1 i_257_76_1454 (.A1(n_257_76_1243), .A2(n_257_76_1451), .ZN(
      n_257_76_1452));
   INV_X1 i_257_76_1455 (.A(n_257_76_1452), .ZN(n_257_76_1453));
   NAND3_X1 i_257_76_1456 (.A1(n_257_76_1250), .A2(n_257_76_1453), .A3(n_257_37), 
      .ZN(n_257_76_1454));
   INV_X1 i_257_76_1457 (.A(n_257_76_1454), .ZN(n_257_76_1455));
   NAND3_X1 i_257_76_1458 (.A1(n_257_76_1449), .A2(n_257_76_1241), .A3(
      n_257_76_1455), .ZN(n_257_76_1456));
   NOR2_X1 i_257_76_1459 (.A1(n_257_76_1456), .A2(n_257_76_1304), .ZN(
      n_257_76_1457));
   NAND4_X1 i_257_76_1460 (.A1(n_257_76_1214), .A2(n_257_76_1302), .A3(
      n_257_76_1233), .A4(n_257_76_1234), .ZN(n_257_76_1458));
   INV_X1 i_257_76_1461 (.A(n_257_76_1458), .ZN(n_257_76_1459));
   NAND3_X1 i_257_76_1462 (.A1(n_257_76_1457), .A2(n_257_76_1232), .A3(
      n_257_76_1459), .ZN(n_257_76_1460));
   INV_X1 i_257_76_1463 (.A(n_257_76_1460), .ZN(n_257_76_1461));
   NAND3_X1 i_257_76_1464 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1461), .ZN(n_257_76_1462));
   INV_X1 i_257_76_1465 (.A(n_257_76_1462), .ZN(n_257_76_1463));
   NAND2_X1 i_257_76_1466 (.A1(n_257_67), .A2(n_257_76_1463), .ZN(n_257_76_1464));
   NAND3_X1 i_257_76_1467 (.A1(n_257_76_1240), .A2(n_257_76_1241), .A3(n_257_449), 
      .ZN(n_257_76_1465));
   NAND2_X1 i_257_76_1468 (.A1(n_257_76_18056), .A2(n_257_1075), .ZN(
      n_257_76_1466));
   INV_X1 i_257_76_1469 (.A(n_257_76_1466), .ZN(n_257_76_1467));
   NAND4_X1 i_257_76_1470 (.A1(n_257_76_1467), .A2(n_257_76_1248), .A3(
      n_257_76_1249), .A4(n_257_76_1250), .ZN(n_257_76_1468));
   NOR2_X1 i_257_76_1471 (.A1(n_257_76_1465), .A2(n_257_76_1468), .ZN(
      n_257_76_1469));
   NAND3_X1 i_257_76_1472 (.A1(n_257_76_1232), .A2(n_257_76_1469), .A3(
      n_257_76_1238), .ZN(n_257_76_1470));
   INV_X1 i_257_76_1473 (.A(n_257_76_1470), .ZN(n_257_76_1471));
   NAND3_X1 i_257_76_1474 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1471), .ZN(n_257_76_1472));
   INV_X1 i_257_76_1475 (.A(n_257_76_1472), .ZN(n_257_76_1473));
   NAND2_X1 i_257_76_1476 (.A1(n_257_27), .A2(n_257_76_1473), .ZN(n_257_76_1474));
   NAND2_X1 i_257_76_1477 (.A1(n_257_76_1307), .A2(n_257_154), .ZN(n_257_76_1475));
   INV_X1 i_257_76_1478 (.A(n_257_76_1475), .ZN(n_257_76_1476));
   NAND2_X1 i_257_76_1479 (.A1(n_257_429), .A2(n_257_76_1226), .ZN(n_257_76_1477));
   INV_X1 i_257_76_1480 (.A(n_257_76_1477), .ZN(n_257_76_1478));
   NAND3_X1 i_257_76_1481 (.A1(n_257_76_1243), .A2(n_257_76_1284), .A3(
      n_257_76_1478), .ZN(n_257_76_1479));
   INV_X1 i_257_76_1482 (.A(n_257_76_1479), .ZN(n_257_76_1480));
   NAND3_X1 i_257_76_1483 (.A1(n_257_76_1480), .A2(n_257_76_1290), .A3(
      n_257_76_1250), .ZN(n_257_76_1481));
   INV_X1 i_257_76_1484 (.A(n_257_76_1481), .ZN(n_257_76_1482));
   NAND3_X1 i_257_76_1485 (.A1(n_257_76_1339), .A2(n_257_76_1482), .A3(
      n_257_76_1241), .ZN(n_257_76_1483));
   NOR2_X1 i_257_76_1486 (.A1(n_257_76_1483), .A2(n_257_76_1304), .ZN(
      n_257_76_1484));
   NOR2_X1 i_257_76_1487 (.A1(n_257_76_1303), .A2(n_257_76_1294), .ZN(
      n_257_76_1485));
   NAND4_X1 i_257_76_1488 (.A1(n_257_76_1476), .A2(n_257_76_1484), .A3(
      n_257_76_1485), .A4(n_257_76_1232), .ZN(n_257_76_1486));
   INV_X1 i_257_76_1489 (.A(n_257_76_1486), .ZN(n_257_76_1487));
   NAND3_X1 i_257_76_1490 (.A1(n_257_76_1487), .A2(n_257_76_1212), .A3(
      n_257_76_1213), .ZN(n_257_76_1488));
   INV_X1 i_257_76_1491 (.A(n_257_76_1488), .ZN(n_257_76_1489));
   NAND2_X1 i_257_76_1492 (.A1(n_257_184), .A2(n_257_76_1489), .ZN(n_257_76_1490));
   NAND3_X1 i_257_76_1493 (.A1(n_257_76_1464), .A2(n_257_76_1474), .A3(
      n_257_76_1490), .ZN(n_257_76_1491));
   INV_X1 i_257_76_1494 (.A(n_257_76_1491), .ZN(n_257_76_1492));
   NAND2_X1 i_257_76_1495 (.A1(n_257_1067), .A2(n_257_76_1226), .ZN(
      n_257_76_1493));
   INV_X1 i_257_76_1496 (.A(n_257_76_1493), .ZN(n_257_76_1494));
   NAND2_X1 i_257_76_1497 (.A1(n_257_438), .A2(n_257_76_1494), .ZN(n_257_76_1495));
   INV_X1 i_257_76_1498 (.A(n_257_76_1495), .ZN(n_257_76_1496));
   NAND3_X1 i_257_76_1499 (.A1(n_257_76_1496), .A2(n_257_76_1248), .A3(
      n_257_76_1250), .ZN(n_257_76_1497));
   INV_X1 i_257_76_1500 (.A(n_257_76_1497), .ZN(n_257_76_1498));
   NAND2_X1 i_257_76_1501 (.A1(n_257_76_1214), .A2(n_257_76_1498), .ZN(
      n_257_76_1499));
   INV_X1 i_257_76_1502 (.A(n_257_76_1499), .ZN(n_257_76_1500));
   NAND3_X1 i_257_76_1503 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1500), .ZN(n_257_76_1501));
   INV_X1 i_257_76_1504 (.A(n_257_76_1501), .ZN(n_257_76_1502));
   NAND2_X1 i_257_76_1505 (.A1(n_257_19), .A2(n_257_76_1502), .ZN(n_257_76_1503));
   NAND4_X1 i_257_76_1506 (.A1(n_257_76_1248), .A2(n_257_76_1249), .A3(
      n_257_76_1290), .A4(n_257_76_1250), .ZN(n_257_76_1504));
   NAND3_X1 i_257_76_1507 (.A1(n_257_442), .A2(n_257_76_1215), .A3(n_257_893), 
      .ZN(n_257_76_1505));
   INV_X1 i_257_76_1508 (.A(n_257_76_1505), .ZN(n_257_76_1506));
   NAND3_X1 i_257_76_1509 (.A1(n_257_420), .A2(n_257_76_1280), .A3(n_257_76_1506), 
      .ZN(n_257_76_1507));
   INV_X1 i_257_76_1510 (.A(n_257_76_1507), .ZN(n_257_76_1508));
   NAND2_X1 i_257_76_1511 (.A1(n_257_76_1288), .A2(n_257_76_1508), .ZN(
      n_257_76_1509));
   INV_X1 i_257_76_1512 (.A(n_257_76_1509), .ZN(n_257_76_1510));
   NAND2_X1 i_257_76_1513 (.A1(n_257_76_1243), .A2(n_257_76_1284), .ZN(
      n_257_76_1511));
   INV_X1 i_257_76_1514 (.A(n_257_76_1511), .ZN(n_257_76_1512));
   NAND2_X1 i_257_76_1515 (.A1(n_257_312), .A2(n_257_422), .ZN(n_257_76_1513));
   NAND4_X1 i_257_76_1516 (.A1(n_257_76_1510), .A2(n_257_76_1512), .A3(
      n_257_76_1513), .A4(n_257_76_1287), .ZN(n_257_76_1514));
   NOR2_X1 i_257_76_1517 (.A1(n_257_76_1504), .A2(n_257_76_1514), .ZN(
      n_257_76_1515));
   NAND2_X1 i_257_76_1518 (.A1(n_257_274), .A2(n_257_423), .ZN(n_257_76_1516));
   NAND4_X1 i_257_76_1519 (.A1(n_257_76_1241), .A2(n_257_76_1516), .A3(
      n_257_76_1296), .A4(n_257_76_1297), .ZN(n_257_76_1517));
   INV_X1 i_257_76_1520 (.A(n_257_76_1517), .ZN(n_257_76_1518));
   NAND3_X1 i_257_76_1521 (.A1(n_257_76_1515), .A2(n_257_76_1518), .A3(
      n_257_76_1386), .ZN(n_257_76_1519));
   NAND3_X1 i_257_76_1522 (.A1(n_257_76_1385), .A2(n_257_76_1307), .A3(
      n_257_76_1295), .ZN(n_257_76_1520));
   NOR2_X1 i_257_76_1523 (.A1(n_257_76_1519), .A2(n_257_76_1520), .ZN(
      n_257_76_1521));
   NAND2_X1 i_257_76_1524 (.A1(n_257_351), .A2(n_257_421), .ZN(n_257_76_1522));
   NAND4_X1 i_257_76_1525 (.A1(n_257_76_1232), .A2(n_257_76_1278), .A3(
      n_257_76_1306), .A4(n_257_76_1522), .ZN(n_257_76_1523));
   INV_X1 i_257_76_1526 (.A(n_257_76_1523), .ZN(n_257_76_1524));
   NAND4_X1 i_257_76_1527 (.A1(n_257_76_1212), .A2(n_257_76_1521), .A3(
      n_257_76_1524), .A4(n_257_76_1213), .ZN(n_257_76_1525));
   INV_X1 i_257_76_1528 (.A(n_257_76_1525), .ZN(n_257_76_1526));
   NAND2_X1 i_257_76_1529 (.A1(n_257_382), .A2(n_257_76_1526), .ZN(n_257_76_1527));
   NAND4_X1 i_257_76_1530 (.A1(n_257_76_1233), .A2(n_257_76_1234), .A3(
      n_257_76_1235), .A4(n_257_76_1239), .ZN(n_257_76_1528));
   NOR2_X1 i_257_76_1531 (.A1(n_257_76_1528), .A2(n_257_76_1303), .ZN(
      n_257_76_1529));
   INV_X1 i_257_76_1532 (.A(n_257_76_1250), .ZN(n_257_76_1530));
   NAND2_X1 i_257_76_1533 (.A1(n_257_430), .A2(n_257_76_1226), .ZN(n_257_76_1531));
   INV_X1 i_257_76_1534 (.A(n_257_76_1531), .ZN(n_257_76_1532));
   NAND3_X1 i_257_76_1535 (.A1(n_257_76_1243), .A2(n_257_76_1284), .A3(
      n_257_76_1532), .ZN(n_257_76_1533));
   NOR2_X1 i_257_76_1536 (.A1(n_257_76_1530), .A2(n_257_76_1533), .ZN(
      n_257_76_1534));
   NAND3_X1 i_257_76_1537 (.A1(n_257_76_1406), .A2(n_257_76_1534), .A3(
      n_257_76_1408), .ZN(n_257_76_1535));
   NAND3_X1 i_257_76_1538 (.A1(n_257_76_1240), .A2(n_257_76_1241), .A3(n_257_115), 
      .ZN(n_257_76_1536));
   NOR2_X1 i_257_76_1539 (.A1(n_257_76_1535), .A2(n_257_76_1536), .ZN(
      n_257_76_1537));
   NAND4_X1 i_257_76_1540 (.A1(n_257_76_1232), .A2(n_257_76_1529), .A3(
      n_257_76_1307), .A4(n_257_76_1537), .ZN(n_257_76_1538));
   INV_X1 i_257_76_1541 (.A(n_257_76_1538), .ZN(n_257_76_1539));
   NAND3_X1 i_257_76_1542 (.A1(n_257_76_1539), .A2(n_257_76_1212), .A3(
      n_257_76_1213), .ZN(n_257_76_1540));
   INV_X1 i_257_76_1543 (.A(n_257_76_1540), .ZN(n_257_76_1541));
   NAND2_X1 i_257_76_1544 (.A1(n_257_145), .A2(n_257_76_1541), .ZN(n_257_76_1542));
   NAND3_X1 i_257_76_1545 (.A1(n_257_76_1503), .A2(n_257_76_1527), .A3(
      n_257_76_1542), .ZN(n_257_76_1543));
   INV_X1 i_257_76_1546 (.A(n_257_76_1543), .ZN(n_257_76_1544));
   INV_X1 i_257_76_1547 (.A(n_257_767), .ZN(n_257_76_1545));
   NOR2_X1 i_257_76_1548 (.A1(n_257_76_1216), .A2(n_257_76_1545), .ZN(
      n_257_76_1546));
   NAND3_X1 i_257_76_1549 (.A1(n_257_76_1249), .A2(n_257_76_1250), .A3(
      n_257_76_1546), .ZN(n_257_76_1547));
   INV_X1 i_257_76_1550 (.A(n_257_76_1547), .ZN(n_257_76_1548));
   NAND2_X1 i_257_76_1551 (.A1(n_257_447), .A2(n_257_76_1248), .ZN(n_257_76_1549));
   INV_X1 i_257_76_1552 (.A(n_257_76_1549), .ZN(n_257_76_1550));
   NAND4_X1 i_257_76_1553 (.A1(n_257_76_1548), .A2(n_257_76_1550), .A3(
      n_257_76_1235), .A4(n_257_76_1241), .ZN(n_257_76_1551));
   NAND2_X1 i_257_76_1554 (.A1(n_257_76_1214), .A2(n_257_76_1234), .ZN(
      n_257_76_1552));
   NOR2_X1 i_257_76_1555 (.A1(n_257_76_1551), .A2(n_257_76_1552), .ZN(
      n_257_76_1553));
   NAND3_X1 i_257_76_1556 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1553), .ZN(n_257_76_1554));
   INV_X1 i_257_76_1557 (.A(n_257_76_1554), .ZN(n_257_76_1555));
   NAND2_X1 i_257_76_1558 (.A1(n_257_77), .A2(n_257_76_1214), .ZN(n_257_76_1556));
   NAND3_X1 i_257_76_1559 (.A1(n_257_76_1302), .A2(n_257_76_1233), .A3(
      n_257_76_1234), .ZN(n_257_76_1557));
   NOR2_X1 i_257_76_1560 (.A1(n_257_76_1556), .A2(n_257_76_1557), .ZN(
      n_257_76_1558));
   NAND2_X1 i_257_76_1561 (.A1(n_257_431), .A2(n_257_76_1226), .ZN(n_257_76_1559));
   INV_X1 i_257_76_1562 (.A(n_257_76_1559), .ZN(n_257_76_1560));
   NAND3_X1 i_257_76_1563 (.A1(n_257_76_1243), .A2(n_257_76_1284), .A3(
      n_257_76_1560), .ZN(n_257_76_1561));
   INV_X1 i_257_76_1564 (.A(n_257_76_1561), .ZN(n_257_76_1562));
   NAND3_X1 i_257_76_1565 (.A1(n_257_76_1562), .A2(n_257_76_1290), .A3(
      n_257_76_1250), .ZN(n_257_76_1563));
   INV_X1 i_257_76_1566 (.A(n_257_76_1563), .ZN(n_257_76_1564));
   NAND3_X1 i_257_76_1567 (.A1(n_257_76_1339), .A2(n_257_76_1564), .A3(
      n_257_76_1241), .ZN(n_257_76_1565));
   NOR2_X1 i_257_76_1568 (.A1(n_257_76_1565), .A2(n_257_76_1304), .ZN(
      n_257_76_1566));
   NAND3_X1 i_257_76_1569 (.A1(n_257_76_1232), .A2(n_257_76_1558), .A3(
      n_257_76_1566), .ZN(n_257_76_1567));
   INV_X1 i_257_76_1570 (.A(n_257_76_1567), .ZN(n_257_76_1568));
   NAND3_X1 i_257_76_1571 (.A1(n_257_76_1212), .A2(n_257_76_1568), .A3(
      n_257_76_1213), .ZN(n_257_76_1569));
   INV_X1 i_257_76_1572 (.A(n_257_76_1569), .ZN(n_257_76_1570));
   AOI22_X1 i_257_76_1573 (.A1(n_257_23), .A2(n_257_76_1555), .B1(n_257_107), 
      .B2(n_257_76_1570), .ZN(n_257_76_1571));
   NAND3_X1 i_257_76_1574 (.A1(n_257_76_1492), .A2(n_257_76_1544), .A3(
      n_257_76_1571), .ZN(n_257_76_1572));
   NAND2_X1 i_257_76_1575 (.A1(n_257_76_1214), .A2(n_257_76_1233), .ZN(
      n_257_76_1573));
   INV_X1 i_257_76_1576 (.A(n_257_76_1573), .ZN(n_257_76_1574));
   NAND3_X1 i_257_76_1577 (.A1(n_257_448), .A2(n_257_76_1250), .A3(
      n_257_76_18056), .ZN(n_257_76_1575));
   INV_X1 i_257_76_1578 (.A(n_257_76_1575), .ZN(n_257_76_1576));
   NAND3_X1 i_257_76_1579 (.A1(n_257_76_1576), .A2(n_257_76_1323), .A3(
      n_257_76_1241), .ZN(n_257_76_1577));
   INV_X1 i_257_76_1580 (.A(n_257_76_1577), .ZN(n_257_76_1578));
   NAND3_X1 i_257_76_1581 (.A1(n_257_76_1234), .A2(n_257_76_1235), .A3(
      n_257_76_1240), .ZN(n_257_76_1579));
   INV_X1 i_257_76_1582 (.A(n_257_76_1579), .ZN(n_257_76_1580));
   NAND4_X1 i_257_76_1583 (.A1(n_257_76_1574), .A2(n_257_76_1578), .A3(n_257_671), 
      .A4(n_257_76_1580), .ZN(n_257_76_1581));
   INV_X1 i_257_76_1584 (.A(n_257_76_1581), .ZN(n_257_76_1582));
   NAND3_X1 i_257_76_1585 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1582), .ZN(n_257_76_1583));
   INV_X1 i_257_76_1586 (.A(n_257_76_1583), .ZN(n_257_76_1584));
   NAND2_X1 i_257_76_1587 (.A1(n_257_26), .A2(n_257_76_1584), .ZN(n_257_76_1585));
   NAND2_X1 i_257_76_1588 (.A1(n_257_76_1212), .A2(n_257_76_1213), .ZN(
      n_257_76_1586));
   NAND2_X1 i_257_76_1589 (.A1(n_257_425), .A2(n_257_76_1226), .ZN(n_257_76_1587));
   NOR2_X1 i_257_76_1590 (.A1(n_257_76_1281), .A2(n_257_76_1587), .ZN(
      n_257_76_1588));
   NAND3_X1 i_257_76_1591 (.A1(n_257_76_1243), .A2(n_257_76_1588), .A3(
      n_257_76_1284), .ZN(n_257_76_1589));
   INV_X1 i_257_76_1592 (.A(n_257_76_1589), .ZN(n_257_76_1590));
   NAND4_X1 i_257_76_1593 (.A1(n_257_76_1590), .A2(n_257_76_1290), .A3(
      n_257_76_1250), .A4(n_257_76_1287), .ZN(n_257_76_1591));
   INV_X1 i_257_76_1594 (.A(n_257_76_1591), .ZN(n_257_76_1592));
   NAND2_X1 i_257_76_1595 (.A1(n_257_76_1592), .A2(n_257_76_1339), .ZN(
      n_257_76_1593));
   NAND3_X1 i_257_76_1596 (.A1(n_257_76_1234), .A2(n_257_76_1235), .A3(
      n_257_76_1239), .ZN(n_257_76_1594));
   NAND3_X1 i_257_76_1597 (.A1(n_257_76_1240), .A2(n_257_76_1241), .A3(
      n_257_76_1296), .ZN(n_257_76_1595));
   NOR3_X1 i_257_76_1598 (.A1(n_257_76_1593), .A2(n_257_76_1594), .A3(
      n_257_76_1595), .ZN(n_257_76_1596));
   INV_X1 i_257_76_1599 (.A(n_257_76_1372), .ZN(n_257_76_1597));
   NAND3_X1 i_257_76_1600 (.A1(n_257_76_1302), .A2(n_257_76_1293), .A3(
      n_257_76_1233), .ZN(n_257_76_1598));
   INV_X1 i_257_76_1601 (.A(n_257_76_1598), .ZN(n_257_76_1599));
   NAND4_X1 i_257_76_1602 (.A1(n_257_76_1599), .A2(n_257_76_1307), .A3(n_257_234), 
      .A4(n_257_76_1214), .ZN(n_257_76_1600));
   INV_X1 i_257_76_1603 (.A(n_257_76_1600), .ZN(n_257_76_1601));
   NAND3_X1 i_257_76_1604 (.A1(n_257_76_1596), .A2(n_257_76_1597), .A3(
      n_257_76_1601), .ZN(n_257_76_1602));
   NOR2_X1 i_257_76_1605 (.A1(n_257_76_1586), .A2(n_257_76_1602), .ZN(
      n_257_76_1603));
   NAND2_X1 i_257_76_1606 (.A1(n_257_264), .A2(n_257_76_1603), .ZN(n_257_76_1604));
   NAND2_X1 i_257_76_1607 (.A1(n_257_421), .A2(n_257_76_1226), .ZN(n_257_76_1605));
   NOR2_X1 i_257_76_1608 (.A1(n_257_76_1281), .A2(n_257_76_1605), .ZN(
      n_257_76_1606));
   NAND3_X1 i_257_76_1609 (.A1(n_257_76_1606), .A2(n_257_76_1243), .A3(
      n_257_76_1284), .ZN(n_257_76_1607));
   INV_X1 i_257_76_1610 (.A(n_257_76_1607), .ZN(n_257_76_1608));
   NAND4_X1 i_257_76_1611 (.A1(n_257_76_1608), .A2(n_257_76_1513), .A3(
      n_257_76_1287), .A4(n_257_76_1288), .ZN(n_257_76_1609));
   NOR2_X1 i_257_76_1612 (.A1(n_257_76_1504), .A2(n_257_76_1609), .ZN(
      n_257_76_1610));
   NAND3_X1 i_257_76_1613 (.A1(n_257_76_1610), .A2(n_257_76_1518), .A3(
      n_257_76_1386), .ZN(n_257_76_1611));
   NAND2_X1 i_257_76_1614 (.A1(n_257_76_1302), .A2(n_257_76_1293), .ZN(
      n_257_76_1612));
   INV_X1 i_257_76_1615 (.A(n_257_76_1612), .ZN(n_257_76_1613));
   INV_X1 i_257_76_1616 (.A(n_257_76_1334), .ZN(n_257_76_1614));
   NAND3_X1 i_257_76_1617 (.A1(n_257_76_1613), .A2(n_257_76_1214), .A3(
      n_257_76_1614), .ZN(n_257_76_1615));
   NOR2_X1 i_257_76_1618 (.A1(n_257_76_1611), .A2(n_257_76_1615), .ZN(
      n_257_76_1616));
   INV_X1 i_257_76_1619 (.A(n_257_76_1279), .ZN(n_257_76_1617));
   INV_X1 i_257_76_1620 (.A(n_257_76_1306), .ZN(n_257_76_1618));
   NAND2_X1 i_257_76_1621 (.A1(n_257_76_1307), .A2(n_257_351), .ZN(n_257_76_1619));
   NOR2_X1 i_257_76_1622 (.A1(n_257_76_1618), .A2(n_257_76_1619), .ZN(
      n_257_76_1620));
   NAND3_X1 i_257_76_1623 (.A1(n_257_76_1616), .A2(n_257_76_1617), .A3(
      n_257_76_1620), .ZN(n_257_76_1621));
   NOR2_X1 i_257_76_1624 (.A1(n_257_76_1621), .A2(n_257_76_1586), .ZN(
      n_257_76_1622));
   NAND2_X1 i_257_76_1625 (.A1(n_257_381), .A2(n_257_76_1622), .ZN(n_257_76_1623));
   NAND3_X1 i_257_76_1626 (.A1(n_257_76_1585), .A2(n_257_76_1604), .A3(
      n_257_76_1623), .ZN(n_257_76_1624));
   INV_X1 i_257_76_1627 (.A(n_257_76_1624), .ZN(n_257_76_1625));
   INV_X1 i_257_76_1628 (.A(n_257_567), .ZN(n_257_76_1626));
   NAND3_X1 i_257_76_1629 (.A1(n_257_76_1626), .A2(n_257_442), .A3(n_257_76_1215), 
      .ZN(n_257_76_1627));
   OAI21_X1 i_257_76_1630 (.A(n_257_76_1627), .B1(n_257_428), .B2(n_257_76_1216), 
      .ZN(n_257_76_1628));
   NAND3_X1 i_257_76_1631 (.A1(n_257_427), .A2(n_257_76_1284), .A3(n_257_76_1628), 
      .ZN(n_257_76_1629));
   INV_X1 i_257_76_1632 (.A(n_257_76_1629), .ZN(n_257_76_1630));
   NAND2_X1 i_257_76_1633 (.A1(n_257_76_1243), .A2(n_257_194), .ZN(n_257_76_1631));
   INV_X1 i_257_76_1634 (.A(n_257_76_1631), .ZN(n_257_76_1632));
   NAND4_X1 i_257_76_1635 (.A1(n_257_76_1297), .A2(n_257_76_1630), .A3(
      n_257_76_1290), .A4(n_257_76_1632), .ZN(n_257_76_1633));
   INV_X1 i_257_76_1636 (.A(n_257_76_1633), .ZN(n_257_76_1634));
   NAND3_X1 i_257_76_1637 (.A1(n_257_76_1634), .A2(n_257_76_1214), .A3(
      n_257_76_1302), .ZN(n_257_76_1635));
   INV_X1 i_257_76_1638 (.A(n_257_76_1635), .ZN(n_257_76_1636));
   NAND3_X1 i_257_76_1639 (.A1(n_257_76_1248), .A2(n_257_76_1249), .A3(
      n_257_76_1250), .ZN(n_257_76_1637));
   INV_X1 i_257_76_1640 (.A(n_257_76_1637), .ZN(n_257_76_1638));
   NAND4_X1 i_257_76_1641 (.A1(n_257_76_1638), .A2(n_257_76_1239), .A3(
      n_257_76_1240), .A4(n_257_76_1241), .ZN(n_257_76_1639));
   INV_X1 i_257_76_1642 (.A(n_257_76_1639), .ZN(n_257_76_1640));
   NAND4_X1 i_257_76_1643 (.A1(n_257_76_1293), .A2(n_257_76_1233), .A3(
      n_257_76_1234), .A4(n_257_76_1235), .ZN(n_257_76_1641));
   INV_X1 i_257_76_1644 (.A(n_257_76_1641), .ZN(n_257_76_1642));
   NAND3_X1 i_257_76_1645 (.A1(n_257_76_1636), .A2(n_257_76_1640), .A3(
      n_257_76_1642), .ZN(n_257_76_1643));
   NOR2_X1 i_257_76_1646 (.A1(n_257_76_1333), .A2(n_257_76_1643), .ZN(
      n_257_76_1644));
   NAND3_X1 i_257_76_1647 (.A1(n_257_76_1644), .A2(n_257_76_1212), .A3(
      n_257_76_1213), .ZN(n_257_76_1645));
   INV_X1 i_257_76_1648 (.A(n_257_76_1645), .ZN(n_257_76_1646));
   NAND2_X1 i_257_76_1649 (.A1(n_257_224), .A2(n_257_76_1646), .ZN(n_257_76_1647));
   NAND2_X1 i_257_76_1650 (.A1(n_257_76_1290), .A2(n_257_76_1250), .ZN(
      n_257_76_1648));
   INV_X1 i_257_76_1651 (.A(n_257_76_1648), .ZN(n_257_76_1649));
   NAND2_X1 i_257_76_1652 (.A1(n_257_76_18056), .A2(n_257_454), .ZN(
      n_257_76_1650));
   INV_X1 i_257_76_1653 (.A(n_257_76_1650), .ZN(n_257_76_1651));
   NAND4_X1 i_257_76_1654 (.A1(n_257_76_1323), .A2(n_257_76_1649), .A3(n_257_451), 
      .A4(n_257_76_1651), .ZN(n_257_76_1652));
   NOR2_X1 i_257_76_1655 (.A1(n_257_76_1652), .A2(n_257_76_1242), .ZN(
      n_257_76_1653));
   NAND3_X1 i_257_76_1656 (.A1(n_257_76_1653), .A2(n_257_76_1232), .A3(
      n_257_76_1238), .ZN(n_257_76_1654));
   INV_X1 i_257_76_1657 (.A(n_257_76_1654), .ZN(n_257_76_1655));
   NAND3_X1 i_257_76_1658 (.A1(n_257_76_1212), .A2(n_257_76_1213), .A3(
      n_257_76_1655), .ZN(n_257_76_1656));
   INV_X1 i_257_76_1659 (.A(n_257_76_1656), .ZN(n_257_76_1657));
   NAND2_X1 i_257_76_1660 (.A1(n_257_434), .A2(n_257_76_1657), .ZN(n_257_76_1658));
   NOR2_X1 i_257_76_1661 (.A1(n_257_76_1294), .A2(n_257_76_1304), .ZN(
      n_257_76_1659));
   NAND2_X1 i_257_76_1662 (.A1(n_257_76_1243), .A2(n_257_503), .ZN(n_257_76_1660));
   INV_X1 i_257_76_1663 (.A(n_257_76_1660), .ZN(n_257_76_1661));
   NAND3_X1 i_257_76_1664 (.A1(n_257_76_1284), .A2(n_257_76_1628), .A3(n_257_424), 
      .ZN(n_257_76_1662));
   INV_X1 i_257_76_1665 (.A(n_257_76_1662), .ZN(n_257_76_1663));
   NAND4_X1 i_257_76_1666 (.A1(n_257_76_1297), .A2(n_257_76_1290), .A3(
      n_257_76_1661), .A4(n_257_76_1663), .ZN(n_257_76_1664));
   INV_X1 i_257_76_1667 (.A(n_257_76_1664), .ZN(n_257_76_1665));
   NAND3_X1 i_257_76_1668 (.A1(n_257_76_1665), .A2(n_257_76_1214), .A3(
      n_257_76_1302), .ZN(n_257_76_1666));
   INV_X1 i_257_76_1669 (.A(n_257_76_1666), .ZN(n_257_76_1667));
   NAND2_X1 i_257_76_1670 (.A1(n_257_76_1241), .A2(n_257_76_1296), .ZN(
      n_257_76_1668));
   NAND4_X1 i_257_76_1671 (.A1(n_257_76_1248), .A2(n_257_76_1249), .A3(
      n_257_76_1250), .A4(n_257_76_1287), .ZN(n_257_76_1669));
   NOR2_X1 i_257_76_1672 (.A1(n_257_76_1668), .A2(n_257_76_1669), .ZN(
      n_257_76_1670));
   NAND4_X1 i_257_76_1673 (.A1(n_257_76_1659), .A2(n_257_76_1667), .A3(
      n_257_76_1307), .A4(n_257_76_1670), .ZN(n_257_76_1671));
   NAND3_X1 i_257_76_1674 (.A1(n_257_76_1232), .A2(n_257_76_1278), .A3(
      n_257_76_1306), .ZN(n_257_76_1672));
   NOR2_X1 i_257_76_1675 (.A1(n_257_76_1671), .A2(n_257_76_1672), .ZN(
      n_257_76_1673));
   NAND3_X1 i_257_76_1676 (.A1(n_257_76_1673), .A2(n_257_76_1212), .A3(
      n_257_76_1213), .ZN(n_257_76_1674));
   INV_X1 i_257_76_1677 (.A(n_257_76_1674), .ZN(n_257_76_1675));
   NAND2_X1 i_257_76_1678 (.A1(n_257_265), .A2(n_257_76_1675), .ZN(n_257_76_1676));
   NAND3_X1 i_257_76_1679 (.A1(n_257_76_1647), .A2(n_257_76_1658), .A3(
      n_257_76_1676), .ZN(n_257_76_1677));
   INV_X1 i_257_76_1680 (.A(n_257_76_1677), .ZN(n_257_76_1678));
   NOR2_X1 i_257_76_1681 (.A1(n_257_76_1598), .A2(n_257_76_1594), .ZN(
      n_257_76_1679));
   NAND2_X1 i_257_76_1682 (.A1(n_257_76_1250), .A2(n_257_76_1287), .ZN(
      n_257_76_1680));
   INV_X1 i_257_76_1683 (.A(n_257_76_1680), .ZN(n_257_76_1681));
   NAND3_X1 i_257_76_1684 (.A1(n_257_76_1323), .A2(n_257_76_1296), .A3(
      n_257_76_1681), .ZN(n_257_76_1682));
   NAND3_X1 i_257_76_1685 (.A1(n_257_76_1240), .A2(n_257_76_1241), .A3(
      n_257_76_1516), .ZN(n_257_76_1683));
   NOR2_X1 i_257_76_1686 (.A1(n_257_76_1682), .A2(n_257_76_1683), .ZN(
      n_257_76_1684));
   NAND3_X1 i_257_76_1687 (.A1(n_257_76_1288), .A2(n_257_312), .A3(n_257_76_1243), 
      .ZN(n_257_76_1685));
   INV_X1 i_257_76_1688 (.A(n_257_76_1685), .ZN(n_257_76_1686));
   NAND3_X1 i_257_76_1689 (.A1(n_257_76_1284), .A2(n_257_76_1628), .A3(n_257_422), 
      .ZN(n_257_76_1687));
   INV_X1 i_257_76_1690 (.A(n_257_76_1687), .ZN(n_257_76_1688));
   NAND4_X1 i_257_76_1691 (.A1(n_257_76_1686), .A2(n_257_76_1297), .A3(
      n_257_76_1290), .A4(n_257_76_1688), .ZN(n_257_76_1689));
   NOR2_X1 i_257_76_1692 (.A1(n_257_76_1237), .A2(n_257_76_1689), .ZN(
      n_257_76_1690));
   NAND4_X1 i_257_76_1693 (.A1(n_257_76_1679), .A2(n_257_76_1684), .A3(
      n_257_76_1307), .A4(n_257_76_1690), .ZN(n_257_76_1691));
   NOR2_X1 i_257_76_1694 (.A1(n_257_76_1691), .A2(n_257_76_1672), .ZN(
      n_257_76_1692));
   NAND3_X1 i_257_76_1695 (.A1(n_257_76_1692), .A2(n_257_76_1212), .A3(
      n_257_76_1213), .ZN(n_257_76_1693));
   INV_X1 i_257_76_1696 (.A(n_257_76_1693), .ZN(n_257_76_1694));
   NAND2_X1 i_257_76_1697 (.A1(n_257_342), .A2(n_257_76_1694), .ZN(n_257_76_1695));
   NAND2_X1 i_257_76_1698 (.A1(n_257_76_1516), .A2(n_257_76_1296), .ZN(
      n_257_76_1696));
   INV_X1 i_257_76_1699 (.A(n_257_76_1696), .ZN(n_257_76_1697));
   INV_X1 i_257_76_1700 (.A(n_257_76_1297), .ZN(n_257_76_1698));
   NOR2_X1 i_257_76_1701 (.A1(n_257_76_1322), .A2(n_257_76_1698), .ZN(
      n_257_76_1699));
   NAND2_X1 i_257_76_1702 (.A1(n_257_76_1697), .A2(n_257_76_1699), .ZN(
      n_257_76_1700));
   NAND2_X1 i_257_76_1703 (.A1(n_257_76_1250), .A2(n_257_76_1513), .ZN(
      n_257_76_1701));
   INV_X1 i_257_76_1704 (.A(n_257_76_1290), .ZN(n_257_76_1702));
   NOR2_X1 i_257_76_1705 (.A1(n_257_76_1701), .A2(n_257_76_1702), .ZN(
      n_257_76_1703));
   NAND2_X1 i_257_76_1706 (.A1(n_257_420), .A2(n_257_893), .ZN(n_257_76_1704));
   NAND2_X1 i_257_76_1707 (.A1(n_257_76_1243), .A2(n_257_76_1704), .ZN(
      n_257_76_1705));
   INV_X1 i_257_76_1708 (.A(n_257_76_1705), .ZN(n_257_76_1706));
   NAND3_X1 i_257_76_1709 (.A1(n_257_484), .A2(n_257_76_1226), .A3(n_257_390), 
      .ZN(n_257_76_1707));
   INV_X1 i_257_76_1710 (.A(n_257_76_1707), .ZN(n_257_76_1708));
   NAND2_X1 i_257_76_1711 (.A1(n_257_76_1280), .A2(n_257_76_1708), .ZN(
      n_257_76_1709));
   INV_X1 i_257_76_1712 (.A(n_257_76_1709), .ZN(n_257_76_1710));
   NAND2_X1 i_257_76_1713 (.A1(n_257_76_1710), .A2(n_257_76_1284), .ZN(
      n_257_76_1711));
   INV_X1 i_257_76_1714 (.A(n_257_76_1711), .ZN(n_257_76_1712));
   NAND2_X1 i_257_76_1715 (.A1(n_257_76_1706), .A2(n_257_76_1712), .ZN(
      n_257_76_1713));
   NAND2_X1 i_257_76_1716 (.A1(n_257_76_1287), .A2(n_257_76_1288), .ZN(
      n_257_76_1714));
   NOR2_X1 i_257_76_1717 (.A1(n_257_76_1713), .A2(n_257_76_1714), .ZN(
      n_257_76_1715));
   NAND2_X1 i_257_76_1718 (.A1(n_257_76_1703), .A2(n_257_76_1715), .ZN(
      n_257_76_1716));
   NOR2_X1 i_257_76_1719 (.A1(n_257_76_1700), .A2(n_257_76_1716), .ZN(
      n_257_76_1717));
   NAND2_X1 i_257_76_1720 (.A1(n_257_76_1235), .A2(n_257_76_1239), .ZN(
      n_257_76_1718));
   NAND2_X1 i_257_76_1721 (.A1(n_257_76_1240), .A2(n_257_76_1241), .ZN(
      n_257_76_1719));
   NOR2_X1 i_257_76_1722 (.A1(n_257_76_1718), .A2(n_257_76_1719), .ZN(
      n_257_76_1720));
   NAND2_X1 i_257_76_1723 (.A1(n_257_76_1717), .A2(n_257_76_1720), .ZN(
      n_257_76_1721));
   NAND2_X1 i_257_76_1724 (.A1(n_257_76_1307), .A2(n_257_76_1214), .ZN(
      n_257_76_1722));
   INV_X1 i_257_76_1725 (.A(n_257_76_1722), .ZN(n_257_76_1723));
   NOR2_X1 i_257_76_1726 (.A1(n_257_76_1612), .A2(n_257_76_1334), .ZN(
      n_257_76_1724));
   NAND2_X1 i_257_76_1727 (.A1(n_257_76_1723), .A2(n_257_76_1724), .ZN(
      n_257_76_1725));
   NOR2_X1 i_257_76_1728 (.A1(n_257_76_1721), .A2(n_257_76_1725), .ZN(
      n_257_76_1726));
   NAND2_X1 i_257_76_1729 (.A1(n_257_76_1306), .A2(n_257_76_1522), .ZN(
      n_257_76_1727));
   NOR2_X1 i_257_76_1730 (.A1(n_257_76_1279), .A2(n_257_76_1727), .ZN(
      n_257_76_1728));
   NAND2_X1 i_257_76_1731 (.A1(n_257_76_1726), .A2(n_257_76_1728), .ZN(
      n_257_76_1729));
   NOR2_X1 i_257_76_1732 (.A1(n_257_76_1729), .A2(n_257_76_1586), .ZN(
      n_257_76_1730));
   NAND2_X1 i_257_76_1733 (.A1(n_257_12), .A2(n_257_76_1730), .ZN(n_257_76_1731));
   NAND2_X1 i_257_76_1734 (.A1(n_257_76_1621), .A2(n_257_76_1602), .ZN(
      n_257_76_1732));
   INV_X1 i_257_76_1735 (.A(n_257_76_1732), .ZN(n_257_76_1733));
   NAND2_X1 i_257_76_1736 (.A1(n_257_76_1300), .A2(n_257_76_1384), .ZN(
      n_257_76_1734));
   NAND2_X1 i_257_76_1737 (.A1(n_257_671), .A2(n_257_76_17958), .ZN(
      n_257_76_1735));
   NAND2_X1 i_257_76_1738 (.A1(n_257_154), .A2(n_257_76_17331), .ZN(
      n_257_76_1736));
   NAND2_X1 i_257_76_1739 (.A1(n_257_76_1735), .A2(n_257_76_1736), .ZN(
      n_257_76_1737));
   NOR2_X1 i_257_76_1740 (.A1(n_257_76_1734), .A2(n_257_76_1737), .ZN(
      n_257_76_1738));
   NAND2_X1 i_257_76_1741 (.A1(n_257_767), .A2(n_257_442), .ZN(n_257_76_1739));
   INV_X1 i_257_76_1742 (.A(n_257_76_1739), .ZN(n_257_76_1740));
   AOI22_X1 i_257_76_1743 (.A1(n_257_449), .A2(n_257_76_9364), .B1(n_257_447), 
      .B2(n_257_76_1740), .ZN(n_257_76_1741));
   AOI22_X1 i_257_76_1744 (.A1(n_257_799), .A2(n_257_76_17952), .B1(n_257_37), 
      .B2(n_257_76_17918), .ZN(n_257_76_1742));
   NAND2_X1 i_257_76_1745 (.A1(n_257_76_1741), .A2(n_257_76_1742), .ZN(
      n_257_76_1743));
   INV_X1 i_257_76_1746 (.A(Small_Packet_Data_Size[2]), .ZN(n_257_76_1744));
   NAND2_X1 i_257_76_1747 (.A1(n_257_76_1707), .A2(n_257_76_18057), .ZN(
      n_257_76_1745));
   INV_X1 i_257_76_1748 (.A(n_257_76_1745), .ZN(n_257_76_1746));
   NAND2_X1 i_257_76_1749 (.A1(n_257_76_1746), .A2(n_257_76_1342), .ZN(
      n_257_76_1747));
   NAND2_X1 i_257_76_1750 (.A1(n_257_599), .A2(n_257_442), .ZN(n_257_76_1748));
   INV_X1 i_257_76_1751 (.A(n_257_76_1748), .ZN(n_257_76_1749));
   NAND2_X1 i_257_76_1752 (.A1(n_257_432), .A2(n_257_76_1749), .ZN(n_257_76_1750));
   INV_X1 i_257_76_1753 (.A(n_257_76_1750), .ZN(n_257_76_1751));
   NOR2_X1 i_257_76_1754 (.A1(n_257_76_1747), .A2(n_257_76_1751), .ZN(
      n_257_76_1752));
   NAND2_X1 i_257_76_1755 (.A1(n_257_76_1752), .A2(n_257_76_1507), .ZN(
      n_257_76_1753));
   NAND3_X1 i_257_76_1756 (.A1(n_257_703), .A2(n_257_435), .A3(n_257_442), 
      .ZN(n_257_76_1754));
   INV_X1 i_257_76_1757 (.A(n_257_631), .ZN(n_257_76_1755));
   OAI21_X1 i_257_76_1758 (.A(n_257_76_1754), .B1(n_257_76_1755), .B2(
      n_257_76_17927), .ZN(n_257_76_1756));
   NOR2_X1 i_257_76_1759 (.A1(n_257_76_1753), .A2(n_257_76_1756), .ZN(
      n_257_76_1757));
   NAND2_X1 i_257_76_1760 (.A1(n_257_442), .A2(n_257_933), .ZN(n_257_76_1758));
   INV_X1 i_257_76_1761 (.A(n_257_76_1758), .ZN(n_257_76_1759));
   NAND2_X1 i_257_76_1762 (.A1(n_257_440), .A2(n_257_76_1759), .ZN(n_257_76_1760));
   NAND2_X1 i_257_76_1763 (.A1(n_257_438), .A2(n_257_76_4949), .ZN(n_257_76_1761));
   NAND2_X1 i_257_76_1764 (.A1(n_257_76_1760), .A2(n_257_76_1761), .ZN(
      n_257_76_1762));
   NAND3_X1 i_257_76_1765 (.A1(n_257_439), .A2(n_257_901), .A3(n_257_442), 
      .ZN(n_257_76_1763));
   INV_X1 i_257_76_1766 (.A(n_257_76_1763), .ZN(n_257_76_1764));
   NOR2_X1 i_257_76_1767 (.A1(n_257_76_1762), .A2(n_257_76_1764), .ZN(
      n_257_76_1765));
   NAND2_X1 i_257_76_1768 (.A1(n_257_76_1757), .A2(n_257_76_1765), .ZN(
      n_257_76_1766));
   NOR2_X1 i_257_76_1769 (.A1(n_257_76_1743), .A2(n_257_76_1766), .ZN(
      n_257_76_1767));
   NAND2_X1 i_257_76_1770 (.A1(n_257_115), .A2(n_257_76_17925), .ZN(
      n_257_76_1768));
   NAND2_X1 i_257_76_1771 (.A1(n_257_735), .A2(n_257_76_17935), .ZN(
      n_257_76_1769));
   NAND2_X1 i_257_76_1772 (.A1(n_257_76_1768), .A2(n_257_76_1769), .ZN(
      n_257_76_1770));
   NAND2_X1 i_257_76_1773 (.A1(n_257_863), .A2(n_257_76_17903), .ZN(
      n_257_76_1771));
   NAND2_X1 i_257_76_1774 (.A1(n_257_831), .A2(n_257_442), .ZN(n_257_76_1772));
   INV_X1 i_257_76_1775 (.A(n_257_76_1772), .ZN(n_257_76_1773));
   NAND2_X1 i_257_76_1776 (.A1(n_257_446), .A2(n_257_76_1773), .ZN(n_257_76_1774));
   NAND2_X1 i_257_76_1777 (.A1(n_257_76_1771), .A2(n_257_76_1774), .ZN(
      n_257_76_1775));
   NOR2_X1 i_257_76_1778 (.A1(n_257_76_1770), .A2(n_257_76_1775), .ZN(
      n_257_76_1776));
   NAND2_X1 i_257_76_1779 (.A1(n_257_76_1767), .A2(n_257_76_1776), .ZN(
      n_257_76_1777));
   NAND2_X1 i_257_76_1780 (.A1(n_257_965), .A2(n_257_442), .ZN(n_257_76_1778));
   INV_X1 i_257_76_1781 (.A(n_257_76_1778), .ZN(n_257_76_1779));
   NAND2_X1 i_257_76_1782 (.A1(n_257_441), .A2(n_257_76_1779), .ZN(n_257_76_1780));
   NAND2_X1 i_257_76_1783 (.A1(n_257_76_1780), .A2(n_257_76_1633), .ZN(
      n_257_76_1781));
   NAND2_X1 i_257_76_1784 (.A1(n_257_454), .A2(n_257_442), .ZN(n_257_76_1782));
   INV_X1 i_257_76_1785 (.A(n_257_76_1782), .ZN(n_257_76_1783));
   NAND2_X1 i_257_76_1786 (.A1(n_257_451), .A2(n_257_76_1783), .ZN(n_257_76_1784));
   NAND2_X1 i_257_76_1787 (.A1(n_257_76_1664), .A2(n_257_76_1784), .ZN(
      n_257_76_1785));
   NOR2_X1 i_257_76_1788 (.A1(n_257_76_1781), .A2(n_257_76_1785), .ZN(
      n_257_76_1786));
   INV_X1 i_257_76_1789 (.A(n_257_76_1689), .ZN(n_257_76_1787));
   AOI21_X1 i_257_76_1790 (.A(n_257_76_1787), .B1(n_257_77), .B2(n_257_76_17932), 
      .ZN(n_257_76_1788));
   NAND2_X1 i_257_76_1791 (.A1(n_257_76_1786), .A2(n_257_76_1788), .ZN(
      n_257_76_1789));
   NOR2_X1 i_257_76_1792 (.A1(n_257_76_1777), .A2(n_257_76_1789), .ZN(
      n_257_76_1790));
   NAND2_X1 i_257_76_1793 (.A1(n_257_76_1738), .A2(n_257_76_1790), .ZN(
      n_257_76_1791));
   NAND2_X1 i_257_76_1794 (.A1(n_257_1029), .A2(n_257_76_17969), .ZN(
      n_257_76_1792));
   NAND2_X1 i_257_76_1795 (.A1(n_257_997), .A2(n_257_76_17964), .ZN(
      n_257_76_1793));
   NAND2_X1 i_257_76_1796 (.A1(n_257_76_1792), .A2(n_257_76_1793), .ZN(
      n_257_76_1794));
   NOR2_X1 i_257_76_1797 (.A1(n_257_76_1791), .A2(n_257_76_1794), .ZN(
      n_257_76_1795));
   NAND2_X1 i_257_76_1798 (.A1(n_257_76_1733), .A2(n_257_76_1795), .ZN(
      n_257_76_1796));
   NAND3_X1 i_257_76_1799 (.A1(n_257_76_1695), .A2(n_257_76_1731), .A3(
      n_257_76_1796), .ZN(n_257_76_1797));
   INV_X1 i_257_76_1800 (.A(n_257_76_1797), .ZN(n_257_76_1798));
   NAND3_X1 i_257_76_1801 (.A1(n_257_76_1625), .A2(n_257_76_1678), .A3(
      n_257_76_1798), .ZN(n_257_76_1799));
   NOR2_X1 i_257_76_1802 (.A1(n_257_76_1572), .A2(n_257_76_1799), .ZN(
      n_257_76_1800));
   NAND2_X1 i_257_76_1803 (.A1(n_257_76_1447), .A2(n_257_76_1800), .ZN(n_2));
   NAND2_X1 i_257_76_1804 (.A1(n_257_998), .A2(n_257_444), .ZN(n_257_76_1801));
   NAND2_X1 i_257_76_1805 (.A1(n_257_441), .A2(n_257_966), .ZN(n_257_76_1802));
   INV_X1 i_257_76_1806 (.A(n_257_1062), .ZN(n_257_76_1803));
   NAND2_X1 i_257_76_1807 (.A1(n_257_76_1803), .A2(n_257_442), .ZN(n_257_76_1804));
   INV_X1 i_257_76_1808 (.A(n_257_934), .ZN(n_257_76_1805));
   NOR2_X1 i_257_76_1809 (.A1(n_257_76_1804), .A2(n_257_76_1805), .ZN(
      n_257_76_1806));
   NAND2_X1 i_257_76_1810 (.A1(n_257_440), .A2(n_257_76_1806), .ZN(n_257_76_1807));
   INV_X1 i_257_76_1811 (.A(n_257_76_1807), .ZN(n_257_76_1808));
   NAND2_X1 i_257_76_1812 (.A1(n_257_76_1802), .A2(n_257_76_1808), .ZN(
      n_257_76_1809));
   INV_X1 i_257_76_1813 (.A(n_257_76_1809), .ZN(n_257_76_1810));
   NAND2_X1 i_257_76_1814 (.A1(n_257_76_1801), .A2(n_257_76_1810), .ZN(
      n_257_76_1811));
   INV_X1 i_257_76_1815 (.A(n_257_76_1811), .ZN(n_257_76_1812));
   NAND2_X1 i_257_76_1816 (.A1(n_257_1030), .A2(n_257_443), .ZN(n_257_76_1813));
   NAND2_X1 i_257_76_1817 (.A1(n_257_76_1812), .A2(n_257_76_1813), .ZN(
      n_257_76_1814));
   INV_X1 i_257_76_1818 (.A(n_257_76_1814), .ZN(n_257_76_1815));
   NAND2_X1 i_257_76_1819 (.A1(n_257_17), .A2(n_257_76_1815), .ZN(n_257_76_1816));
   INV_X1 i_257_76_1820 (.A(n_257_76_1804), .ZN(n_257_76_1817));
   NAND2_X1 i_257_76_1821 (.A1(n_257_443), .A2(n_257_76_1817), .ZN(n_257_76_1818));
   INV_X1 i_257_76_1822 (.A(n_257_76_1818), .ZN(n_257_76_1819));
   NAND2_X1 i_257_76_1823 (.A1(n_257_1030), .A2(n_257_76_1819), .ZN(
      n_257_76_1820));
   INV_X1 i_257_76_1824 (.A(n_257_76_1820), .ZN(n_257_76_1821));
   NAND2_X1 i_257_76_1825 (.A1(n_257_14), .A2(n_257_76_1821), .ZN(n_257_76_1822));
   NAND2_X1 i_257_76_1826 (.A1(n_257_736), .A2(n_257_436), .ZN(n_257_76_1823));
   NAND2_X1 i_257_76_1827 (.A1(n_257_76_1802), .A2(n_257_76_1823), .ZN(
      n_257_76_1824));
   NAND2_X1 i_257_76_1828 (.A1(n_257_864), .A2(n_257_445), .ZN(n_257_76_1825));
   NAND2_X1 i_257_76_1829 (.A1(n_257_800), .A2(n_257_437), .ZN(n_257_76_1826));
   NAND2_X1 i_257_76_1830 (.A1(n_257_446), .A2(n_257_832), .ZN(n_257_76_1827));
   NAND3_X1 i_257_76_1831 (.A1(n_257_76_1825), .A2(n_257_76_1826), .A3(
      n_257_76_1827), .ZN(n_257_76_1828));
   NOR2_X1 i_257_76_1832 (.A1(n_257_76_1824), .A2(n_257_76_1828), .ZN(
      n_257_76_1829));
   NAND2_X1 i_257_76_1833 (.A1(n_257_672), .A2(n_257_448), .ZN(n_257_76_1830));
   NAND2_X1 i_257_76_1834 (.A1(n_257_704), .A2(n_257_435), .ZN(n_257_76_1831));
   NAND2_X1 i_257_76_1835 (.A1(n_257_450), .A2(n_257_76_1817), .ZN(n_257_76_1832));
   INV_X1 i_257_76_1836 (.A(n_257_76_1832), .ZN(n_257_76_1833));
   NAND3_X1 i_257_76_1837 (.A1(n_257_632), .A2(n_257_76_1831), .A3(n_257_76_1833), 
      .ZN(n_257_76_1834));
   INV_X1 i_257_76_1838 (.A(n_257_76_1834), .ZN(n_257_76_1835));
   NAND2_X1 i_257_76_1839 (.A1(n_257_440), .A2(n_257_934), .ZN(n_257_76_1836));
   NAND2_X1 i_257_76_1840 (.A1(n_257_438), .A2(n_257_1068), .ZN(n_257_76_1837));
   NAND2_X1 i_257_76_1841 (.A1(n_257_439), .A2(n_257_902), .ZN(n_257_76_1838));
   NAND4_X1 i_257_76_1842 (.A1(n_257_76_1835), .A2(n_257_76_1836), .A3(
      n_257_76_1837), .A4(n_257_76_1838), .ZN(n_257_76_1839));
   NAND2_X1 i_257_76_1843 (.A1(n_257_449), .A2(n_257_1076), .ZN(n_257_76_1840));
   NAND2_X1 i_257_76_1844 (.A1(n_257_447), .A2(n_257_768), .ZN(n_257_76_1841));
   NAND2_X1 i_257_76_1845 (.A1(n_257_76_1840), .A2(n_257_76_1841), .ZN(
      n_257_76_1842));
   NOR2_X1 i_257_76_1846 (.A1(n_257_76_1839), .A2(n_257_76_1842), .ZN(
      n_257_76_1843));
   NAND3_X1 i_257_76_1847 (.A1(n_257_76_1829), .A2(n_257_76_1830), .A3(
      n_257_76_1843), .ZN(n_257_76_1844));
   INV_X1 i_257_76_1848 (.A(n_257_76_1844), .ZN(n_257_76_1845));
   NAND2_X1 i_257_76_1849 (.A1(n_257_76_1845), .A2(n_257_76_1801), .ZN(
      n_257_76_1846));
   INV_X1 i_257_76_1850 (.A(n_257_76_1813), .ZN(n_257_76_1847));
   NOR2_X1 i_257_76_1851 (.A1(n_257_76_1846), .A2(n_257_76_1847), .ZN(
      n_257_76_1848));
   NAND2_X1 i_257_76_1852 (.A1(n_257_28), .A2(n_257_76_1848), .ZN(n_257_76_1849));
   NAND3_X1 i_257_76_1853 (.A1(n_257_76_1816), .A2(n_257_76_1822), .A3(
      n_257_76_1849), .ZN(n_257_76_1850));
   NAND3_X1 i_257_76_1854 (.A1(n_257_446), .A2(n_257_76_1836), .A3(n_257_76_1837), 
      .ZN(n_257_76_1851));
   INV_X1 i_257_76_1855 (.A(n_257_76_1851), .ZN(n_257_76_1852));
   NAND2_X1 i_257_76_1856 (.A1(n_257_832), .A2(n_257_76_1817), .ZN(n_257_76_1853));
   INV_X1 i_257_76_1857 (.A(n_257_76_1853), .ZN(n_257_76_1854));
   NAND2_X1 i_257_76_1858 (.A1(n_257_76_1838), .A2(n_257_76_1854), .ZN(
      n_257_76_1855));
   INV_X1 i_257_76_1859 (.A(n_257_76_1855), .ZN(n_257_76_1856));
   NAND4_X1 i_257_76_1860 (.A1(n_257_76_1802), .A2(n_257_76_1852), .A3(
      n_257_76_1825), .A4(n_257_76_1856), .ZN(n_257_76_1857));
   INV_X1 i_257_76_1861 (.A(n_257_76_1857), .ZN(n_257_76_1858));
   NAND2_X1 i_257_76_1862 (.A1(n_257_76_1801), .A2(n_257_76_1858), .ZN(
      n_257_76_1859));
   INV_X1 i_257_76_1863 (.A(n_257_76_1859), .ZN(n_257_76_1860));
   NAND2_X1 i_257_76_1864 (.A1(n_257_76_1860), .A2(n_257_76_1813), .ZN(
      n_257_76_1861));
   INV_X1 i_257_76_1865 (.A(n_257_76_1861), .ZN(n_257_76_1862));
   NAND2_X1 i_257_76_1866 (.A1(n_257_21), .A2(n_257_76_1862), .ZN(n_257_76_1863));
   INV_X1 i_257_76_1867 (.A(n_257_76_1836), .ZN(n_257_76_1864));
   NAND3_X1 i_257_76_1868 (.A1(n_257_439), .A2(n_257_902), .A3(n_257_76_1817), 
      .ZN(n_257_76_1865));
   NOR2_X1 i_257_76_1869 (.A1(n_257_76_1864), .A2(n_257_76_1865), .ZN(
      n_257_76_1866));
   NAND2_X1 i_257_76_1870 (.A1(n_257_76_1802), .A2(n_257_76_1866), .ZN(
      n_257_76_1867));
   INV_X1 i_257_76_1871 (.A(n_257_76_1867), .ZN(n_257_76_1868));
   NAND2_X1 i_257_76_1872 (.A1(n_257_76_1801), .A2(n_257_76_1868), .ZN(
      n_257_76_1869));
   INV_X1 i_257_76_1873 (.A(n_257_76_1869), .ZN(n_257_76_1870));
   NAND2_X1 i_257_76_1874 (.A1(n_257_76_1870), .A2(n_257_76_1813), .ZN(
      n_257_76_1871));
   INV_X1 i_257_76_1875 (.A(n_257_76_1871), .ZN(n_257_76_1872));
   NAND2_X1 i_257_76_1876 (.A1(n_257_18), .A2(n_257_76_1872), .ZN(n_257_76_1873));
   NAND2_X1 i_257_76_1877 (.A1(n_257_536), .A2(n_257_426), .ZN(n_257_76_1874));
   NAND2_X1 i_257_76_1878 (.A1(n_257_38), .A2(n_257_433), .ZN(n_257_76_1875));
   NAND3_X1 i_257_76_1879 (.A1(n_257_76_1874), .A2(n_257_275), .A3(n_257_76_1875), 
      .ZN(n_257_76_1876));
   INV_X1 i_257_76_1880 (.A(n_257_76_1826), .ZN(n_257_76_1877));
   NOR2_X1 i_257_76_1881 (.A1(n_257_76_1876), .A2(n_257_76_1877), .ZN(
      n_257_76_1878));
   NAND2_X1 i_257_76_1882 (.A1(n_257_76_1823), .A2(n_257_76_1825), .ZN(
      n_257_76_1879));
   INV_X1 i_257_76_1883 (.A(n_257_76_1879), .ZN(n_257_76_1880));
   NAND2_X1 i_257_76_1884 (.A1(n_257_504), .A2(n_257_424), .ZN(n_257_76_1881));
   NAND2_X1 i_257_76_1885 (.A1(n_257_76_1881), .A2(n_257_76_1831), .ZN(
      n_257_76_1882));
   INV_X1 i_257_76_1886 (.A(n_257_76_1882), .ZN(n_257_76_1883));
   NAND2_X1 i_257_76_1887 (.A1(n_257_632), .A2(n_257_450), .ZN(n_257_76_1884));
   NAND2_X1 i_257_76_1888 (.A1(n_257_195), .A2(n_257_427), .ZN(n_257_76_1885));
   NAND2_X1 i_257_76_1889 (.A1(n_257_432), .A2(n_257_600), .ZN(n_257_76_1886));
   NAND2_X1 i_257_76_1890 (.A1(n_257_428), .A2(n_257_568), .ZN(n_257_76_1887));
   NAND2_X1 i_257_76_1891 (.A1(n_257_423), .A2(n_257_76_1817), .ZN(n_257_76_1888));
   INV_X1 i_257_76_1892 (.A(n_257_76_1888), .ZN(n_257_76_1889));
   NAND3_X1 i_257_76_1893 (.A1(n_257_76_1886), .A2(n_257_76_1887), .A3(
      n_257_76_1889), .ZN(n_257_76_1890));
   INV_X1 i_257_76_1894 (.A(n_257_76_1890), .ZN(n_257_76_1891));
   NAND4_X1 i_257_76_1895 (.A1(n_257_76_1883), .A2(n_257_76_1884), .A3(
      n_257_76_1885), .A4(n_257_76_1891), .ZN(n_257_76_1892));
   NAND3_X1 i_257_76_1896 (.A1(n_257_76_1836), .A2(n_257_76_1837), .A3(
      n_257_76_1838), .ZN(n_257_76_1893));
   NOR2_X1 i_257_76_1897 (.A1(n_257_76_1892), .A2(n_257_76_1893), .ZN(
      n_257_76_1894));
   NAND2_X1 i_257_76_1898 (.A1(n_257_116), .A2(n_257_430), .ZN(n_257_76_1895));
   NAND4_X1 i_257_76_1899 (.A1(n_257_76_1878), .A2(n_257_76_1880), .A3(
      n_257_76_1894), .A4(n_257_76_1895), .ZN(n_257_76_1896));
   INV_X1 i_257_76_1900 (.A(n_257_76_1896), .ZN(n_257_76_1897));
   NAND2_X1 i_257_76_1901 (.A1(n_257_76_1801), .A2(n_257_76_1897), .ZN(
      n_257_76_1898));
   INV_X1 i_257_76_1902 (.A(n_257_76_1898), .ZN(n_257_76_1899));
   NAND2_X1 i_257_76_1903 (.A1(n_257_78), .A2(n_257_431), .ZN(n_257_76_1900));
   NAND2_X1 i_257_76_1904 (.A1(n_257_451), .A2(n_257_455), .ZN(n_257_76_1901));
   NAND2_X1 i_257_76_1905 (.A1(n_257_76_1802), .A2(n_257_76_1901), .ZN(
      n_257_76_1902));
   INV_X1 i_257_76_1906 (.A(n_257_76_1902), .ZN(n_257_76_1903));
   NAND3_X1 i_257_76_1907 (.A1(n_257_76_1827), .A2(n_257_76_1840), .A3(
      n_257_76_1841), .ZN(n_257_76_1904));
   INV_X1 i_257_76_1908 (.A(n_257_76_1904), .ZN(n_257_76_1905));
   NAND3_X1 i_257_76_1909 (.A1(n_257_76_1900), .A2(n_257_76_1903), .A3(
      n_257_76_1905), .ZN(n_257_76_1906));
   INV_X1 i_257_76_1910 (.A(n_257_76_1906), .ZN(n_257_76_1907));
   NAND2_X1 i_257_76_1911 (.A1(n_257_155), .A2(n_257_429), .ZN(n_257_76_1908));
   NAND3_X1 i_257_76_1912 (.A1(n_257_76_1907), .A2(n_257_76_1908), .A3(
      n_257_76_1830), .ZN(n_257_76_1909));
   INV_X1 i_257_76_1913 (.A(n_257_76_1909), .ZN(n_257_76_1910));
   NAND2_X1 i_257_76_1914 (.A1(n_257_235), .A2(n_257_425), .ZN(n_257_76_1911));
   NAND4_X1 i_257_76_1915 (.A1(n_257_76_1899), .A2(n_257_76_1813), .A3(
      n_257_76_1910), .A4(n_257_76_1911), .ZN(n_257_76_1912));
   INV_X1 i_257_76_1916 (.A(n_257_76_1912), .ZN(n_257_76_1913));
   NAND2_X1 i_257_76_1917 (.A1(n_257_304), .A2(n_257_76_1913), .ZN(n_257_76_1914));
   NAND3_X1 i_257_76_1918 (.A1(n_257_76_1863), .A2(n_257_76_1873), .A3(
      n_257_76_1914), .ZN(n_257_76_1915));
   NOR2_X1 i_257_76_1919 (.A1(n_257_76_1850), .A2(n_257_76_1915), .ZN(
      n_257_76_1916));
   NAND2_X1 i_257_76_1920 (.A1(n_257_966), .A2(n_257_76_1817), .ZN(n_257_76_1917));
   INV_X1 i_257_76_1921 (.A(n_257_76_1917), .ZN(n_257_76_1918));
   NAND2_X1 i_257_76_1922 (.A1(n_257_441), .A2(n_257_76_1918), .ZN(n_257_76_1919));
   INV_X1 i_257_76_1923 (.A(n_257_76_1919), .ZN(n_257_76_1920));
   NAND2_X1 i_257_76_1924 (.A1(n_257_76_1801), .A2(n_257_76_1920), .ZN(
      n_257_76_1921));
   INV_X1 i_257_76_1925 (.A(n_257_76_1921), .ZN(n_257_76_1922));
   NAND2_X1 i_257_76_1926 (.A1(n_257_76_1922), .A2(n_257_76_1813), .ZN(
      n_257_76_1923));
   INV_X1 i_257_76_1927 (.A(n_257_76_1923), .ZN(n_257_76_1924));
   NAND2_X1 i_257_76_1928 (.A1(n_257_16), .A2(n_257_76_1924), .ZN(n_257_76_1925));
   INV_X1 i_257_76_1929 (.A(n_257_704), .ZN(n_257_76_1926));
   NAND2_X1 i_257_76_1930 (.A1(n_257_435), .A2(n_257_76_1817), .ZN(n_257_76_1927));
   NOR2_X1 i_257_76_1931 (.A1(n_257_76_1926), .A2(n_257_76_1927), .ZN(
      n_257_76_1928));
   NAND4_X1 i_257_76_1932 (.A1(n_257_76_1836), .A2(n_257_76_1837), .A3(
      n_257_76_1838), .A4(n_257_76_1928), .ZN(n_257_76_1929));
   INV_X1 i_257_76_1933 (.A(n_257_76_1929), .ZN(n_257_76_1930));
   NAND4_X1 i_257_76_1934 (.A1(n_257_76_1930), .A2(n_257_76_1826), .A3(
      n_257_76_1827), .A4(n_257_76_1841), .ZN(n_257_76_1931));
   NAND3_X1 i_257_76_1935 (.A1(n_257_76_1802), .A2(n_257_76_1823), .A3(
      n_257_76_1825), .ZN(n_257_76_1932));
   NOR2_X1 i_257_76_1936 (.A1(n_257_76_1931), .A2(n_257_76_1932), .ZN(
      n_257_76_1933));
   NAND2_X1 i_257_76_1937 (.A1(n_257_76_1801), .A2(n_257_76_1933), .ZN(
      n_257_76_1934));
   INV_X1 i_257_76_1938 (.A(n_257_76_1934), .ZN(n_257_76_1935));
   NAND2_X1 i_257_76_1939 (.A1(n_257_76_1935), .A2(n_257_76_1813), .ZN(
      n_257_76_1936));
   INV_X1 i_257_76_1940 (.A(n_257_76_1936), .ZN(n_257_76_1937));
   NAND2_X1 i_257_76_1941 (.A1(n_257_25), .A2(n_257_76_1937), .ZN(n_257_76_1938));
   NAND3_X1 i_257_76_1942 (.A1(n_257_76_1895), .A2(n_257_76_1802), .A3(
      n_257_76_1901), .ZN(n_257_76_1939));
   INV_X1 i_257_76_1943 (.A(n_257_76_1939), .ZN(n_257_76_1940));
   NAND3_X1 i_257_76_1944 (.A1(n_257_76_1826), .A2(n_257_76_1827), .A3(
      n_257_76_1840), .ZN(n_257_76_1941));
   NOR2_X1 i_257_76_1945 (.A1(n_257_76_1941), .A2(n_257_76_1879), .ZN(
      n_257_76_1942));
   NAND3_X1 i_257_76_1946 (.A1(n_257_76_1841), .A2(n_257_76_1875), .A3(
      n_257_76_1836), .ZN(n_257_76_1943));
   INV_X1 i_257_76_1947 (.A(n_257_76_1831), .ZN(n_257_76_1944));
   NAND3_X1 i_257_76_1948 (.A1(n_257_76_1803), .A2(n_257_442), .A3(n_257_568), 
      .ZN(n_257_76_1945));
   INV_X1 i_257_76_1949 (.A(n_257_76_1945), .ZN(n_257_76_1946));
   NAND2_X1 i_257_76_1950 (.A1(n_257_428), .A2(n_257_76_1946), .ZN(n_257_76_1947));
   INV_X1 i_257_76_1951 (.A(n_257_76_1947), .ZN(n_257_76_1948));
   NAND2_X1 i_257_76_1952 (.A1(n_257_76_1886), .A2(n_257_76_1948), .ZN(
      n_257_76_1949));
   NOR2_X1 i_257_76_1953 (.A1(n_257_76_1944), .A2(n_257_76_1949), .ZN(
      n_257_76_1950));
   NAND4_X1 i_257_76_1954 (.A1(n_257_76_1950), .A2(n_257_76_1837), .A3(
      n_257_76_1838), .A4(n_257_76_1884), .ZN(n_257_76_1951));
   NOR2_X1 i_257_76_1955 (.A1(n_257_76_1943), .A2(n_257_76_1951), .ZN(
      n_257_76_1952));
   NAND4_X1 i_257_76_1956 (.A1(n_257_76_1940), .A2(n_257_76_1942), .A3(
      n_257_76_1900), .A4(n_257_76_1952), .ZN(n_257_76_1953));
   INV_X1 i_257_76_1957 (.A(n_257_76_1953), .ZN(n_257_76_1954));
   NAND2_X1 i_257_76_1958 (.A1(n_257_76_1908), .A2(n_257_76_1830), .ZN(
      n_257_76_1955));
   INV_X1 i_257_76_1959 (.A(n_257_76_1955), .ZN(n_257_76_1956));
   NAND3_X1 i_257_76_1960 (.A1(n_257_76_1954), .A2(n_257_76_1956), .A3(
      n_257_76_1801), .ZN(n_257_76_1957));
   NOR2_X1 i_257_76_1961 (.A1(n_257_76_1957), .A2(n_257_76_1847), .ZN(
      n_257_76_1958));
   NAND2_X1 i_257_76_1962 (.A1(n_257_185), .A2(n_257_76_1958), .ZN(n_257_76_1959));
   NAND3_X1 i_257_76_1963 (.A1(n_257_76_1925), .A2(n_257_76_1938), .A3(
      n_257_76_1959), .ZN(n_257_76_1960));
   NAND2_X1 i_257_76_1964 (.A1(n_257_442), .A2(n_257_1062), .ZN(n_257_76_1961));
   INV_X1 i_257_76_1965 (.A(n_257_76_1961), .ZN(n_257_76_1962));
   NAND2_X1 i_257_76_1966 (.A1(n_257_13), .A2(n_257_76_1962), .ZN(n_257_76_1963));
   NAND2_X1 i_257_76_1967 (.A1(n_257_864), .A2(n_257_76_1836), .ZN(n_257_76_1964));
   INV_X1 i_257_76_1968 (.A(n_257_76_1964), .ZN(n_257_76_1965));
   NAND2_X1 i_257_76_1969 (.A1(n_257_445), .A2(n_257_76_1817), .ZN(n_257_76_1966));
   INV_X1 i_257_76_1970 (.A(n_257_76_1966), .ZN(n_257_76_1967));
   NAND3_X1 i_257_76_1971 (.A1(n_257_76_1837), .A2(n_257_76_1838), .A3(
      n_257_76_1967), .ZN(n_257_76_1968));
   INV_X1 i_257_76_1972 (.A(n_257_76_1968), .ZN(n_257_76_1969));
   NAND3_X1 i_257_76_1973 (.A1(n_257_76_1802), .A2(n_257_76_1965), .A3(
      n_257_76_1969), .ZN(n_257_76_1970));
   INV_X1 i_257_76_1974 (.A(n_257_76_1970), .ZN(n_257_76_1971));
   NAND2_X1 i_257_76_1975 (.A1(n_257_76_1801), .A2(n_257_76_1971), .ZN(
      n_257_76_1972));
   INV_X1 i_257_76_1976 (.A(n_257_76_1972), .ZN(n_257_76_1973));
   NAND2_X1 i_257_76_1977 (.A1(n_257_76_1973), .A2(n_257_76_1813), .ZN(
      n_257_76_1974));
   INV_X1 i_257_76_1978 (.A(n_257_76_1974), .ZN(n_257_76_1975));
   NAND2_X1 i_257_76_1979 (.A1(n_257_20), .A2(n_257_76_1975), .ZN(n_257_76_1976));
   NAND2_X1 i_257_76_1980 (.A1(n_257_76_1963), .A2(n_257_76_1976), .ZN(
      n_257_76_1977));
   NOR2_X1 i_257_76_1981 (.A1(n_257_76_1960), .A2(n_257_76_1977), .ZN(
      n_257_76_1978));
   INV_X1 i_257_76_1982 (.A(n_257_76_1801), .ZN(n_257_76_1979));
   NAND4_X1 i_257_76_1983 (.A1(n_257_76_1875), .A2(n_257_76_1836), .A3(
      n_257_76_1837), .A4(n_257_536), .ZN(n_257_76_1980));
   INV_X1 i_257_76_1984 (.A(n_257_76_1887), .ZN(n_257_76_1981));
   NAND2_X1 i_257_76_1985 (.A1(n_257_426), .A2(n_257_76_1817), .ZN(n_257_76_1982));
   NOR2_X1 i_257_76_1986 (.A1(n_257_76_1981), .A2(n_257_76_1982), .ZN(
      n_257_76_1983));
   NAND3_X1 i_257_76_1987 (.A1(n_257_76_1831), .A2(n_257_76_1983), .A3(
      n_257_76_1886), .ZN(n_257_76_1984));
   INV_X1 i_257_76_1988 (.A(n_257_76_1984), .ZN(n_257_76_1985));
   NAND4_X1 i_257_76_1989 (.A1(n_257_76_1985), .A2(n_257_76_1838), .A3(
      n_257_76_1884), .A4(n_257_76_1885), .ZN(n_257_76_1986));
   NOR2_X1 i_257_76_1990 (.A1(n_257_76_1980), .A2(n_257_76_1986), .ZN(
      n_257_76_1987));
   NAND3_X1 i_257_76_1991 (.A1(n_257_76_1823), .A2(n_257_76_1825), .A3(
      n_257_76_1826), .ZN(n_257_76_1988));
   INV_X1 i_257_76_1992 (.A(n_257_76_1988), .ZN(n_257_76_1989));
   NAND3_X1 i_257_76_1993 (.A1(n_257_76_1987), .A2(n_257_76_1989), .A3(
      n_257_76_1895), .ZN(n_257_76_1990));
   NOR2_X1 i_257_76_1994 (.A1(n_257_76_1979), .A2(n_257_76_1990), .ZN(
      n_257_76_1991));
   NAND3_X1 i_257_76_1995 (.A1(n_257_76_1991), .A2(n_257_76_1813), .A3(
      n_257_76_1910), .ZN(n_257_76_1992));
   INV_X1 i_257_76_1996 (.A(n_257_76_1992), .ZN(n_257_76_1993));
   NAND2_X1 i_257_76_1997 (.A1(n_257_225), .A2(n_257_76_1993), .ZN(n_257_76_1994));
   NAND2_X1 i_257_76_1998 (.A1(n_257_736), .A2(n_257_76_1836), .ZN(n_257_76_1995));
   INV_X1 i_257_76_1999 (.A(n_257_76_1995), .ZN(n_257_76_1996));
   NAND2_X1 i_257_76_2000 (.A1(n_257_436), .A2(n_257_76_1817), .ZN(n_257_76_1997));
   INV_X1 i_257_76_2001 (.A(n_257_76_1997), .ZN(n_257_76_1998));
   NAND3_X1 i_257_76_2002 (.A1(n_257_76_1837), .A2(n_257_76_1838), .A3(
      n_257_76_1998), .ZN(n_257_76_1999));
   INV_X1 i_257_76_2003 (.A(n_257_76_1999), .ZN(n_257_76_2000));
   NAND4_X1 i_257_76_2004 (.A1(n_257_76_1996), .A2(n_257_76_2000), .A3(
      n_257_76_1827), .A4(n_257_76_1841), .ZN(n_257_76_2001));
   NAND3_X1 i_257_76_2005 (.A1(n_257_76_1802), .A2(n_257_76_1825), .A3(
      n_257_76_1826), .ZN(n_257_76_2002));
   NOR2_X1 i_257_76_2006 (.A1(n_257_76_2001), .A2(n_257_76_2002), .ZN(
      n_257_76_2003));
   NAND2_X1 i_257_76_2007 (.A1(n_257_76_1801), .A2(n_257_76_2003), .ZN(
      n_257_76_2004));
   INV_X1 i_257_76_2008 (.A(n_257_76_2004), .ZN(n_257_76_2005));
   NAND2_X1 i_257_76_2009 (.A1(n_257_76_2005), .A2(n_257_76_1813), .ZN(
      n_257_76_2006));
   INV_X1 i_257_76_2010 (.A(n_257_76_2006), .ZN(n_257_76_2007));
   NAND2_X1 i_257_76_2011 (.A1(n_257_24), .A2(n_257_76_2007), .ZN(n_257_76_2008));
   NOR2_X1 i_257_76_2012 (.A1(n_257_76_1902), .A2(n_257_76_1988), .ZN(
      n_257_76_2009));
   INV_X1 i_257_76_2013 (.A(n_257_600), .ZN(n_257_76_2010));
   NOR2_X1 i_257_76_2014 (.A1(n_257_76_1804), .A2(n_257_76_2010), .ZN(
      n_257_76_2011));
   NAND2_X1 i_257_76_2015 (.A1(n_257_432), .A2(n_257_76_2011), .ZN(n_257_76_2012));
   INV_X1 i_257_76_2016 (.A(n_257_76_2012), .ZN(n_257_76_2013));
   NAND2_X1 i_257_76_2017 (.A1(n_257_76_1831), .A2(n_257_76_2013), .ZN(
      n_257_76_2014));
   INV_X1 i_257_76_2018 (.A(n_257_76_2014), .ZN(n_257_76_2015));
   NAND3_X1 i_257_76_2019 (.A1(n_257_76_2015), .A2(n_257_76_1838), .A3(
      n_257_76_1884), .ZN(n_257_76_2016));
   INV_X1 i_257_76_2020 (.A(n_257_76_2016), .ZN(n_257_76_2017));
   NAND2_X1 i_257_76_2021 (.A1(n_257_76_1836), .A2(n_257_76_1837), .ZN(
      n_257_76_2018));
   INV_X1 i_257_76_2022 (.A(n_257_76_2018), .ZN(n_257_76_2019));
   NAND3_X1 i_257_76_2023 (.A1(n_257_76_2017), .A2(n_257_76_2019), .A3(
      n_257_76_1875), .ZN(n_257_76_2020));
   NOR2_X1 i_257_76_2024 (.A1(n_257_76_2020), .A2(n_257_76_1904), .ZN(
      n_257_76_2021));
   NAND3_X1 i_257_76_2025 (.A1(n_257_76_2009), .A2(n_257_76_1830), .A3(
      n_257_76_2021), .ZN(n_257_76_2022));
   INV_X1 i_257_76_2026 (.A(n_257_76_2022), .ZN(n_257_76_2023));
   NAND2_X1 i_257_76_2027 (.A1(n_257_76_2023), .A2(n_257_76_1801), .ZN(
      n_257_76_2024));
   NOR2_X1 i_257_76_2028 (.A1(n_257_76_2024), .A2(n_257_76_1847), .ZN(
      n_257_76_2025));
   NAND2_X1 i_257_76_2029 (.A1(n_257_68), .A2(n_257_76_2025), .ZN(n_257_76_2026));
   NAND3_X1 i_257_76_2030 (.A1(n_257_76_1994), .A2(n_257_76_2008), .A3(
      n_257_76_2026), .ZN(n_257_76_2027));
   NAND2_X1 i_257_76_2031 (.A1(n_257_437), .A2(n_257_76_1817), .ZN(n_257_76_2028));
   INV_X1 i_257_76_2032 (.A(n_257_76_2028), .ZN(n_257_76_2029));
   NAND2_X1 i_257_76_2033 (.A1(n_257_76_1838), .A2(n_257_76_2029), .ZN(
      n_257_76_2030));
   INV_X1 i_257_76_2034 (.A(n_257_76_2030), .ZN(n_257_76_2031));
   NAND4_X1 i_257_76_2035 (.A1(n_257_76_2019), .A2(n_257_76_1827), .A3(
      n_257_76_2031), .A4(n_257_800), .ZN(n_257_76_2032));
   NAND2_X1 i_257_76_2036 (.A1(n_257_76_1802), .A2(n_257_76_1825), .ZN(
      n_257_76_2033));
   NOR2_X1 i_257_76_2037 (.A1(n_257_76_2032), .A2(n_257_76_2033), .ZN(
      n_257_76_2034));
   NAND2_X1 i_257_76_2038 (.A1(n_257_76_1801), .A2(n_257_76_2034), .ZN(
      n_257_76_2035));
   INV_X1 i_257_76_2039 (.A(n_257_76_2035), .ZN(n_257_76_2036));
   NAND2_X1 i_257_76_2040 (.A1(n_257_76_2036), .A2(n_257_76_1813), .ZN(
      n_257_76_2037));
   INV_X1 i_257_76_2041 (.A(n_257_76_2037), .ZN(n_257_76_2038));
   NAND2_X1 i_257_76_2042 (.A1(n_257_22), .A2(n_257_76_2038), .ZN(n_257_76_2039));
   NAND2_X1 i_257_76_2043 (.A1(n_257_444), .A2(n_257_76_1817), .ZN(n_257_76_2040));
   INV_X1 i_257_76_2044 (.A(n_257_76_2040), .ZN(n_257_76_2041));
   NAND2_X1 i_257_76_2045 (.A1(n_257_998), .A2(n_257_76_2041), .ZN(n_257_76_2042));
   INV_X1 i_257_76_2046 (.A(n_257_76_2042), .ZN(n_257_76_2043));
   NAND2_X1 i_257_76_2047 (.A1(n_257_76_1813), .A2(n_257_76_2043), .ZN(
      n_257_76_2044));
   INV_X1 i_257_76_2048 (.A(n_257_76_2044), .ZN(n_257_76_2045));
   NAND2_X1 i_257_76_2049 (.A1(n_257_15), .A2(n_257_76_2045), .ZN(n_257_76_2046));
   NAND2_X1 i_257_76_2050 (.A1(n_257_76_2039), .A2(n_257_76_2046), .ZN(
      n_257_76_2047));
   NOR2_X1 i_257_76_2051 (.A1(n_257_76_2027), .A2(n_257_76_2047), .ZN(
      n_257_76_2048));
   NAND3_X1 i_257_76_2052 (.A1(n_257_76_1916), .A2(n_257_76_1978), .A3(
      n_257_76_2048), .ZN(n_257_76_2049));
   INV_X1 i_257_76_2053 (.A(n_257_76_2049), .ZN(n_257_76_2050));
   INV_X1 i_257_76_2054 (.A(n_257_38), .ZN(n_257_76_2051));
   NAND2_X1 i_257_76_2055 (.A1(n_257_433), .A2(n_257_76_1817), .ZN(n_257_76_2052));
   INV_X1 i_257_76_2056 (.A(n_257_76_2052), .ZN(n_257_76_2053));
   NAND2_X1 i_257_76_2057 (.A1(n_257_76_1831), .A2(n_257_76_2053), .ZN(
      n_257_76_2054));
   NOR2_X1 i_257_76_2058 (.A1(n_257_76_2051), .A2(n_257_76_2054), .ZN(
      n_257_76_2055));
   NAND2_X1 i_257_76_2059 (.A1(n_257_76_1838), .A2(n_257_76_1884), .ZN(
      n_257_76_2056));
   INV_X1 i_257_76_2060 (.A(n_257_76_2056), .ZN(n_257_76_2057));
   NAND3_X1 i_257_76_2061 (.A1(n_257_76_2055), .A2(n_257_76_2019), .A3(
      n_257_76_2057), .ZN(n_257_76_2058));
   NOR2_X1 i_257_76_2062 (.A1(n_257_76_2058), .A2(n_257_76_1904), .ZN(
      n_257_76_2059));
   NAND3_X1 i_257_76_2063 (.A1(n_257_76_2009), .A2(n_257_76_1830), .A3(
      n_257_76_2059), .ZN(n_257_76_2060));
   INV_X1 i_257_76_2064 (.A(n_257_76_2060), .ZN(n_257_76_2061));
   NAND2_X1 i_257_76_2065 (.A1(n_257_76_2061), .A2(n_257_76_1801), .ZN(
      n_257_76_2062));
   NOR2_X1 i_257_76_2066 (.A1(n_257_76_2062), .A2(n_257_76_1847), .ZN(
      n_257_76_2063));
   NAND2_X1 i_257_76_2067 (.A1(n_257_67), .A2(n_257_76_2063), .ZN(n_257_76_2064));
   NAND2_X1 i_257_76_2068 (.A1(n_257_76_1841), .A2(n_257_449), .ZN(n_257_76_2065));
   NAND2_X1 i_257_76_2069 (.A1(n_257_1076), .A2(n_257_76_1817), .ZN(
      n_257_76_2066));
   INV_X1 i_257_76_2070 (.A(n_257_76_2066), .ZN(n_257_76_2067));
   NAND2_X1 i_257_76_2071 (.A1(n_257_76_1831), .A2(n_257_76_2067), .ZN(
      n_257_76_2068));
   INV_X1 i_257_76_2072 (.A(n_257_76_2068), .ZN(n_257_76_2069));
   NAND4_X1 i_257_76_2073 (.A1(n_257_76_2069), .A2(n_257_76_1836), .A3(
      n_257_76_1837), .A4(n_257_76_1838), .ZN(n_257_76_2070));
   NOR2_X1 i_257_76_2074 (.A1(n_257_76_2065), .A2(n_257_76_2070), .ZN(
      n_257_76_2071));
   INV_X1 i_257_76_2075 (.A(n_257_76_1824), .ZN(n_257_76_2072));
   INV_X1 i_257_76_2076 (.A(n_257_76_1828), .ZN(n_257_76_2073));
   NAND3_X1 i_257_76_2077 (.A1(n_257_76_2071), .A2(n_257_76_2072), .A3(
      n_257_76_2073), .ZN(n_257_76_2074));
   INV_X1 i_257_76_2078 (.A(n_257_76_1830), .ZN(n_257_76_2075));
   NOR2_X1 i_257_76_2079 (.A1(n_257_76_2074), .A2(n_257_76_2075), .ZN(
      n_257_76_2076));
   NAND2_X1 i_257_76_2080 (.A1(n_257_76_1801), .A2(n_257_76_2076), .ZN(
      n_257_76_2077));
   NOR2_X1 i_257_76_2081 (.A1(n_257_76_2077), .A2(n_257_76_1847), .ZN(
      n_257_76_2078));
   NAND2_X1 i_257_76_2082 (.A1(n_257_27), .A2(n_257_76_2078), .ZN(n_257_76_2079));
   NAND2_X1 i_257_76_2083 (.A1(n_257_429), .A2(n_257_76_1817), .ZN(n_257_76_2080));
   INV_X1 i_257_76_2084 (.A(n_257_76_2080), .ZN(n_257_76_2081));
   NAND2_X1 i_257_76_2085 (.A1(n_257_76_1886), .A2(n_257_76_2081), .ZN(
      n_257_76_2082));
   NOR2_X1 i_257_76_2086 (.A1(n_257_76_1944), .A2(n_257_76_2082), .ZN(
      n_257_76_2083));
   NAND4_X1 i_257_76_2087 (.A1(n_257_76_2083), .A2(n_257_76_1837), .A3(
      n_257_76_1838), .A4(n_257_76_1884), .ZN(n_257_76_2084));
   NOR2_X1 i_257_76_2088 (.A1(n_257_76_1943), .A2(n_257_76_2084), .ZN(
      n_257_76_2085));
   NAND4_X1 i_257_76_2089 (.A1(n_257_76_1940), .A2(n_257_76_1942), .A3(
      n_257_76_1900), .A4(n_257_76_2085), .ZN(n_257_76_2086));
   NAND2_X1 i_257_76_2090 (.A1(n_257_76_1830), .A2(n_257_155), .ZN(n_257_76_2087));
   NOR2_X1 i_257_76_2091 (.A1(n_257_76_2086), .A2(n_257_76_2087), .ZN(
      n_257_76_2088));
   NAND3_X1 i_257_76_2092 (.A1(n_257_76_2088), .A2(n_257_76_1813), .A3(
      n_257_76_1801), .ZN(n_257_76_2089));
   INV_X1 i_257_76_2093 (.A(n_257_76_2089), .ZN(n_257_76_2090));
   NAND2_X1 i_257_76_2094 (.A1(n_257_184), .A2(n_257_76_2090), .ZN(n_257_76_2091));
   NAND3_X1 i_257_76_2095 (.A1(n_257_76_2064), .A2(n_257_76_2079), .A3(
      n_257_76_2091), .ZN(n_257_76_2092));
   INV_X1 i_257_76_2096 (.A(n_257_76_2092), .ZN(n_257_76_2093));
   NAND2_X1 i_257_76_2097 (.A1(n_257_1068), .A2(n_257_76_1817), .ZN(
      n_257_76_2094));
   INV_X1 i_257_76_2098 (.A(n_257_76_2094), .ZN(n_257_76_2095));
   NAND2_X1 i_257_76_2099 (.A1(n_257_438), .A2(n_257_76_2095), .ZN(n_257_76_2096));
   INV_X1 i_257_76_2100 (.A(n_257_76_2096), .ZN(n_257_76_2097));
   NAND3_X1 i_257_76_2101 (.A1(n_257_76_2097), .A2(n_257_76_1836), .A3(
      n_257_76_1838), .ZN(n_257_76_2098));
   INV_X1 i_257_76_2102 (.A(n_257_76_2098), .ZN(n_257_76_2099));
   NAND2_X1 i_257_76_2103 (.A1(n_257_76_1802), .A2(n_257_76_2099), .ZN(
      n_257_76_2100));
   INV_X1 i_257_76_2104 (.A(n_257_76_2100), .ZN(n_257_76_2101));
   NAND2_X1 i_257_76_2105 (.A1(n_257_76_1801), .A2(n_257_76_2101), .ZN(
      n_257_76_2102));
   INV_X1 i_257_76_2106 (.A(n_257_76_2102), .ZN(n_257_76_2103));
   NAND2_X1 i_257_76_2107 (.A1(n_257_76_2103), .A2(n_257_76_1813), .ZN(
      n_257_76_2104));
   INV_X1 i_257_76_2108 (.A(n_257_76_2104), .ZN(n_257_76_2105));
   NAND2_X1 i_257_76_2109 (.A1(n_257_19), .A2(n_257_76_2105), .ZN(n_257_76_2106));
   INV_X1 i_257_76_2110 (.A(n_257_76_1881), .ZN(n_257_76_2107));
   NAND3_X1 i_257_76_2111 (.A1(n_257_76_1803), .A2(n_257_442), .A3(n_257_894), 
      .ZN(n_257_76_2108));
   INV_X1 i_257_76_2112 (.A(n_257_76_2108), .ZN(n_257_76_2109));
   NAND3_X1 i_257_76_2113 (.A1(n_257_420), .A2(n_257_76_1887), .A3(n_257_76_2109), 
      .ZN(n_257_76_2110));
   NOR2_X1 i_257_76_2114 (.A1(n_257_76_2107), .A2(n_257_76_2110), .ZN(
      n_257_76_2111));
   NAND2_X1 i_257_76_2115 (.A1(n_257_76_1831), .A2(n_257_76_1886), .ZN(
      n_257_76_2112));
   INV_X1 i_257_76_2116 (.A(n_257_76_2112), .ZN(n_257_76_2113));
   NAND4_X1 i_257_76_2117 (.A1(n_257_76_2111), .A2(n_257_76_2113), .A3(
      n_257_76_1884), .A4(n_257_76_1885), .ZN(n_257_76_2114));
   NAND2_X1 i_257_76_2118 (.A1(n_257_313), .A2(n_257_422), .ZN(n_257_76_2115));
   NAND4_X1 i_257_76_2119 (.A1(n_257_76_1836), .A2(n_257_76_2115), .A3(
      n_257_76_1837), .A4(n_257_76_1838), .ZN(n_257_76_2116));
   NOR2_X1 i_257_76_2120 (.A1(n_257_76_2114), .A2(n_257_76_2116), .ZN(
      n_257_76_2117));
   NAND4_X1 i_257_76_2121 (.A1(n_257_76_1840), .A2(n_257_76_1841), .A3(
      n_257_76_1874), .A4(n_257_76_1875), .ZN(n_257_76_2118));
   INV_X1 i_257_76_2122 (.A(n_257_76_2118), .ZN(n_257_76_2119));
   NAND3_X1 i_257_76_2123 (.A1(n_257_76_2117), .A2(n_257_76_2073), .A3(
      n_257_76_2119), .ZN(n_257_76_2120));
   NAND2_X1 i_257_76_2124 (.A1(n_257_275), .A2(n_257_423), .ZN(n_257_76_2121));
   NAND3_X1 i_257_76_2125 (.A1(n_257_76_1901), .A2(n_257_76_1823), .A3(
      n_257_76_2121), .ZN(n_257_76_2122));
   INV_X1 i_257_76_2126 (.A(n_257_76_2122), .ZN(n_257_76_2123));
   NAND2_X1 i_257_76_2127 (.A1(n_257_76_1895), .A2(n_257_76_1802), .ZN(
      n_257_76_2124));
   INV_X1 i_257_76_2128 (.A(n_257_76_2124), .ZN(n_257_76_2125));
   NAND3_X1 i_257_76_2129 (.A1(n_257_76_2123), .A2(n_257_76_2125), .A3(
      n_257_76_1900), .ZN(n_257_76_2126));
   NOR2_X1 i_257_76_2130 (.A1(n_257_76_2120), .A2(n_257_76_2126), .ZN(
      n_257_76_2127));
   NAND2_X1 i_257_76_2131 (.A1(n_257_352), .A2(n_257_421), .ZN(n_257_76_2128));
   NAND2_X1 i_257_76_2132 (.A1(n_257_76_1830), .A2(n_257_76_2128), .ZN(
      n_257_76_2129));
   INV_X1 i_257_76_2133 (.A(n_257_76_2129), .ZN(n_257_76_2130));
   NAND4_X1 i_257_76_2134 (.A1(n_257_76_2127), .A2(n_257_76_1801), .A3(
      n_257_76_2130), .A4(n_257_76_1908), .ZN(n_257_76_2131));
   NAND2_X1 i_257_76_2135 (.A1(n_257_76_1813), .A2(n_257_76_1911), .ZN(
      n_257_76_2132));
   NOR2_X1 i_257_76_2136 (.A1(n_257_76_2131), .A2(n_257_76_2132), .ZN(
      n_257_76_2133));
   NAND2_X1 i_257_76_2137 (.A1(n_257_382), .A2(n_257_76_2133), .ZN(n_257_76_2134));
   NAND4_X1 i_257_76_2138 (.A1(n_257_76_1827), .A2(n_257_116), .A3(n_257_76_1840), 
      .A4(n_257_76_1841), .ZN(n_257_76_2135));
   NAND2_X1 i_257_76_2139 (.A1(n_257_430), .A2(n_257_76_1817), .ZN(n_257_76_2136));
   INV_X1 i_257_76_2140 (.A(n_257_76_2136), .ZN(n_257_76_2137));
   NAND2_X1 i_257_76_2141 (.A1(n_257_76_1886), .A2(n_257_76_2137), .ZN(
      n_257_76_2138));
   NOR2_X1 i_257_76_2142 (.A1(n_257_76_1944), .A2(n_257_76_2138), .ZN(
      n_257_76_2139));
   NAND4_X1 i_257_76_2143 (.A1(n_257_76_2019), .A2(n_257_76_2057), .A3(
      n_257_76_1875), .A4(n_257_76_2139), .ZN(n_257_76_2140));
   NOR2_X1 i_257_76_2144 (.A1(n_257_76_2135), .A2(n_257_76_2140), .ZN(
      n_257_76_2141));
   NAND4_X1 i_257_76_2145 (.A1(n_257_76_1830), .A2(n_257_76_2141), .A3(
      n_257_76_2009), .A4(n_257_76_1900), .ZN(n_257_76_2142));
   INV_X1 i_257_76_2146 (.A(n_257_76_2142), .ZN(n_257_76_2143));
   NAND3_X1 i_257_76_2147 (.A1(n_257_76_2143), .A2(n_257_76_1813), .A3(
      n_257_76_1801), .ZN(n_257_76_2144));
   INV_X1 i_257_76_2148 (.A(n_257_76_2144), .ZN(n_257_76_2145));
   NAND2_X1 i_257_76_2149 (.A1(n_257_145), .A2(n_257_76_2145), .ZN(n_257_76_2146));
   NAND3_X1 i_257_76_2150 (.A1(n_257_76_2106), .A2(n_257_76_2134), .A3(
      n_257_76_2146), .ZN(n_257_76_2147));
   INV_X1 i_257_76_2151 (.A(n_257_76_2147), .ZN(n_257_76_2148));
   INV_X1 i_257_76_2152 (.A(n_257_768), .ZN(n_257_76_2149));
   NOR2_X1 i_257_76_2153 (.A1(n_257_76_1804), .A2(n_257_76_2149), .ZN(
      n_257_76_2150));
   NAND3_X1 i_257_76_2154 (.A1(n_257_76_1837), .A2(n_257_76_1838), .A3(
      n_257_76_2150), .ZN(n_257_76_2151));
   INV_X1 i_257_76_2155 (.A(n_257_76_2151), .ZN(n_257_76_2152));
   NAND2_X1 i_257_76_2156 (.A1(n_257_447), .A2(n_257_76_1836), .ZN(n_257_76_2153));
   INV_X1 i_257_76_2157 (.A(n_257_76_2153), .ZN(n_257_76_2154));
   NAND4_X1 i_257_76_2158 (.A1(n_257_76_2152), .A2(n_257_76_2154), .A3(
      n_257_76_1826), .A4(n_257_76_1827), .ZN(n_257_76_2155));
   NOR2_X1 i_257_76_2159 (.A1(n_257_76_2155), .A2(n_257_76_2033), .ZN(
      n_257_76_2156));
   NAND2_X1 i_257_76_2160 (.A1(n_257_76_1801), .A2(n_257_76_2156), .ZN(
      n_257_76_2157));
   INV_X1 i_257_76_2161 (.A(n_257_76_2157), .ZN(n_257_76_2158));
   NAND2_X1 i_257_76_2162 (.A1(n_257_76_2158), .A2(n_257_76_1813), .ZN(
      n_257_76_2159));
   INV_X1 i_257_76_2163 (.A(n_257_76_2159), .ZN(n_257_76_2160));
   NAND3_X1 i_257_76_2164 (.A1(n_257_76_1875), .A2(n_257_76_1836), .A3(
      n_257_76_1837), .ZN(n_257_76_2161));
   NAND2_X1 i_257_76_2165 (.A1(n_257_431), .A2(n_257_76_1817), .ZN(n_257_76_2162));
   INV_X1 i_257_76_2166 (.A(n_257_76_2162), .ZN(n_257_76_2163));
   NAND2_X1 i_257_76_2167 (.A1(n_257_76_1886), .A2(n_257_76_2163), .ZN(
      n_257_76_2164));
   INV_X1 i_257_76_2168 (.A(n_257_76_2164), .ZN(n_257_76_2165));
   NAND4_X1 i_257_76_2169 (.A1(n_257_76_1838), .A2(n_257_76_1884), .A3(
      n_257_76_1831), .A4(n_257_76_2165), .ZN(n_257_76_2166));
   NOR2_X1 i_257_76_2170 (.A1(n_257_76_2161), .A2(n_257_76_2166), .ZN(
      n_257_76_2167));
   NAND2_X1 i_257_76_2171 (.A1(n_257_76_1825), .A2(n_257_76_1826), .ZN(
      n_257_76_2168));
   INV_X1 i_257_76_2172 (.A(n_257_76_2168), .ZN(n_257_76_2169));
   NAND3_X1 i_257_76_2173 (.A1(n_257_76_2167), .A2(n_257_76_1905), .A3(
      n_257_76_2169), .ZN(n_257_76_2170));
   NAND4_X1 i_257_76_2174 (.A1(n_257_78), .A2(n_257_76_1802), .A3(n_257_76_1901), 
      .A4(n_257_76_1823), .ZN(n_257_76_2171));
   NOR2_X1 i_257_76_2175 (.A1(n_257_76_2170), .A2(n_257_76_2171), .ZN(
      n_257_76_2172));
   NAND3_X1 i_257_76_2176 (.A1(n_257_76_2172), .A2(n_257_76_1801), .A3(
      n_257_76_1830), .ZN(n_257_76_2173));
   NOR2_X1 i_257_76_2177 (.A1(n_257_76_2173), .A2(n_257_76_1847), .ZN(
      n_257_76_2174));
   AOI22_X1 i_257_76_2178 (.A1(n_257_23), .A2(n_257_76_2160), .B1(n_257_107), 
      .B2(n_257_76_2174), .ZN(n_257_76_2175));
   NAND3_X1 i_257_76_2179 (.A1(n_257_76_2093), .A2(n_257_76_2148), .A3(
      n_257_76_2175), .ZN(n_257_76_2176));
   NAND3_X1 i_257_76_2180 (.A1(n_257_76_1826), .A2(n_257_76_1827), .A3(
      n_257_76_1841), .ZN(n_257_76_2177));
   NAND3_X1 i_257_76_2181 (.A1(n_257_448), .A2(n_257_76_1838), .A3(
      n_257_76_18054), .ZN(n_257_76_2178));
   INV_X1 i_257_76_2182 (.A(n_257_76_2178), .ZN(n_257_76_2179));
   NAND2_X1 i_257_76_2183 (.A1(n_257_76_2179), .A2(n_257_76_2019), .ZN(
      n_257_76_2180));
   NOR2_X1 i_257_76_2184 (.A1(n_257_76_2177), .A2(n_257_76_2180), .ZN(
      n_257_76_2181));
   INV_X1 i_257_76_2185 (.A(n_257_76_1932), .ZN(n_257_76_2182));
   NAND3_X1 i_257_76_2186 (.A1(n_257_76_2181), .A2(n_257_76_2182), .A3(n_257_672), 
      .ZN(n_257_76_2183));
   INV_X1 i_257_76_2187 (.A(n_257_76_2183), .ZN(n_257_76_2184));
   NAND2_X1 i_257_76_2188 (.A1(n_257_76_1801), .A2(n_257_76_2184), .ZN(
      n_257_76_2185));
   NOR2_X1 i_257_76_2189 (.A1(n_257_76_1847), .A2(n_257_76_2185), .ZN(
      n_257_76_2186));
   NAND2_X1 i_257_76_2190 (.A1(n_257_26), .A2(n_257_76_2186), .ZN(n_257_76_2187));
   NAND2_X1 i_257_76_2191 (.A1(n_257_425), .A2(n_257_76_1817), .ZN(n_257_76_2188));
   INV_X1 i_257_76_2192 (.A(n_257_76_2188), .ZN(n_257_76_2189));
   NAND3_X1 i_257_76_2193 (.A1(n_257_76_1886), .A2(n_257_76_1887), .A3(
      n_257_76_2189), .ZN(n_257_76_2190));
   INV_X1 i_257_76_2194 (.A(n_257_76_2190), .ZN(n_257_76_2191));
   NAND3_X1 i_257_76_2195 (.A1(n_257_76_1885), .A2(n_257_76_2191), .A3(
      n_257_76_1831), .ZN(n_257_76_2192));
   INV_X1 i_257_76_2196 (.A(n_257_76_2192), .ZN(n_257_76_2193));
   NAND3_X1 i_257_76_2197 (.A1(n_257_76_2019), .A2(n_257_76_2193), .A3(
      n_257_76_2057), .ZN(n_257_76_2194));
   NAND3_X1 i_257_76_2198 (.A1(n_257_76_1841), .A2(n_257_76_1874), .A3(
      n_257_76_1875), .ZN(n_257_76_2195));
   NOR2_X1 i_257_76_2199 (.A1(n_257_76_2194), .A2(n_257_76_2195), .ZN(
      n_257_76_2196));
   NAND3_X1 i_257_76_2200 (.A1(n_257_76_1940), .A2(n_257_76_1942), .A3(
      n_257_76_2196), .ZN(n_257_76_2197));
   INV_X1 i_257_76_2201 (.A(n_257_76_2197), .ZN(n_257_76_2198));
   NAND2_X1 i_257_76_2202 (.A1(n_257_76_1830), .A2(n_257_76_1900), .ZN(
      n_257_76_2199));
   INV_X1 i_257_76_2203 (.A(n_257_76_2199), .ZN(n_257_76_2200));
   NAND4_X1 i_257_76_2204 (.A1(n_257_76_2198), .A2(n_257_76_2200), .A3(n_257_235), 
      .A4(n_257_76_1908), .ZN(n_257_76_2201));
   NAND2_X1 i_257_76_2205 (.A1(n_257_76_1813), .A2(n_257_76_1801), .ZN(
      n_257_76_2202));
   NOR2_X1 i_257_76_2206 (.A1(n_257_76_2201), .A2(n_257_76_2202), .ZN(
      n_257_76_2203));
   NAND2_X1 i_257_76_2207 (.A1(n_257_264), .A2(n_257_76_2203), .ZN(n_257_76_2204));
   NAND2_X1 i_257_76_2208 (.A1(n_257_76_1900), .A2(n_257_352), .ZN(n_257_76_2205));
   INV_X1 i_257_76_2209 (.A(n_257_76_2205), .ZN(n_257_76_2206));
   NAND4_X1 i_257_76_2210 (.A1(n_257_76_1823), .A2(n_257_76_2121), .A3(
      n_257_76_1825), .A4(n_257_76_1826), .ZN(n_257_76_2207));
   NOR2_X1 i_257_76_2211 (.A1(n_257_76_1939), .A2(n_257_76_2207), .ZN(
      n_257_76_2208));
   NAND2_X1 i_257_76_2212 (.A1(n_257_421), .A2(n_257_76_1817), .ZN(n_257_76_2209));
   NOR2_X1 i_257_76_2213 (.A1(n_257_76_1981), .A2(n_257_76_2209), .ZN(
      n_257_76_2210));
   NAND4_X1 i_257_76_2214 (.A1(n_257_76_1881), .A2(n_257_76_1831), .A3(
      n_257_76_2210), .A4(n_257_76_1886), .ZN(n_257_76_2211));
   NAND2_X1 i_257_76_2215 (.A1(n_257_76_1884), .A2(n_257_76_1885), .ZN(
      n_257_76_2212));
   NOR2_X1 i_257_76_2216 (.A1(n_257_76_2211), .A2(n_257_76_2212), .ZN(
      n_257_76_2213));
   NAND2_X1 i_257_76_2217 (.A1(n_257_76_1875), .A2(n_257_76_1836), .ZN(
      n_257_76_2214));
   INV_X1 i_257_76_2218 (.A(n_257_76_2214), .ZN(n_257_76_2215));
   NAND3_X1 i_257_76_2219 (.A1(n_257_76_2115), .A2(n_257_76_1837), .A3(
      n_257_76_1838), .ZN(n_257_76_2216));
   INV_X1 i_257_76_2220 (.A(n_257_76_2216), .ZN(n_257_76_2217));
   NAND3_X1 i_257_76_2221 (.A1(n_257_76_2213), .A2(n_257_76_2215), .A3(
      n_257_76_2217), .ZN(n_257_76_2218));
   NAND4_X1 i_257_76_2222 (.A1(n_257_76_1827), .A2(n_257_76_1840), .A3(
      n_257_76_1841), .A4(n_257_76_1874), .ZN(n_257_76_2219));
   NOR2_X1 i_257_76_2223 (.A1(n_257_76_2218), .A2(n_257_76_2219), .ZN(
      n_257_76_2220));
   NAND4_X1 i_257_76_2224 (.A1(n_257_76_2206), .A2(n_257_76_2208), .A3(
      n_257_76_1830), .A4(n_257_76_2220), .ZN(n_257_76_2221));
   INV_X1 i_257_76_2225 (.A(n_257_76_2221), .ZN(n_257_76_2222));
   NAND2_X1 i_257_76_2226 (.A1(n_257_76_1801), .A2(n_257_76_1908), .ZN(
      n_257_76_2223));
   INV_X1 i_257_76_2227 (.A(n_257_76_2223), .ZN(n_257_76_2224));
   NAND4_X1 i_257_76_2228 (.A1(n_257_76_2222), .A2(n_257_76_2224), .A3(
      n_257_76_1813), .A4(n_257_76_1911), .ZN(n_257_76_2225));
   INV_X1 i_257_76_2229 (.A(n_257_76_2225), .ZN(n_257_76_2226));
   NAND2_X1 i_257_76_2230 (.A1(n_257_381), .A2(n_257_76_2226), .ZN(n_257_76_2227));
   NAND3_X1 i_257_76_2231 (.A1(n_257_76_2187), .A2(n_257_76_2204), .A3(
      n_257_76_2227), .ZN(n_257_76_2228));
   INV_X1 i_257_76_2232 (.A(n_257_76_2228), .ZN(n_257_76_2229));
   NAND2_X1 i_257_76_2233 (.A1(n_257_76_1831), .A2(n_257_195), .ZN(n_257_76_2230));
   INV_X1 i_257_76_2234 (.A(n_257_76_2230), .ZN(n_257_76_2231));
   INV_X1 i_257_76_2235 (.A(n_257_568), .ZN(n_257_76_2232));
   NAND3_X1 i_257_76_2236 (.A1(n_257_76_1803), .A2(n_257_76_2232), .A3(n_257_442), 
      .ZN(n_257_76_2233));
   OAI21_X1 i_257_76_2237 (.A(n_257_76_2233), .B1(n_257_428), .B2(n_257_76_1804), 
      .ZN(n_257_76_2234));
   NAND3_X1 i_257_76_2238 (.A1(n_257_427), .A2(n_257_76_1886), .A3(n_257_76_2234), 
      .ZN(n_257_76_2235));
   INV_X1 i_257_76_2239 (.A(n_257_76_2235), .ZN(n_257_76_2236));
   NAND4_X1 i_257_76_2240 (.A1(n_257_76_1875), .A2(n_257_76_1884), .A3(
      n_257_76_2231), .A4(n_257_76_2236), .ZN(n_257_76_2237));
   INV_X1 i_257_76_2241 (.A(n_257_76_2237), .ZN(n_257_76_2238));
   NAND3_X1 i_257_76_2242 (.A1(n_257_76_2238), .A2(n_257_76_1895), .A3(
      n_257_76_1802), .ZN(n_257_76_2239));
   INV_X1 i_257_76_2243 (.A(n_257_76_2239), .ZN(n_257_76_2240));
   NAND4_X1 i_257_76_2244 (.A1(n_257_76_1901), .A2(n_257_76_1823), .A3(
      n_257_76_1825), .A4(n_257_76_1826), .ZN(n_257_76_2241));
   INV_X1 i_257_76_2245 (.A(n_257_76_2241), .ZN(n_257_76_2242));
   INV_X1 i_257_76_2246 (.A(n_257_76_1893), .ZN(n_257_76_2243));
   NAND4_X1 i_257_76_2247 (.A1(n_257_76_2243), .A2(n_257_76_1827), .A3(
      n_257_76_1840), .A4(n_257_76_1841), .ZN(n_257_76_2244));
   INV_X1 i_257_76_2248 (.A(n_257_76_2244), .ZN(n_257_76_2245));
   NAND4_X1 i_257_76_2249 (.A1(n_257_76_2240), .A2(n_257_76_2242), .A3(
      n_257_76_2245), .A4(n_257_76_1900), .ZN(n_257_76_2246));
   INV_X1 i_257_76_2250 (.A(n_257_76_2246), .ZN(n_257_76_2247));
   NAND3_X1 i_257_76_2251 (.A1(n_257_76_2247), .A2(n_257_76_1956), .A3(
      n_257_76_1801), .ZN(n_257_76_2248));
   NOR2_X1 i_257_76_2252 (.A1(n_257_76_2248), .A2(n_257_76_1847), .ZN(
      n_257_76_2249));
   NAND2_X1 i_257_76_2253 (.A1(n_257_224), .A2(n_257_76_2249), .ZN(n_257_76_2250));
   NAND2_X1 i_257_76_2254 (.A1(n_257_76_1838), .A2(n_257_76_18054), .ZN(
      n_257_76_2251));
   INV_X1 i_257_76_2255 (.A(n_257_76_2251), .ZN(n_257_76_2252));
   NAND2_X1 i_257_76_2256 (.A1(n_257_76_1884), .A2(n_257_455), .ZN(n_257_76_2253));
   INV_X1 i_257_76_2257 (.A(n_257_76_2253), .ZN(n_257_76_2254));
   NAND3_X1 i_257_76_2258 (.A1(n_257_76_2019), .A2(n_257_76_2252), .A3(
      n_257_76_2254), .ZN(n_257_76_2255));
   NAND3_X1 i_257_76_2259 (.A1(n_257_76_1840), .A2(n_257_76_1841), .A3(n_257_451), 
      .ZN(n_257_76_2256));
   NOR2_X1 i_257_76_2260 (.A1(n_257_76_2255), .A2(n_257_76_2256), .ZN(
      n_257_76_2257));
   NAND3_X1 i_257_76_2261 (.A1(n_257_76_1829), .A2(n_257_76_1830), .A3(
      n_257_76_2257), .ZN(n_257_76_2258));
   INV_X1 i_257_76_2262 (.A(n_257_76_2258), .ZN(n_257_76_2259));
   NAND2_X1 i_257_76_2263 (.A1(n_257_76_2259), .A2(n_257_76_1801), .ZN(
      n_257_76_2260));
   NOR2_X1 i_257_76_2264 (.A1(n_257_76_2260), .A2(n_257_76_1847), .ZN(
      n_257_76_2261));
   NAND2_X1 i_257_76_2265 (.A1(n_257_434), .A2(n_257_76_2261), .ZN(n_257_76_2262));
   NOR2_X1 i_257_76_2266 (.A1(n_257_76_1988), .A2(n_257_76_1904), .ZN(
      n_257_76_2263));
   NAND3_X1 i_257_76_2267 (.A1(n_257_504), .A2(n_257_76_2234), .A3(n_257_424), 
      .ZN(n_257_76_2264));
   NOR2_X1 i_257_76_2268 (.A1(n_257_76_2112), .A2(n_257_76_2264), .ZN(
      n_257_76_2265));
   INV_X1 i_257_76_2269 (.A(n_257_76_2212), .ZN(n_257_76_2266));
   NAND3_X1 i_257_76_2270 (.A1(n_257_76_2265), .A2(n_257_76_2266), .A3(
      n_257_76_1838), .ZN(n_257_76_2267));
   NAND4_X1 i_257_76_2271 (.A1(n_257_76_1874), .A2(n_257_76_1875), .A3(
      n_257_76_1836), .A4(n_257_76_1837), .ZN(n_257_76_2268));
   NOR2_X1 i_257_76_2272 (.A1(n_257_76_2267), .A2(n_257_76_2268), .ZN(
      n_257_76_2269));
   NAND4_X1 i_257_76_2273 (.A1(n_257_76_1940), .A2(n_257_76_2263), .A3(
      n_257_76_1900), .A4(n_257_76_2269), .ZN(n_257_76_2270));
   NOR2_X1 i_257_76_2274 (.A1(n_257_76_2270), .A2(n_257_76_1955), .ZN(
      n_257_76_2271));
   NAND2_X1 i_257_76_2275 (.A1(n_257_76_1911), .A2(n_257_76_1801), .ZN(
      n_257_76_2272));
   INV_X1 i_257_76_2276 (.A(n_257_76_2272), .ZN(n_257_76_2273));
   NAND3_X1 i_257_76_2277 (.A1(n_257_76_2271), .A2(n_257_76_2273), .A3(
      n_257_76_1813), .ZN(n_257_76_2274));
   INV_X1 i_257_76_2278 (.A(n_257_76_2274), .ZN(n_257_76_2275));
   NAND2_X1 i_257_76_2279 (.A1(n_257_265), .A2(n_257_76_2275), .ZN(n_257_76_2276));
   NAND3_X1 i_257_76_2280 (.A1(n_257_76_2250), .A2(n_257_76_2262), .A3(
      n_257_76_2276), .ZN(n_257_76_2277));
   INV_X1 i_257_76_2281 (.A(n_257_76_2277), .ZN(n_257_76_2278));
   NAND3_X1 i_257_76_2282 (.A1(n_257_76_1886), .A2(n_257_76_2234), .A3(n_257_422), 
      .ZN(n_257_76_2279));
   NOR2_X1 i_257_76_2283 (.A1(n_257_76_2279), .A2(n_257_76_1944), .ZN(
      n_257_76_2280));
   NAND2_X1 i_257_76_2284 (.A1(n_257_313), .A2(n_257_76_1881), .ZN(n_257_76_2281));
   INV_X1 i_257_76_2285 (.A(n_257_76_2281), .ZN(n_257_76_2282));
   NAND4_X1 i_257_76_2286 (.A1(n_257_76_2280), .A2(n_257_76_1875), .A3(
      n_257_76_2282), .A4(n_257_76_1884), .ZN(n_257_76_2283));
   INV_X1 i_257_76_2287 (.A(n_257_76_1895), .ZN(n_257_76_2284));
   NOR2_X1 i_257_76_2288 (.A1(n_257_76_2283), .A2(n_257_76_2284), .ZN(
      n_257_76_2285));
   NAND3_X1 i_257_76_2289 (.A1(n_257_76_2285), .A2(n_257_76_1900), .A3(
      n_257_76_1903), .ZN(n_257_76_2286));
   INV_X1 i_257_76_2290 (.A(n_257_76_2286), .ZN(n_257_76_2287));
   NAND2_X1 i_257_76_2291 (.A1(n_257_76_1841), .A2(n_257_76_1874), .ZN(
      n_257_76_2288));
   NAND4_X1 i_257_76_2292 (.A1(n_257_76_1836), .A2(n_257_76_1837), .A3(
      n_257_76_1838), .A4(n_257_76_1885), .ZN(n_257_76_2289));
   NOR2_X1 i_257_76_2293 (.A1(n_257_76_2288), .A2(n_257_76_2289), .ZN(
      n_257_76_2290));
   NAND3_X1 i_257_76_2294 (.A1(n_257_76_1823), .A2(n_257_76_2121), .A3(
      n_257_76_1825), .ZN(n_257_76_2291));
   INV_X1 i_257_76_2295 (.A(n_257_76_2291), .ZN(n_257_76_2292));
   INV_X1 i_257_76_2296 (.A(n_257_76_1941), .ZN(n_257_76_2293));
   NAND3_X1 i_257_76_2297 (.A1(n_257_76_2290), .A2(n_257_76_2292), .A3(
      n_257_76_2293), .ZN(n_257_76_2294));
   INV_X1 i_257_76_2298 (.A(n_257_76_2294), .ZN(n_257_76_2295));
   NAND4_X1 i_257_76_2299 (.A1(n_257_76_2287), .A2(n_257_76_1908), .A3(
      n_257_76_2295), .A4(n_257_76_1830), .ZN(n_257_76_2296));
   INV_X1 i_257_76_2300 (.A(n_257_76_2296), .ZN(n_257_76_2297));
   NAND3_X1 i_257_76_2301 (.A1(n_257_76_2297), .A2(n_257_76_2273), .A3(
      n_257_76_1813), .ZN(n_257_76_2298));
   INV_X1 i_257_76_2302 (.A(n_257_76_2298), .ZN(n_257_76_2299));
   NAND2_X1 i_257_76_2303 (.A1(n_257_342), .A2(n_257_76_2299), .ZN(n_257_76_2300));
   NOR2_X1 i_257_76_2304 (.A1(n_257_76_1979), .A2(n_257_76_1955), .ZN(
      n_257_76_2301));
   NAND2_X1 i_257_76_2305 (.A1(n_257_76_2121), .A2(n_257_76_1825), .ZN(
      n_257_76_2302));
   INV_X1 i_257_76_2306 (.A(n_257_76_2302), .ZN(n_257_76_2303));
   NAND2_X1 i_257_76_2307 (.A1(n_257_76_1826), .A2(n_257_76_1827), .ZN(
      n_257_76_2304));
   INV_X1 i_257_76_2308 (.A(n_257_76_2304), .ZN(n_257_76_2305));
   NAND2_X1 i_257_76_2309 (.A1(n_257_76_2303), .A2(n_257_76_2305), .ZN(
      n_257_76_2306));
   NAND2_X1 i_257_76_2310 (.A1(n_257_76_1901), .A2(n_257_76_1823), .ZN(
      n_257_76_2307));
   NOR2_X1 i_257_76_2311 (.A1(n_257_76_2306), .A2(n_257_76_2307), .ZN(
      n_257_76_2308));
   INV_X1 i_257_76_2312 (.A(n_257_76_1842), .ZN(n_257_76_2309));
   INV_X1 i_257_76_2313 (.A(n_257_76_1874), .ZN(n_257_76_2310));
   NOR2_X1 i_257_76_2314 (.A1(n_257_76_2214), .A2(n_257_76_2310), .ZN(
      n_257_76_2311));
   NAND2_X1 i_257_76_2315 (.A1(n_257_76_2309), .A2(n_257_76_2311), .ZN(
      n_257_76_2312));
   NAND2_X1 i_257_76_2316 (.A1(n_257_76_2115), .A2(n_257_76_1837), .ZN(
      n_257_76_2313));
   NOR2_X1 i_257_76_2317 (.A1(n_257_76_2313), .A2(n_257_76_2056), .ZN(
      n_257_76_2314));
   NAND2_X1 i_257_76_2318 (.A1(n_257_420), .A2(n_257_894), .ZN(n_257_76_2315));
   NAND2_X1 i_257_76_2319 (.A1(n_257_76_1831), .A2(n_257_76_2315), .ZN(
      n_257_76_2316));
   INV_X1 i_257_76_2320 (.A(n_257_76_2316), .ZN(n_257_76_2317));
   NAND2_X1 i_257_76_2321 (.A1(n_257_76_1817), .A2(n_257_484), .ZN(n_257_76_2318));
   INV_X1 i_257_76_2322 (.A(n_257_76_2318), .ZN(n_257_76_2319));
   NAND2_X1 i_257_76_2323 (.A1(n_257_76_2319), .A2(n_257_391), .ZN(n_257_76_2320));
   INV_X1 i_257_76_2324 (.A(n_257_76_2320), .ZN(n_257_76_2321));
   NAND2_X1 i_257_76_2325 (.A1(n_257_76_2321), .A2(n_257_76_1887), .ZN(
      n_257_76_2322));
   INV_X1 i_257_76_2326 (.A(n_257_76_1886), .ZN(n_257_76_2323));
   NOR2_X1 i_257_76_2327 (.A1(n_257_76_2322), .A2(n_257_76_2323), .ZN(
      n_257_76_2324));
   NAND2_X1 i_257_76_2328 (.A1(n_257_76_2317), .A2(n_257_76_2324), .ZN(
      n_257_76_2325));
   NAND2_X1 i_257_76_2329 (.A1(n_257_76_1885), .A2(n_257_76_1881), .ZN(
      n_257_76_2326));
   NOR2_X1 i_257_76_2330 (.A1(n_257_76_2325), .A2(n_257_76_2326), .ZN(
      n_257_76_2327));
   NAND2_X1 i_257_76_2331 (.A1(n_257_76_2314), .A2(n_257_76_2327), .ZN(
      n_257_76_2328));
   NOR2_X1 i_257_76_2332 (.A1(n_257_76_2312), .A2(n_257_76_2328), .ZN(
      n_257_76_2329));
   NAND2_X1 i_257_76_2333 (.A1(n_257_76_2308), .A2(n_257_76_2329), .ZN(
      n_257_76_2330));
   NAND2_X1 i_257_76_2334 (.A1(n_257_76_2125), .A2(n_257_76_1900), .ZN(
      n_257_76_2331));
   INV_X1 i_257_76_2335 (.A(n_257_76_2331), .ZN(n_257_76_2332));
   NAND2_X1 i_257_76_2336 (.A1(n_257_76_2332), .A2(n_257_76_2128), .ZN(
      n_257_76_2333));
   NOR2_X1 i_257_76_2337 (.A1(n_257_76_2330), .A2(n_257_76_2333), .ZN(
      n_257_76_2334));
   NAND2_X1 i_257_76_2338 (.A1(n_257_76_2301), .A2(n_257_76_2334), .ZN(
      n_257_76_2335));
   NOR2_X1 i_257_76_2339 (.A1(n_257_76_2335), .A2(n_257_76_2132), .ZN(
      n_257_76_2336));
   NAND2_X1 i_257_76_2340 (.A1(n_257_12), .A2(n_257_76_2336), .ZN(n_257_76_2337));
   INV_X1 i_257_76_2341 (.A(n_257_1030), .ZN(n_257_76_2338));
   OAI21_X1 i_257_76_2342 (.A(n_257_76_2221), .B1(n_257_76_2338), .B2(
      n_257_76_17968), .ZN(n_257_76_2339));
   INV_X1 i_257_76_2343 (.A(n_257_76_2201), .ZN(n_257_76_2340));
   NOR2_X1 i_257_76_2344 (.A1(n_257_76_2339), .A2(n_257_76_2340), .ZN(
      n_257_76_2341));
   NAND2_X1 i_257_76_2345 (.A1(n_257_155), .A2(n_257_76_17331), .ZN(
      n_257_76_2342));
   AOI22_X1 i_257_76_2346 (.A1(n_257_672), .A2(n_257_76_17958), .B1(n_257_78), 
      .B2(n_257_76_17932), .ZN(n_257_76_2343));
   NAND2_X1 i_257_76_2347 (.A1(n_257_76_2342), .A2(n_257_76_2343), .ZN(
      n_257_76_2344));
   INV_X1 i_257_76_2348 (.A(n_257_76_2344), .ZN(n_257_76_2345));
   NAND2_X1 i_257_76_2349 (.A1(n_257_116), .A2(n_257_76_17925), .ZN(
      n_257_76_2346));
   NAND2_X1 i_257_76_2350 (.A1(n_257_76_2237), .A2(n_257_76_2346), .ZN(
      n_257_76_2347));
   INV_X1 i_257_76_2351 (.A(n_257_76_2283), .ZN(n_257_76_2348));
   NOR2_X1 i_257_76_2352 (.A1(n_257_76_2347), .A2(n_257_76_2348), .ZN(
      n_257_76_2349));
   NAND2_X1 i_257_76_2353 (.A1(n_257_966), .A2(n_257_442), .ZN(n_257_76_2350));
   INV_X1 i_257_76_2354 (.A(n_257_76_2350), .ZN(n_257_76_2351));
   NAND2_X1 i_257_76_2355 (.A1(n_257_441), .A2(n_257_76_2351), .ZN(n_257_76_2352));
   NAND2_X1 i_257_76_2356 (.A1(n_257_455), .A2(n_257_442), .ZN(n_257_76_2353));
   INV_X1 i_257_76_2357 (.A(n_257_76_2353), .ZN(n_257_76_2354));
   NAND2_X1 i_257_76_2358 (.A1(n_257_451), .A2(n_257_76_2354), .ZN(n_257_76_2355));
   NAND2_X1 i_257_76_2359 (.A1(n_257_76_2352), .A2(n_257_76_2355), .ZN(
      n_257_76_2356));
   NAND2_X1 i_257_76_2360 (.A1(n_257_736), .A2(n_257_76_17935), .ZN(
      n_257_76_2357));
   NAND2_X1 i_257_76_2361 (.A1(n_257_864), .A2(n_257_76_17903), .ZN(
      n_257_76_2358));
   NAND2_X1 i_257_76_2362 (.A1(n_257_76_2357), .A2(n_257_76_2358), .ZN(
      n_257_76_2359));
   NOR2_X1 i_257_76_2363 (.A1(n_257_76_2356), .A2(n_257_76_2359), .ZN(
      n_257_76_2360));
   NAND2_X1 i_257_76_2364 (.A1(n_257_76_2349), .A2(n_257_76_2360), .ZN(
      n_257_76_2361));
   NAND2_X1 i_257_76_2365 (.A1(n_257_38), .A2(n_257_76_17918), .ZN(n_257_76_2362));
   NAND3_X1 i_257_76_2366 (.A1(n_257_439), .A2(n_257_902), .A3(n_257_442), 
      .ZN(n_257_76_2363));
   NAND2_X1 i_257_76_2367 (.A1(n_257_76_2362), .A2(n_257_76_2363), .ZN(
      n_257_76_2364));
   NAND2_X1 i_257_76_2368 (.A1(n_257_442), .A2(n_257_934), .ZN(n_257_76_2365));
   INV_X1 i_257_76_2369 (.A(n_257_76_2365), .ZN(n_257_76_2366));
   NAND2_X1 i_257_76_2370 (.A1(n_257_440), .A2(n_257_76_2366), .ZN(n_257_76_2367));
   NAND2_X1 i_257_76_2371 (.A1(n_257_438), .A2(n_257_76_5502), .ZN(n_257_76_2368));
   NAND2_X1 i_257_76_2372 (.A1(n_257_76_2367), .A2(n_257_76_2368), .ZN(
      n_257_76_2369));
   NOR2_X1 i_257_76_2373 (.A1(n_257_76_2364), .A2(n_257_76_2369), .ZN(
      n_257_76_2370));
   NAND3_X1 i_257_76_2374 (.A1(n_257_704), .A2(n_257_435), .A3(n_257_442), 
      .ZN(n_257_76_2371));
   NAND2_X1 i_257_76_2375 (.A1(n_257_76_2371), .A2(n_257_76_2110), .ZN(
      n_257_76_2372));
   INV_X1 i_257_76_2376 (.A(n_257_76_2372), .ZN(n_257_76_2373));
   NAND2_X1 i_257_76_2377 (.A1(n_257_600), .A2(n_257_442), .ZN(n_257_76_2374));
   INV_X1 i_257_76_2378 (.A(n_257_76_2374), .ZN(n_257_76_2375));
   NAND2_X1 i_257_76_2379 (.A1(n_257_432), .A2(n_257_76_2375), .ZN(n_257_76_2376));
   NAND2_X1 i_257_76_2380 (.A1(n_257_76_2376), .A2(n_257_76_2320), .ZN(
      n_257_76_2377));
   INV_X1 i_257_76_2381 (.A(Small_Packet_Data_Size[3]), .ZN(n_257_76_2378));
   NAND2_X1 i_257_76_2382 (.A1(n_257_76_1947), .A2(n_257_76_18055), .ZN(
      n_257_76_2379));
   NOR2_X1 i_257_76_2383 (.A1(n_257_76_2377), .A2(n_257_76_2379), .ZN(
      n_257_76_2380));
   NAND2_X1 i_257_76_2384 (.A1(n_257_76_2373), .A2(n_257_76_2380), .ZN(
      n_257_76_2381));
   INV_X1 i_257_76_2385 (.A(n_257_632), .ZN(n_257_76_2382));
   OAI21_X1 i_257_76_2386 (.A(n_257_76_2264), .B1(n_257_76_2382), .B2(
      n_257_76_17927), .ZN(n_257_76_2383));
   NOR2_X1 i_257_76_2387 (.A1(n_257_76_2381), .A2(n_257_76_2383), .ZN(
      n_257_76_2384));
   NAND2_X1 i_257_76_2388 (.A1(n_257_76_2370), .A2(n_257_76_2384), .ZN(
      n_257_76_2385));
   INV_X1 i_257_76_2389 (.A(n_257_76_2385), .ZN(n_257_76_2386));
   NAND2_X1 i_257_76_2390 (.A1(n_257_800), .A2(n_257_76_17952), .ZN(
      n_257_76_2387));
   NAND2_X1 i_257_76_2391 (.A1(n_257_832), .A2(n_257_442), .ZN(n_257_76_2388));
   INV_X1 i_257_76_2392 (.A(n_257_76_2388), .ZN(n_257_76_2389));
   NAND2_X1 i_257_76_2393 (.A1(n_257_446), .A2(n_257_76_2389), .ZN(n_257_76_2390));
   NAND2_X1 i_257_76_2394 (.A1(n_257_76_2387), .A2(n_257_76_2390), .ZN(
      n_257_76_2391));
   NAND2_X1 i_257_76_2395 (.A1(n_257_449), .A2(n_257_76_9900), .ZN(n_257_76_2392));
   NAND2_X1 i_257_76_2396 (.A1(n_257_768), .A2(n_257_442), .ZN(n_257_76_2393));
   INV_X1 i_257_76_2397 (.A(n_257_76_2393), .ZN(n_257_76_2394));
   NAND2_X1 i_257_76_2398 (.A1(n_257_447), .A2(n_257_76_2394), .ZN(n_257_76_2395));
   NAND2_X1 i_257_76_2399 (.A1(n_257_76_2392), .A2(n_257_76_2395), .ZN(
      n_257_76_2396));
   NOR2_X1 i_257_76_2400 (.A1(n_257_76_2391), .A2(n_257_76_2396), .ZN(
      n_257_76_2397));
   NAND2_X1 i_257_76_2401 (.A1(n_257_76_2386), .A2(n_257_76_2397), .ZN(
      n_257_76_2398));
   NOR2_X1 i_257_76_2402 (.A1(n_257_76_2361), .A2(n_257_76_2398), .ZN(
      n_257_76_2399));
   NAND2_X1 i_257_76_2403 (.A1(n_257_76_2345), .A2(n_257_76_2399), .ZN(
      n_257_76_2400));
   NAND2_X1 i_257_76_2404 (.A1(n_257_76_1896), .A2(n_257_76_1990), .ZN(
      n_257_76_2401));
   INV_X1 i_257_76_2405 (.A(n_257_76_2401), .ZN(n_257_76_2402));
   NAND2_X1 i_257_76_2406 (.A1(n_257_998), .A2(n_257_76_17964), .ZN(
      n_257_76_2403));
   NAND2_X1 i_257_76_2407 (.A1(n_257_76_2402), .A2(n_257_76_2403), .ZN(
      n_257_76_2404));
   NOR2_X1 i_257_76_2408 (.A1(n_257_76_2400), .A2(n_257_76_2404), .ZN(
      n_257_76_2405));
   NAND2_X1 i_257_76_2409 (.A1(n_257_76_2341), .A2(n_257_76_2405), .ZN(
      n_257_76_2406));
   NAND3_X1 i_257_76_2410 (.A1(n_257_76_2300), .A2(n_257_76_2337), .A3(
      n_257_76_2406), .ZN(n_257_76_2407));
   INV_X1 i_257_76_2411 (.A(n_257_76_2407), .ZN(n_257_76_2408));
   NAND3_X1 i_257_76_2412 (.A1(n_257_76_2229), .A2(n_257_76_2278), .A3(
      n_257_76_2408), .ZN(n_257_76_2409));
   NOR2_X1 i_257_76_2413 (.A1(n_257_76_2176), .A2(n_257_76_2409), .ZN(
      n_257_76_2410));
   NAND2_X1 i_257_76_2414 (.A1(n_257_76_2050), .A2(n_257_76_2410), .ZN(n_3));
   NAND2_X1 i_257_76_2415 (.A1(n_257_1031), .A2(n_257_443), .ZN(n_257_76_2411));
   NAND2_X1 i_257_76_2416 (.A1(n_257_999), .A2(n_257_444), .ZN(n_257_76_2412));
   NAND2_X1 i_257_76_2417 (.A1(n_257_441), .A2(n_257_967), .ZN(n_257_76_2413));
   INV_X1 i_257_76_2418 (.A(n_257_1063), .ZN(n_257_76_2414));
   NAND2_X1 i_257_76_2419 (.A1(n_257_442), .A2(n_257_76_2414), .ZN(n_257_76_2415));
   INV_X1 i_257_76_2420 (.A(n_257_935), .ZN(n_257_76_2416));
   NOR2_X1 i_257_76_2421 (.A1(n_257_76_2415), .A2(n_257_76_2416), .ZN(
      n_257_76_2417));
   NAND2_X1 i_257_76_2422 (.A1(n_257_440), .A2(n_257_76_2417), .ZN(n_257_76_2418));
   INV_X1 i_257_76_2423 (.A(n_257_76_2418), .ZN(n_257_76_2419));
   NAND2_X1 i_257_76_2424 (.A1(n_257_76_2413), .A2(n_257_76_2419), .ZN(
      n_257_76_2420));
   INV_X1 i_257_76_2425 (.A(n_257_76_2420), .ZN(n_257_76_2421));
   NAND2_X1 i_257_76_2426 (.A1(n_257_76_2412), .A2(n_257_76_2421), .ZN(
      n_257_76_2422));
   INV_X1 i_257_76_2427 (.A(n_257_76_2422), .ZN(n_257_76_2423));
   NAND2_X1 i_257_76_2428 (.A1(n_257_76_2411), .A2(n_257_76_2423), .ZN(
      n_257_76_2424));
   INV_X1 i_257_76_2429 (.A(n_257_76_2424), .ZN(n_257_76_2425));
   NAND2_X1 i_257_76_2430 (.A1(n_257_17), .A2(n_257_76_2425), .ZN(n_257_76_2426));
   INV_X1 i_257_76_2431 (.A(n_257_76_2415), .ZN(n_257_76_2427));
   NAND2_X1 i_257_76_2432 (.A1(n_257_443), .A2(n_257_76_2427), .ZN(n_257_76_2428));
   INV_X1 i_257_76_2433 (.A(n_257_76_2428), .ZN(n_257_76_2429));
   NAND2_X1 i_257_76_2434 (.A1(n_257_1031), .A2(n_257_76_2429), .ZN(
      n_257_76_2430));
   INV_X1 i_257_76_2435 (.A(n_257_76_2430), .ZN(n_257_76_2431));
   NAND2_X1 i_257_76_2436 (.A1(n_257_14), .A2(n_257_76_2431), .ZN(n_257_76_2432));
   INV_X1 i_257_76_2437 (.A(n_257_76_2411), .ZN(n_257_76_2433));
   NAND2_X1 i_257_76_2438 (.A1(n_257_440), .A2(n_257_935), .ZN(n_257_76_2434));
   NAND2_X1 i_257_76_2439 (.A1(n_257_438), .A2(n_257_1069), .ZN(n_257_76_2435));
   NAND2_X1 i_257_76_2440 (.A1(n_257_865), .A2(n_257_445), .ZN(n_257_76_2436));
   NAND3_X1 i_257_76_2441 (.A1(n_257_76_2434), .A2(n_257_76_2435), .A3(
      n_257_76_2436), .ZN(n_257_76_2437));
   INV_X1 i_257_76_2442 (.A(n_257_76_2437), .ZN(n_257_76_2438));
   NAND2_X1 i_257_76_2443 (.A1(n_257_737), .A2(n_257_436), .ZN(n_257_76_2439));
   NAND2_X1 i_257_76_2444 (.A1(n_257_801), .A2(n_257_437), .ZN(n_257_76_2440));
   NAND2_X1 i_257_76_2445 (.A1(n_257_76_2439), .A2(n_257_76_2440), .ZN(
      n_257_76_2441));
   INV_X1 i_257_76_2446 (.A(n_257_76_2441), .ZN(n_257_76_2442));
   NAND2_X1 i_257_76_2447 (.A1(n_257_439), .A2(n_257_903), .ZN(n_257_76_2443));
   NAND2_X1 i_257_76_2448 (.A1(n_257_435), .A2(n_257_705), .ZN(n_257_76_2444));
   NAND3_X1 i_257_76_2449 (.A1(n_257_76_2444), .A2(n_257_450), .A3(n_257_76_2427), 
      .ZN(n_257_76_2445));
   INV_X1 i_257_76_2450 (.A(n_257_76_2445), .ZN(n_257_76_2446));
   NAND3_X1 i_257_76_2451 (.A1(n_257_76_2443), .A2(n_257_633), .A3(n_257_76_2446), 
      .ZN(n_257_76_2447));
   INV_X1 i_257_76_2452 (.A(n_257_76_2447), .ZN(n_257_76_2448));
   NAND3_X1 i_257_76_2453 (.A1(n_257_76_2438), .A2(n_257_76_2442), .A3(
      n_257_76_2448), .ZN(n_257_76_2449));
   NAND2_X1 i_257_76_2454 (.A1(n_257_446), .A2(n_257_833), .ZN(n_257_76_2450));
   NAND2_X1 i_257_76_2455 (.A1(n_257_449), .A2(n_257_1077), .ZN(n_257_76_2451));
   NAND2_X1 i_257_76_2456 (.A1(n_257_447), .A2(n_257_769), .ZN(n_257_76_2452));
   NAND3_X1 i_257_76_2457 (.A1(n_257_76_2450), .A2(n_257_76_2451), .A3(
      n_257_76_2452), .ZN(n_257_76_2453));
   NOR2_X1 i_257_76_2458 (.A1(n_257_76_2449), .A2(n_257_76_2453), .ZN(
      n_257_76_2454));
   NAND2_X1 i_257_76_2459 (.A1(n_257_673), .A2(n_257_448), .ZN(n_257_76_2455));
   NAND2_X1 i_257_76_2460 (.A1(n_257_76_2455), .A2(n_257_76_2413), .ZN(
      n_257_76_2456));
   INV_X1 i_257_76_2461 (.A(n_257_76_2456), .ZN(n_257_76_2457));
   NAND3_X1 i_257_76_2462 (.A1(n_257_76_2454), .A2(n_257_76_2457), .A3(
      n_257_76_2412), .ZN(n_257_76_2458));
   NOR2_X1 i_257_76_2463 (.A1(n_257_76_2433), .A2(n_257_76_2458), .ZN(
      n_257_76_2459));
   NAND2_X1 i_257_76_2464 (.A1(n_257_28), .A2(n_257_76_2459), .ZN(n_257_76_2460));
   NAND3_X1 i_257_76_2465 (.A1(n_257_76_2426), .A2(n_257_76_2432), .A3(
      n_257_76_2460), .ZN(n_257_76_2461));
   NAND3_X1 i_257_76_2466 (.A1(n_257_446), .A2(n_257_76_2434), .A3(n_257_76_2435), 
      .ZN(n_257_76_2462));
   INV_X1 i_257_76_2467 (.A(n_257_76_2462), .ZN(n_257_76_2463));
   INV_X1 i_257_76_2468 (.A(n_257_833), .ZN(n_257_76_2464));
   NOR2_X1 i_257_76_2469 (.A1(n_257_76_2464), .A2(n_257_76_2415), .ZN(
      n_257_76_2465));
   NAND3_X1 i_257_76_2470 (.A1(n_257_76_2436), .A2(n_257_76_2443), .A3(
      n_257_76_2465), .ZN(n_257_76_2466));
   INV_X1 i_257_76_2471 (.A(n_257_76_2466), .ZN(n_257_76_2467));
   NAND3_X1 i_257_76_2472 (.A1(n_257_76_2413), .A2(n_257_76_2463), .A3(
      n_257_76_2467), .ZN(n_257_76_2468));
   INV_X1 i_257_76_2473 (.A(n_257_76_2468), .ZN(n_257_76_2469));
   NAND2_X1 i_257_76_2474 (.A1(n_257_76_2412), .A2(n_257_76_2469), .ZN(
      n_257_76_2470));
   INV_X1 i_257_76_2475 (.A(n_257_76_2470), .ZN(n_257_76_2471));
   NAND2_X1 i_257_76_2476 (.A1(n_257_76_2411), .A2(n_257_76_2471), .ZN(
      n_257_76_2472));
   INV_X1 i_257_76_2477 (.A(n_257_76_2472), .ZN(n_257_76_2473));
   NAND2_X1 i_257_76_2478 (.A1(n_257_21), .A2(n_257_76_2473), .ZN(n_257_76_2474));
   INV_X1 i_257_76_2479 (.A(n_257_76_2434), .ZN(n_257_76_2475));
   NAND3_X1 i_257_76_2480 (.A1(n_257_439), .A2(n_257_903), .A3(n_257_76_2427), 
      .ZN(n_257_76_2476));
   NOR2_X1 i_257_76_2481 (.A1(n_257_76_2475), .A2(n_257_76_2476), .ZN(
      n_257_76_2477));
   NAND2_X1 i_257_76_2482 (.A1(n_257_76_2413), .A2(n_257_76_2477), .ZN(
      n_257_76_2478));
   INV_X1 i_257_76_2483 (.A(n_257_76_2478), .ZN(n_257_76_2479));
   NAND2_X1 i_257_76_2484 (.A1(n_257_76_2412), .A2(n_257_76_2479), .ZN(
      n_257_76_2480));
   INV_X1 i_257_76_2485 (.A(n_257_76_2480), .ZN(n_257_76_2481));
   NAND2_X1 i_257_76_2486 (.A1(n_257_76_2411), .A2(n_257_76_2481), .ZN(
      n_257_76_2482));
   INV_X1 i_257_76_2487 (.A(n_257_76_2482), .ZN(n_257_76_2483));
   NAND2_X1 i_257_76_2488 (.A1(n_257_18), .A2(n_257_76_2483), .ZN(n_257_76_2484));
   NAND2_X1 i_257_76_2489 (.A1(n_257_505), .A2(n_257_424), .ZN(n_257_76_2485));
   NAND2_X1 i_257_76_2490 (.A1(n_257_76_2485), .A2(n_257_276), .ZN(n_257_76_2486));
   NAND2_X1 i_257_76_2491 (.A1(n_257_428), .A2(n_257_569), .ZN(n_257_76_2487));
   INV_X1 i_257_76_2492 (.A(n_257_76_2487), .ZN(n_257_76_2488));
   NAND2_X1 i_257_76_2493 (.A1(n_257_423), .A2(n_257_76_2427), .ZN(n_257_76_2489));
   NOR2_X1 i_257_76_2494 (.A1(n_257_76_2488), .A2(n_257_76_2489), .ZN(
      n_257_76_2490));
   NAND2_X1 i_257_76_2495 (.A1(n_257_432), .A2(n_257_601), .ZN(n_257_76_2491));
   NAND3_X1 i_257_76_2496 (.A1(n_257_76_2490), .A2(n_257_76_2444), .A3(
      n_257_76_2491), .ZN(n_257_76_2492));
   NOR2_X1 i_257_76_2497 (.A1(n_257_76_2486), .A2(n_257_76_2492), .ZN(
      n_257_76_2493));
   NAND2_X1 i_257_76_2498 (.A1(n_257_633), .A2(n_257_450), .ZN(n_257_76_2494));
   NAND2_X1 i_257_76_2499 (.A1(n_257_39), .A2(n_257_433), .ZN(n_257_76_2495));
   NAND2_X1 i_257_76_2500 (.A1(n_257_76_2494), .A2(n_257_76_2495), .ZN(
      n_257_76_2496));
   INV_X1 i_257_76_2501 (.A(n_257_76_2496), .ZN(n_257_76_2497));
   NAND2_X1 i_257_76_2502 (.A1(n_257_117), .A2(n_257_430), .ZN(n_257_76_2498));
   NAND3_X1 i_257_76_2503 (.A1(n_257_76_2493), .A2(n_257_76_2497), .A3(
      n_257_76_2498), .ZN(n_257_76_2499));
   INV_X1 i_257_76_2504 (.A(n_257_76_2499), .ZN(n_257_76_2500));
   NAND2_X1 i_257_76_2505 (.A1(n_257_156), .A2(n_257_429), .ZN(n_257_76_2501));
   NAND3_X1 i_257_76_2506 (.A1(n_257_76_2500), .A2(n_257_76_2455), .A3(
      n_257_76_2501), .ZN(n_257_76_2502));
   INV_X1 i_257_76_2507 (.A(n_257_76_2412), .ZN(n_257_76_2503));
   NOR2_X1 i_257_76_2508 (.A1(n_257_76_2502), .A2(n_257_76_2503), .ZN(
      n_257_76_2504));
   NAND3_X1 i_257_76_2509 (.A1(n_257_76_2440), .A2(n_257_76_2434), .A3(
      n_257_76_2435), .ZN(n_257_76_2505));
   NAND2_X1 i_257_76_2510 (.A1(n_257_427), .A2(n_257_196), .ZN(n_257_76_2506));
   NAND3_X1 i_257_76_2511 (.A1(n_257_76_2436), .A2(n_257_76_2443), .A3(
      n_257_76_2506), .ZN(n_257_76_2507));
   NOR2_X1 i_257_76_2512 (.A1(n_257_76_2505), .A2(n_257_76_2507), .ZN(
      n_257_76_2508));
   INV_X1 i_257_76_2513 (.A(n_257_76_2453), .ZN(n_257_76_2509));
   NAND2_X1 i_257_76_2514 (.A1(n_257_451), .A2(n_257_456), .ZN(n_257_76_2510));
   NAND2_X1 i_257_76_2515 (.A1(n_257_537), .A2(n_257_426), .ZN(n_257_76_2511));
   NAND3_X1 i_257_76_2516 (.A1(n_257_76_2510), .A2(n_257_76_2511), .A3(
      n_257_76_2439), .ZN(n_257_76_2512));
   INV_X1 i_257_76_2517 (.A(n_257_76_2512), .ZN(n_257_76_2513));
   NAND3_X1 i_257_76_2518 (.A1(n_257_76_2508), .A2(n_257_76_2509), .A3(
      n_257_76_2513), .ZN(n_257_76_2514));
   NAND2_X1 i_257_76_2519 (.A1(n_257_236), .A2(n_257_425), .ZN(n_257_76_2515));
   NAND2_X1 i_257_76_2520 (.A1(n_257_79), .A2(n_257_431), .ZN(n_257_76_2516));
   NAND3_X1 i_257_76_2521 (.A1(n_257_76_2515), .A2(n_257_76_2413), .A3(
      n_257_76_2516), .ZN(n_257_76_2517));
   NOR2_X1 i_257_76_2522 (.A1(n_257_76_2514), .A2(n_257_76_2517), .ZN(
      n_257_76_2518));
   NAND3_X1 i_257_76_2523 (.A1(n_257_76_2504), .A2(n_257_76_2411), .A3(
      n_257_76_2518), .ZN(n_257_76_2519));
   INV_X1 i_257_76_2524 (.A(n_257_76_2519), .ZN(n_257_76_2520));
   NAND2_X1 i_257_76_2525 (.A1(n_257_304), .A2(n_257_76_2520), .ZN(n_257_76_2521));
   NAND3_X1 i_257_76_2526 (.A1(n_257_76_2474), .A2(n_257_76_2484), .A3(
      n_257_76_2521), .ZN(n_257_76_2522));
   NOR2_X1 i_257_76_2527 (.A1(n_257_76_2461), .A2(n_257_76_2522), .ZN(
      n_257_76_2523));
   NAND2_X1 i_257_76_2528 (.A1(n_257_967), .A2(n_257_76_2427), .ZN(n_257_76_2524));
   INV_X1 i_257_76_2529 (.A(n_257_76_2524), .ZN(n_257_76_2525));
   NAND2_X1 i_257_76_2530 (.A1(n_257_441), .A2(n_257_76_2525), .ZN(n_257_76_2526));
   INV_X1 i_257_76_2531 (.A(n_257_76_2526), .ZN(n_257_76_2527));
   NAND2_X1 i_257_76_2532 (.A1(n_257_76_2412), .A2(n_257_76_2527), .ZN(
      n_257_76_2528));
   INV_X1 i_257_76_2533 (.A(n_257_76_2528), .ZN(n_257_76_2529));
   NAND2_X1 i_257_76_2534 (.A1(n_257_76_2411), .A2(n_257_76_2529), .ZN(
      n_257_76_2530));
   INV_X1 i_257_76_2535 (.A(n_257_76_2530), .ZN(n_257_76_2531));
   NAND2_X1 i_257_76_2536 (.A1(n_257_16), .A2(n_257_76_2531), .ZN(n_257_76_2532));
   NAND2_X1 i_257_76_2537 (.A1(n_257_76_2450), .A2(n_257_76_2452), .ZN(
      n_257_76_2533));
   INV_X1 i_257_76_2538 (.A(n_257_76_2533), .ZN(n_257_76_2534));
   NAND3_X1 i_257_76_2539 (.A1(n_257_435), .A2(n_257_705), .A3(n_257_76_2427), 
      .ZN(n_257_76_2535));
   INV_X1 i_257_76_2540 (.A(n_257_76_2535), .ZN(n_257_76_2536));
   NAND4_X1 i_257_76_2541 (.A1(n_257_76_2435), .A2(n_257_76_2436), .A3(
      n_257_76_2443), .A4(n_257_76_2536), .ZN(n_257_76_2537));
   INV_X1 i_257_76_2542 (.A(n_257_76_2537), .ZN(n_257_76_2538));
   NAND3_X1 i_257_76_2543 (.A1(n_257_76_2439), .A2(n_257_76_2440), .A3(
      n_257_76_2434), .ZN(n_257_76_2539));
   INV_X1 i_257_76_2544 (.A(n_257_76_2539), .ZN(n_257_76_2540));
   NAND4_X1 i_257_76_2545 (.A1(n_257_76_2534), .A2(n_257_76_2538), .A3(
      n_257_76_2413), .A4(n_257_76_2540), .ZN(n_257_76_2541));
   INV_X1 i_257_76_2546 (.A(n_257_76_2541), .ZN(n_257_76_2542));
   NAND2_X1 i_257_76_2547 (.A1(n_257_76_2542), .A2(n_257_76_2412), .ZN(
      n_257_76_2543));
   NOR2_X1 i_257_76_2548 (.A1(n_257_76_2433), .A2(n_257_76_2543), .ZN(
      n_257_76_2544));
   NAND2_X1 i_257_76_2549 (.A1(n_257_25), .A2(n_257_76_2544), .ZN(n_257_76_2545));
   NAND3_X1 i_257_76_2550 (.A1(n_257_442), .A2(n_257_569), .A3(n_257_76_2414), 
      .ZN(n_257_76_2546));
   INV_X1 i_257_76_2551 (.A(n_257_76_2546), .ZN(n_257_76_2547));
   NAND2_X1 i_257_76_2552 (.A1(n_257_428), .A2(n_257_76_2547), .ZN(n_257_76_2548));
   INV_X1 i_257_76_2553 (.A(n_257_76_2548), .ZN(n_257_76_2549));
   NAND3_X1 i_257_76_2554 (.A1(n_257_76_2444), .A2(n_257_76_2491), .A3(
      n_257_76_2549), .ZN(n_257_76_2550));
   INV_X1 i_257_76_2555 (.A(n_257_76_2550), .ZN(n_257_76_2551));
   NAND3_X1 i_257_76_2556 (.A1(n_257_76_2494), .A2(n_257_76_2551), .A3(
      n_257_76_2495), .ZN(n_257_76_2552));
   INV_X1 i_257_76_2557 (.A(n_257_76_2552), .ZN(n_257_76_2553));
   NAND2_X1 i_257_76_2558 (.A1(n_257_76_2436), .A2(n_257_76_2443), .ZN(
      n_257_76_2554));
   INV_X1 i_257_76_2559 (.A(n_257_76_2554), .ZN(n_257_76_2555));
   NAND2_X1 i_257_76_2560 (.A1(n_257_76_2553), .A2(n_257_76_2555), .ZN(
      n_257_76_2556));
   NAND4_X1 i_257_76_2561 (.A1(n_257_76_2439), .A2(n_257_76_2440), .A3(
      n_257_76_2434), .A4(n_257_76_2435), .ZN(n_257_76_2557));
   NOR2_X1 i_257_76_2562 (.A1(n_257_76_2556), .A2(n_257_76_2557), .ZN(
      n_257_76_2558));
   NAND3_X1 i_257_76_2563 (.A1(n_257_76_2413), .A2(n_257_76_2516), .A3(
      n_257_76_2450), .ZN(n_257_76_2559));
   INV_X1 i_257_76_2564 (.A(n_257_76_2559), .ZN(n_257_76_2560));
   NAND4_X1 i_257_76_2565 (.A1(n_257_76_2451), .A2(n_257_76_2452), .A3(
      n_257_76_2510), .A4(n_257_76_2498), .ZN(n_257_76_2561));
   INV_X1 i_257_76_2566 (.A(n_257_76_2561), .ZN(n_257_76_2562));
   NAND4_X1 i_257_76_2567 (.A1(n_257_76_2558), .A2(n_257_76_2560), .A3(
      n_257_76_2501), .A4(n_257_76_2562), .ZN(n_257_76_2563));
   INV_X1 i_257_76_2568 (.A(n_257_76_2563), .ZN(n_257_76_2564));
   NAND2_X1 i_257_76_2569 (.A1(n_257_76_2412), .A2(n_257_76_2455), .ZN(
      n_257_76_2565));
   INV_X1 i_257_76_2570 (.A(n_257_76_2565), .ZN(n_257_76_2566));
   NAND3_X1 i_257_76_2571 (.A1(n_257_76_2564), .A2(n_257_76_2411), .A3(
      n_257_76_2566), .ZN(n_257_76_2567));
   INV_X1 i_257_76_2572 (.A(n_257_76_2567), .ZN(n_257_76_2568));
   NAND2_X1 i_257_76_2573 (.A1(n_257_185), .A2(n_257_76_2568), .ZN(n_257_76_2569));
   NAND3_X1 i_257_76_2574 (.A1(n_257_76_2532), .A2(n_257_76_2545), .A3(
      n_257_76_2569), .ZN(n_257_76_2570));
   NAND2_X1 i_257_76_2575 (.A1(n_257_442), .A2(n_257_1063), .ZN(n_257_76_2571));
   INV_X1 i_257_76_2576 (.A(n_257_76_2571), .ZN(n_257_76_2572));
   NAND2_X1 i_257_76_2577 (.A1(n_257_13), .A2(n_257_76_2572), .ZN(n_257_76_2573));
   INV_X1 i_257_76_2578 (.A(n_257_76_2413), .ZN(n_257_76_2574));
   NAND2_X1 i_257_76_2579 (.A1(n_257_445), .A2(n_257_76_2427), .ZN(n_257_76_2575));
   INV_X1 i_257_76_2580 (.A(n_257_76_2575), .ZN(n_257_76_2576));
   NAND2_X1 i_257_76_2581 (.A1(n_257_76_2576), .A2(n_257_865), .ZN(n_257_76_2577));
   INV_X1 i_257_76_2582 (.A(n_257_76_2577), .ZN(n_257_76_2578));
   NAND4_X1 i_257_76_2583 (.A1(n_257_76_2578), .A2(n_257_76_2434), .A3(
      n_257_76_2435), .A4(n_257_76_2443), .ZN(n_257_76_2579));
   NOR2_X1 i_257_76_2584 (.A1(n_257_76_2574), .A2(n_257_76_2579), .ZN(
      n_257_76_2580));
   NAND2_X1 i_257_76_2585 (.A1(n_257_76_2412), .A2(n_257_76_2580), .ZN(
      n_257_76_2581));
   INV_X1 i_257_76_2586 (.A(n_257_76_2581), .ZN(n_257_76_2582));
   NAND2_X1 i_257_76_2587 (.A1(n_257_76_2411), .A2(n_257_76_2582), .ZN(
      n_257_76_2583));
   INV_X1 i_257_76_2588 (.A(n_257_76_2583), .ZN(n_257_76_2584));
   NAND2_X1 i_257_76_2589 (.A1(n_257_20), .A2(n_257_76_2584), .ZN(n_257_76_2585));
   NAND2_X1 i_257_76_2590 (.A1(n_257_76_2573), .A2(n_257_76_2585), .ZN(
      n_257_76_2586));
   NOR2_X1 i_257_76_2591 (.A1(n_257_76_2570), .A2(n_257_76_2586), .ZN(
      n_257_76_2587));
   NAND2_X1 i_257_76_2592 (.A1(n_257_426), .A2(n_257_76_2427), .ZN(n_257_76_2588));
   NOR2_X1 i_257_76_2593 (.A1(n_257_76_2488), .A2(n_257_76_2588), .ZN(
      n_257_76_2589));
   NAND3_X1 i_257_76_2594 (.A1(n_257_76_2589), .A2(n_257_76_2444), .A3(
      n_257_76_2491), .ZN(n_257_76_2590));
   INV_X1 i_257_76_2595 (.A(n_257_76_2590), .ZN(n_257_76_2591));
   NAND3_X1 i_257_76_2596 (.A1(n_257_76_2591), .A2(n_257_76_2495), .A3(
      n_257_76_2506), .ZN(n_257_76_2592));
   NAND3_X1 i_257_76_2597 (.A1(n_257_537), .A2(n_257_76_2443), .A3(n_257_76_2494), 
      .ZN(n_257_76_2593));
   NOR2_X1 i_257_76_2598 (.A1(n_257_76_2592), .A2(n_257_76_2593), .ZN(
      n_257_76_2594));
   NAND3_X1 i_257_76_2599 (.A1(n_257_76_2498), .A2(n_257_76_2439), .A3(
      n_257_76_2440), .ZN(n_257_76_2595));
   INV_X1 i_257_76_2600 (.A(n_257_76_2595), .ZN(n_257_76_2596));
   NAND4_X1 i_257_76_2601 (.A1(n_257_76_2594), .A2(n_257_76_2596), .A3(
      n_257_76_2516), .A4(n_257_76_2438), .ZN(n_257_76_2597));
   INV_X1 i_257_76_2602 (.A(n_257_76_2597), .ZN(n_257_76_2598));
   NAND2_X1 i_257_76_2603 (.A1(n_257_76_2455), .A2(n_257_76_2501), .ZN(
      n_257_76_2599));
   INV_X1 i_257_76_2604 (.A(n_257_76_2599), .ZN(n_257_76_2600));
   NAND2_X1 i_257_76_2605 (.A1(n_257_76_2450), .A2(n_257_76_2451), .ZN(
      n_257_76_2601));
   INV_X1 i_257_76_2606 (.A(n_257_76_2601), .ZN(n_257_76_2602));
   NAND2_X1 i_257_76_2607 (.A1(n_257_76_2452), .A2(n_257_76_2510), .ZN(
      n_257_76_2603));
   INV_X1 i_257_76_2608 (.A(n_257_76_2603), .ZN(n_257_76_2604));
   NAND3_X1 i_257_76_2609 (.A1(n_257_76_2602), .A2(n_257_76_2604), .A3(
      n_257_76_2413), .ZN(n_257_76_2605));
   INV_X1 i_257_76_2610 (.A(n_257_76_2605), .ZN(n_257_76_2606));
   NAND4_X1 i_257_76_2611 (.A1(n_257_76_2598), .A2(n_257_76_2600), .A3(
      n_257_76_2412), .A4(n_257_76_2606), .ZN(n_257_76_2607));
   NOR2_X1 i_257_76_2612 (.A1(n_257_76_2607), .A2(n_257_76_2433), .ZN(
      n_257_76_2608));
   NAND2_X1 i_257_76_2613 (.A1(n_257_225), .A2(n_257_76_2608), .ZN(n_257_76_2609));
   NAND2_X1 i_257_76_2614 (.A1(n_257_436), .A2(n_257_76_2427), .ZN(n_257_76_2610));
   INV_X1 i_257_76_2615 (.A(n_257_76_2610), .ZN(n_257_76_2611));
   NAND4_X1 i_257_76_2616 (.A1(n_257_76_2436), .A2(n_257_76_2443), .A3(n_257_737), 
      .A4(n_257_76_2611), .ZN(n_257_76_2612));
   NOR2_X1 i_257_76_2617 (.A1(n_257_76_2612), .A2(n_257_76_2505), .ZN(
      n_257_76_2613));
   NAND3_X1 i_257_76_2618 (.A1(n_257_76_2613), .A2(n_257_76_2534), .A3(
      n_257_76_2413), .ZN(n_257_76_2614));
   INV_X1 i_257_76_2619 (.A(n_257_76_2614), .ZN(n_257_76_2615));
   NAND2_X1 i_257_76_2620 (.A1(n_257_76_2615), .A2(n_257_76_2412), .ZN(
      n_257_76_2616));
   NOR2_X1 i_257_76_2621 (.A1(n_257_76_2433), .A2(n_257_76_2616), .ZN(
      n_257_76_2617));
   NAND2_X1 i_257_76_2622 (.A1(n_257_24), .A2(n_257_76_2617), .ZN(n_257_76_2618));
   NOR2_X1 i_257_76_2623 (.A1(n_257_76_2453), .A2(n_257_76_2574), .ZN(
      n_257_76_2619));
   NAND3_X1 i_257_76_2624 (.A1(n_257_76_2435), .A2(n_257_76_2436), .A3(
      n_257_76_2443), .ZN(n_257_76_2620));
   INV_X1 i_257_76_2625 (.A(n_257_76_2620), .ZN(n_257_76_2621));
   INV_X1 i_257_76_2626 (.A(n_257_76_2444), .ZN(n_257_76_2622));
   INV_X1 i_257_76_2627 (.A(n_257_601), .ZN(n_257_76_2623));
   NOR2_X1 i_257_76_2628 (.A1(n_257_76_2415), .A2(n_257_76_2623), .ZN(
      n_257_76_2624));
   NAND2_X1 i_257_76_2629 (.A1(n_257_432), .A2(n_257_76_2624), .ZN(n_257_76_2625));
   NOR2_X1 i_257_76_2630 (.A1(n_257_76_2622), .A2(n_257_76_2625), .ZN(
      n_257_76_2626));
   NAND3_X1 i_257_76_2631 (.A1(n_257_76_2494), .A2(n_257_76_2626), .A3(
      n_257_76_2495), .ZN(n_257_76_2627));
   INV_X1 i_257_76_2632 (.A(n_257_76_2627), .ZN(n_257_76_2628));
   NAND4_X1 i_257_76_2633 (.A1(n_257_76_2540), .A2(n_257_76_2621), .A3(
      n_257_76_2510), .A4(n_257_76_2628), .ZN(n_257_76_2629));
   INV_X1 i_257_76_2634 (.A(n_257_76_2629), .ZN(n_257_76_2630));
   NAND4_X1 i_257_76_2635 (.A1(n_257_76_2412), .A2(n_257_76_2619), .A3(
      n_257_76_2630), .A4(n_257_76_2455), .ZN(n_257_76_2631));
   NOR2_X1 i_257_76_2636 (.A1(n_257_76_2631), .A2(n_257_76_2433), .ZN(
      n_257_76_2632));
   NAND2_X1 i_257_76_2637 (.A1(n_257_68), .A2(n_257_76_2632), .ZN(n_257_76_2633));
   NAND3_X1 i_257_76_2638 (.A1(n_257_76_2609), .A2(n_257_76_2618), .A3(
      n_257_76_2633), .ZN(n_257_76_2634));
   NAND2_X1 i_257_76_2639 (.A1(n_257_437), .A2(n_257_76_2427), .ZN(n_257_76_2635));
   INV_X1 i_257_76_2640 (.A(n_257_76_2635), .ZN(n_257_76_2636));
   NAND3_X1 i_257_76_2641 (.A1(n_257_76_2443), .A2(n_257_801), .A3(n_257_76_2636), 
      .ZN(n_257_76_2637));
   INV_X1 i_257_76_2642 (.A(n_257_76_2637), .ZN(n_257_76_2638));
   NAND4_X1 i_257_76_2643 (.A1(n_257_76_2413), .A2(n_257_76_2438), .A3(
      n_257_76_2450), .A4(n_257_76_2638), .ZN(n_257_76_2639));
   INV_X1 i_257_76_2644 (.A(n_257_76_2639), .ZN(n_257_76_2640));
   NAND2_X1 i_257_76_2645 (.A1(n_257_76_2412), .A2(n_257_76_2640), .ZN(
      n_257_76_2641));
   INV_X1 i_257_76_2646 (.A(n_257_76_2641), .ZN(n_257_76_2642));
   NAND2_X1 i_257_76_2647 (.A1(n_257_76_2411), .A2(n_257_76_2642), .ZN(
      n_257_76_2643));
   INV_X1 i_257_76_2648 (.A(n_257_76_2643), .ZN(n_257_76_2644));
   NAND2_X1 i_257_76_2649 (.A1(n_257_22), .A2(n_257_76_2644), .ZN(n_257_76_2645));
   NAND2_X1 i_257_76_2650 (.A1(n_257_444), .A2(n_257_76_2427), .ZN(n_257_76_2646));
   INV_X1 i_257_76_2651 (.A(n_257_76_2646), .ZN(n_257_76_2647));
   NAND2_X1 i_257_76_2652 (.A1(n_257_999), .A2(n_257_76_2647), .ZN(n_257_76_2648));
   INV_X1 i_257_76_2653 (.A(n_257_76_2648), .ZN(n_257_76_2649));
   NAND2_X1 i_257_76_2654 (.A1(n_257_76_2411), .A2(n_257_76_2649), .ZN(
      n_257_76_2650));
   INV_X1 i_257_76_2655 (.A(n_257_76_2650), .ZN(n_257_76_2651));
   NAND2_X1 i_257_76_2656 (.A1(n_257_15), .A2(n_257_76_2651), .ZN(n_257_76_2652));
   NAND2_X1 i_257_76_2657 (.A1(n_257_76_2645), .A2(n_257_76_2652), .ZN(
      n_257_76_2653));
   NOR2_X1 i_257_76_2658 (.A1(n_257_76_2634), .A2(n_257_76_2653), .ZN(
      n_257_76_2654));
   NAND3_X1 i_257_76_2659 (.A1(n_257_76_2523), .A2(n_257_76_2587), .A3(
      n_257_76_2654), .ZN(n_257_76_2655));
   INV_X1 i_257_76_2660 (.A(n_257_76_2655), .ZN(n_257_76_2656));
   INV_X1 i_257_76_2661 (.A(n_257_76_2494), .ZN(n_257_76_2657));
   NAND2_X1 i_257_76_2662 (.A1(n_257_433), .A2(n_257_76_2427), .ZN(n_257_76_2658));
   INV_X1 i_257_76_2663 (.A(n_257_76_2658), .ZN(n_257_76_2659));
   NAND3_X1 i_257_76_2664 (.A1(n_257_39), .A2(n_257_76_2444), .A3(n_257_76_2659), 
      .ZN(n_257_76_2660));
   NOR2_X1 i_257_76_2665 (.A1(n_257_76_2657), .A2(n_257_76_2660), .ZN(
      n_257_76_2661));
   NAND4_X1 i_257_76_2666 (.A1(n_257_76_2540), .A2(n_257_76_2621), .A3(
      n_257_76_2510), .A4(n_257_76_2661), .ZN(n_257_76_2662));
   INV_X1 i_257_76_2667 (.A(n_257_76_2662), .ZN(n_257_76_2663));
   NAND4_X1 i_257_76_2668 (.A1(n_257_76_2412), .A2(n_257_76_2619), .A3(
      n_257_76_2663), .A4(n_257_76_2455), .ZN(n_257_76_2664));
   NOR2_X1 i_257_76_2669 (.A1(n_257_76_2664), .A2(n_257_76_2433), .ZN(
      n_257_76_2665));
   NAND2_X1 i_257_76_2670 (.A1(n_257_67), .A2(n_257_76_2665), .ZN(n_257_76_2666));
   NAND2_X1 i_257_76_2671 (.A1(n_257_1077), .A2(n_257_76_2427), .ZN(
      n_257_76_2667));
   INV_X1 i_257_76_2672 (.A(n_257_76_2667), .ZN(n_257_76_2668));
   NAND2_X1 i_257_76_2673 (.A1(n_257_76_2668), .A2(n_257_76_2444), .ZN(
      n_257_76_2669));
   INV_X1 i_257_76_2674 (.A(n_257_76_2669), .ZN(n_257_76_2670));
   NAND3_X1 i_257_76_2675 (.A1(n_257_76_2436), .A2(n_257_76_2443), .A3(
      n_257_76_2670), .ZN(n_257_76_2671));
   NAND2_X1 i_257_76_2676 (.A1(n_257_76_2434), .A2(n_257_76_2435), .ZN(
      n_257_76_2672));
   NOR2_X1 i_257_76_2677 (.A1(n_257_76_2671), .A2(n_257_76_2672), .ZN(
      n_257_76_2673));
   NAND3_X1 i_257_76_2678 (.A1(n_257_76_2439), .A2(n_257_449), .A3(n_257_76_2440), 
      .ZN(n_257_76_2674));
   INV_X1 i_257_76_2679 (.A(n_257_76_2674), .ZN(n_257_76_2675));
   NAND3_X1 i_257_76_2680 (.A1(n_257_76_2673), .A2(n_257_76_2534), .A3(
      n_257_76_2675), .ZN(n_257_76_2676));
   INV_X1 i_257_76_2681 (.A(n_257_76_2676), .ZN(n_257_76_2677));
   NAND3_X1 i_257_76_2682 (.A1(n_257_76_2677), .A2(n_257_76_2457), .A3(
      n_257_76_2412), .ZN(n_257_76_2678));
   NOR2_X1 i_257_76_2683 (.A1(n_257_76_2433), .A2(n_257_76_2678), .ZN(
      n_257_76_2679));
   NAND2_X1 i_257_76_2684 (.A1(n_257_27), .A2(n_257_76_2679), .ZN(n_257_76_2680));
   NAND4_X1 i_257_76_2685 (.A1(n_257_76_2602), .A2(n_257_76_2413), .A3(n_257_156), 
      .A4(n_257_76_2516), .ZN(n_257_76_2681));
   NAND2_X1 i_257_76_2686 (.A1(n_257_429), .A2(n_257_76_2427), .ZN(n_257_76_2682));
   INV_X1 i_257_76_2687 (.A(n_257_76_2682), .ZN(n_257_76_2683));
   NAND3_X1 i_257_76_2688 (.A1(n_257_76_2444), .A2(n_257_76_2491), .A3(
      n_257_76_2683), .ZN(n_257_76_2684));
   INV_X1 i_257_76_2689 (.A(n_257_76_2684), .ZN(n_257_76_2685));
   NAND3_X1 i_257_76_2690 (.A1(n_257_76_2494), .A2(n_257_76_2685), .A3(
      n_257_76_2495), .ZN(n_257_76_2686));
   NOR2_X1 i_257_76_2691 (.A1(n_257_76_2620), .A2(n_257_76_2686), .ZN(
      n_257_76_2687));
   NAND4_X1 i_257_76_2692 (.A1(n_257_76_2498), .A2(n_257_76_2439), .A3(
      n_257_76_2440), .A4(n_257_76_2434), .ZN(n_257_76_2688));
   INV_X1 i_257_76_2693 (.A(n_257_76_2688), .ZN(n_257_76_2689));
   NAND3_X1 i_257_76_2694 (.A1(n_257_76_2687), .A2(n_257_76_2604), .A3(
      n_257_76_2689), .ZN(n_257_76_2690));
   NOR2_X1 i_257_76_2695 (.A1(n_257_76_2681), .A2(n_257_76_2690), .ZN(
      n_257_76_2691));
   NAND3_X1 i_257_76_2696 (.A1(n_257_76_2691), .A2(n_257_76_2411), .A3(
      n_257_76_2566), .ZN(n_257_76_2692));
   INV_X1 i_257_76_2697 (.A(n_257_76_2692), .ZN(n_257_76_2693));
   NAND2_X1 i_257_76_2698 (.A1(n_257_184), .A2(n_257_76_2693), .ZN(n_257_76_2694));
   NAND3_X1 i_257_76_2699 (.A1(n_257_76_2666), .A2(n_257_76_2680), .A3(
      n_257_76_2694), .ZN(n_257_76_2695));
   INV_X1 i_257_76_2700 (.A(n_257_76_2695), .ZN(n_257_76_2696));
   NAND2_X1 i_257_76_2701 (.A1(n_257_1069), .A2(n_257_76_2427), .ZN(
      n_257_76_2697));
   INV_X1 i_257_76_2702 (.A(n_257_76_2697), .ZN(n_257_76_2698));
   NAND2_X1 i_257_76_2703 (.A1(n_257_438), .A2(n_257_76_2698), .ZN(n_257_76_2699));
   INV_X1 i_257_76_2704 (.A(n_257_76_2699), .ZN(n_257_76_2700));
   NAND3_X1 i_257_76_2705 (.A1(n_257_76_2700), .A2(n_257_76_2434), .A3(
      n_257_76_2443), .ZN(n_257_76_2701));
   INV_X1 i_257_76_2706 (.A(n_257_76_2701), .ZN(n_257_76_2702));
   NAND2_X1 i_257_76_2707 (.A1(n_257_76_2413), .A2(n_257_76_2702), .ZN(
      n_257_76_2703));
   INV_X1 i_257_76_2708 (.A(n_257_76_2703), .ZN(n_257_76_2704));
   NAND2_X1 i_257_76_2709 (.A1(n_257_76_2412), .A2(n_257_76_2704), .ZN(
      n_257_76_2705));
   INV_X1 i_257_76_2710 (.A(n_257_76_2705), .ZN(n_257_76_2706));
   NAND2_X1 i_257_76_2711 (.A1(n_257_76_2411), .A2(n_257_76_2706), .ZN(
      n_257_76_2707));
   INV_X1 i_257_76_2712 (.A(n_257_76_2707), .ZN(n_257_76_2708));
   NAND2_X1 i_257_76_2713 (.A1(n_257_19), .A2(n_257_76_2708), .ZN(n_257_76_2709));
   NAND2_X1 i_257_76_2714 (.A1(n_257_76_2413), .A2(n_257_76_2516), .ZN(
      n_257_76_2710));
   INV_X1 i_257_76_2715 (.A(n_257_76_2710), .ZN(n_257_76_2711));
   NAND2_X1 i_257_76_2716 (.A1(n_257_353), .A2(n_257_421), .ZN(n_257_76_2712));
   NAND2_X1 i_257_76_2717 (.A1(n_257_76_2712), .A2(n_257_76_2450), .ZN(
      n_257_76_2713));
   INV_X1 i_257_76_2718 (.A(n_257_76_2713), .ZN(n_257_76_2714));
   NAND2_X1 i_257_76_2719 (.A1(n_257_76_2711), .A2(n_257_76_2714), .ZN(
      n_257_76_2715));
   NAND2_X1 i_257_76_2720 (.A1(n_257_76_2501), .A2(n_257_76_2515), .ZN(
      n_257_76_2716));
   NOR2_X1 i_257_76_2721 (.A1(n_257_76_2715), .A2(n_257_76_2716), .ZN(
      n_257_76_2717));
   NAND2_X1 i_257_76_2722 (.A1(n_257_76_2506), .A2(n_257_76_2485), .ZN(
      n_257_76_2718));
   INV_X1 i_257_76_2723 (.A(n_257_76_2718), .ZN(n_257_76_2719));
   INV_X1 i_257_76_2724 (.A(n_257_895), .ZN(n_257_76_2720));
   NOR2_X1 i_257_76_2725 (.A1(n_257_1063), .A2(n_257_76_2720), .ZN(n_257_76_2721));
   NAND2_X1 i_257_76_2726 (.A1(n_257_442), .A2(n_257_76_2721), .ZN(n_257_76_2722));
   INV_X1 i_257_76_2727 (.A(n_257_76_2722), .ZN(n_257_76_2723));
   NAND2_X1 i_257_76_2728 (.A1(n_257_420), .A2(n_257_76_2723), .ZN(n_257_76_2724));
   NOR2_X1 i_257_76_2729 (.A1(n_257_76_2724), .A2(n_257_76_2488), .ZN(
      n_257_76_2725));
   NAND2_X1 i_257_76_2730 (.A1(n_257_76_2725), .A2(n_257_76_2491), .ZN(
      n_257_76_2726));
   NAND2_X1 i_257_76_2731 (.A1(n_257_314), .A2(n_257_422), .ZN(n_257_76_2727));
   NAND2_X1 i_257_76_2732 (.A1(n_257_76_2727), .A2(n_257_76_2444), .ZN(
      n_257_76_2728));
   NOR2_X1 i_257_76_2733 (.A1(n_257_76_2726), .A2(n_257_76_2728), .ZN(
      n_257_76_2729));
   NAND2_X1 i_257_76_2734 (.A1(n_257_76_2719), .A2(n_257_76_2729), .ZN(
      n_257_76_2730));
   NAND2_X1 i_257_76_2735 (.A1(n_257_276), .A2(n_257_423), .ZN(n_257_76_2731));
   NAND2_X1 i_257_76_2736 (.A1(n_257_76_2731), .A2(n_257_76_2495), .ZN(
      n_257_76_2732));
   INV_X1 i_257_76_2737 (.A(n_257_76_2732), .ZN(n_257_76_2733));
   NAND2_X1 i_257_76_2738 (.A1(n_257_76_2733), .A2(n_257_76_2494), .ZN(
      n_257_76_2734));
   NOR2_X1 i_257_76_2739 (.A1(n_257_76_2730), .A2(n_257_76_2734), .ZN(
      n_257_76_2735));
   NOR2_X1 i_257_76_2740 (.A1(n_257_76_2672), .A2(n_257_76_2554), .ZN(
      n_257_76_2736));
   NAND2_X1 i_257_76_2741 (.A1(n_257_76_2735), .A2(n_257_76_2736), .ZN(
      n_257_76_2737));
   INV_X1 i_257_76_2742 (.A(n_257_76_2451), .ZN(n_257_76_2738));
   NOR2_X1 i_257_76_2743 (.A1(n_257_76_2603), .A2(n_257_76_2738), .ZN(
      n_257_76_2739));
   NAND2_X1 i_257_76_2744 (.A1(n_257_76_2511), .A2(n_257_76_2498), .ZN(
      n_257_76_2740));
   NOR2_X1 i_257_76_2745 (.A1(n_257_76_2740), .A2(n_257_76_2441), .ZN(
      n_257_76_2741));
   NAND2_X1 i_257_76_2746 (.A1(n_257_76_2739), .A2(n_257_76_2741), .ZN(
      n_257_76_2742));
   NOR2_X1 i_257_76_2747 (.A1(n_257_76_2737), .A2(n_257_76_2742), .ZN(
      n_257_76_2743));
   NAND2_X1 i_257_76_2748 (.A1(n_257_76_2717), .A2(n_257_76_2743), .ZN(
      n_257_76_2744));
   NAND2_X1 i_257_76_2749 (.A1(n_257_76_2411), .A2(n_257_76_2566), .ZN(
      n_257_76_2745));
   NOR2_X1 i_257_76_2750 (.A1(n_257_76_2744), .A2(n_257_76_2745), .ZN(
      n_257_76_2746));
   NAND2_X1 i_257_76_2751 (.A1(n_257_382), .A2(n_257_76_2746), .ZN(n_257_76_2747));
   NAND2_X1 i_257_76_2752 (.A1(n_257_430), .A2(n_257_76_2427), .ZN(n_257_76_2748));
   INV_X1 i_257_76_2753 (.A(n_257_76_2748), .ZN(n_257_76_2749));
   NAND3_X1 i_257_76_2754 (.A1(n_257_76_2444), .A2(n_257_76_2491), .A3(
      n_257_76_2749), .ZN(n_257_76_2750));
   INV_X1 i_257_76_2755 (.A(n_257_76_2750), .ZN(n_257_76_2751));
   NAND4_X1 i_257_76_2756 (.A1(n_257_76_2494), .A2(n_257_117), .A3(n_257_76_2751), 
      .A4(n_257_76_2495), .ZN(n_257_76_2752));
   INV_X1 i_257_76_2757 (.A(n_257_76_2752), .ZN(n_257_76_2753));
   NAND3_X1 i_257_76_2758 (.A1(n_257_76_2540), .A2(n_257_76_2753), .A3(
      n_257_76_2621), .ZN(n_257_76_2754));
   NAND4_X1 i_257_76_2759 (.A1(n_257_76_2450), .A2(n_257_76_2451), .A3(
      n_257_76_2452), .A4(n_257_76_2510), .ZN(n_257_76_2755));
   NOR2_X1 i_257_76_2760 (.A1(n_257_76_2754), .A2(n_257_76_2755), .ZN(
      n_257_76_2756));
   INV_X1 i_257_76_2761 (.A(n_257_76_2455), .ZN(n_257_76_2757));
   NOR2_X1 i_257_76_2762 (.A1(n_257_76_2757), .A2(n_257_76_2710), .ZN(
      n_257_76_2758));
   NAND3_X1 i_257_76_2763 (.A1(n_257_76_2756), .A2(n_257_76_2758), .A3(
      n_257_76_2412), .ZN(n_257_76_2759));
   NOR2_X1 i_257_76_2764 (.A1(n_257_76_2759), .A2(n_257_76_2433), .ZN(
      n_257_76_2760));
   NAND2_X1 i_257_76_2765 (.A1(n_257_145), .A2(n_257_76_2760), .ZN(n_257_76_2761));
   NAND3_X1 i_257_76_2766 (.A1(n_257_76_2709), .A2(n_257_76_2747), .A3(
      n_257_76_2761), .ZN(n_257_76_2762));
   INV_X1 i_257_76_2767 (.A(n_257_76_2762), .ZN(n_257_76_2763));
   NAND2_X1 i_257_76_2768 (.A1(n_257_769), .A2(n_257_76_2414), .ZN(n_257_76_2764));
   NOR2_X1 i_257_76_2769 (.A1(n_257_76_17412), .A2(n_257_76_2764), .ZN(
      n_257_76_2765));
   NAND4_X1 i_257_76_2770 (.A1(n_257_76_2435), .A2(n_257_76_2436), .A3(
      n_257_76_2443), .A4(n_257_76_2765), .ZN(n_257_76_2766));
   INV_X1 i_257_76_2771 (.A(n_257_76_2766), .ZN(n_257_76_2767));
   NAND3_X1 i_257_76_2772 (.A1(n_257_76_2440), .A2(n_257_447), .A3(n_257_76_2434), 
      .ZN(n_257_76_2768));
   INV_X1 i_257_76_2773 (.A(n_257_76_2768), .ZN(n_257_76_2769));
   NAND4_X1 i_257_76_2774 (.A1(n_257_76_2767), .A2(n_257_76_2413), .A3(
      n_257_76_2769), .A4(n_257_76_2450), .ZN(n_257_76_2770));
   INV_X1 i_257_76_2775 (.A(n_257_76_2770), .ZN(n_257_76_2771));
   NAND2_X1 i_257_76_2776 (.A1(n_257_76_2412), .A2(n_257_76_2771), .ZN(
      n_257_76_2772));
   INV_X1 i_257_76_2777 (.A(n_257_76_2772), .ZN(n_257_76_2773));
   NAND2_X1 i_257_76_2778 (.A1(n_257_76_2411), .A2(n_257_76_2773), .ZN(
      n_257_76_2774));
   INV_X1 i_257_76_2779 (.A(n_257_76_2774), .ZN(n_257_76_2775));
   NAND3_X1 i_257_76_2780 (.A1(n_257_76_2510), .A2(n_257_79), .A3(n_257_76_2439), 
      .ZN(n_257_76_2776));
   NAND4_X1 i_257_76_2781 (.A1(n_257_76_2440), .A2(n_257_76_2434), .A3(
      n_257_76_2435), .A4(n_257_76_2436), .ZN(n_257_76_2777));
   NAND2_X1 i_257_76_2782 (.A1(n_257_431), .A2(n_257_76_2427), .ZN(n_257_76_2778));
   INV_X1 i_257_76_2783 (.A(n_257_76_2778), .ZN(n_257_76_2779));
   NAND3_X1 i_257_76_2784 (.A1(n_257_76_2444), .A2(n_257_76_2491), .A3(
      n_257_76_2779), .ZN(n_257_76_2780));
   INV_X1 i_257_76_2785 (.A(n_257_76_2780), .ZN(n_257_76_2781));
   NAND4_X1 i_257_76_2786 (.A1(n_257_76_2443), .A2(n_257_76_2494), .A3(
      n_257_76_2781), .A4(n_257_76_2495), .ZN(n_257_76_2782));
   NOR3_X1 i_257_76_2787 (.A1(n_257_76_2776), .A2(n_257_76_2777), .A3(
      n_257_76_2782), .ZN(n_257_76_2783));
   NAND4_X1 i_257_76_2788 (.A1(n_257_76_2783), .A2(n_257_76_2412), .A3(
      n_257_76_2455), .A4(n_257_76_2619), .ZN(n_257_76_2784));
   NOR2_X1 i_257_76_2789 (.A1(n_257_76_2784), .A2(n_257_76_2433), .ZN(
      n_257_76_2785));
   AOI22_X1 i_257_76_2790 (.A1(n_257_23), .A2(n_257_76_2775), .B1(n_257_107), 
      .B2(n_257_76_2785), .ZN(n_257_76_2786));
   NAND3_X1 i_257_76_2791 (.A1(n_257_76_2696), .A2(n_257_76_2763), .A3(
      n_257_76_2786), .ZN(n_257_76_2787));
   NAND3_X1 i_257_76_2792 (.A1(n_257_448), .A2(n_257_76_2443), .A3(
      n_257_76_18053), .ZN(n_257_76_2788));
   INV_X1 i_257_76_2793 (.A(n_257_76_2788), .ZN(n_257_76_2789));
   NAND4_X1 i_257_76_2794 (.A1(n_257_76_2438), .A2(n_257_76_2442), .A3(
      n_257_76_2789), .A4(n_257_76_2452), .ZN(n_257_76_2790));
   INV_X1 i_257_76_2795 (.A(n_257_76_2790), .ZN(n_257_76_2791));
   NAND3_X1 i_257_76_2796 (.A1(n_257_673), .A2(n_257_76_2413), .A3(n_257_76_2450), 
      .ZN(n_257_76_2792));
   INV_X1 i_257_76_2797 (.A(n_257_76_2792), .ZN(n_257_76_2793));
   NAND3_X1 i_257_76_2798 (.A1(n_257_76_2412), .A2(n_257_76_2791), .A3(
      n_257_76_2793), .ZN(n_257_76_2794));
   INV_X1 i_257_76_2799 (.A(n_257_76_2794), .ZN(n_257_76_2795));
   NAND2_X1 i_257_76_2800 (.A1(n_257_76_2795), .A2(n_257_76_2411), .ZN(
      n_257_76_2796));
   INV_X1 i_257_76_2801 (.A(n_257_76_2796), .ZN(n_257_76_2797));
   NAND2_X1 i_257_76_2802 (.A1(n_257_26), .A2(n_257_76_2797), .ZN(n_257_76_2798));
   NAND2_X1 i_257_76_2803 (.A1(n_257_76_2411), .A2(n_257_76_2412), .ZN(
      n_257_76_2799));
   NAND3_X1 i_257_76_2804 (.A1(n_257_76_2413), .A2(n_257_76_2516), .A3(n_257_236), 
      .ZN(n_257_76_2800));
   NOR2_X1 i_257_76_2805 (.A1(n_257_76_2800), .A2(n_257_76_2755), .ZN(
      n_257_76_2801));
   NAND2_X1 i_257_76_2806 (.A1(n_257_425), .A2(n_257_76_2427), .ZN(n_257_76_2802));
   NOR2_X1 i_257_76_2807 (.A1(n_257_76_2488), .A2(n_257_76_2802), .ZN(
      n_257_76_2803));
   NAND3_X1 i_257_76_2808 (.A1(n_257_76_2803), .A2(n_257_76_2444), .A3(
      n_257_76_2491), .ZN(n_257_76_2804));
   INV_X1 i_257_76_2809 (.A(n_257_76_2804), .ZN(n_257_76_2805));
   NAND3_X1 i_257_76_2810 (.A1(n_257_76_2805), .A2(n_257_76_2495), .A3(
      n_257_76_2506), .ZN(n_257_76_2806));
   INV_X1 i_257_76_2811 (.A(n_257_76_2806), .ZN(n_257_76_2807));
   NAND3_X1 i_257_76_2812 (.A1(n_257_76_2436), .A2(n_257_76_2443), .A3(
      n_257_76_2494), .ZN(n_257_76_2808));
   INV_X1 i_257_76_2813 (.A(n_257_76_2808), .ZN(n_257_76_2809));
   INV_X1 i_257_76_2814 (.A(n_257_76_2672), .ZN(n_257_76_2810));
   NAND3_X1 i_257_76_2815 (.A1(n_257_76_2807), .A2(n_257_76_2809), .A3(
      n_257_76_2810), .ZN(n_257_76_2811));
   NAND4_X1 i_257_76_2816 (.A1(n_257_76_2511), .A2(n_257_76_2498), .A3(
      n_257_76_2439), .A4(n_257_76_2440), .ZN(n_257_76_2812));
   NOR2_X1 i_257_76_2817 (.A1(n_257_76_2811), .A2(n_257_76_2812), .ZN(
      n_257_76_2813));
   NAND3_X1 i_257_76_2818 (.A1(n_257_76_2801), .A2(n_257_76_2600), .A3(
      n_257_76_2813), .ZN(n_257_76_2814));
   NOR2_X1 i_257_76_2819 (.A1(n_257_76_2799), .A2(n_257_76_2814), .ZN(
      n_257_76_2815));
   NAND2_X1 i_257_76_2820 (.A1(n_257_264), .A2(n_257_76_2815), .ZN(n_257_76_2816));
   INV_X1 i_257_76_2821 (.A(n_257_76_2728), .ZN(n_257_76_2817));
   INV_X1 i_257_76_2822 (.A(n_257_76_2491), .ZN(n_257_76_2818));
   NAND3_X1 i_257_76_2823 (.A1(n_257_76_2487), .A2(n_257_421), .A3(n_257_76_2427), 
      .ZN(n_257_76_2819));
   NOR2_X1 i_257_76_2824 (.A1(n_257_76_2818), .A2(n_257_76_2819), .ZN(
      n_257_76_2820));
   NAND4_X1 i_257_76_2825 (.A1(n_257_76_2817), .A2(n_257_76_2820), .A3(
      n_257_76_2506), .A4(n_257_76_2485), .ZN(n_257_76_2821));
   NAND3_X1 i_257_76_2826 (.A1(n_257_76_2494), .A2(n_257_76_2731), .A3(
      n_257_76_2495), .ZN(n_257_76_2822));
   NOR2_X1 i_257_76_2827 (.A1(n_257_76_2821), .A2(n_257_76_2822), .ZN(
      n_257_76_2823));
   NAND3_X1 i_257_76_2828 (.A1(n_257_353), .A2(n_257_76_2440), .A3(n_257_76_2434), 
      .ZN(n_257_76_2824));
   NOR2_X1 i_257_76_2829 (.A1(n_257_76_2824), .A2(n_257_76_2620), .ZN(
      n_257_76_2825));
   NAND3_X1 i_257_76_2830 (.A1(n_257_76_2511), .A2(n_257_76_2498), .A3(
      n_257_76_2439), .ZN(n_257_76_2826));
   INV_X1 i_257_76_2831 (.A(n_257_76_2826), .ZN(n_257_76_2827));
   NAND4_X1 i_257_76_2832 (.A1(n_257_76_2823), .A2(n_257_76_2825), .A3(
      n_257_76_2827), .A4(n_257_76_2516), .ZN(n_257_76_2828));
   NOR2_X1 i_257_76_2833 (.A1(n_257_76_2828), .A2(n_257_76_2503), .ZN(
      n_257_76_2829));
   NAND4_X1 i_257_76_2834 (.A1(n_257_76_2515), .A2(n_257_76_2602), .A3(
      n_257_76_2604), .A4(n_257_76_2413), .ZN(n_257_76_2830));
   NOR2_X1 i_257_76_2835 (.A1(n_257_76_2830), .A2(n_257_76_2599), .ZN(
      n_257_76_2831));
   NAND3_X1 i_257_76_2836 (.A1(n_257_76_2829), .A2(n_257_76_2411), .A3(
      n_257_76_2831), .ZN(n_257_76_2832));
   INV_X1 i_257_76_2837 (.A(n_257_76_2832), .ZN(n_257_76_2833));
   NAND2_X1 i_257_76_2838 (.A1(n_257_381), .A2(n_257_76_2833), .ZN(n_257_76_2834));
   NAND3_X1 i_257_76_2839 (.A1(n_257_76_2798), .A2(n_257_76_2816), .A3(
      n_257_76_2834), .ZN(n_257_76_2835));
   INV_X1 i_257_76_2840 (.A(n_257_76_2835), .ZN(n_257_76_2836));
   NAND4_X1 i_257_76_2841 (.A1(n_257_76_2413), .A2(n_257_76_2516), .A3(
      n_257_76_2450), .A4(n_257_76_2451), .ZN(n_257_76_2837));
   NAND4_X1 i_257_76_2842 (.A1(n_257_76_2540), .A2(n_257_76_2621), .A3(
      n_257_76_2452), .A4(n_257_76_2510), .ZN(n_257_76_2838));
   NOR2_X1 i_257_76_2843 (.A1(n_257_76_2837), .A2(n_257_76_2838), .ZN(
      n_257_76_2839));
   INV_X1 i_257_76_2844 (.A(n_257_569), .ZN(n_257_76_2840));
   NAND3_X1 i_257_76_2845 (.A1(n_257_76_2840), .A2(n_257_442), .A3(n_257_76_2414), 
      .ZN(n_257_76_2841));
   OAI21_X1 i_257_76_2846 (.A(n_257_76_2841), .B1(n_257_428), .B2(n_257_76_2415), 
      .ZN(n_257_76_2842));
   NAND2_X1 i_257_76_2847 (.A1(n_257_196), .A2(n_257_76_2842), .ZN(n_257_76_2843));
   INV_X1 i_257_76_2848 (.A(n_257_76_2843), .ZN(n_257_76_2844));
   NAND4_X1 i_257_76_2849 (.A1(n_257_76_2844), .A2(n_257_427), .A3(n_257_76_2444), 
      .A4(n_257_76_2491), .ZN(n_257_76_2845));
   INV_X1 i_257_76_2850 (.A(n_257_76_2845), .ZN(n_257_76_2846));
   NAND4_X1 i_257_76_2851 (.A1(n_257_76_2846), .A2(n_257_76_2498), .A3(
      n_257_76_2494), .A4(n_257_76_2495), .ZN(n_257_76_2847));
   INV_X1 i_257_76_2852 (.A(n_257_76_2847), .ZN(n_257_76_2848));
   NAND3_X1 i_257_76_2853 (.A1(n_257_76_2455), .A2(n_257_76_2501), .A3(
      n_257_76_2848), .ZN(n_257_76_2849));
   INV_X1 i_257_76_2854 (.A(n_257_76_2849), .ZN(n_257_76_2850));
   NAND3_X1 i_257_76_2855 (.A1(n_257_76_2839), .A2(n_257_76_2850), .A3(
      n_257_76_2412), .ZN(n_257_76_2851));
   NOR2_X1 i_257_76_2856 (.A1(n_257_76_2851), .A2(n_257_76_2433), .ZN(
      n_257_76_2852));
   NAND2_X1 i_257_76_2857 (.A1(n_257_224), .A2(n_257_76_2852), .ZN(n_257_76_2853));
   NAND4_X1 i_257_76_2858 (.A1(n_257_76_2442), .A2(n_257_76_2450), .A3(
      n_257_76_2451), .A4(n_257_76_2452), .ZN(n_257_76_2854));
   NAND2_X1 i_257_76_2859 (.A1(n_257_76_18053), .A2(n_257_456), .ZN(
      n_257_76_2855));
   INV_X1 i_257_76_2860 (.A(n_257_76_2855), .ZN(n_257_76_2856));
   NAND3_X1 i_257_76_2861 (.A1(n_257_76_2856), .A2(n_257_76_2443), .A3(
      n_257_76_2494), .ZN(n_257_76_2857));
   INV_X1 i_257_76_2862 (.A(n_257_76_2857), .ZN(n_257_76_2858));
   NAND2_X1 i_257_76_2863 (.A1(n_257_451), .A2(n_257_76_2434), .ZN(n_257_76_2859));
   INV_X1 i_257_76_2864 (.A(n_257_76_2859), .ZN(n_257_76_2860));
   NAND2_X1 i_257_76_2865 (.A1(n_257_76_2435), .A2(n_257_76_2436), .ZN(
      n_257_76_2861));
   INV_X1 i_257_76_2866 (.A(n_257_76_2861), .ZN(n_257_76_2862));
   NAND3_X1 i_257_76_2867 (.A1(n_257_76_2858), .A2(n_257_76_2860), .A3(
      n_257_76_2862), .ZN(n_257_76_2863));
   NOR2_X1 i_257_76_2868 (.A1(n_257_76_2854), .A2(n_257_76_2863), .ZN(
      n_257_76_2864));
   NAND3_X1 i_257_76_2869 (.A1(n_257_76_2864), .A2(n_257_76_2457), .A3(
      n_257_76_2412), .ZN(n_257_76_2865));
   NOR2_X1 i_257_76_2870 (.A1(n_257_76_2865), .A2(n_257_76_2433), .ZN(
      n_257_76_2866));
   NAND2_X1 i_257_76_2871 (.A1(n_257_434), .A2(n_257_76_2866), .ZN(n_257_76_2867));
   NAND3_X1 i_257_76_2872 (.A1(n_257_76_2455), .A2(n_257_76_2501), .A3(
      n_257_76_2515), .ZN(n_257_76_2868));
   NOR2_X1 i_257_76_2873 (.A1(n_257_76_2503), .A2(n_257_76_2868), .ZN(
      n_257_76_2869));
   NAND2_X1 i_257_76_2874 (.A1(n_257_424), .A2(n_257_76_2427), .ZN(n_257_76_2870));
   INV_X1 i_257_76_2875 (.A(n_257_76_2870), .ZN(n_257_76_2871));
   NAND3_X1 i_257_76_2876 (.A1(n_257_505), .A2(n_257_76_2487), .A3(n_257_76_2871), 
      .ZN(n_257_76_2872));
   INV_X1 i_257_76_2877 (.A(n_257_76_2872), .ZN(n_257_76_2873));
   NAND2_X1 i_257_76_2878 (.A1(n_257_76_2444), .A2(n_257_76_2491), .ZN(
      n_257_76_2874));
   INV_X1 i_257_76_2879 (.A(n_257_76_2874), .ZN(n_257_76_2875));
   NAND4_X1 i_257_76_2880 (.A1(n_257_76_2873), .A2(n_257_76_2495), .A3(
      n_257_76_2506), .A4(n_257_76_2875), .ZN(n_257_76_2876));
   NOR2_X1 i_257_76_2881 (.A1(n_257_76_2876), .A2(n_257_76_2808), .ZN(
      n_257_76_2877));
   NAND3_X1 i_257_76_2882 (.A1(n_257_76_2510), .A2(n_257_76_2511), .A3(
      n_257_76_2498), .ZN(n_257_76_2878));
   INV_X1 i_257_76_2883 (.A(n_257_76_2878), .ZN(n_257_76_2879));
   INV_X1 i_257_76_2884 (.A(n_257_76_2557), .ZN(n_257_76_2880));
   NAND3_X1 i_257_76_2885 (.A1(n_257_76_2877), .A2(n_257_76_2879), .A3(
      n_257_76_2880), .ZN(n_257_76_2881));
   NAND2_X1 i_257_76_2886 (.A1(n_257_76_2451), .A2(n_257_76_2452), .ZN(
      n_257_76_2882));
   INV_X1 i_257_76_2887 (.A(n_257_76_2882), .ZN(n_257_76_2883));
   NAND4_X1 i_257_76_2888 (.A1(n_257_76_2883), .A2(n_257_76_2413), .A3(
      n_257_76_2516), .A4(n_257_76_2450), .ZN(n_257_76_2884));
   NOR2_X1 i_257_76_2889 (.A1(n_257_76_2881), .A2(n_257_76_2884), .ZN(
      n_257_76_2885));
   NAND3_X1 i_257_76_2890 (.A1(n_257_76_2869), .A2(n_257_76_2411), .A3(
      n_257_76_2885), .ZN(n_257_76_2886));
   INV_X1 i_257_76_2891 (.A(n_257_76_2886), .ZN(n_257_76_2887));
   NAND2_X1 i_257_76_2892 (.A1(n_257_265), .A2(n_257_76_2887), .ZN(n_257_76_2888));
   NAND3_X1 i_257_76_2893 (.A1(n_257_76_2853), .A2(n_257_76_2867), .A3(
      n_257_76_2888), .ZN(n_257_76_2889));
   INV_X1 i_257_76_2894 (.A(n_257_76_2889), .ZN(n_257_76_2890));
   NAND4_X1 i_257_76_2895 (.A1(n_257_76_2602), .A2(n_257_76_2604), .A3(
      n_257_76_2413), .A4(n_257_76_2516), .ZN(n_257_76_2891));
   NAND4_X1 i_257_76_2896 (.A1(n_257_76_2731), .A2(n_257_76_2495), .A3(
      n_257_76_2506), .A4(n_257_76_2875), .ZN(n_257_76_2892));
   NOR2_X1 i_257_76_2897 (.A1(n_257_76_2892), .A2(n_257_76_2808), .ZN(
      n_257_76_2893));
   NAND3_X1 i_257_76_2898 (.A1(n_257_76_2487), .A2(n_257_422), .A3(n_257_76_2427), 
      .ZN(n_257_76_2894));
   INV_X1 i_257_76_2899 (.A(n_257_76_2894), .ZN(n_257_76_2895));
   NAND3_X1 i_257_76_2900 (.A1(n_257_76_2485), .A2(n_257_314), .A3(n_257_76_2895), 
      .ZN(n_257_76_2896));
   INV_X1 i_257_76_2901 (.A(n_257_76_2896), .ZN(n_257_76_2897));
   NAND3_X1 i_257_76_2902 (.A1(n_257_76_2511), .A2(n_257_76_2498), .A3(
      n_257_76_2897), .ZN(n_257_76_2898));
   INV_X1 i_257_76_2903 (.A(n_257_76_2898), .ZN(n_257_76_2899));
   NAND3_X1 i_257_76_2904 (.A1(n_257_76_2893), .A2(n_257_76_2899), .A3(
      n_257_76_2880), .ZN(n_257_76_2900));
   NOR2_X1 i_257_76_2905 (.A1(n_257_76_2891), .A2(n_257_76_2900), .ZN(
      n_257_76_2901));
   NAND3_X1 i_257_76_2906 (.A1(n_257_76_2411), .A2(n_257_76_2869), .A3(
      n_257_76_2901), .ZN(n_257_76_2902));
   INV_X1 i_257_76_2907 (.A(n_257_76_2902), .ZN(n_257_76_2903));
   NAND2_X1 i_257_76_2908 (.A1(n_257_342), .A2(n_257_76_2903), .ZN(n_257_76_2904));
   NAND2_X1 i_257_76_2909 (.A1(n_257_76_2516), .A2(n_257_76_2712), .ZN(
      n_257_76_2905));
   INV_X1 i_257_76_2910 (.A(n_257_76_2905), .ZN(n_257_76_2906));
   NAND2_X1 i_257_76_2911 (.A1(n_257_76_2906), .A2(n_257_76_2413), .ZN(
      n_257_76_2907));
   NOR2_X1 i_257_76_2912 (.A1(n_257_76_2907), .A2(n_257_76_2716), .ZN(
      n_257_76_2908));
   NAND3_X1 i_257_76_2913 (.A1(n_257_442), .A2(n_257_392), .A3(n_257_76_2414), 
      .ZN(n_257_76_2909));
   INV_X1 i_257_76_2914 (.A(n_257_76_2909), .ZN(n_257_76_2910));
   NAND2_X1 i_257_76_2915 (.A1(n_257_76_2910), .A2(n_257_484), .ZN(n_257_76_2911));
   INV_X1 i_257_76_2916 (.A(n_257_76_2911), .ZN(n_257_76_2912));
   NAND2_X1 i_257_76_2917 (.A1(n_257_76_2487), .A2(n_257_76_2912), .ZN(
      n_257_76_2913));
   NAND2_X1 i_257_76_2918 (.A1(n_257_420), .A2(n_257_895), .ZN(n_257_76_2914));
   INV_X1 i_257_76_2919 (.A(n_257_76_2914), .ZN(n_257_76_2915));
   NOR2_X1 i_257_76_2920 (.A1(n_257_76_2913), .A2(n_257_76_2915), .ZN(
      n_257_76_2916));
   NAND2_X1 i_257_76_2921 (.A1(n_257_76_2916), .A2(n_257_76_2491), .ZN(
      n_257_76_2917));
   NOR2_X1 i_257_76_2922 (.A1(n_257_76_2917), .A2(n_257_76_2728), .ZN(
      n_257_76_2918));
   NAND2_X1 i_257_76_2923 (.A1(n_257_76_2719), .A2(n_257_76_2918), .ZN(
      n_257_76_2919));
   NAND2_X1 i_257_76_2924 (.A1(n_257_76_2443), .A2(n_257_76_2494), .ZN(
      n_257_76_2920));
   INV_X1 i_257_76_2925 (.A(n_257_76_2920), .ZN(n_257_76_2921));
   NAND2_X1 i_257_76_2926 (.A1(n_257_76_2921), .A2(n_257_76_2733), .ZN(
      n_257_76_2922));
   NOR2_X1 i_257_76_2927 (.A1(n_257_76_2919), .A2(n_257_76_2922), .ZN(
      n_257_76_2923));
   NAND2_X1 i_257_76_2928 (.A1(n_257_76_2440), .A2(n_257_76_2434), .ZN(
      n_257_76_2924));
   NOR2_X1 i_257_76_2929 (.A1(n_257_76_2924), .A2(n_257_76_2861), .ZN(
      n_257_76_2925));
   NAND2_X1 i_257_76_2930 (.A1(n_257_76_2923), .A2(n_257_76_2925), .ZN(
      n_257_76_2926));
   INV_X1 i_257_76_2931 (.A(n_257_76_2450), .ZN(n_257_76_2927));
   NOR2_X1 i_257_76_2932 (.A1(n_257_76_2882), .A2(n_257_76_2927), .ZN(
      n_257_76_2928));
   NAND2_X1 i_257_76_2933 (.A1(n_257_76_2510), .A2(n_257_76_2511), .ZN(
      n_257_76_2929));
   NAND2_X1 i_257_76_2934 (.A1(n_257_76_2498), .A2(n_257_76_2439), .ZN(
      n_257_76_2930));
   NOR2_X1 i_257_76_2935 (.A1(n_257_76_2929), .A2(n_257_76_2930), .ZN(
      n_257_76_2931));
   NAND2_X1 i_257_76_2936 (.A1(n_257_76_2928), .A2(n_257_76_2931), .ZN(
      n_257_76_2932));
   NOR2_X1 i_257_76_2937 (.A1(n_257_76_2926), .A2(n_257_76_2932), .ZN(
      n_257_76_2933));
   NAND2_X1 i_257_76_2938 (.A1(n_257_76_2908), .A2(n_257_76_2933), .ZN(
      n_257_76_2934));
   NOR2_X1 i_257_76_2939 (.A1(n_257_76_2934), .A2(n_257_76_2745), .ZN(
      n_257_76_2935));
   NAND2_X1 i_257_76_2940 (.A1(n_257_12), .A2(n_257_76_2935), .ZN(n_257_76_2936));
   NAND2_X1 i_257_76_2941 (.A1(n_257_999), .A2(n_257_76_17964), .ZN(
      n_257_76_2937));
   NAND2_X1 i_257_76_2942 (.A1(n_257_76_2597), .A2(n_257_76_2937), .ZN(
      n_257_76_2938));
   NAND2_X1 i_257_76_2943 (.A1(n_257_673), .A2(n_257_76_17958), .ZN(
      n_257_76_2939));
   NAND2_X1 i_257_76_2944 (.A1(n_257_156), .A2(n_257_76_17331), .ZN(
      n_257_76_2940));
   NAND2_X1 i_257_76_2945 (.A1(n_257_76_2939), .A2(n_257_76_2940), .ZN(
      n_257_76_2941));
   NOR2_X1 i_257_76_2946 (.A1(n_257_76_2938), .A2(n_257_76_2941), .ZN(
      n_257_76_2942));
   NAND2_X1 i_257_76_2947 (.A1(n_257_76_2499), .A2(n_257_76_2847), .ZN(
      n_257_76_2943));
   INV_X1 i_257_76_2948 (.A(n_257_76_2943), .ZN(n_257_76_2944));
   NAND2_X1 i_257_76_2949 (.A1(n_257_967), .A2(n_257_442), .ZN(n_257_76_2945));
   INV_X1 i_257_76_2950 (.A(n_257_76_2945), .ZN(n_257_76_2946));
   NAND2_X1 i_257_76_2951 (.A1(n_257_441), .A2(n_257_76_2946), .ZN(n_257_76_2947));
   NAND2_X1 i_257_76_2952 (.A1(n_257_79), .A2(n_257_76_17932), .ZN(n_257_76_2948));
   NAND2_X1 i_257_76_2953 (.A1(n_257_76_2947), .A2(n_257_76_2948), .ZN(
      n_257_76_2949));
   NAND2_X1 i_257_76_2954 (.A1(n_257_833), .A2(n_257_442), .ZN(n_257_76_2950));
   INV_X1 i_257_76_2955 (.A(n_257_76_2950), .ZN(n_257_76_2951));
   NAND2_X1 i_257_76_2956 (.A1(n_257_446), .A2(n_257_76_2951), .ZN(n_257_76_2952));
   NAND2_X1 i_257_76_2957 (.A1(n_257_449), .A2(n_257_76_10424), .ZN(
      n_257_76_2953));
   NAND2_X1 i_257_76_2958 (.A1(n_257_76_2952), .A2(n_257_76_2953), .ZN(
      n_257_76_2954));
   NOR2_X1 i_257_76_2959 (.A1(n_257_76_2949), .A2(n_257_76_2954), .ZN(
      n_257_76_2955));
   NAND2_X1 i_257_76_2960 (.A1(n_257_76_2944), .A2(n_257_76_2955), .ZN(
      n_257_76_2956));
   NAND3_X1 i_257_76_2961 (.A1(n_257_435), .A2(n_257_705), .A3(n_257_442), 
      .ZN(n_257_76_2957));
   NAND2_X1 i_257_76_2962 (.A1(n_257_601), .A2(n_257_442), .ZN(n_257_76_2958));
   INV_X1 i_257_76_2963 (.A(n_257_76_2958), .ZN(n_257_76_2959));
   NAND2_X1 i_257_76_2964 (.A1(n_257_432), .A2(n_257_76_2959), .ZN(n_257_76_2960));
   NAND2_X1 i_257_76_2965 (.A1(n_257_76_2957), .A2(n_257_76_2960), .ZN(
      n_257_76_2961));
   INV_X1 i_257_76_2966 (.A(n_257_76_2961), .ZN(n_257_76_2962));
   NAND2_X1 i_257_76_2967 (.A1(n_257_76_2724), .A2(n_257_76_2548), .ZN(
      n_257_76_2963));
   NAND2_X1 i_257_76_2968 (.A1(n_257_76_2414), .A2(Small_Packet_Data_Size[4]), 
      .ZN(n_257_76_2964));
   INV_X1 i_257_76_2969 (.A(Small_Packet_Data_Size[4]), .ZN(n_257_76_2965));
   OAI21_X1 i_257_76_2970 (.A(n_257_76_2964), .B1(n_257_442), .B2(n_257_76_2965), 
      .ZN(n_257_76_2966));
   NAND2_X1 i_257_76_2971 (.A1(n_257_76_2911), .A2(n_257_76_2966), .ZN(
      n_257_76_2967));
   NOR2_X1 i_257_76_2972 (.A1(n_257_76_2963), .A2(n_257_76_2967), .ZN(
      n_257_76_2968));
   NAND2_X1 i_257_76_2973 (.A1(n_257_76_2962), .A2(n_257_76_2968), .ZN(
      n_257_76_2969));
   NAND2_X1 i_257_76_2974 (.A1(n_257_39), .A2(n_257_76_17918), .ZN(n_257_76_2970));
   NAND2_X1 i_257_76_2975 (.A1(n_257_76_2970), .A2(n_257_76_2872), .ZN(
      n_257_76_2971));
   NOR2_X1 i_257_76_2976 (.A1(n_257_76_2969), .A2(n_257_76_2971), .ZN(
      n_257_76_2972));
   AOI22_X1 i_257_76_2977 (.A1(n_257_438), .A2(n_257_76_6054), .B1(n_257_633), 
      .B2(n_257_76_17928), .ZN(n_257_76_2973));
   NAND2_X1 i_257_76_2978 (.A1(n_257_76_2972), .A2(n_257_76_2973), .ZN(
      n_257_76_2974));
   NAND2_X1 i_257_76_2979 (.A1(n_257_76_17903), .A2(n_257_865), .ZN(
      n_257_76_2975));
   NAND2_X1 i_257_76_2980 (.A1(n_257_76_2975), .A2(n_257_76_2896), .ZN(
      n_257_76_2976));
   INV_X1 i_257_76_2981 (.A(n_257_76_2976), .ZN(n_257_76_2977));
   NAND3_X1 i_257_76_2982 (.A1(n_257_439), .A2(n_257_903), .A3(n_257_442), 
      .ZN(n_257_76_2978));
   NAND2_X1 i_257_76_2983 (.A1(n_257_935), .A2(n_257_442), .ZN(n_257_76_2979));
   INV_X1 i_257_76_2984 (.A(n_257_76_2979), .ZN(n_257_76_2980));
   NAND2_X1 i_257_76_2985 (.A1(n_257_440), .A2(n_257_76_2980), .ZN(n_257_76_2981));
   NAND2_X1 i_257_76_2986 (.A1(n_257_76_2978), .A2(n_257_76_2981), .ZN(
      n_257_76_2982));
   INV_X1 i_257_76_2987 (.A(n_257_76_2982), .ZN(n_257_76_2983));
   NAND2_X1 i_257_76_2988 (.A1(n_257_76_2977), .A2(n_257_76_2983), .ZN(
      n_257_76_2984));
   NOR2_X1 i_257_76_2989 (.A1(n_257_76_2974), .A2(n_257_76_2984), .ZN(
      n_257_76_2985));
   AOI22_X1 i_257_76_2990 (.A1(n_257_737), .A2(n_257_76_17935), .B1(n_257_801), 
      .B2(n_257_76_17952), .ZN(n_257_76_2986));
   NAND2_X1 i_257_76_2991 (.A1(n_257_117), .A2(n_257_76_17925), .ZN(
      n_257_76_2987));
   NAND2_X1 i_257_76_2992 (.A1(n_257_76_2986), .A2(n_257_76_2987), .ZN(
      n_257_76_2988));
   NAND2_X1 i_257_76_2993 (.A1(n_257_442), .A2(n_257_769), .ZN(n_257_76_2989));
   INV_X1 i_257_76_2994 (.A(n_257_76_2989), .ZN(n_257_76_2990));
   NAND2_X1 i_257_76_2995 (.A1(n_257_447), .A2(n_257_76_2990), .ZN(n_257_76_2991));
   NAND2_X1 i_257_76_2996 (.A1(n_257_456), .A2(n_257_442), .ZN(n_257_76_2992));
   INV_X1 i_257_76_2997 (.A(n_257_76_2992), .ZN(n_257_76_2993));
   NAND2_X1 i_257_76_2998 (.A1(n_257_451), .A2(n_257_76_2993), .ZN(n_257_76_2994));
   NAND2_X1 i_257_76_2999 (.A1(n_257_76_2991), .A2(n_257_76_2994), .ZN(
      n_257_76_2995));
   NOR2_X1 i_257_76_3000 (.A1(n_257_76_2988), .A2(n_257_76_2995), .ZN(
      n_257_76_2996));
   NAND2_X1 i_257_76_3001 (.A1(n_257_76_2985), .A2(n_257_76_2996), .ZN(
      n_257_76_2997));
   NOR2_X1 i_257_76_3002 (.A1(n_257_76_2956), .A2(n_257_76_2997), .ZN(
      n_257_76_2998));
   NAND2_X1 i_257_76_3003 (.A1(n_257_76_2942), .A2(n_257_76_2998), .ZN(
      n_257_76_2999));
   INV_X1 i_257_76_3004 (.A(n_257_76_2999), .ZN(n_257_76_3000));
   INV_X1 i_257_76_3005 (.A(n_257_1031), .ZN(n_257_76_3001));
   OAI21_X1 i_257_76_3006 (.A(n_257_76_2828), .B1(n_257_76_3001), .B2(
      n_257_76_17968), .ZN(n_257_76_3002));
   INV_X1 i_257_76_3007 (.A(n_257_76_2814), .ZN(n_257_76_3003));
   NOR2_X1 i_257_76_3008 (.A1(n_257_76_3002), .A2(n_257_76_3003), .ZN(
      n_257_76_3004));
   NAND2_X1 i_257_76_3009 (.A1(n_257_76_3000), .A2(n_257_76_3004), .ZN(
      n_257_76_3005));
   NAND3_X1 i_257_76_3010 (.A1(n_257_76_2904), .A2(n_257_76_2936), .A3(
      n_257_76_3005), .ZN(n_257_76_3006));
   INV_X1 i_257_76_3011 (.A(n_257_76_3006), .ZN(n_257_76_3007));
   NAND3_X1 i_257_76_3012 (.A1(n_257_76_2836), .A2(n_257_76_2890), .A3(
      n_257_76_3007), .ZN(n_257_76_3008));
   NOR2_X1 i_257_76_3013 (.A1(n_257_76_2787), .A2(n_257_76_3008), .ZN(
      n_257_76_3009));
   NAND2_X1 i_257_76_3014 (.A1(n_257_76_2656), .A2(n_257_76_3009), .ZN(n_4));
   NAND2_X1 i_257_76_3015 (.A1(n_257_1000), .A2(n_257_444), .ZN(n_257_76_3010));
   NAND2_X1 i_257_76_3016 (.A1(n_257_441), .A2(n_257_968), .ZN(n_257_76_3011));
   INV_X1 i_257_76_3017 (.A(n_257_1064), .ZN(n_257_76_3012));
   NAND2_X1 i_257_76_3018 (.A1(n_257_442), .A2(n_257_76_3012), .ZN(n_257_76_3013));
   INV_X1 i_257_76_3019 (.A(n_257_936), .ZN(n_257_76_3014));
   NOR2_X1 i_257_76_3020 (.A1(n_257_76_3013), .A2(n_257_76_3014), .ZN(
      n_257_76_3015));
   NAND2_X1 i_257_76_3021 (.A1(n_257_440), .A2(n_257_76_3015), .ZN(n_257_76_3016));
   INV_X1 i_257_76_3022 (.A(n_257_76_3016), .ZN(n_257_76_3017));
   NAND2_X1 i_257_76_3023 (.A1(n_257_76_3011), .A2(n_257_76_3017), .ZN(
      n_257_76_3018));
   INV_X1 i_257_76_3024 (.A(n_257_76_3018), .ZN(n_257_76_3019));
   NAND2_X1 i_257_76_3025 (.A1(n_257_76_3010), .A2(n_257_76_3019), .ZN(
      n_257_76_3020));
   INV_X1 i_257_76_3026 (.A(n_257_76_3020), .ZN(n_257_76_3021));
   NAND2_X1 i_257_76_3027 (.A1(n_257_1032), .A2(n_257_443), .ZN(n_257_76_3022));
   NAND2_X1 i_257_76_3028 (.A1(n_257_76_3021), .A2(n_257_76_3022), .ZN(
      n_257_76_3023));
   INV_X1 i_257_76_3029 (.A(n_257_76_3023), .ZN(n_257_76_3024));
   NAND2_X1 i_257_76_3030 (.A1(n_257_17), .A2(n_257_76_3024), .ZN(n_257_76_3025));
   INV_X1 i_257_76_3031 (.A(n_257_76_3013), .ZN(n_257_76_3026));
   NAND2_X1 i_257_76_3032 (.A1(n_257_443), .A2(n_257_76_3026), .ZN(n_257_76_3027));
   INV_X1 i_257_76_3033 (.A(n_257_76_3027), .ZN(n_257_76_3028));
   NAND2_X1 i_257_76_3034 (.A1(n_257_1032), .A2(n_257_76_3028), .ZN(
      n_257_76_3029));
   INV_X1 i_257_76_3035 (.A(n_257_76_3029), .ZN(n_257_76_3030));
   NAND2_X1 i_257_76_3036 (.A1(n_257_76_18072), .A2(n_257_76_3030), .ZN(
      n_257_76_3031));
   INV_X1 i_257_76_3037 (.A(n_257_634), .ZN(n_257_76_3032));
   NAND2_X1 i_257_76_3038 (.A1(n_257_435), .A2(n_257_706), .ZN(n_257_76_3033));
   NAND3_X1 i_257_76_3039 (.A1(n_257_76_3033), .A2(n_257_450), .A3(n_257_76_3026), 
      .ZN(n_257_76_3034));
   NOR2_X1 i_257_76_3040 (.A1(n_257_76_3032), .A2(n_257_76_3034), .ZN(
      n_257_76_3035));
   NAND2_X1 i_257_76_3041 (.A1(n_257_440), .A2(n_257_936), .ZN(n_257_76_3036));
   NAND2_X1 i_257_76_3042 (.A1(n_257_438), .A2(n_257_1070), .ZN(n_257_76_3037));
   NAND2_X1 i_257_76_3043 (.A1(n_257_439), .A2(n_257_904), .ZN(n_257_76_3038));
   NAND4_X1 i_257_76_3044 (.A1(n_257_76_3035), .A2(n_257_76_3036), .A3(
      n_257_76_3037), .A4(n_257_76_3038), .ZN(n_257_76_3039));
   NAND2_X1 i_257_76_3045 (.A1(n_257_738), .A2(n_257_436), .ZN(n_257_76_3040));
   NAND2_X1 i_257_76_3046 (.A1(n_257_866), .A2(n_257_445), .ZN(n_257_76_3041));
   NAND2_X1 i_257_76_3047 (.A1(n_257_802), .A2(n_257_437), .ZN(n_257_76_3042));
   NAND3_X1 i_257_76_3048 (.A1(n_257_76_3040), .A2(n_257_76_3041), .A3(
      n_257_76_3042), .ZN(n_257_76_3043));
   NOR2_X1 i_257_76_3049 (.A1(n_257_76_3039), .A2(n_257_76_3043), .ZN(
      n_257_76_3044));
   NAND2_X1 i_257_76_3050 (.A1(n_257_674), .A2(n_257_448), .ZN(n_257_76_3045));
   NAND2_X1 i_257_76_3051 (.A1(n_257_446), .A2(n_257_834), .ZN(n_257_76_3046));
   NAND2_X1 i_257_76_3052 (.A1(n_257_449), .A2(n_257_1078), .ZN(n_257_76_3047));
   NAND2_X1 i_257_76_3053 (.A1(n_257_447), .A2(n_257_770), .ZN(n_257_76_3048));
   NAND3_X1 i_257_76_3054 (.A1(n_257_76_3046), .A2(n_257_76_3047), .A3(
      n_257_76_3048), .ZN(n_257_76_3049));
   INV_X1 i_257_76_3055 (.A(n_257_76_3049), .ZN(n_257_76_3050));
   NAND4_X1 i_257_76_3056 (.A1(n_257_76_3044), .A2(n_257_76_3045), .A3(
      n_257_76_3011), .A4(n_257_76_3050), .ZN(n_257_76_3051));
   INV_X1 i_257_76_3057 (.A(n_257_76_3051), .ZN(n_257_76_3052));
   NAND3_X1 i_257_76_3058 (.A1(n_257_76_3052), .A2(n_257_76_3022), .A3(
      n_257_76_3010), .ZN(n_257_76_3053));
   INV_X1 i_257_76_3059 (.A(n_257_76_3053), .ZN(n_257_76_3054));
   NAND2_X1 i_257_76_3060 (.A1(n_257_28), .A2(n_257_76_3054), .ZN(n_257_76_3055));
   NAND3_X1 i_257_76_3061 (.A1(n_257_76_3025), .A2(n_257_76_3031), .A3(
      n_257_76_3055), .ZN(n_257_76_3056));
   NAND3_X1 i_257_76_3062 (.A1(n_257_76_3041), .A2(n_257_446), .A3(n_257_76_3036), 
      .ZN(n_257_76_3057));
   INV_X1 i_257_76_3063 (.A(n_257_76_3057), .ZN(n_257_76_3058));
   NAND2_X1 i_257_76_3064 (.A1(n_257_76_3026), .A2(n_257_834), .ZN(n_257_76_3059));
   INV_X1 i_257_76_3065 (.A(n_257_76_3059), .ZN(n_257_76_3060));
   NAND3_X1 i_257_76_3066 (.A1(n_257_76_3037), .A2(n_257_76_3038), .A3(
      n_257_76_3060), .ZN(n_257_76_3061));
   INV_X1 i_257_76_3067 (.A(n_257_76_3061), .ZN(n_257_76_3062));
   NAND3_X1 i_257_76_3068 (.A1(n_257_76_3011), .A2(n_257_76_3058), .A3(
      n_257_76_3062), .ZN(n_257_76_3063));
   INV_X1 i_257_76_3069 (.A(n_257_76_3063), .ZN(n_257_76_3064));
   NAND2_X1 i_257_76_3070 (.A1(n_257_76_3010), .A2(n_257_76_3064), .ZN(
      n_257_76_3065));
   INV_X1 i_257_76_3071 (.A(n_257_76_3065), .ZN(n_257_76_3066));
   NAND2_X1 i_257_76_3072 (.A1(n_257_76_3066), .A2(n_257_76_3022), .ZN(
      n_257_76_3067));
   INV_X1 i_257_76_3073 (.A(n_257_76_3067), .ZN(n_257_76_3068));
   NAND2_X1 i_257_76_3074 (.A1(n_257_76_18070), .A2(n_257_76_3068), .ZN(
      n_257_76_3069));
   INV_X1 i_257_76_3075 (.A(n_257_76_3036), .ZN(n_257_76_3070));
   NAND3_X1 i_257_76_3076 (.A1(n_257_439), .A2(n_257_904), .A3(n_257_76_3026), 
      .ZN(n_257_76_3071));
   NOR2_X1 i_257_76_3077 (.A1(n_257_76_3070), .A2(n_257_76_3071), .ZN(
      n_257_76_3072));
   NAND2_X1 i_257_76_3078 (.A1(n_257_76_3011), .A2(n_257_76_3072), .ZN(
      n_257_76_3073));
   INV_X1 i_257_76_3079 (.A(n_257_76_3073), .ZN(n_257_76_3074));
   NAND2_X1 i_257_76_3080 (.A1(n_257_76_3010), .A2(n_257_76_3074), .ZN(
      n_257_76_3075));
   INV_X1 i_257_76_3081 (.A(n_257_76_3075), .ZN(n_257_76_3076));
   NAND2_X1 i_257_76_3082 (.A1(n_257_76_3076), .A2(n_257_76_3022), .ZN(
      n_257_76_3077));
   INV_X1 i_257_76_3083 (.A(n_257_76_3077), .ZN(n_257_76_3078));
   NAND2_X1 i_257_76_3084 (.A1(n_257_18), .A2(n_257_76_3078), .ZN(n_257_76_3079));
   INV_X1 i_257_76_3085 (.A(n_257_76_3010), .ZN(n_257_76_3080));
   NAND2_X1 i_257_76_3086 (.A1(n_257_634), .A2(n_257_450), .ZN(n_257_76_3081));
   NAND2_X1 i_257_76_3087 (.A1(n_257_40), .A2(n_257_433), .ZN(n_257_76_3082));
   NAND3_X1 i_257_76_3088 (.A1(n_257_76_3081), .A2(n_257_277), .A3(n_257_76_3082), 
      .ZN(n_257_76_3083));
   INV_X1 i_257_76_3089 (.A(n_257_76_3083), .ZN(n_257_76_3084));
   NAND2_X1 i_257_76_3090 (.A1(n_257_427), .A2(n_257_197), .ZN(n_257_76_3085));
   NAND2_X1 i_257_76_3091 (.A1(n_257_432), .A2(n_257_602), .ZN(n_257_76_3086));
   NAND2_X1 i_257_76_3092 (.A1(n_257_76_3033), .A2(n_257_76_3086), .ZN(
      n_257_76_3087));
   INV_X1 i_257_76_3093 (.A(n_257_76_3087), .ZN(n_257_76_3088));
   NAND2_X1 i_257_76_3094 (.A1(n_257_506), .A2(n_257_424), .ZN(n_257_76_3089));
   NAND2_X1 i_257_76_3095 (.A1(n_257_428), .A2(n_257_570), .ZN(n_257_76_3090));
   INV_X1 i_257_76_3096 (.A(n_257_76_3090), .ZN(n_257_76_3091));
   NAND2_X1 i_257_76_3097 (.A1(n_257_423), .A2(n_257_76_3026), .ZN(n_257_76_3092));
   NOR2_X1 i_257_76_3098 (.A1(n_257_76_3091), .A2(n_257_76_3092), .ZN(
      n_257_76_3093));
   NAND4_X1 i_257_76_3099 (.A1(n_257_76_3085), .A2(n_257_76_3088), .A3(
      n_257_76_3089), .A4(n_257_76_3093), .ZN(n_257_76_3094));
   INV_X1 i_257_76_3100 (.A(n_257_76_3094), .ZN(n_257_76_3095));
   NAND2_X1 i_257_76_3101 (.A1(n_257_538), .A2(n_257_426), .ZN(n_257_76_3096));
   NAND2_X1 i_257_76_3102 (.A1(n_257_118), .A2(n_257_430), .ZN(n_257_76_3097));
   NAND4_X1 i_257_76_3103 (.A1(n_257_76_3084), .A2(n_257_76_3095), .A3(
      n_257_76_3096), .A4(n_257_76_3097), .ZN(n_257_76_3098));
   INV_X1 i_257_76_3104 (.A(n_257_76_3098), .ZN(n_257_76_3099));
   NAND2_X1 i_257_76_3105 (.A1(n_257_76_3045), .A2(n_257_76_3099), .ZN(
      n_257_76_3100));
   NOR2_X1 i_257_76_3106 (.A1(n_257_76_3080), .A2(n_257_76_3100), .ZN(
      n_257_76_3101));
   NAND2_X1 i_257_76_3107 (.A1(n_257_237), .A2(n_257_425), .ZN(n_257_76_3102));
   NAND2_X1 i_257_76_3108 (.A1(n_257_157), .A2(n_257_429), .ZN(n_257_76_3103));
   NAND2_X1 i_257_76_3109 (.A1(n_257_80), .A2(n_257_431), .ZN(n_257_76_3104));
   NAND3_X1 i_257_76_3110 (.A1(n_257_76_3102), .A2(n_257_76_3103), .A3(
      n_257_76_3104), .ZN(n_257_76_3105));
   NAND2_X1 i_257_76_3111 (.A1(n_257_451), .A2(n_257_457), .ZN(n_257_76_3106));
   NAND3_X1 i_257_76_3112 (.A1(n_257_76_3106), .A2(n_257_76_3040), .A3(
      n_257_76_3041), .ZN(n_257_76_3107));
   INV_X1 i_257_76_3113 (.A(n_257_76_3107), .ZN(n_257_76_3108));
   NAND4_X1 i_257_76_3114 (.A1(n_257_76_3042), .A2(n_257_76_3036), .A3(
      n_257_76_3037), .A4(n_257_76_3038), .ZN(n_257_76_3109));
   INV_X1 i_257_76_3115 (.A(n_257_76_3109), .ZN(n_257_76_3110));
   NAND4_X1 i_257_76_3116 (.A1(n_257_76_3050), .A2(n_257_76_3108), .A3(
      n_257_76_3011), .A4(n_257_76_3110), .ZN(n_257_76_3111));
   NOR2_X1 i_257_76_3117 (.A1(n_257_76_3105), .A2(n_257_76_3111), .ZN(
      n_257_76_3112));
   NAND3_X1 i_257_76_3118 (.A1(n_257_76_3101), .A2(n_257_76_3022), .A3(
      n_257_76_3112), .ZN(n_257_76_3113));
   INV_X1 i_257_76_3119 (.A(n_257_76_3113), .ZN(n_257_76_3114));
   NAND2_X1 i_257_76_3120 (.A1(n_257_76_18066), .A2(n_257_76_3114), .ZN(
      n_257_76_3115));
   NAND3_X1 i_257_76_3121 (.A1(n_257_76_3069), .A2(n_257_76_3079), .A3(
      n_257_76_3115), .ZN(n_257_76_3116));
   NOR2_X1 i_257_76_3122 (.A1(n_257_76_3056), .A2(n_257_76_3116), .ZN(
      n_257_76_3117));
   NAND2_X1 i_257_76_3123 (.A1(n_257_968), .A2(n_257_76_3026), .ZN(n_257_76_3118));
   INV_X1 i_257_76_3124 (.A(n_257_76_3118), .ZN(n_257_76_3119));
   NAND2_X1 i_257_76_3125 (.A1(n_257_441), .A2(n_257_76_3119), .ZN(n_257_76_3120));
   INV_X1 i_257_76_3126 (.A(n_257_76_3120), .ZN(n_257_76_3121));
   NAND2_X1 i_257_76_3127 (.A1(n_257_76_3010), .A2(n_257_76_3121), .ZN(
      n_257_76_3122));
   INV_X1 i_257_76_3128 (.A(n_257_76_3122), .ZN(n_257_76_3123));
   NAND2_X1 i_257_76_3129 (.A1(n_257_76_3123), .A2(n_257_76_3022), .ZN(
      n_257_76_3124));
   INV_X1 i_257_76_3130 (.A(n_257_76_3124), .ZN(n_257_76_3125));
   NAND2_X1 i_257_76_3131 (.A1(n_257_76_18071), .A2(n_257_76_3125), .ZN(
      n_257_76_3126));
   INV_X1 i_257_76_3132 (.A(n_257_76_3022), .ZN(n_257_76_3127));
   NAND2_X1 i_257_76_3133 (.A1(n_257_76_3046), .A2(n_257_76_3048), .ZN(
      n_257_76_3128));
   INV_X1 i_257_76_3134 (.A(n_257_76_3128), .ZN(n_257_76_3129));
   NAND3_X1 i_257_76_3135 (.A1(n_257_435), .A2(n_257_706), .A3(n_257_76_3026), 
      .ZN(n_257_76_3130));
   INV_X1 i_257_76_3136 (.A(n_257_76_3130), .ZN(n_257_76_3131));
   NAND4_X1 i_257_76_3137 (.A1(n_257_76_3036), .A2(n_257_76_3037), .A3(
      n_257_76_3038), .A4(n_257_76_3131), .ZN(n_257_76_3132));
   INV_X1 i_257_76_3138 (.A(n_257_76_3132), .ZN(n_257_76_3133));
   INV_X1 i_257_76_3139 (.A(n_257_76_3043), .ZN(n_257_76_3134));
   NAND4_X1 i_257_76_3140 (.A1(n_257_76_3129), .A2(n_257_76_3133), .A3(
      n_257_76_3134), .A4(n_257_76_3011), .ZN(n_257_76_3135));
   INV_X1 i_257_76_3141 (.A(n_257_76_3135), .ZN(n_257_76_3136));
   NAND2_X1 i_257_76_3142 (.A1(n_257_76_3010), .A2(n_257_76_3136), .ZN(
      n_257_76_3137));
   NOR2_X1 i_257_76_3143 (.A1(n_257_76_3127), .A2(n_257_76_3137), .ZN(
      n_257_76_3138));
   NAND2_X1 i_257_76_3144 (.A1(n_257_76_18078), .A2(n_257_76_3138), .ZN(
      n_257_76_3139));
   NAND3_X1 i_257_76_3145 (.A1(n_257_76_3036), .A2(n_257_76_3037), .A3(
      n_257_76_3081), .ZN(n_257_76_3140));
   NAND3_X1 i_257_76_3146 (.A1(n_257_442), .A2(n_257_570), .A3(n_257_76_3012), 
      .ZN(n_257_76_3141));
   INV_X1 i_257_76_3147 (.A(n_257_76_3141), .ZN(n_257_76_3142));
   NAND2_X1 i_257_76_3148 (.A1(n_257_428), .A2(n_257_76_3142), .ZN(n_257_76_3143));
   INV_X1 i_257_76_3149 (.A(n_257_76_3143), .ZN(n_257_76_3144));
   NAND3_X1 i_257_76_3150 (.A1(n_257_76_3033), .A2(n_257_76_3086), .A3(
      n_257_76_3144), .ZN(n_257_76_3145));
   INV_X1 i_257_76_3151 (.A(n_257_76_3145), .ZN(n_257_76_3146));
   NAND3_X1 i_257_76_3152 (.A1(n_257_76_3038), .A2(n_257_76_3146), .A3(
      n_257_76_3082), .ZN(n_257_76_3147));
   NOR2_X1 i_257_76_3153 (.A1(n_257_76_3140), .A2(n_257_76_3147), .ZN(
      n_257_76_3148));
   NAND2_X1 i_257_76_3154 (.A1(n_257_76_3106), .A2(n_257_76_3097), .ZN(
      n_257_76_3149));
   INV_X1 i_257_76_3155 (.A(n_257_76_3149), .ZN(n_257_76_3150));
   NAND3_X1 i_257_76_3156 (.A1(n_257_76_3148), .A2(n_257_76_3150), .A3(
      n_257_76_3134), .ZN(n_257_76_3151));
   NAND4_X1 i_257_76_3157 (.A1(n_257_76_3011), .A2(n_257_76_3046), .A3(
      n_257_76_3047), .A4(n_257_76_3048), .ZN(n_257_76_3152));
   NOR2_X1 i_257_76_3158 (.A1(n_257_76_3151), .A2(n_257_76_3152), .ZN(
      n_257_76_3153));
   NAND3_X1 i_257_76_3159 (.A1(n_257_76_3045), .A2(n_257_76_3103), .A3(
      n_257_76_3104), .ZN(n_257_76_3154));
   INV_X1 i_257_76_3160 (.A(n_257_76_3154), .ZN(n_257_76_3155));
   NAND3_X1 i_257_76_3161 (.A1(n_257_76_3153), .A2(n_257_76_3155), .A3(
      n_257_76_3010), .ZN(n_257_76_3156));
   NOR2_X1 i_257_76_3162 (.A1(n_257_76_3156), .A2(n_257_76_3127), .ZN(
      n_257_76_3157));
   NAND2_X1 i_257_76_3163 (.A1(n_257_76_18074), .A2(n_257_76_3157), .ZN(
      n_257_76_3158));
   NAND3_X1 i_257_76_3164 (.A1(n_257_76_3126), .A2(n_257_76_3139), .A3(
      n_257_76_3158), .ZN(n_257_76_3159));
   NAND2_X1 i_257_76_3165 (.A1(n_257_442), .A2(n_257_1064), .ZN(n_257_76_3160));
   INV_X1 i_257_76_3166 (.A(n_257_76_3160), .ZN(n_257_76_3161));
   NAND2_X1 i_257_76_3167 (.A1(n_257_13), .A2(n_257_76_3161), .ZN(n_257_76_3162));
   INV_X1 i_257_76_3168 (.A(n_257_76_3011), .ZN(n_257_76_3163));
   NAND2_X1 i_257_76_3169 (.A1(n_257_76_3036), .A2(n_257_76_3037), .ZN(
      n_257_76_3164));
   INV_X1 i_257_76_3170 (.A(n_257_76_3164), .ZN(n_257_76_3165));
   NAND2_X1 i_257_76_3171 (.A1(n_257_445), .A2(n_257_76_3026), .ZN(n_257_76_3166));
   INV_X1 i_257_76_3172 (.A(n_257_76_3166), .ZN(n_257_76_3167));
   NAND3_X1 i_257_76_3173 (.A1(n_257_76_3038), .A2(n_257_866), .A3(n_257_76_3167), 
      .ZN(n_257_76_3168));
   INV_X1 i_257_76_3174 (.A(n_257_76_3168), .ZN(n_257_76_3169));
   NAND2_X1 i_257_76_3175 (.A1(n_257_76_3165), .A2(n_257_76_3169), .ZN(
      n_257_76_3170));
   NOR2_X1 i_257_76_3176 (.A1(n_257_76_3163), .A2(n_257_76_3170), .ZN(
      n_257_76_3171));
   NAND2_X1 i_257_76_3177 (.A1(n_257_76_3010), .A2(n_257_76_3171), .ZN(
      n_257_76_3172));
   INV_X1 i_257_76_3178 (.A(n_257_76_3172), .ZN(n_257_76_3173));
   NAND2_X1 i_257_76_3179 (.A1(n_257_76_3173), .A2(n_257_76_3022), .ZN(
      n_257_76_3174));
   INV_X1 i_257_76_3180 (.A(n_257_76_3174), .ZN(n_257_76_3175));
   NAND2_X1 i_257_76_3181 (.A1(n_257_76_18077), .A2(n_257_76_3175), .ZN(
      n_257_76_3176));
   NAND2_X1 i_257_76_3182 (.A1(n_257_76_3162), .A2(n_257_76_3176), .ZN(
      n_257_76_3177));
   NOR2_X1 i_257_76_3183 (.A1(n_257_76_3159), .A2(n_257_76_3177), .ZN(
      n_257_76_3178));
   NAND2_X1 i_257_76_3184 (.A1(n_257_76_3046), .A2(n_257_76_3047), .ZN(
      n_257_76_3179));
   INV_X1 i_257_76_3185 (.A(n_257_76_3179), .ZN(n_257_76_3180));
   NAND3_X1 i_257_76_3186 (.A1(n_257_76_3180), .A2(n_257_76_3104), .A3(
      n_257_76_3011), .ZN(n_257_76_3181));
   NAND3_X1 i_257_76_3187 (.A1(n_257_76_3036), .A2(n_257_76_3037), .A3(
      n_257_76_3038), .ZN(n_257_76_3182));
   INV_X1 i_257_76_3188 (.A(n_257_76_3182), .ZN(n_257_76_3183));
   NAND4_X1 i_257_76_3189 (.A1(n_257_76_3134), .A2(n_257_76_3048), .A3(
      n_257_76_3183), .A4(n_257_76_3106), .ZN(n_257_76_3184));
   NOR2_X1 i_257_76_3190 (.A1(n_257_76_3181), .A2(n_257_76_3184), .ZN(
      n_257_76_3185));
   NAND2_X1 i_257_76_3191 (.A1(n_257_426), .A2(n_257_76_3026), .ZN(n_257_76_3186));
   NOR2_X1 i_257_76_3192 (.A1(n_257_76_3091), .A2(n_257_76_3186), .ZN(
      n_257_76_3187));
   NAND3_X1 i_257_76_3193 (.A1(n_257_76_3187), .A2(n_257_76_3033), .A3(
      n_257_76_3086), .ZN(n_257_76_3188));
   INV_X1 i_257_76_3194 (.A(n_257_76_3188), .ZN(n_257_76_3189));
   NAND3_X1 i_257_76_3195 (.A1(n_257_76_3189), .A2(n_257_76_3082), .A3(
      n_257_76_3085), .ZN(n_257_76_3190));
   INV_X1 i_257_76_3196 (.A(n_257_76_3190), .ZN(n_257_76_3191));
   NAND2_X1 i_257_76_3197 (.A1(n_257_538), .A2(n_257_76_3081), .ZN(n_257_76_3192));
   INV_X1 i_257_76_3198 (.A(n_257_76_3192), .ZN(n_257_76_3193));
   NAND3_X1 i_257_76_3199 (.A1(n_257_76_3191), .A2(n_257_76_3193), .A3(
      n_257_76_3097), .ZN(n_257_76_3194));
   INV_X1 i_257_76_3200 (.A(n_257_76_3194), .ZN(n_257_76_3195));
   NAND3_X1 i_257_76_3201 (.A1(n_257_76_3195), .A2(n_257_76_3045), .A3(
      n_257_76_3103), .ZN(n_257_76_3196));
   INV_X1 i_257_76_3202 (.A(n_257_76_3196), .ZN(n_257_76_3197));
   NAND3_X1 i_257_76_3203 (.A1(n_257_76_3185), .A2(n_257_76_3197), .A3(
      n_257_76_3010), .ZN(n_257_76_3198));
   NOR2_X1 i_257_76_3204 (.A1(n_257_76_3198), .A2(n_257_76_3127), .ZN(
      n_257_76_3199));
   NAND2_X1 i_257_76_3205 (.A1(n_257_76_18076), .A2(n_257_76_3199), .ZN(
      n_257_76_3200));
   NAND3_X1 i_257_76_3206 (.A1(n_257_76_3041), .A2(n_257_76_3042), .A3(
      n_257_76_3036), .ZN(n_257_76_3201));
   INV_X1 i_257_76_3207 (.A(n_257_76_3201), .ZN(n_257_76_3202));
   NAND2_X1 i_257_76_3208 (.A1(n_257_436), .A2(n_257_76_3026), .ZN(n_257_76_3203));
   INV_X1 i_257_76_3209 (.A(n_257_76_3203), .ZN(n_257_76_3204));
   NAND4_X1 i_257_76_3210 (.A1(n_257_76_3037), .A2(n_257_76_3038), .A3(n_257_738), 
      .A4(n_257_76_3204), .ZN(n_257_76_3205));
   INV_X1 i_257_76_3211 (.A(n_257_76_3205), .ZN(n_257_76_3206));
   NAND4_X1 i_257_76_3212 (.A1(n_257_76_3129), .A2(n_257_76_3202), .A3(
      n_257_76_3206), .A4(n_257_76_3011), .ZN(n_257_76_3207));
   INV_X1 i_257_76_3213 (.A(n_257_76_3207), .ZN(n_257_76_3208));
   NAND2_X1 i_257_76_3214 (.A1(n_257_76_3010), .A2(n_257_76_3208), .ZN(
      n_257_76_3209));
   INV_X1 i_257_76_3215 (.A(n_257_76_3209), .ZN(n_257_76_3210));
   NAND2_X1 i_257_76_3216 (.A1(n_257_76_3210), .A2(n_257_76_3022), .ZN(
      n_257_76_3211));
   INV_X1 i_257_76_3217 (.A(n_257_76_3211), .ZN(n_257_76_3212));
   NAND2_X1 i_257_76_3218 (.A1(n_257_24), .A2(n_257_76_3212), .ZN(n_257_76_3213));
   NOR2_X1 i_257_76_3219 (.A1(n_257_76_3163), .A2(n_257_76_3179), .ZN(
      n_257_76_3214));
   NAND4_X1 i_257_76_3220 (.A1(n_257_76_3048), .A2(n_257_76_3106), .A3(
      n_257_76_3040), .A4(n_257_76_3041), .ZN(n_257_76_3215));
   INV_X1 i_257_76_3221 (.A(n_257_76_3215), .ZN(n_257_76_3216));
   INV_X1 i_257_76_3222 (.A(n_257_76_3033), .ZN(n_257_76_3217));
   INV_X1 i_257_76_3223 (.A(n_257_602), .ZN(n_257_76_3218));
   NOR2_X1 i_257_76_3224 (.A1(n_257_76_3013), .A2(n_257_76_3218), .ZN(
      n_257_76_3219));
   NAND2_X1 i_257_76_3225 (.A1(n_257_432), .A2(n_257_76_3219), .ZN(n_257_76_3220));
   NOR2_X1 i_257_76_3226 (.A1(n_257_76_3217), .A2(n_257_76_3220), .ZN(
      n_257_76_3221));
   NAND4_X1 i_257_76_3227 (.A1(n_257_76_3081), .A2(n_257_76_3038), .A3(
      n_257_76_3221), .A4(n_257_76_3082), .ZN(n_257_76_3222));
   NAND3_X1 i_257_76_3228 (.A1(n_257_76_3042), .A2(n_257_76_3036), .A3(
      n_257_76_3037), .ZN(n_257_76_3223));
   NOR2_X1 i_257_76_3229 (.A1(n_257_76_3222), .A2(n_257_76_3223), .ZN(
      n_257_76_3224));
   NAND4_X1 i_257_76_3230 (.A1(n_257_76_3214), .A2(n_257_76_3045), .A3(
      n_257_76_3216), .A4(n_257_76_3224), .ZN(n_257_76_3225));
   INV_X1 i_257_76_3231 (.A(n_257_76_3225), .ZN(n_257_76_3226));
   NAND3_X1 i_257_76_3232 (.A1(n_257_76_3226), .A2(n_257_76_3022), .A3(
      n_257_76_3010), .ZN(n_257_76_3227));
   INV_X1 i_257_76_3233 (.A(n_257_76_3227), .ZN(n_257_76_3228));
   NAND2_X1 i_257_76_3234 (.A1(n_257_68), .A2(n_257_76_3228), .ZN(n_257_76_3229));
   NAND3_X1 i_257_76_3235 (.A1(n_257_76_3200), .A2(n_257_76_3213), .A3(
      n_257_76_3229), .ZN(n_257_76_3230));
   NAND2_X1 i_257_76_3236 (.A1(n_257_437), .A2(n_257_76_3026), .ZN(n_257_76_3231));
   INV_X1 i_257_76_3237 (.A(n_257_76_3231), .ZN(n_257_76_3232));
   NAND4_X1 i_257_76_3238 (.A1(n_257_76_3037), .A2(n_257_76_3038), .A3(n_257_802), 
      .A4(n_257_76_3232), .ZN(n_257_76_3233));
   INV_X1 i_257_76_3239 (.A(n_257_76_3233), .ZN(n_257_76_3234));
   NAND2_X1 i_257_76_3240 (.A1(n_257_76_3041), .A2(n_257_76_3036), .ZN(
      n_257_76_3235));
   INV_X1 i_257_76_3241 (.A(n_257_76_3235), .ZN(n_257_76_3236));
   NAND4_X1 i_257_76_3242 (.A1(n_257_76_3011), .A2(n_257_76_3234), .A3(
      n_257_76_3046), .A4(n_257_76_3236), .ZN(n_257_76_3237));
   INV_X1 i_257_76_3243 (.A(n_257_76_3237), .ZN(n_257_76_3238));
   NAND2_X1 i_257_76_3244 (.A1(n_257_76_3010), .A2(n_257_76_3238), .ZN(
      n_257_76_3239));
   INV_X1 i_257_76_3245 (.A(n_257_76_3239), .ZN(n_257_76_3240));
   NAND2_X1 i_257_76_3246 (.A1(n_257_76_3240), .A2(n_257_76_3022), .ZN(
      n_257_76_3241));
   INV_X1 i_257_76_3247 (.A(n_257_76_3241), .ZN(n_257_76_3242));
   NAND2_X1 i_257_76_3248 (.A1(n_257_22), .A2(n_257_76_3242), .ZN(n_257_76_3243));
   NAND2_X1 i_257_76_3249 (.A1(n_257_444), .A2(n_257_76_3026), .ZN(n_257_76_3244));
   INV_X1 i_257_76_3250 (.A(n_257_76_3244), .ZN(n_257_76_3245));
   NAND2_X1 i_257_76_3251 (.A1(n_257_1000), .A2(n_257_76_3245), .ZN(
      n_257_76_3246));
   INV_X1 i_257_76_3252 (.A(n_257_76_3246), .ZN(n_257_76_3247));
   NAND2_X1 i_257_76_3253 (.A1(n_257_76_3022), .A2(n_257_76_3247), .ZN(
      n_257_76_3248));
   INV_X1 i_257_76_3254 (.A(n_257_76_3248), .ZN(n_257_76_3249));
   NAND2_X1 i_257_76_3255 (.A1(n_257_76_18075), .A2(n_257_76_3249), .ZN(
      n_257_76_3250));
   NAND2_X1 i_257_76_3256 (.A1(n_257_76_3243), .A2(n_257_76_3250), .ZN(
      n_257_76_3251));
   NOR2_X1 i_257_76_3257 (.A1(n_257_76_3230), .A2(n_257_76_3251), .ZN(
      n_257_76_3252));
   NAND3_X1 i_257_76_3258 (.A1(n_257_76_3117), .A2(n_257_76_3178), .A3(
      n_257_76_3252), .ZN(n_257_76_3253));
   INV_X1 i_257_76_3259 (.A(n_257_76_3253), .ZN(n_257_76_3254));
   NAND2_X1 i_257_76_3260 (.A1(n_257_433), .A2(n_257_76_3026), .ZN(n_257_76_3255));
   INV_X1 i_257_76_3261 (.A(n_257_76_3255), .ZN(n_257_76_3256));
   NAND3_X1 i_257_76_3262 (.A1(n_257_40), .A2(n_257_76_3033), .A3(n_257_76_3256), 
      .ZN(n_257_76_3257));
   INV_X1 i_257_76_3263 (.A(n_257_76_3257), .ZN(n_257_76_3258));
   NAND3_X1 i_257_76_3264 (.A1(n_257_76_3258), .A2(n_257_76_3081), .A3(
      n_257_76_3038), .ZN(n_257_76_3259));
   NOR2_X1 i_257_76_3265 (.A1(n_257_76_3223), .A2(n_257_76_3259), .ZN(
      n_257_76_3260));
   NAND4_X1 i_257_76_3266 (.A1(n_257_76_3214), .A2(n_257_76_3045), .A3(
      n_257_76_3216), .A4(n_257_76_3260), .ZN(n_257_76_3261));
   INV_X1 i_257_76_3267 (.A(n_257_76_3261), .ZN(n_257_76_3262));
   NAND3_X1 i_257_76_3268 (.A1(n_257_76_3262), .A2(n_257_76_3022), .A3(
      n_257_76_3010), .ZN(n_257_76_3263));
   INV_X1 i_257_76_3269 (.A(n_257_76_3263), .ZN(n_257_76_3264));
   NAND2_X1 i_257_76_3270 (.A1(n_257_76_18081), .A2(n_257_76_3264), .ZN(
      n_257_76_3265));
   NAND3_X1 i_257_76_3271 (.A1(n_257_76_3011), .A2(n_257_76_3046), .A3(
      n_257_76_3048), .ZN(n_257_76_3266));
   NAND3_X1 i_257_76_3272 (.A1(n_257_76_3042), .A2(n_257_449), .A3(n_257_76_3036), 
      .ZN(n_257_76_3267));
   INV_X1 i_257_76_3273 (.A(n_257_76_3267), .ZN(n_257_76_3268));
   NAND2_X1 i_257_76_3274 (.A1(n_257_76_3040), .A2(n_257_76_3041), .ZN(
      n_257_76_3269));
   INV_X1 i_257_76_3275 (.A(n_257_76_3269), .ZN(n_257_76_3270));
   NAND3_X1 i_257_76_3276 (.A1(n_257_76_3033), .A2(n_257_1078), .A3(
      n_257_76_3026), .ZN(n_257_76_3271));
   INV_X1 i_257_76_3277 (.A(n_257_76_3271), .ZN(n_257_76_3272));
   NAND3_X1 i_257_76_3278 (.A1(n_257_76_3037), .A2(n_257_76_3038), .A3(
      n_257_76_3272), .ZN(n_257_76_3273));
   INV_X1 i_257_76_3279 (.A(n_257_76_3273), .ZN(n_257_76_3274));
   NAND3_X1 i_257_76_3280 (.A1(n_257_76_3268), .A2(n_257_76_3270), .A3(
      n_257_76_3274), .ZN(n_257_76_3275));
   NOR2_X1 i_257_76_3281 (.A1(n_257_76_3266), .A2(n_257_76_3275), .ZN(
      n_257_76_3276));
   NAND3_X1 i_257_76_3282 (.A1(n_257_76_3276), .A2(n_257_76_3010), .A3(
      n_257_76_3045), .ZN(n_257_76_3277));
   NOR2_X1 i_257_76_3283 (.A1(n_257_76_3277), .A2(n_257_76_3127), .ZN(
      n_257_76_3278));
   NAND2_X1 i_257_76_3284 (.A1(n_257_27), .A2(n_257_76_3278), .ZN(n_257_76_3279));
   INV_X1 i_257_76_3285 (.A(n_257_76_3045), .ZN(n_257_76_3280));
   NAND3_X1 i_257_76_3286 (.A1(n_257_76_3104), .A2(n_257_157), .A3(n_257_76_3011), 
      .ZN(n_257_76_3281));
   NOR2_X1 i_257_76_3287 (.A1(n_257_76_3280), .A2(n_257_76_3281), .ZN(
      n_257_76_3282));
   NAND2_X1 i_257_76_3288 (.A1(n_257_429), .A2(n_257_76_3026), .ZN(n_257_76_3283));
   INV_X1 i_257_76_3289 (.A(n_257_76_3283), .ZN(n_257_76_3284));
   NAND3_X1 i_257_76_3290 (.A1(n_257_76_3033), .A2(n_257_76_3086), .A3(
      n_257_76_3284), .ZN(n_257_76_3285));
   INV_X1 i_257_76_3291 (.A(n_257_76_3285), .ZN(n_257_76_3286));
   NAND3_X1 i_257_76_3292 (.A1(n_257_76_3038), .A2(n_257_76_3286), .A3(
      n_257_76_3082), .ZN(n_257_76_3287));
   NAND2_X1 i_257_76_3293 (.A1(n_257_76_3037), .A2(n_257_76_3081), .ZN(
      n_257_76_3288));
   NOR2_X1 i_257_76_3294 (.A1(n_257_76_3287), .A2(n_257_76_3288), .ZN(
      n_257_76_3289));
   NAND2_X1 i_257_76_3295 (.A1(n_257_76_3097), .A2(n_257_76_3040), .ZN(
      n_257_76_3290));
   INV_X1 i_257_76_3296 (.A(n_257_76_3290), .ZN(n_257_76_3291));
   NAND3_X1 i_257_76_3297 (.A1(n_257_76_3289), .A2(n_257_76_3291), .A3(
      n_257_76_3202), .ZN(n_257_76_3292));
   NAND4_X1 i_257_76_3298 (.A1(n_257_76_3046), .A2(n_257_76_3047), .A3(
      n_257_76_3048), .A4(n_257_76_3106), .ZN(n_257_76_3293));
   NOR2_X1 i_257_76_3299 (.A1(n_257_76_3292), .A2(n_257_76_3293), .ZN(
      n_257_76_3294));
   NAND3_X1 i_257_76_3300 (.A1(n_257_76_3010), .A2(n_257_76_3282), .A3(
      n_257_76_3294), .ZN(n_257_76_3295));
   NOR2_X1 i_257_76_3301 (.A1(n_257_76_3295), .A2(n_257_76_3127), .ZN(
      n_257_76_3296));
   NAND2_X1 i_257_76_3302 (.A1(n_257_76_18061), .A2(n_257_76_3296), .ZN(
      n_257_76_3297));
   NAND3_X1 i_257_76_3303 (.A1(n_257_76_3265), .A2(n_257_76_3279), .A3(
      n_257_76_3297), .ZN(n_257_76_3298));
   INV_X1 i_257_76_3304 (.A(n_257_76_3298), .ZN(n_257_76_3299));
   NAND2_X1 i_257_76_3305 (.A1(n_257_1070), .A2(n_257_76_3026), .ZN(
      n_257_76_3300));
   INV_X1 i_257_76_3306 (.A(n_257_76_3300), .ZN(n_257_76_3301));
   NAND2_X1 i_257_76_3307 (.A1(n_257_438), .A2(n_257_76_3301), .ZN(n_257_76_3302));
   INV_X1 i_257_76_3308 (.A(n_257_76_3302), .ZN(n_257_76_3303));
   NAND3_X1 i_257_76_3309 (.A1(n_257_76_3303), .A2(n_257_76_3036), .A3(
      n_257_76_3038), .ZN(n_257_76_3304));
   INV_X1 i_257_76_3310 (.A(n_257_76_3304), .ZN(n_257_76_3305));
   NAND2_X1 i_257_76_3311 (.A1(n_257_76_3011), .A2(n_257_76_3305), .ZN(
      n_257_76_3306));
   INV_X1 i_257_76_3312 (.A(n_257_76_3306), .ZN(n_257_76_3307));
   NAND2_X1 i_257_76_3313 (.A1(n_257_76_3010), .A2(n_257_76_3307), .ZN(
      n_257_76_3308));
   INV_X1 i_257_76_3314 (.A(n_257_76_3308), .ZN(n_257_76_3309));
   NAND2_X1 i_257_76_3315 (.A1(n_257_76_3309), .A2(n_257_76_3022), .ZN(
      n_257_76_3310));
   INV_X1 i_257_76_3316 (.A(n_257_76_3310), .ZN(n_257_76_3311));
   NAND2_X1 i_257_76_3317 (.A1(n_257_76_18067), .A2(n_257_76_3311), .ZN(
      n_257_76_3312));
   NAND2_X1 i_257_76_3318 (.A1(n_257_354), .A2(n_257_421), .ZN(n_257_76_3313));
   NAND2_X1 i_257_76_3319 (.A1(n_257_76_3011), .A2(n_257_76_3313), .ZN(
      n_257_76_3314));
   INV_X1 i_257_76_3320 (.A(n_257_76_3314), .ZN(n_257_76_3315));
   NAND2_X1 i_257_76_3321 (.A1(n_257_76_3315), .A2(n_257_76_3104), .ZN(
      n_257_76_3316));
   NAND2_X1 i_257_76_3322 (.A1(n_257_76_3102), .A2(n_257_76_3103), .ZN(
      n_257_76_3317));
   NOR2_X1 i_257_76_3323 (.A1(n_257_76_3316), .A2(n_257_76_3317), .ZN(
      n_257_76_3318));
   NAND2_X1 i_257_76_3324 (.A1(n_257_76_3089), .A2(n_257_76_3033), .ZN(
      n_257_76_3319));
   INV_X1 i_257_76_3325 (.A(n_257_896), .ZN(n_257_76_3320));
   NOR2_X1 i_257_76_3326 (.A1(n_257_1064), .A2(n_257_76_3320), .ZN(n_257_76_3321));
   NAND2_X1 i_257_76_3327 (.A1(n_257_442), .A2(n_257_76_3321), .ZN(n_257_76_3322));
   INV_X1 i_257_76_3328 (.A(n_257_76_3322), .ZN(n_257_76_3323));
   NAND2_X1 i_257_76_3329 (.A1(n_257_420), .A2(n_257_76_3323), .ZN(n_257_76_3324));
   NOR2_X1 i_257_76_3330 (.A1(n_257_76_3324), .A2(n_257_76_3091), .ZN(
      n_257_76_3325));
   NAND2_X1 i_257_76_3331 (.A1(n_257_76_3325), .A2(n_257_76_3086), .ZN(
      n_257_76_3326));
   NOR2_X1 i_257_76_3332 (.A1(n_257_76_3319), .A2(n_257_76_3326), .ZN(
      n_257_76_3327));
   NAND2_X1 i_257_76_3333 (.A1(n_257_315), .A2(n_257_422), .ZN(n_257_76_3328));
   NAND2_X1 i_257_76_3334 (.A1(n_257_76_3085), .A2(n_257_76_3328), .ZN(
      n_257_76_3329));
   INV_X1 i_257_76_3335 (.A(n_257_76_3329), .ZN(n_257_76_3330));
   NAND2_X1 i_257_76_3336 (.A1(n_257_76_3327), .A2(n_257_76_3330), .ZN(
      n_257_76_3331));
   NAND2_X1 i_257_76_3337 (.A1(n_257_76_3038), .A2(n_257_76_3082), .ZN(
      n_257_76_3332));
   INV_X1 i_257_76_3338 (.A(n_257_76_3332), .ZN(n_257_76_3333));
   NAND2_X1 i_257_76_3339 (.A1(n_257_76_3333), .A2(n_257_76_3081), .ZN(
      n_257_76_3334));
   NOR2_X1 i_257_76_3340 (.A1(n_257_76_3331), .A2(n_257_76_3334), .ZN(
      n_257_76_3335));
   NAND2_X1 i_257_76_3341 (.A1(n_257_76_3041), .A2(n_257_76_3042), .ZN(
      n_257_76_3336));
   NOR2_X1 i_257_76_3342 (.A1(n_257_76_3336), .A2(n_257_76_3164), .ZN(
      n_257_76_3337));
   NAND2_X1 i_257_76_3343 (.A1(n_257_76_3335), .A2(n_257_76_3337), .ZN(
      n_257_76_3338));
   NAND2_X1 i_257_76_3344 (.A1(n_257_76_3048), .A2(n_257_76_3106), .ZN(
      n_257_76_3339));
   NOR2_X1 i_257_76_3345 (.A1(n_257_76_3179), .A2(n_257_76_3339), .ZN(
      n_257_76_3340));
   NAND2_X1 i_257_76_3346 (.A1(n_257_76_3096), .A2(n_257_76_3097), .ZN(
      n_257_76_3341));
   NAND2_X1 i_257_76_3347 (.A1(n_257_277), .A2(n_257_423), .ZN(n_257_76_3342));
   NAND2_X1 i_257_76_3348 (.A1(n_257_76_3342), .A2(n_257_76_3040), .ZN(
      n_257_76_3343));
   NOR2_X1 i_257_76_3349 (.A1(n_257_76_3341), .A2(n_257_76_3343), .ZN(
      n_257_76_3344));
   NAND2_X1 i_257_76_3350 (.A1(n_257_76_3340), .A2(n_257_76_3344), .ZN(
      n_257_76_3345));
   NOR2_X1 i_257_76_3351 (.A1(n_257_76_3338), .A2(n_257_76_3345), .ZN(
      n_257_76_3346));
   NAND2_X1 i_257_76_3352 (.A1(n_257_76_3318), .A2(n_257_76_3346), .ZN(
      n_257_76_3347));
   NAND2_X1 i_257_76_3353 (.A1(n_257_76_3010), .A2(n_257_76_3045), .ZN(
      n_257_76_3348));
   INV_X1 i_257_76_3354 (.A(n_257_76_3348), .ZN(n_257_76_3349));
   NAND2_X1 i_257_76_3355 (.A1(n_257_76_3349), .A2(n_257_76_3022), .ZN(
      n_257_76_3350));
   NOR2_X1 i_257_76_3356 (.A1(n_257_76_3347), .A2(n_257_76_3350), .ZN(
      n_257_76_3351));
   NAND2_X1 i_257_76_3357 (.A1(n_257_76_18073), .A2(n_257_76_3351), .ZN(
      n_257_76_3352));
   NAND2_X1 i_257_76_3358 (.A1(n_257_76_3104), .A2(n_257_76_3011), .ZN(
      n_257_76_3353));
   NOR2_X1 i_257_76_3359 (.A1(n_257_76_3280), .A2(n_257_76_3353), .ZN(
      n_257_76_3354));
   NAND2_X1 i_257_76_3360 (.A1(n_257_430), .A2(n_257_76_3026), .ZN(n_257_76_3355));
   INV_X1 i_257_76_3361 (.A(n_257_76_3355), .ZN(n_257_76_3356));
   NAND3_X1 i_257_76_3362 (.A1(n_257_76_3033), .A2(n_257_76_3086), .A3(
      n_257_76_3356), .ZN(n_257_76_3357));
   INV_X1 i_257_76_3363 (.A(n_257_76_3357), .ZN(n_257_76_3358));
   NAND4_X1 i_257_76_3364 (.A1(n_257_118), .A2(n_257_76_3038), .A3(n_257_76_3358), 
      .A4(n_257_76_3082), .ZN(n_257_76_3359));
   INV_X1 i_257_76_3365 (.A(n_257_76_3359), .ZN(n_257_76_3360));
   INV_X1 i_257_76_3366 (.A(n_257_76_3140), .ZN(n_257_76_3361));
   NAND3_X1 i_257_76_3367 (.A1(n_257_76_3134), .A2(n_257_76_3360), .A3(
      n_257_76_3361), .ZN(n_257_76_3362));
   NOR2_X1 i_257_76_3368 (.A1(n_257_76_3362), .A2(n_257_76_3293), .ZN(
      n_257_76_3363));
   NAND3_X1 i_257_76_3369 (.A1(n_257_76_3010), .A2(n_257_76_3354), .A3(
      n_257_76_3363), .ZN(n_257_76_3364));
   NOR2_X1 i_257_76_3370 (.A1(n_257_76_3364), .A2(n_257_76_3127), .ZN(
      n_257_76_3365));
   NAND2_X1 i_257_76_3371 (.A1(n_257_76_18068), .A2(n_257_76_3365), .ZN(
      n_257_76_3366));
   NAND3_X1 i_257_76_3372 (.A1(n_257_76_3312), .A2(n_257_76_3352), .A3(
      n_257_76_3366), .ZN(n_257_76_3367));
   INV_X1 i_257_76_3373 (.A(n_257_76_3367), .ZN(n_257_76_3368));
   INV_X1 i_257_76_3374 (.A(n_257_770), .ZN(n_257_76_3369));
   NOR2_X1 i_257_76_3375 (.A1(n_257_76_3013), .A2(n_257_76_3369), .ZN(
      n_257_76_3370));
   NAND4_X1 i_257_76_3376 (.A1(n_257_76_3036), .A2(n_257_76_3037), .A3(
      n_257_76_3038), .A4(n_257_76_3370), .ZN(n_257_76_3371));
   INV_X1 i_257_76_3377 (.A(n_257_76_3371), .ZN(n_257_76_3372));
   NAND3_X1 i_257_76_3378 (.A1(n_257_76_3041), .A2(n_257_76_3042), .A3(n_257_447), 
      .ZN(n_257_76_3373));
   INV_X1 i_257_76_3379 (.A(n_257_76_3373), .ZN(n_257_76_3374));
   NAND4_X1 i_257_76_3380 (.A1(n_257_76_3011), .A2(n_257_76_3372), .A3(
      n_257_76_3374), .A4(n_257_76_3046), .ZN(n_257_76_3375));
   INV_X1 i_257_76_3381 (.A(n_257_76_3375), .ZN(n_257_76_3376));
   NAND2_X1 i_257_76_3382 (.A1(n_257_76_3010), .A2(n_257_76_3376), .ZN(
      n_257_76_3377));
   INV_X1 i_257_76_3383 (.A(n_257_76_3377), .ZN(n_257_76_3378));
   NAND2_X1 i_257_76_3384 (.A1(n_257_76_3378), .A2(n_257_76_3022), .ZN(
      n_257_76_3379));
   INV_X1 i_257_76_3385 (.A(n_257_76_3379), .ZN(n_257_76_3380));
   NAND3_X1 i_257_76_3386 (.A1(n_257_76_3011), .A2(n_257_80), .A3(n_257_76_3046), 
      .ZN(n_257_76_3381));
   INV_X1 i_257_76_3387 (.A(n_257_76_3381), .ZN(n_257_76_3382));
   NAND4_X1 i_257_76_3388 (.A1(n_257_76_3041), .A2(n_257_76_3042), .A3(
      n_257_76_3036), .A4(n_257_76_3037), .ZN(n_257_76_3383));
   NAND2_X1 i_257_76_3389 (.A1(n_257_431), .A2(n_257_76_3026), .ZN(n_257_76_3384));
   INV_X1 i_257_76_3390 (.A(n_257_76_3384), .ZN(n_257_76_3385));
   NAND3_X1 i_257_76_3391 (.A1(n_257_76_3033), .A2(n_257_76_3086), .A3(
      n_257_76_3385), .ZN(n_257_76_3386));
   INV_X1 i_257_76_3392 (.A(n_257_76_3386), .ZN(n_257_76_3387));
   NAND4_X1 i_257_76_3393 (.A1(n_257_76_3081), .A2(n_257_76_3038), .A3(
      n_257_76_3387), .A4(n_257_76_3082), .ZN(n_257_76_3388));
   NOR2_X1 i_257_76_3394 (.A1(n_257_76_3383), .A2(n_257_76_3388), .ZN(
      n_257_76_3389));
   NAND4_X1 i_257_76_3395 (.A1(n_257_76_3047), .A2(n_257_76_3048), .A3(
      n_257_76_3106), .A4(n_257_76_3040), .ZN(n_257_76_3390));
   INV_X1 i_257_76_3396 (.A(n_257_76_3390), .ZN(n_257_76_3391));
   NAND4_X1 i_257_76_3397 (.A1(n_257_76_3382), .A2(n_257_76_3389), .A3(
      n_257_76_3045), .A4(n_257_76_3391), .ZN(n_257_76_3392));
   INV_X1 i_257_76_3398 (.A(n_257_76_3392), .ZN(n_257_76_3393));
   NAND3_X1 i_257_76_3399 (.A1(n_257_76_3393), .A2(n_257_76_3022), .A3(
      n_257_76_3010), .ZN(n_257_76_3394));
   INV_X1 i_257_76_3400 (.A(n_257_76_3394), .ZN(n_257_76_3395));
   AOI22_X1 i_257_76_3401 (.A1(n_257_76_18085), .A2(n_257_76_3380), .B1(
      n_257_76_18080), .B2(n_257_76_3395), .ZN(n_257_76_3396));
   NAND3_X1 i_257_76_3402 (.A1(n_257_76_3299), .A2(n_257_76_3368), .A3(
      n_257_76_3396), .ZN(n_257_76_3397));
   NAND3_X1 i_257_76_3403 (.A1(n_257_448), .A2(n_257_76_3038), .A3(
      n_257_76_18052), .ZN(n_257_76_3398));
   NOR2_X1 i_257_76_3404 (.A1(n_257_76_3398), .A2(n_257_76_3164), .ZN(
      n_257_76_3399));
   NAND3_X1 i_257_76_3405 (.A1(n_257_76_3399), .A2(n_257_76_3129), .A3(
      n_257_76_3134), .ZN(n_257_76_3400));
   NAND2_X1 i_257_76_3406 (.A1(n_257_674), .A2(n_257_76_3011), .ZN(n_257_76_3401));
   NOR2_X1 i_257_76_3407 (.A1(n_257_76_3400), .A2(n_257_76_3401), .ZN(
      n_257_76_3402));
   NAND2_X1 i_257_76_3408 (.A1(n_257_76_3402), .A2(n_257_76_3010), .ZN(
      n_257_76_3403));
   NOR2_X1 i_257_76_3409 (.A1(n_257_76_3403), .A2(n_257_76_3127), .ZN(
      n_257_76_3404));
   NAND2_X1 i_257_76_3410 (.A1(n_257_76_18079), .A2(n_257_76_3404), .ZN(
      n_257_76_3405));
   NAND2_X1 i_257_76_3411 (.A1(n_257_76_3022), .A2(n_257_76_3010), .ZN(
      n_257_76_3406));
   NAND2_X1 i_257_76_3412 (.A1(n_257_425), .A2(n_257_76_3026), .ZN(n_257_76_3407));
   NOR2_X1 i_257_76_3413 (.A1(n_257_76_3091), .A2(n_257_76_3407), .ZN(
      n_257_76_3408));
   NAND3_X1 i_257_76_3414 (.A1(n_257_76_3408), .A2(n_257_76_3033), .A3(
      n_257_76_3086), .ZN(n_257_76_3409));
   INV_X1 i_257_76_3415 (.A(n_257_76_3409), .ZN(n_257_76_3410));
   NAND4_X1 i_257_76_3416 (.A1(n_257_76_3410), .A2(n_257_76_3038), .A3(
      n_257_76_3082), .A4(n_257_76_3085), .ZN(n_257_76_3411));
   NOR2_X1 i_257_76_3417 (.A1(n_257_76_3411), .A2(n_257_76_3140), .ZN(
      n_257_76_3412));
   NAND3_X1 i_257_76_3418 (.A1(n_257_76_3048), .A2(n_257_76_3106), .A3(
      n_257_76_3096), .ZN(n_257_76_3413));
   INV_X1 i_257_76_3419 (.A(n_257_76_3413), .ZN(n_257_76_3414));
   NAND4_X1 i_257_76_3420 (.A1(n_257_76_3097), .A2(n_257_76_3040), .A3(
      n_257_76_3041), .A4(n_257_76_3042), .ZN(n_257_76_3415));
   INV_X1 i_257_76_3421 (.A(n_257_76_3415), .ZN(n_257_76_3416));
   NAND3_X1 i_257_76_3422 (.A1(n_257_76_3412), .A2(n_257_76_3414), .A3(
      n_257_76_3416), .ZN(n_257_76_3417));
   INV_X1 i_257_76_3423 (.A(n_257_76_3417), .ZN(n_257_76_3418));
   NAND2_X1 i_257_76_3424 (.A1(n_257_76_3045), .A2(n_257_76_3103), .ZN(
      n_257_76_3419));
   INV_X1 i_257_76_3425 (.A(n_257_76_3419), .ZN(n_257_76_3420));
   NAND4_X1 i_257_76_3426 (.A1(n_257_76_3180), .A2(n_257_76_3104), .A3(n_257_237), 
      .A4(n_257_76_3011), .ZN(n_257_76_3421));
   INV_X1 i_257_76_3427 (.A(n_257_76_3421), .ZN(n_257_76_3422));
   NAND3_X1 i_257_76_3428 (.A1(n_257_76_3418), .A2(n_257_76_3420), .A3(
      n_257_76_3422), .ZN(n_257_76_3423));
   NOR2_X1 i_257_76_3429 (.A1(n_257_76_3406), .A2(n_257_76_3423), .ZN(
      n_257_76_3424));
   NAND2_X1 i_257_76_3430 (.A1(n_257_76_18064), .A2(n_257_76_3424), .ZN(
      n_257_76_3425));
   NAND3_X1 i_257_76_3431 (.A1(n_257_76_3045), .A2(n_257_76_3102), .A3(
      n_257_76_3103), .ZN(n_257_76_3426));
   INV_X1 i_257_76_3432 (.A(n_257_76_3339), .ZN(n_257_76_3427));
   NAND3_X1 i_257_76_3433 (.A1(n_257_76_3180), .A2(n_257_76_3427), .A3(
      n_257_76_3011), .ZN(n_257_76_3428));
   NOR2_X1 i_257_76_3434 (.A1(n_257_76_3426), .A2(n_257_76_3428), .ZN(
      n_257_76_3429));
   NAND3_X1 i_257_76_3435 (.A1(n_257_76_3040), .A2(n_257_76_3041), .A3(n_257_354), 
      .ZN(n_257_76_3430));
   NOR2_X1 i_257_76_3436 (.A1(n_257_76_3430), .A2(n_257_76_3223), .ZN(
      n_257_76_3431));
   NAND2_X1 i_257_76_3437 (.A1(n_257_421), .A2(n_257_76_3026), .ZN(n_257_76_3432));
   NOR2_X1 i_257_76_3438 (.A1(n_257_76_3091), .A2(n_257_76_3432), .ZN(
      n_257_76_3433));
   NAND3_X1 i_257_76_3439 (.A1(n_257_76_3433), .A2(n_257_76_3033), .A3(
      n_257_76_3086), .ZN(n_257_76_3434));
   INV_X1 i_257_76_3440 (.A(n_257_76_3434), .ZN(n_257_76_3435));
   NAND4_X1 i_257_76_3441 (.A1(n_257_76_3435), .A2(n_257_76_3085), .A3(
      n_257_76_3328), .A4(n_257_76_3089), .ZN(n_257_76_3436));
   NAND3_X1 i_257_76_3442 (.A1(n_257_76_3081), .A2(n_257_76_3038), .A3(
      n_257_76_3082), .ZN(n_257_76_3437));
   NOR2_X1 i_257_76_3443 (.A1(n_257_76_3436), .A2(n_257_76_3437), .ZN(
      n_257_76_3438));
   NAND3_X1 i_257_76_3444 (.A1(n_257_76_3096), .A2(n_257_76_3097), .A3(
      n_257_76_3342), .ZN(n_257_76_3439));
   INV_X1 i_257_76_3445 (.A(n_257_76_3439), .ZN(n_257_76_3440));
   NAND4_X1 i_257_76_3446 (.A1(n_257_76_3431), .A2(n_257_76_3438), .A3(
      n_257_76_3440), .A4(n_257_76_3104), .ZN(n_257_76_3441));
   INV_X1 i_257_76_3447 (.A(n_257_76_3441), .ZN(n_257_76_3442));
   NAND4_X1 i_257_76_3448 (.A1(n_257_76_3429), .A2(n_257_76_3022), .A3(
      n_257_76_3442), .A4(n_257_76_3010), .ZN(n_257_76_3443));
   INV_X1 i_257_76_3449 (.A(n_257_76_3443), .ZN(n_257_76_3444));
   NAND2_X1 i_257_76_3450 (.A1(n_257_76_18082), .A2(n_257_76_3444), .ZN(
      n_257_76_3445));
   NAND3_X1 i_257_76_3451 (.A1(n_257_76_3405), .A2(n_257_76_3425), .A3(
      n_257_76_3445), .ZN(n_257_76_3446));
   INV_X1 i_257_76_3452 (.A(n_257_76_3446), .ZN(n_257_76_3447));
   NAND3_X1 i_257_76_3453 (.A1(n_257_76_3038), .A2(n_257_76_3082), .A3(
      n_257_76_3033), .ZN(n_257_76_3448));
   NOR2_X1 i_257_76_3454 (.A1(n_257_76_3448), .A2(n_257_76_3288), .ZN(
      n_257_76_3449));
   NAND3_X1 i_257_76_3455 (.A1(n_257_76_3097), .A2(n_257_76_3040), .A3(
      n_257_76_3041), .ZN(n_257_76_3450));
   INV_X1 i_257_76_3456 (.A(n_257_76_3450), .ZN(n_257_76_3451));
   INV_X1 i_257_76_3457 (.A(n_257_570), .ZN(n_257_76_3452));
   NAND3_X1 i_257_76_3458 (.A1(n_257_76_3452), .A2(n_257_442), .A3(n_257_76_3012), 
      .ZN(n_257_76_3453));
   OAI21_X1 i_257_76_3459 (.A(n_257_76_3453), .B1(n_257_428), .B2(n_257_76_3013), 
      .ZN(n_257_76_3454));
   NAND4_X1 i_257_76_3460 (.A1(n_257_427), .A2(n_257_197), .A3(n_257_76_3086), 
      .A4(n_257_76_3454), .ZN(n_257_76_3455));
   INV_X1 i_257_76_3461 (.A(n_257_76_3455), .ZN(n_257_76_3456));
   NAND3_X1 i_257_76_3462 (.A1(n_257_76_3042), .A2(n_257_76_3456), .A3(
      n_257_76_3036), .ZN(n_257_76_3457));
   INV_X1 i_257_76_3463 (.A(n_257_76_3457), .ZN(n_257_76_3458));
   NAND3_X1 i_257_76_3464 (.A1(n_257_76_3449), .A2(n_257_76_3451), .A3(
      n_257_76_3458), .ZN(n_257_76_3459));
   NOR2_X1 i_257_76_3465 (.A1(n_257_76_3459), .A2(n_257_76_3428), .ZN(
      n_257_76_3460));
   NAND3_X1 i_257_76_3466 (.A1(n_257_76_3460), .A2(n_257_76_3155), .A3(
      n_257_76_3010), .ZN(n_257_76_3461));
   NOR2_X1 i_257_76_3467 (.A1(n_257_76_3461), .A2(n_257_76_3127), .ZN(
      n_257_76_3462));
   NAND2_X1 i_257_76_3468 (.A1(n_257_76_18065), .A2(n_257_76_3462), .ZN(
      n_257_76_3463));
   NAND3_X1 i_257_76_3469 (.A1(n_257_451), .A2(n_257_76_3036), .A3(n_257_76_3037), 
      .ZN(n_257_76_3464));
   NAND3_X1 i_257_76_3470 (.A1(n_257_457), .A2(n_257_76_3033), .A3(n_257_76_3026), 
      .ZN(n_257_76_3465));
   INV_X1 i_257_76_3471 (.A(n_257_76_3465), .ZN(n_257_76_3466));
   NAND3_X1 i_257_76_3472 (.A1(n_257_76_3081), .A2(n_257_76_3038), .A3(
      n_257_76_3466), .ZN(n_257_76_3467));
   NOR3_X1 i_257_76_3473 (.A1(n_257_76_3043), .A2(n_257_76_3464), .A3(
      n_257_76_3467), .ZN(n_257_76_3468));
   NOR2_X1 i_257_76_3474 (.A1(n_257_76_3049), .A2(n_257_76_3163), .ZN(
      n_257_76_3469));
   NAND3_X1 i_257_76_3475 (.A1(n_257_76_3468), .A2(n_257_76_3045), .A3(
      n_257_76_3469), .ZN(n_257_76_3470));
   INV_X1 i_257_76_3476 (.A(n_257_76_3470), .ZN(n_257_76_3471));
   NAND3_X1 i_257_76_3477 (.A1(n_257_76_3471), .A2(n_257_76_3022), .A3(
      n_257_76_3010), .ZN(n_257_76_3472));
   INV_X1 i_257_76_3478 (.A(n_257_76_3472), .ZN(n_257_76_3473));
   NAND2_X1 i_257_76_3479 (.A1(n_257_76_18063), .A2(n_257_76_3473), .ZN(
      n_257_76_3474));
   NAND4_X1 i_257_76_3480 (.A1(n_257_76_3038), .A2(n_257_76_3082), .A3(
      n_257_76_3085), .A4(n_257_76_3033), .ZN(n_257_76_3475));
   NAND3_X1 i_257_76_3481 (.A1(n_257_76_3090), .A2(n_257_424), .A3(n_257_76_3026), 
      .ZN(n_257_76_3476));
   INV_X1 i_257_76_3482 (.A(n_257_76_3476), .ZN(n_257_76_3477));
   NAND3_X1 i_257_76_3483 (.A1(n_257_76_3477), .A2(n_257_506), .A3(n_257_76_3086), 
      .ZN(n_257_76_3478));
   INV_X1 i_257_76_3484 (.A(n_257_76_3478), .ZN(n_257_76_3479));
   NAND3_X1 i_257_76_3485 (.A1(n_257_76_3037), .A2(n_257_76_3081), .A3(
      n_257_76_3479), .ZN(n_257_76_3480));
   NOR2_X1 i_257_76_3486 (.A1(n_257_76_3475), .A2(n_257_76_3480), .ZN(
      n_257_76_3481));
   NAND3_X1 i_257_76_3487 (.A1(n_257_76_3106), .A2(n_257_76_3096), .A3(
      n_257_76_3097), .ZN(n_257_76_3482));
   INV_X1 i_257_76_3488 (.A(n_257_76_3482), .ZN(n_257_76_3483));
   NAND4_X1 i_257_76_3489 (.A1(n_257_76_3040), .A2(n_257_76_3041), .A3(
      n_257_76_3042), .A4(n_257_76_3036), .ZN(n_257_76_3484));
   INV_X1 i_257_76_3490 (.A(n_257_76_3484), .ZN(n_257_76_3485));
   NAND4_X1 i_257_76_3491 (.A1(n_257_76_3481), .A2(n_257_76_3050), .A3(
      n_257_76_3483), .A4(n_257_76_3485), .ZN(n_257_76_3486));
   NAND3_X1 i_257_76_3492 (.A1(n_257_76_3103), .A2(n_257_76_3104), .A3(
      n_257_76_3011), .ZN(n_257_76_3487));
   NOR2_X1 i_257_76_3493 (.A1(n_257_76_3486), .A2(n_257_76_3487), .ZN(
      n_257_76_3488));
   NAND2_X1 i_257_76_3494 (.A1(n_257_76_3045), .A2(n_257_76_3102), .ZN(
      n_257_76_3489));
   INV_X1 i_257_76_3495 (.A(n_257_76_3489), .ZN(n_257_76_3490));
   NAND2_X1 i_257_76_3496 (.A1(n_257_76_3010), .A2(n_257_76_3490), .ZN(
      n_257_76_3491));
   INV_X1 i_257_76_3497 (.A(n_257_76_3491), .ZN(n_257_76_3492));
   NAND3_X1 i_257_76_3498 (.A1(n_257_76_3488), .A2(n_257_76_3492), .A3(
      n_257_76_3022), .ZN(n_257_76_3493));
   INV_X1 i_257_76_3499 (.A(n_257_76_3493), .ZN(n_257_76_3494));
   NAND2_X1 i_257_76_3500 (.A1(n_257_76_18062), .A2(n_257_76_3494), .ZN(
      n_257_76_3495));
   NAND3_X1 i_257_76_3501 (.A1(n_257_76_3463), .A2(n_257_76_3474), .A3(
      n_257_76_3495), .ZN(n_257_76_3496));
   INV_X1 i_257_76_3502 (.A(n_257_76_3496), .ZN(n_257_76_3497));
   NOR2_X1 i_257_76_3503 (.A1(n_257_76_3140), .A2(n_257_76_3475), .ZN(
      n_257_76_3498));
   NAND3_X1 i_257_76_3504 (.A1(n_257_76_3090), .A2(n_257_422), .A3(n_257_76_3026), 
      .ZN(n_257_76_3499));
   INV_X1 i_257_76_3505 (.A(n_257_76_3499), .ZN(n_257_76_3500));
   NAND4_X1 i_257_76_3506 (.A1(n_257_76_3089), .A2(n_257_315), .A3(n_257_76_3086), 
      .A4(n_257_76_3500), .ZN(n_257_76_3501));
   INV_X1 i_257_76_3507 (.A(n_257_76_3501), .ZN(n_257_76_3502));
   NAND4_X1 i_257_76_3508 (.A1(n_257_76_3106), .A2(n_257_76_3502), .A3(
      n_257_76_3096), .A4(n_257_76_3097), .ZN(n_257_76_3503));
   INV_X1 i_257_76_3509 (.A(n_257_76_3503), .ZN(n_257_76_3504));
   NAND4_X1 i_257_76_3510 (.A1(n_257_76_3342), .A2(n_257_76_3040), .A3(
      n_257_76_3041), .A4(n_257_76_3042), .ZN(n_257_76_3505));
   INV_X1 i_257_76_3511 (.A(n_257_76_3505), .ZN(n_257_76_3506));
   NAND4_X1 i_257_76_3512 (.A1(n_257_76_3498), .A2(n_257_76_3504), .A3(
      n_257_76_3050), .A4(n_257_76_3506), .ZN(n_257_76_3507));
   NOR2_X1 i_257_76_3513 (.A1(n_257_76_3507), .A2(n_257_76_3487), .ZN(
      n_257_76_3508));
   NAND3_X1 i_257_76_3514 (.A1(n_257_76_3508), .A2(n_257_76_3492), .A3(
      n_257_76_3022), .ZN(n_257_76_3509));
   INV_X1 i_257_76_3515 (.A(n_257_76_3509), .ZN(n_257_76_3510));
   NAND2_X1 i_257_76_3516 (.A1(n_257_342), .A2(n_257_76_3510), .ZN(n_257_76_3511));
   NAND2_X1 i_257_76_3517 (.A1(n_257_76_3081), .A2(n_257_76_3038), .ZN(
      n_257_76_3512));
   NAND2_X1 i_257_76_3518 (.A1(n_257_76_3082), .A2(n_257_76_3085), .ZN(
      n_257_76_3513));
   NOR2_X1 i_257_76_3519 (.A1(n_257_76_3512), .A2(n_257_76_3513), .ZN(
      n_257_76_3514));
   NAND2_X1 i_257_76_3520 (.A1(n_257_420), .A2(n_257_896), .ZN(n_257_76_3515));
   INV_X1 i_257_76_3521 (.A(n_257_76_3515), .ZN(n_257_76_3516));
   NAND3_X1 i_257_76_3522 (.A1(n_257_484), .A2(n_257_76_3026), .A3(n_257_393), 
      .ZN(n_257_76_3517));
   INV_X1 i_257_76_3523 (.A(n_257_76_3517), .ZN(n_257_76_3518));
   NAND2_X1 i_257_76_3524 (.A1(n_257_76_3090), .A2(n_257_76_3518), .ZN(
      n_257_76_3519));
   NOR2_X1 i_257_76_3525 (.A1(n_257_76_3516), .A2(n_257_76_3519), .ZN(
      n_257_76_3520));
   NAND2_X1 i_257_76_3526 (.A1(n_257_76_3088), .A2(n_257_76_3520), .ZN(
      n_257_76_3521));
   NAND2_X1 i_257_76_3527 (.A1(n_257_76_3328), .A2(n_257_76_3089), .ZN(
      n_257_76_3522));
   NOR2_X1 i_257_76_3528 (.A1(n_257_76_3521), .A2(n_257_76_3522), .ZN(
      n_257_76_3523));
   NAND2_X1 i_257_76_3529 (.A1(n_257_76_3514), .A2(n_257_76_3523), .ZN(
      n_257_76_3524));
   INV_X1 i_257_76_3530 (.A(n_257_76_3524), .ZN(n_257_76_3525));
   NAND2_X1 i_257_76_3531 (.A1(n_257_76_3525), .A2(n_257_76_3337), .ZN(
      n_257_76_3526));
   NOR2_X1 i_257_76_3532 (.A1(n_257_76_3345), .A2(n_257_76_3526), .ZN(
      n_257_76_3527));
   NAND2_X1 i_257_76_3533 (.A1(n_257_76_3318), .A2(n_257_76_3527), .ZN(
      n_257_76_3528));
   NOR2_X1 i_257_76_3534 (.A1(n_257_76_3528), .A2(n_257_76_3350), .ZN(
      n_257_76_3529));
   NAND2_X1 i_257_76_3535 (.A1(n_257_76_18060), .A2(n_257_76_3529), .ZN(
      n_257_76_3530));
   INV_X1 i_257_76_3536 (.A(n_257_1032), .ZN(n_257_76_3531));
   OAI21_X1 i_257_76_3537 (.A(n_257_76_3441), .B1(n_257_76_3531), .B2(
      n_257_76_17968), .ZN(n_257_76_3532));
   INV_X1 i_257_76_3538 (.A(n_257_76_3423), .ZN(n_257_76_3533));
   NOR2_X1 i_257_76_3539 (.A1(n_257_76_3532), .A2(n_257_76_3533), .ZN(
      n_257_76_3534));
   NAND2_X1 i_257_76_3540 (.A1(n_257_968), .A2(n_257_442), .ZN(n_257_76_3535));
   INV_X1 i_257_76_3541 (.A(n_257_76_3535), .ZN(n_257_76_3536));
   NAND2_X1 i_257_76_3542 (.A1(n_257_441), .A2(n_257_76_3536), .ZN(n_257_76_3537));
   NAND2_X1 i_257_76_3543 (.A1(n_257_834), .A2(n_257_442), .ZN(n_257_76_3538));
   INV_X1 i_257_76_3544 (.A(n_257_76_3538), .ZN(n_257_76_3539));
   AOI22_X1 i_257_76_3545 (.A1(n_257_446), .A2(n_257_76_3539), .B1(n_257_449), 
      .B2(n_257_76_10974), .ZN(n_257_76_3540));
   NAND2_X1 i_257_76_3546 (.A1(n_257_76_3537), .A2(n_257_76_3540), .ZN(
      n_257_76_3541));
   NAND2_X1 i_257_76_3547 (.A1(n_257_80), .A2(n_257_76_17932), .ZN(n_257_76_3542));
   NAND2_X1 i_257_76_3548 (.A1(n_257_76_3194), .A2(n_257_76_3542), .ZN(
      n_257_76_3543));
   NOR2_X1 i_257_76_3549 (.A1(n_257_76_3541), .A2(n_257_76_3543), .ZN(
      n_257_76_3544));
   NAND2_X1 i_257_76_3550 (.A1(n_257_40), .A2(n_257_76_17918), .ZN(n_257_76_3545));
   NAND2_X1 i_257_76_3551 (.A1(n_257_76_3478), .A2(n_257_76_3545), .ZN(
      n_257_76_3546));
   INV_X1 i_257_76_3552 (.A(n_257_76_3546), .ZN(n_257_76_3547));
   NAND2_X1 i_257_76_3553 (.A1(n_257_76_3012), .A2(Small_Packet_Data_Size[5]), 
      .ZN(n_257_76_3548));
   INV_X1 i_257_76_3554 (.A(Small_Packet_Data_Size[5]), .ZN(n_257_76_3549));
   OAI21_X1 i_257_76_3555 (.A(n_257_76_3548), .B1(n_257_442), .B2(n_257_76_3549), 
      .ZN(n_257_76_3550));
   NAND2_X1 i_257_76_3556 (.A1(n_257_76_3517), .A2(n_257_76_3550), .ZN(
      n_257_76_3551));
   NOR2_X1 i_257_76_3557 (.A1(n_257_76_3551), .A2(n_257_76_3144), .ZN(
      n_257_76_3552));
   NAND2_X1 i_257_76_3558 (.A1(n_257_76_3552), .A2(n_257_76_3324), .ZN(
      n_257_76_3553));
   NAND3_X1 i_257_76_3559 (.A1(n_257_435), .A2(n_257_706), .A3(n_257_442), 
      .ZN(n_257_76_3554));
   NAND2_X1 i_257_76_3560 (.A1(n_257_602), .A2(n_257_442), .ZN(n_257_76_3555));
   INV_X1 i_257_76_3561 (.A(n_257_76_3555), .ZN(n_257_76_3556));
   NAND2_X1 i_257_76_3562 (.A1(n_257_432), .A2(n_257_76_3556), .ZN(n_257_76_3557));
   NAND2_X1 i_257_76_3563 (.A1(n_257_76_3554), .A2(n_257_76_3557), .ZN(
      n_257_76_3558));
   NOR2_X1 i_257_76_3564 (.A1(n_257_76_3553), .A2(n_257_76_3558), .ZN(
      n_257_76_3559));
   NAND2_X1 i_257_76_3565 (.A1(n_257_76_3547), .A2(n_257_76_3559), .ZN(
      n_257_76_3560));
   NAND2_X1 i_257_76_3566 (.A1(n_257_634), .A2(n_257_76_17928), .ZN(
      n_257_76_3561));
   NAND2_X1 i_257_76_3567 (.A1(n_257_76_3455), .A2(n_257_76_3561), .ZN(
      n_257_76_3562));
   NOR2_X1 i_257_76_3568 (.A1(n_257_76_3560), .A2(n_257_76_3562), .ZN(
      n_257_76_3563));
   NAND2_X1 i_257_76_3569 (.A1(n_257_802), .A2(n_257_76_17952), .ZN(
      n_257_76_3564));
   NAND3_X1 i_257_76_3570 (.A1(n_257_439), .A2(n_257_904), .A3(n_257_442), 
      .ZN(n_257_76_3565));
   NAND2_X1 i_257_76_3571 (.A1(n_257_76_3564), .A2(n_257_76_3565), .ZN(
      n_257_76_3566));
   NAND2_X1 i_257_76_3572 (.A1(n_257_442), .A2(n_257_936), .ZN(n_257_76_3567));
   INV_X1 i_257_76_3573 (.A(n_257_76_3567), .ZN(n_257_76_3568));
   NAND2_X1 i_257_76_3574 (.A1(n_257_440), .A2(n_257_76_3568), .ZN(n_257_76_3569));
   NAND2_X1 i_257_76_3575 (.A1(n_257_438), .A2(n_257_76_6607), .ZN(n_257_76_3570));
   NAND2_X1 i_257_76_3576 (.A1(n_257_76_3569), .A2(n_257_76_3570), .ZN(
      n_257_76_3571));
   NOR2_X1 i_257_76_3577 (.A1(n_257_76_3566), .A2(n_257_76_3571), .ZN(
      n_257_76_3572));
   NAND2_X1 i_257_76_3578 (.A1(n_257_76_3563), .A2(n_257_76_3572), .ZN(
      n_257_76_3573));
   NAND2_X1 i_257_76_3579 (.A1(n_257_118), .A2(n_257_76_17925), .ZN(
      n_257_76_3574));
   NAND2_X1 i_257_76_3580 (.A1(n_257_738), .A2(n_257_76_17935), .ZN(
      n_257_76_3575));
   NAND2_X1 i_257_76_3581 (.A1(n_257_76_3574), .A2(n_257_76_3575), .ZN(
      n_257_76_3576));
   NAND2_X1 i_257_76_3582 (.A1(n_257_866), .A2(n_257_76_17903), .ZN(
      n_257_76_3577));
   NAND2_X1 i_257_76_3583 (.A1(n_257_76_3501), .A2(n_257_76_3577), .ZN(
      n_257_76_3578));
   NOR2_X1 i_257_76_3584 (.A1(n_257_76_3576), .A2(n_257_76_3578), .ZN(
      n_257_76_3579));
   NAND2_X1 i_257_76_3585 (.A1(n_257_442), .A2(n_257_770), .ZN(n_257_76_3580));
   INV_X1 i_257_76_3586 (.A(n_257_76_3580), .ZN(n_257_76_3581));
   NAND2_X1 i_257_76_3587 (.A1(n_257_457), .A2(n_257_442), .ZN(n_257_76_3582));
   INV_X1 i_257_76_3588 (.A(n_257_76_3582), .ZN(n_257_76_3583));
   AOI22_X1 i_257_76_3589 (.A1(n_257_447), .A2(n_257_76_3581), .B1(n_257_451), 
      .B2(n_257_76_3583), .ZN(n_257_76_3584));
   NAND2_X1 i_257_76_3590 (.A1(n_257_76_3579), .A2(n_257_76_3584), .ZN(
      n_257_76_3585));
   NOR2_X1 i_257_76_3591 (.A1(n_257_76_3573), .A2(n_257_76_3585), .ZN(
      n_257_76_3586));
   NAND2_X1 i_257_76_3592 (.A1(n_257_76_3544), .A2(n_257_76_3586), .ZN(
      n_257_76_3587));
   NAND2_X1 i_257_76_3593 (.A1(n_257_674), .A2(n_257_76_17958), .ZN(
      n_257_76_3588));
   NAND2_X1 i_257_76_3594 (.A1(n_257_157), .A2(n_257_76_17331), .ZN(
      n_257_76_3589));
   NAND2_X1 i_257_76_3595 (.A1(n_257_76_3588), .A2(n_257_76_3589), .ZN(
      n_257_76_3590));
   NOR2_X1 i_257_76_3596 (.A1(n_257_76_3590), .A2(n_257_76_3099), .ZN(
      n_257_76_3591));
   NAND2_X1 i_257_76_3597 (.A1(n_257_1000), .A2(n_257_76_17964), .ZN(
      n_257_76_3592));
   NAND2_X1 i_257_76_3598 (.A1(n_257_76_3591), .A2(n_257_76_3592), .ZN(
      n_257_76_3593));
   NOR2_X1 i_257_76_3599 (.A1(n_257_76_3587), .A2(n_257_76_3593), .ZN(
      n_257_76_3594));
   NAND2_X1 i_257_76_3600 (.A1(n_257_76_3534), .A2(n_257_76_3594), .ZN(
      n_257_76_3595));
   NAND3_X1 i_257_76_3601 (.A1(n_257_76_3511), .A2(n_257_76_3530), .A3(
      n_257_76_3595), .ZN(n_257_76_3596));
   INV_X1 i_257_76_3602 (.A(n_257_76_3596), .ZN(n_257_76_3597));
   NAND3_X1 i_257_76_3603 (.A1(n_257_76_3447), .A2(n_257_76_3497), .A3(
      n_257_76_3597), .ZN(n_257_76_3598));
   NOR2_X1 i_257_76_3604 (.A1(n_257_76_3397), .A2(n_257_76_3598), .ZN(
      n_257_76_3599));
   NAND2_X1 i_257_76_3605 (.A1(n_257_76_3254), .A2(n_257_76_3599), .ZN(n_5));
   NAND2_X1 i_257_76_3606 (.A1(n_257_1033), .A2(n_257_443), .ZN(n_257_76_3600));
   NAND2_X1 i_257_76_3607 (.A1(n_257_1001), .A2(n_257_444), .ZN(n_257_76_3601));
   NAND2_X1 i_257_76_3608 (.A1(n_257_441), .A2(n_257_969), .ZN(n_257_76_3602));
   INV_X1 i_257_76_3609 (.A(n_257_1065), .ZN(n_257_76_3603));
   NAND2_X1 i_257_76_3610 (.A1(n_257_76_3603), .A2(n_257_442), .ZN(n_257_76_3604));
   INV_X1 i_257_76_3611 (.A(n_257_937), .ZN(n_257_76_3605));
   NOR2_X1 i_257_76_3612 (.A1(n_257_76_3604), .A2(n_257_76_3605), .ZN(
      n_257_76_3606));
   NAND2_X1 i_257_76_3613 (.A1(n_257_440), .A2(n_257_76_3606), .ZN(n_257_76_3607));
   INV_X1 i_257_76_3614 (.A(n_257_76_3607), .ZN(n_257_76_3608));
   NAND2_X1 i_257_76_3615 (.A1(n_257_76_3602), .A2(n_257_76_3608), .ZN(
      n_257_76_3609));
   INV_X1 i_257_76_3616 (.A(n_257_76_3609), .ZN(n_257_76_3610));
   NAND2_X1 i_257_76_3617 (.A1(n_257_76_3601), .A2(n_257_76_3610), .ZN(
      n_257_76_3611));
   INV_X1 i_257_76_3618 (.A(n_257_76_3611), .ZN(n_257_76_3612));
   NAND2_X1 i_257_76_3619 (.A1(n_257_76_3600), .A2(n_257_76_3612), .ZN(
      n_257_76_3613));
   INV_X1 i_257_76_3620 (.A(n_257_76_3613), .ZN(n_257_76_3614));
   NAND2_X1 i_257_76_3621 (.A1(n_257_17), .A2(n_257_76_3614), .ZN(n_257_76_3615));
   INV_X1 i_257_76_3622 (.A(n_257_76_3604), .ZN(n_257_76_3616));
   NAND2_X1 i_257_76_3623 (.A1(n_257_443), .A2(n_257_76_3616), .ZN(n_257_76_3617));
   INV_X1 i_257_76_3624 (.A(n_257_76_3617), .ZN(n_257_76_3618));
   NAND2_X1 i_257_76_3625 (.A1(n_257_1033), .A2(n_257_76_3618), .ZN(
      n_257_76_3619));
   INV_X1 i_257_76_3626 (.A(n_257_76_3619), .ZN(n_257_76_3620));
   NAND2_X1 i_257_76_3627 (.A1(n_257_76_18072), .A2(n_257_76_3620), .ZN(
      n_257_76_3621));
   INV_X1 i_257_76_3628 (.A(n_257_76_3600), .ZN(n_257_76_3622));
   NAND2_X1 i_257_76_3629 (.A1(n_257_803), .A2(n_257_437), .ZN(n_257_76_3623));
   NAND2_X1 i_257_76_3630 (.A1(n_257_76_3602), .A2(n_257_76_3623), .ZN(
      n_257_76_3624));
   NAND2_X1 i_257_76_3631 (.A1(n_257_739), .A2(n_257_436), .ZN(n_257_76_3625));
   NAND2_X1 i_257_76_3632 (.A1(n_257_867), .A2(n_257_445), .ZN(n_257_76_3626));
   NAND2_X1 i_257_76_3633 (.A1(n_257_446), .A2(n_257_835), .ZN(n_257_76_3627));
   NAND3_X1 i_257_76_3634 (.A1(n_257_76_3625), .A2(n_257_76_3626), .A3(
      n_257_76_3627), .ZN(n_257_76_3628));
   NOR2_X1 i_257_76_3635 (.A1(n_257_76_3624), .A2(n_257_76_3628), .ZN(
      n_257_76_3629));
   NAND2_X1 i_257_76_3636 (.A1(n_257_675), .A2(n_257_448), .ZN(n_257_76_3630));
   NAND2_X1 i_257_76_3637 (.A1(n_257_905), .A2(n_257_439), .ZN(n_257_76_3631));
   NAND2_X1 i_257_76_3638 (.A1(n_257_707), .A2(n_257_435), .ZN(n_257_76_3632));
   NAND2_X1 i_257_76_3639 (.A1(n_257_450), .A2(n_257_76_3616), .ZN(n_257_76_3633));
   INV_X1 i_257_76_3640 (.A(n_257_76_3633), .ZN(n_257_76_3634));
   NAND3_X1 i_257_76_3641 (.A1(n_257_76_3632), .A2(n_257_635), .A3(n_257_76_3634), 
      .ZN(n_257_76_3635));
   INV_X1 i_257_76_3642 (.A(n_257_76_3635), .ZN(n_257_76_3636));
   NAND2_X1 i_257_76_3643 (.A1(n_257_440), .A2(n_257_937), .ZN(n_257_76_3637));
   NAND2_X1 i_257_76_3644 (.A1(n_257_438), .A2(n_257_1071), .ZN(n_257_76_3638));
   NAND4_X1 i_257_76_3645 (.A1(n_257_76_3631), .A2(n_257_76_3636), .A3(
      n_257_76_3637), .A4(n_257_76_3638), .ZN(n_257_76_3639));
   NAND2_X1 i_257_76_3646 (.A1(n_257_449), .A2(n_257_1079), .ZN(n_257_76_3640));
   NAND2_X1 i_257_76_3647 (.A1(n_257_447), .A2(n_257_771), .ZN(n_257_76_3641));
   NAND2_X1 i_257_76_3648 (.A1(n_257_76_3640), .A2(n_257_76_3641), .ZN(
      n_257_76_3642));
   NOR2_X1 i_257_76_3649 (.A1(n_257_76_3639), .A2(n_257_76_3642), .ZN(
      n_257_76_3643));
   NAND3_X1 i_257_76_3650 (.A1(n_257_76_3629), .A2(n_257_76_3630), .A3(
      n_257_76_3643), .ZN(n_257_76_3644));
   INV_X1 i_257_76_3651 (.A(n_257_76_3644), .ZN(n_257_76_3645));
   NAND2_X1 i_257_76_3652 (.A1(n_257_76_3645), .A2(n_257_76_3601), .ZN(
      n_257_76_3646));
   NOR2_X1 i_257_76_3653 (.A1(n_257_76_3622), .A2(n_257_76_3646), .ZN(
      n_257_76_3647));
   NAND2_X1 i_257_76_3654 (.A1(n_257_28), .A2(n_257_76_3647), .ZN(n_257_76_3648));
   NAND3_X1 i_257_76_3655 (.A1(n_257_76_3615), .A2(n_257_76_3621), .A3(
      n_257_76_3648), .ZN(n_257_76_3649));
   NAND2_X1 i_257_76_3656 (.A1(n_257_76_3631), .A2(n_257_446), .ZN(n_257_76_3650));
   INV_X1 i_257_76_3657 (.A(n_257_76_3650), .ZN(n_257_76_3651));
   NAND2_X1 i_257_76_3658 (.A1(n_257_835), .A2(n_257_76_3616), .ZN(n_257_76_3652));
   INV_X1 i_257_76_3659 (.A(n_257_76_3652), .ZN(n_257_76_3653));
   NAND3_X1 i_257_76_3660 (.A1(n_257_76_3637), .A2(n_257_76_3638), .A3(
      n_257_76_3653), .ZN(n_257_76_3654));
   INV_X1 i_257_76_3661 (.A(n_257_76_3654), .ZN(n_257_76_3655));
   NAND4_X1 i_257_76_3662 (.A1(n_257_76_3602), .A2(n_257_76_3651), .A3(
      n_257_76_3655), .A4(n_257_76_3626), .ZN(n_257_76_3656));
   INV_X1 i_257_76_3663 (.A(n_257_76_3656), .ZN(n_257_76_3657));
   NAND2_X1 i_257_76_3664 (.A1(n_257_76_3601), .A2(n_257_76_3657), .ZN(
      n_257_76_3658));
   INV_X1 i_257_76_3665 (.A(n_257_76_3658), .ZN(n_257_76_3659));
   NAND2_X1 i_257_76_3666 (.A1(n_257_76_3600), .A2(n_257_76_3659), .ZN(
      n_257_76_3660));
   INV_X1 i_257_76_3667 (.A(n_257_76_3660), .ZN(n_257_76_3661));
   NAND2_X1 i_257_76_3668 (.A1(n_257_76_18070), .A2(n_257_76_3661), .ZN(
      n_257_76_3662));
   NAND2_X1 i_257_76_3669 (.A1(n_257_439), .A2(n_257_76_3616), .ZN(n_257_76_3663));
   INV_X1 i_257_76_3670 (.A(n_257_76_3663), .ZN(n_257_76_3664));
   NAND3_X1 i_257_76_3671 (.A1(n_257_76_3664), .A2(n_257_76_3637), .A3(n_257_905), 
      .ZN(n_257_76_3665));
   INV_X1 i_257_76_3672 (.A(n_257_76_3665), .ZN(n_257_76_3666));
   NAND2_X1 i_257_76_3673 (.A1(n_257_76_3602), .A2(n_257_76_3666), .ZN(
      n_257_76_3667));
   INV_X1 i_257_76_3674 (.A(n_257_76_3667), .ZN(n_257_76_3668));
   NAND2_X1 i_257_76_3675 (.A1(n_257_76_3601), .A2(n_257_76_3668), .ZN(
      n_257_76_3669));
   INV_X1 i_257_76_3676 (.A(n_257_76_3669), .ZN(n_257_76_3670));
   NAND2_X1 i_257_76_3677 (.A1(n_257_76_3600), .A2(n_257_76_3670), .ZN(
      n_257_76_3671));
   INV_X1 i_257_76_3678 (.A(n_257_76_3671), .ZN(n_257_76_3672));
   NAND2_X1 i_257_76_3679 (.A1(n_257_76_18084), .A2(n_257_76_3672), .ZN(
      n_257_76_3673));
   NAND2_X1 i_257_76_3680 (.A1(n_257_451), .A2(n_257_458), .ZN(n_257_76_3674));
   NAND2_X1 i_257_76_3681 (.A1(n_257_76_3602), .A2(n_257_76_3674), .ZN(
      n_257_76_3675));
   NAND3_X1 i_257_76_3682 (.A1(n_257_76_3627), .A2(n_257_76_3640), .A3(
      n_257_76_3641), .ZN(n_257_76_3676));
   NOR2_X1 i_257_76_3683 (.A1(n_257_76_3675), .A2(n_257_76_3676), .ZN(
      n_257_76_3677));
   NAND2_X1 i_257_76_3684 (.A1(n_257_238), .A2(n_257_425), .ZN(n_257_76_3678));
   NAND2_X1 i_257_76_3685 (.A1(n_257_81), .A2(n_257_431), .ZN(n_257_76_3679));
   NAND3_X1 i_257_76_3686 (.A1(n_257_76_3677), .A2(n_257_76_3678), .A3(
      n_257_76_3679), .ZN(n_257_76_3680));
   NAND2_X1 i_257_76_3687 (.A1(n_257_158), .A2(n_257_429), .ZN(n_257_76_3681));
   NAND2_X1 i_257_76_3688 (.A1(n_257_76_3681), .A2(n_257_76_3630), .ZN(
      n_257_76_3682));
   NOR2_X1 i_257_76_3689 (.A1(n_257_76_3680), .A2(n_257_76_3682), .ZN(
      n_257_76_3683));
   NAND2_X1 i_257_76_3690 (.A1(n_257_119), .A2(n_257_430), .ZN(n_257_76_3684));
   NAND2_X1 i_257_76_3691 (.A1(n_257_76_3684), .A2(n_257_76_3623), .ZN(
      n_257_76_3685));
   INV_X1 i_257_76_3692 (.A(n_257_76_3685), .ZN(n_257_76_3686));
   NAND2_X1 i_257_76_3693 (.A1(n_257_41), .A2(n_257_433), .ZN(n_257_76_3687));
   NAND2_X1 i_257_76_3694 (.A1(n_257_539), .A2(n_257_426), .ZN(n_257_76_3688));
   NAND4_X1 i_257_76_3695 (.A1(n_257_76_3625), .A2(n_257_76_3626), .A3(
      n_257_76_3687), .A4(n_257_76_3688), .ZN(n_257_76_3689));
   INV_X1 i_257_76_3696 (.A(n_257_76_3689), .ZN(n_257_76_3690));
   NAND2_X1 i_257_76_3697 (.A1(n_257_198), .A2(n_257_427), .ZN(n_257_76_3691));
   NAND4_X1 i_257_76_3698 (.A1(n_257_76_3631), .A2(n_257_278), .A3(n_257_76_3691), 
      .A4(n_257_76_3637), .ZN(n_257_76_3692));
   NAND2_X1 i_257_76_3699 (.A1(n_257_507), .A2(n_257_424), .ZN(n_257_76_3693));
   NAND2_X1 i_257_76_3700 (.A1(n_257_76_3693), .A2(n_257_76_3632), .ZN(
      n_257_76_3694));
   INV_X1 i_257_76_3701 (.A(n_257_76_3694), .ZN(n_257_76_3695));
   NAND2_X1 i_257_76_3702 (.A1(n_257_635), .A2(n_257_450), .ZN(n_257_76_3696));
   NAND2_X1 i_257_76_3703 (.A1(n_257_432), .A2(n_257_603), .ZN(n_257_76_3697));
   NAND2_X1 i_257_76_3704 (.A1(n_257_428), .A2(n_257_571), .ZN(n_257_76_3698));
   NAND2_X1 i_257_76_3705 (.A1(n_257_423), .A2(n_257_76_3616), .ZN(n_257_76_3699));
   INV_X1 i_257_76_3706 (.A(n_257_76_3699), .ZN(n_257_76_3700));
   NAND3_X1 i_257_76_3707 (.A1(n_257_76_3697), .A2(n_257_76_3698), .A3(
      n_257_76_3700), .ZN(n_257_76_3701));
   INV_X1 i_257_76_3708 (.A(n_257_76_3701), .ZN(n_257_76_3702));
   NAND4_X1 i_257_76_3709 (.A1(n_257_76_3695), .A2(n_257_76_3638), .A3(
      n_257_76_3696), .A4(n_257_76_3702), .ZN(n_257_76_3703));
   NOR2_X1 i_257_76_3710 (.A1(n_257_76_3692), .A2(n_257_76_3703), .ZN(
      n_257_76_3704));
   NAND3_X1 i_257_76_3711 (.A1(n_257_76_3686), .A2(n_257_76_3690), .A3(
      n_257_76_3704), .ZN(n_257_76_3705));
   INV_X1 i_257_76_3712 (.A(n_257_76_3705), .ZN(n_257_76_3706));
   NAND2_X1 i_257_76_3713 (.A1(n_257_76_3601), .A2(n_257_76_3706), .ZN(
      n_257_76_3707));
   INV_X1 i_257_76_3714 (.A(n_257_76_3707), .ZN(n_257_76_3708));
   NAND3_X1 i_257_76_3715 (.A1(n_257_76_3683), .A2(n_257_76_3600), .A3(
      n_257_76_3708), .ZN(n_257_76_3709));
   INV_X1 i_257_76_3716 (.A(n_257_76_3709), .ZN(n_257_76_3710));
   NAND2_X1 i_257_76_3717 (.A1(n_257_76_18066), .A2(n_257_76_3710), .ZN(
      n_257_76_3711));
   NAND3_X1 i_257_76_3718 (.A1(n_257_76_3662), .A2(n_257_76_3673), .A3(
      n_257_76_3711), .ZN(n_257_76_3712));
   NOR2_X1 i_257_76_3719 (.A1(n_257_76_3649), .A2(n_257_76_3712), .ZN(
      n_257_76_3713));
   NAND2_X1 i_257_76_3720 (.A1(n_257_969), .A2(n_257_76_3616), .ZN(n_257_76_3714));
   INV_X1 i_257_76_3721 (.A(n_257_76_3714), .ZN(n_257_76_3715));
   NAND2_X1 i_257_76_3722 (.A1(n_257_441), .A2(n_257_76_3715), .ZN(n_257_76_3716));
   INV_X1 i_257_76_3723 (.A(n_257_76_3716), .ZN(n_257_76_3717));
   NAND2_X1 i_257_76_3724 (.A1(n_257_76_3601), .A2(n_257_76_3717), .ZN(
      n_257_76_3718));
   INV_X1 i_257_76_3725 (.A(n_257_76_3718), .ZN(n_257_76_3719));
   NAND2_X1 i_257_76_3726 (.A1(n_257_76_3600), .A2(n_257_76_3719), .ZN(
      n_257_76_3720));
   INV_X1 i_257_76_3727 (.A(n_257_76_3720), .ZN(n_257_76_3721));
   NAND2_X1 i_257_76_3728 (.A1(n_257_76_18071), .A2(n_257_76_3721), .ZN(
      n_257_76_3722));
   NAND4_X1 i_257_76_3729 (.A1(n_257_76_3602), .A2(n_257_76_3623), .A3(
      n_257_76_3625), .A4(n_257_76_3626), .ZN(n_257_76_3723));
   INV_X1 i_257_76_3730 (.A(n_257_707), .ZN(n_257_76_3724));
   NAND2_X1 i_257_76_3731 (.A1(n_257_435), .A2(n_257_76_3616), .ZN(n_257_76_3725));
   NOR2_X1 i_257_76_3732 (.A1(n_257_76_3724), .A2(n_257_76_3725), .ZN(
      n_257_76_3726));
   NAND3_X1 i_257_76_3733 (.A1(n_257_76_3637), .A2(n_257_76_3638), .A3(
      n_257_76_3726), .ZN(n_257_76_3727));
   INV_X1 i_257_76_3734 (.A(n_257_76_3727), .ZN(n_257_76_3728));
   NAND4_X1 i_257_76_3735 (.A1(n_257_76_3728), .A2(n_257_76_3627), .A3(
      n_257_76_3641), .A4(n_257_76_3631), .ZN(n_257_76_3729));
   NOR2_X1 i_257_76_3736 (.A1(n_257_76_3723), .A2(n_257_76_3729), .ZN(
      n_257_76_3730));
   NAND2_X1 i_257_76_3737 (.A1(n_257_76_3601), .A2(n_257_76_3730), .ZN(
      n_257_76_3731));
   INV_X1 i_257_76_3738 (.A(n_257_76_3731), .ZN(n_257_76_3732));
   NAND2_X1 i_257_76_3739 (.A1(n_257_76_3600), .A2(n_257_76_3732), .ZN(
      n_257_76_3733));
   INV_X1 i_257_76_3740 (.A(n_257_76_3733), .ZN(n_257_76_3734));
   NAND2_X1 i_257_76_3741 (.A1(n_257_76_18078), .A2(n_257_76_3734), .ZN(
      n_257_76_3735));
   NAND3_X1 i_257_76_3742 (.A1(n_257_76_3626), .A2(n_257_76_3627), .A3(
      n_257_76_3640), .ZN(n_257_76_3736));
   NAND2_X1 i_257_76_3743 (.A1(n_257_76_3623), .A2(n_257_76_3625), .ZN(
      n_257_76_3737));
   NOR2_X1 i_257_76_3744 (.A1(n_257_76_3736), .A2(n_257_76_3737), .ZN(
      n_257_76_3738));
   NAND3_X1 i_257_76_3745 (.A1(n_257_76_3684), .A2(n_257_76_3602), .A3(
      n_257_76_3674), .ZN(n_257_76_3739));
   INV_X1 i_257_76_3746 (.A(n_257_76_3739), .ZN(n_257_76_3740));
   NAND3_X1 i_257_76_3747 (.A1(n_257_76_3641), .A2(n_257_76_3687), .A3(
      n_257_76_3631), .ZN(n_257_76_3741));
   NAND3_X1 i_257_76_3748 (.A1(n_257_76_3603), .A2(n_257_442), .A3(n_257_571), 
      .ZN(n_257_76_3742));
   INV_X1 i_257_76_3749 (.A(n_257_76_3742), .ZN(n_257_76_3743));
   NAND2_X1 i_257_76_3750 (.A1(n_257_428), .A2(n_257_76_3743), .ZN(n_257_76_3744));
   INV_X1 i_257_76_3751 (.A(n_257_76_3744), .ZN(n_257_76_3745));
   NAND2_X1 i_257_76_3752 (.A1(n_257_76_3697), .A2(n_257_76_3745), .ZN(
      n_257_76_3746));
   INV_X1 i_257_76_3753 (.A(n_257_76_3746), .ZN(n_257_76_3747));
   NAND2_X1 i_257_76_3754 (.A1(n_257_76_3747), .A2(n_257_76_3632), .ZN(
      n_257_76_3748));
   INV_X1 i_257_76_3755 (.A(n_257_76_3748), .ZN(n_257_76_3749));
   NAND4_X1 i_257_76_3756 (.A1(n_257_76_3749), .A2(n_257_76_3637), .A3(
      n_257_76_3638), .A4(n_257_76_3696), .ZN(n_257_76_3750));
   NOR2_X1 i_257_76_3757 (.A1(n_257_76_3741), .A2(n_257_76_3750), .ZN(
      n_257_76_3751));
   NAND4_X1 i_257_76_3758 (.A1(n_257_76_3738), .A2(n_257_76_3740), .A3(
      n_257_76_3679), .A4(n_257_76_3751), .ZN(n_257_76_3752));
   INV_X1 i_257_76_3759 (.A(n_257_76_3752), .ZN(n_257_76_3753));
   INV_X1 i_257_76_3760 (.A(n_257_76_3682), .ZN(n_257_76_3754));
   NAND3_X1 i_257_76_3761 (.A1(n_257_76_3753), .A2(n_257_76_3754), .A3(
      n_257_76_3601), .ZN(n_257_76_3755));
   NOR2_X1 i_257_76_3762 (.A1(n_257_76_3755), .A2(n_257_76_3622), .ZN(
      n_257_76_3756));
   NAND2_X1 i_257_76_3763 (.A1(n_257_76_18074), .A2(n_257_76_3756), .ZN(
      n_257_76_3757));
   NAND3_X1 i_257_76_3764 (.A1(n_257_76_3722), .A2(n_257_76_3735), .A3(
      n_257_76_3757), .ZN(n_257_76_3758));
   NAND2_X1 i_257_76_3765 (.A1(n_257_1065), .A2(n_257_442), .ZN(n_257_76_3759));
   INV_X1 i_257_76_3766 (.A(n_257_76_3759), .ZN(n_257_76_3760));
   NAND2_X1 i_257_76_3767 (.A1(n_257_13), .A2(n_257_76_3760), .ZN(n_257_76_3761));
   NAND2_X1 i_257_76_3768 (.A1(n_257_867), .A2(n_257_76_3631), .ZN(n_257_76_3762));
   INV_X1 i_257_76_3769 (.A(n_257_76_3762), .ZN(n_257_76_3763));
   NAND2_X1 i_257_76_3770 (.A1(n_257_445), .A2(n_257_76_3616), .ZN(n_257_76_3764));
   INV_X1 i_257_76_3771 (.A(n_257_76_3764), .ZN(n_257_76_3765));
   NAND3_X1 i_257_76_3772 (.A1(n_257_76_3637), .A2(n_257_76_3638), .A3(
      n_257_76_3765), .ZN(n_257_76_3766));
   INV_X1 i_257_76_3773 (.A(n_257_76_3766), .ZN(n_257_76_3767));
   NAND3_X1 i_257_76_3774 (.A1(n_257_76_3602), .A2(n_257_76_3763), .A3(
      n_257_76_3767), .ZN(n_257_76_3768));
   INV_X1 i_257_76_3775 (.A(n_257_76_3768), .ZN(n_257_76_3769));
   NAND2_X1 i_257_76_3776 (.A1(n_257_76_3601), .A2(n_257_76_3769), .ZN(
      n_257_76_3770));
   INV_X1 i_257_76_3777 (.A(n_257_76_3770), .ZN(n_257_76_3771));
   NAND2_X1 i_257_76_3778 (.A1(n_257_76_3600), .A2(n_257_76_3771), .ZN(
      n_257_76_3772));
   INV_X1 i_257_76_3779 (.A(n_257_76_3772), .ZN(n_257_76_3773));
   NAND2_X1 i_257_76_3780 (.A1(n_257_76_18077), .A2(n_257_76_3773), .ZN(
      n_257_76_3774));
   NAND2_X1 i_257_76_3781 (.A1(n_257_76_3761), .A2(n_257_76_3774), .ZN(
      n_257_76_3775));
   NOR2_X1 i_257_76_3782 (.A1(n_257_76_3758), .A2(n_257_76_3775), .ZN(
      n_257_76_3776));
   INV_X1 i_257_76_3783 (.A(n_257_76_3601), .ZN(n_257_76_3777));
   INV_X1 i_257_76_3784 (.A(n_257_76_3632), .ZN(n_257_76_3778));
   NAND2_X1 i_257_76_3785 (.A1(n_257_426), .A2(n_257_76_3616), .ZN(n_257_76_3779));
   INV_X1 i_257_76_3786 (.A(n_257_76_3779), .ZN(n_257_76_3780));
   NAND3_X1 i_257_76_3787 (.A1(n_257_76_3697), .A2(n_257_76_3698), .A3(
      n_257_76_3780), .ZN(n_257_76_3781));
   NOR2_X1 i_257_76_3788 (.A1(n_257_76_3778), .A2(n_257_76_3781), .ZN(
      n_257_76_3782));
   NAND4_X1 i_257_76_3789 (.A1(n_257_76_3782), .A2(n_257_539), .A3(n_257_76_3638), 
      .A4(n_257_76_3696), .ZN(n_257_76_3783));
   NAND3_X1 i_257_76_3790 (.A1(n_257_76_3631), .A2(n_257_76_3691), .A3(
      n_257_76_3637), .ZN(n_257_76_3784));
   NOR2_X1 i_257_76_3791 (.A1(n_257_76_3783), .A2(n_257_76_3784), .ZN(
      n_257_76_3785));
   NAND3_X1 i_257_76_3792 (.A1(n_257_76_3625), .A2(n_257_76_3626), .A3(
      n_257_76_3687), .ZN(n_257_76_3786));
   INV_X1 i_257_76_3793 (.A(n_257_76_3786), .ZN(n_257_76_3787));
   NAND3_X1 i_257_76_3794 (.A1(n_257_76_3785), .A2(n_257_76_3686), .A3(
      n_257_76_3787), .ZN(n_257_76_3788));
   NOR2_X1 i_257_76_3795 (.A1(n_257_76_3777), .A2(n_257_76_3788), .ZN(
      n_257_76_3789));
   NAND4_X1 i_257_76_3796 (.A1(n_257_76_3681), .A2(n_257_76_3630), .A3(
      n_257_76_3677), .A4(n_257_76_3679), .ZN(n_257_76_3790));
   INV_X1 i_257_76_3797 (.A(n_257_76_3790), .ZN(n_257_76_3791));
   NAND3_X1 i_257_76_3798 (.A1(n_257_76_3789), .A2(n_257_76_3600), .A3(
      n_257_76_3791), .ZN(n_257_76_3792));
   INV_X1 i_257_76_3799 (.A(n_257_76_3792), .ZN(n_257_76_3793));
   NAND2_X1 i_257_76_3800 (.A1(n_257_76_18076), .A2(n_257_76_3793), .ZN(
      n_257_76_3794));
   NAND4_X1 i_257_76_3801 (.A1(n_257_76_3602), .A2(n_257_76_3623), .A3(
      n_257_76_3626), .A4(n_257_76_3627), .ZN(n_257_76_3795));
   NAND2_X1 i_257_76_3802 (.A1(n_257_436), .A2(n_257_76_3616), .ZN(n_257_76_3796));
   INV_X1 i_257_76_3803 (.A(n_257_76_3796), .ZN(n_257_76_3797));
   NAND3_X1 i_257_76_3804 (.A1(n_257_76_3637), .A2(n_257_76_3638), .A3(
      n_257_76_3797), .ZN(n_257_76_3798));
   INV_X1 i_257_76_3805 (.A(n_257_76_3798), .ZN(n_257_76_3799));
   NAND4_X1 i_257_76_3806 (.A1(n_257_76_3799), .A2(n_257_76_3641), .A3(n_257_739), 
      .A4(n_257_76_3631), .ZN(n_257_76_3800));
   NOR2_X1 i_257_76_3807 (.A1(n_257_76_3795), .A2(n_257_76_3800), .ZN(
      n_257_76_3801));
   NAND2_X1 i_257_76_3808 (.A1(n_257_76_3601), .A2(n_257_76_3801), .ZN(
      n_257_76_3802));
   INV_X1 i_257_76_3809 (.A(n_257_76_3802), .ZN(n_257_76_3803));
   NAND2_X1 i_257_76_3810 (.A1(n_257_76_3600), .A2(n_257_76_3803), .ZN(
      n_257_76_3804));
   INV_X1 i_257_76_3811 (.A(n_257_76_3804), .ZN(n_257_76_3805));
   NAND2_X1 i_257_76_3812 (.A1(n_257_76_18069), .A2(n_257_76_3805), .ZN(
      n_257_76_3806));
   NAND4_X1 i_257_76_3813 (.A1(n_257_76_3626), .A2(n_257_76_3627), .A3(
      n_257_76_3640), .A4(n_257_76_3641), .ZN(n_257_76_3807));
   INV_X1 i_257_76_3814 (.A(n_257_76_3696), .ZN(n_257_76_3808));
   INV_X1 i_257_76_3815 (.A(n_257_603), .ZN(n_257_76_3809));
   NOR2_X1 i_257_76_3816 (.A1(n_257_76_3604), .A2(n_257_76_3809), .ZN(
      n_257_76_3810));
   NAND2_X1 i_257_76_3817 (.A1(n_257_432), .A2(n_257_76_3810), .ZN(n_257_76_3811));
   INV_X1 i_257_76_3818 (.A(n_257_76_3811), .ZN(n_257_76_3812));
   NAND2_X1 i_257_76_3819 (.A1(n_257_76_3632), .A2(n_257_76_3812), .ZN(
      n_257_76_3813));
   NOR2_X1 i_257_76_3820 (.A1(n_257_76_3808), .A2(n_257_76_3813), .ZN(
      n_257_76_3814));
   NAND2_X1 i_257_76_3821 (.A1(n_257_76_3637), .A2(n_257_76_3638), .ZN(
      n_257_76_3815));
   INV_X1 i_257_76_3822 (.A(n_257_76_3815), .ZN(n_257_76_3816));
   NAND4_X1 i_257_76_3823 (.A1(n_257_76_3814), .A2(n_257_76_3816), .A3(
      n_257_76_3687), .A4(n_257_76_3631), .ZN(n_257_76_3817));
   NOR2_X1 i_257_76_3824 (.A1(n_257_76_3807), .A2(n_257_76_3817), .ZN(
      n_257_76_3818));
   NAND4_X1 i_257_76_3825 (.A1(n_257_76_3602), .A2(n_257_76_3674), .A3(
      n_257_76_3623), .A4(n_257_76_3625), .ZN(n_257_76_3819));
   INV_X1 i_257_76_3826 (.A(n_257_76_3819), .ZN(n_257_76_3820));
   NAND3_X1 i_257_76_3827 (.A1(n_257_76_3818), .A2(n_257_76_3630), .A3(
      n_257_76_3820), .ZN(n_257_76_3821));
   NOR2_X1 i_257_76_3828 (.A1(n_257_76_3821), .A2(n_257_76_3777), .ZN(
      n_257_76_3822));
   NAND2_X1 i_257_76_3829 (.A1(n_257_76_3600), .A2(n_257_76_3822), .ZN(
      n_257_76_3823));
   INV_X1 i_257_76_3830 (.A(n_257_76_3823), .ZN(n_257_76_3824));
   NAND2_X1 i_257_76_3831 (.A1(n_257_68), .A2(n_257_76_3824), .ZN(n_257_76_3825));
   NAND3_X1 i_257_76_3832 (.A1(n_257_76_3794), .A2(n_257_76_3806), .A3(
      n_257_76_3825), .ZN(n_257_76_3826));
   NAND2_X1 i_257_76_3833 (.A1(n_257_437), .A2(n_257_76_3616), .ZN(n_257_76_3827));
   INV_X1 i_257_76_3834 (.A(n_257_76_3827), .ZN(n_257_76_3828));
   NAND3_X1 i_257_76_3835 (.A1(n_257_76_3637), .A2(n_257_76_3638), .A3(
      n_257_76_3828), .ZN(n_257_76_3829));
   INV_X1 i_257_76_3836 (.A(n_257_76_3829), .ZN(n_257_76_3830));
   NAND4_X1 i_257_76_3837 (.A1(n_257_76_3830), .A2(n_257_76_3627), .A3(n_257_803), 
      .A4(n_257_76_3631), .ZN(n_257_76_3831));
   NAND2_X1 i_257_76_3838 (.A1(n_257_76_3602), .A2(n_257_76_3626), .ZN(
      n_257_76_3832));
   NOR2_X1 i_257_76_3839 (.A1(n_257_76_3831), .A2(n_257_76_3832), .ZN(
      n_257_76_3833));
   NAND2_X1 i_257_76_3840 (.A1(n_257_76_3601), .A2(n_257_76_3833), .ZN(
      n_257_76_3834));
   INV_X1 i_257_76_3841 (.A(n_257_76_3834), .ZN(n_257_76_3835));
   NAND2_X1 i_257_76_3842 (.A1(n_257_76_3600), .A2(n_257_76_3835), .ZN(
      n_257_76_3836));
   INV_X1 i_257_76_3843 (.A(n_257_76_3836), .ZN(n_257_76_3837));
   NAND2_X1 i_257_76_3844 (.A1(n_257_22), .A2(n_257_76_3837), .ZN(n_257_76_3838));
   NAND2_X1 i_257_76_3845 (.A1(n_257_444), .A2(n_257_76_3616), .ZN(n_257_76_3839));
   INV_X1 i_257_76_3846 (.A(n_257_76_3839), .ZN(n_257_76_3840));
   NAND2_X1 i_257_76_3847 (.A1(n_257_1001), .A2(n_257_76_3840), .ZN(
      n_257_76_3841));
   INV_X1 i_257_76_3848 (.A(n_257_76_3841), .ZN(n_257_76_3842));
   NAND2_X1 i_257_76_3849 (.A1(n_257_76_3600), .A2(n_257_76_3842), .ZN(
      n_257_76_3843));
   INV_X1 i_257_76_3850 (.A(n_257_76_3843), .ZN(n_257_76_3844));
   NAND2_X1 i_257_76_3851 (.A1(n_257_76_18075), .A2(n_257_76_3844), .ZN(
      n_257_76_3845));
   NAND2_X1 i_257_76_3852 (.A1(n_257_76_3838), .A2(n_257_76_3845), .ZN(
      n_257_76_3846));
   NOR2_X1 i_257_76_3853 (.A1(n_257_76_3826), .A2(n_257_76_3846), .ZN(
      n_257_76_3847));
   NAND3_X1 i_257_76_3854 (.A1(n_257_76_3713), .A2(n_257_76_3776), .A3(
      n_257_76_3847), .ZN(n_257_76_3848));
   INV_X1 i_257_76_3855 (.A(n_257_76_3848), .ZN(n_257_76_3849));
   NAND2_X1 i_257_76_3856 (.A1(n_257_433), .A2(n_257_76_3616), .ZN(n_257_76_3850));
   INV_X1 i_257_76_3857 (.A(n_257_76_3850), .ZN(n_257_76_3851));
   NAND2_X1 i_257_76_3858 (.A1(n_257_76_3632), .A2(n_257_76_3851), .ZN(
      n_257_76_3852));
   NOR2_X1 i_257_76_3859 (.A1(n_257_76_3808), .A2(n_257_76_3852), .ZN(
      n_257_76_3853));
   NAND2_X1 i_257_76_3860 (.A1(n_257_41), .A2(n_257_76_3638), .ZN(n_257_76_3854));
   INV_X1 i_257_76_3861 (.A(n_257_76_3854), .ZN(n_257_76_3855));
   NAND4_X1 i_257_76_3862 (.A1(n_257_76_3853), .A2(n_257_76_3855), .A3(
      n_257_76_3631), .A4(n_257_76_3637), .ZN(n_257_76_3856));
   NOR2_X1 i_257_76_3863 (.A1(n_257_76_3807), .A2(n_257_76_3856), .ZN(
      n_257_76_3857));
   NAND3_X1 i_257_76_3864 (.A1(n_257_76_3857), .A2(n_257_76_3630), .A3(
      n_257_76_3820), .ZN(n_257_76_3858));
   NOR2_X1 i_257_76_3865 (.A1(n_257_76_3858), .A2(n_257_76_3777), .ZN(
      n_257_76_3859));
   NAND2_X1 i_257_76_3866 (.A1(n_257_76_3600), .A2(n_257_76_3859), .ZN(
      n_257_76_3860));
   INV_X1 i_257_76_3867 (.A(n_257_76_3860), .ZN(n_257_76_3861));
   NAND2_X1 i_257_76_3868 (.A1(n_257_76_18081), .A2(n_257_76_3861), .ZN(
      n_257_76_3862));
   NAND3_X1 i_257_76_3869 (.A1(n_257_76_3641), .A2(n_257_76_3631), .A3(n_257_449), 
      .ZN(n_257_76_3863));
   NAND2_X1 i_257_76_3870 (.A1(n_257_76_17760), .A2(n_257_76_3616), .ZN(
      n_257_76_3864));
   OAI21_X1 i_257_76_3871 (.A(n_257_76_3864), .B1(n_257_707), .B2(n_257_76_3604), 
      .ZN(n_257_76_3865));
   NAND4_X1 i_257_76_3872 (.A1(n_257_76_3637), .A2(n_257_76_3638), .A3(
      n_257_76_3865), .A4(n_257_1079), .ZN(n_257_76_3866));
   NOR2_X1 i_257_76_3873 (.A1(n_257_76_3863), .A2(n_257_76_3866), .ZN(
      n_257_76_3867));
   NAND3_X1 i_257_76_3874 (.A1(n_257_76_3629), .A2(n_257_76_3630), .A3(
      n_257_76_3867), .ZN(n_257_76_3868));
   INV_X1 i_257_76_3875 (.A(n_257_76_3868), .ZN(n_257_76_3869));
   NAND2_X1 i_257_76_3876 (.A1(n_257_76_3869), .A2(n_257_76_3601), .ZN(
      n_257_76_3870));
   NOR2_X1 i_257_76_3877 (.A1(n_257_76_3622), .A2(n_257_76_3870), .ZN(
      n_257_76_3871));
   NAND2_X1 i_257_76_3878 (.A1(n_257_76_18083), .A2(n_257_76_3871), .ZN(
      n_257_76_3872));
   NAND2_X1 i_257_76_3879 (.A1(n_257_429), .A2(n_257_76_3616), .ZN(n_257_76_3873));
   INV_X1 i_257_76_3880 (.A(n_257_76_3873), .ZN(n_257_76_3874));
   NAND2_X1 i_257_76_3881 (.A1(n_257_76_3697), .A2(n_257_76_3874), .ZN(
      n_257_76_3875));
   INV_X1 i_257_76_3882 (.A(n_257_76_3875), .ZN(n_257_76_3876));
   NAND2_X1 i_257_76_3883 (.A1(n_257_76_3876), .A2(n_257_76_3632), .ZN(
      n_257_76_3877));
   INV_X1 i_257_76_3884 (.A(n_257_76_3877), .ZN(n_257_76_3878));
   NAND4_X1 i_257_76_3885 (.A1(n_257_76_3878), .A2(n_257_76_3637), .A3(
      n_257_76_3638), .A4(n_257_76_3696), .ZN(n_257_76_3879));
   NOR2_X1 i_257_76_3886 (.A1(n_257_76_3741), .A2(n_257_76_3879), .ZN(
      n_257_76_3880));
   NAND4_X1 i_257_76_3887 (.A1(n_257_76_3738), .A2(n_257_76_3740), .A3(
      n_257_76_3679), .A4(n_257_76_3880), .ZN(n_257_76_3881));
   INV_X1 i_257_76_3888 (.A(n_257_76_3881), .ZN(n_257_76_3882));
   NAND2_X1 i_257_76_3889 (.A1(n_257_76_3630), .A2(n_257_158), .ZN(n_257_76_3883));
   INV_X1 i_257_76_3890 (.A(n_257_76_3883), .ZN(n_257_76_3884));
   NAND3_X1 i_257_76_3891 (.A1(n_257_76_3882), .A2(n_257_76_3601), .A3(
      n_257_76_3884), .ZN(n_257_76_3885));
   NOR2_X1 i_257_76_3892 (.A1(n_257_76_3885), .A2(n_257_76_3622), .ZN(
      n_257_76_3886));
   NAND2_X1 i_257_76_3893 (.A1(n_257_76_18061), .A2(n_257_76_3886), .ZN(
      n_257_76_3887));
   NAND3_X1 i_257_76_3894 (.A1(n_257_76_3862), .A2(n_257_76_3872), .A3(
      n_257_76_3887), .ZN(n_257_76_3888));
   INV_X1 i_257_76_3895 (.A(n_257_76_3888), .ZN(n_257_76_3889));
   NAND2_X1 i_257_76_3896 (.A1(n_257_1071), .A2(n_257_76_3616), .ZN(
      n_257_76_3890));
   INV_X1 i_257_76_3897 (.A(n_257_76_3890), .ZN(n_257_76_3891));
   NAND2_X1 i_257_76_3898 (.A1(n_257_438), .A2(n_257_76_3891), .ZN(n_257_76_3892));
   INV_X1 i_257_76_3899 (.A(n_257_76_3892), .ZN(n_257_76_3893));
   NAND3_X1 i_257_76_3900 (.A1(n_257_76_3631), .A2(n_257_76_3893), .A3(
      n_257_76_3637), .ZN(n_257_76_3894));
   INV_X1 i_257_76_3901 (.A(n_257_76_3894), .ZN(n_257_76_3895));
   NAND2_X1 i_257_76_3902 (.A1(n_257_76_3602), .A2(n_257_76_3895), .ZN(
      n_257_76_3896));
   INV_X1 i_257_76_3903 (.A(n_257_76_3896), .ZN(n_257_76_3897));
   NAND2_X1 i_257_76_3904 (.A1(n_257_76_3601), .A2(n_257_76_3897), .ZN(
      n_257_76_3898));
   INV_X1 i_257_76_3905 (.A(n_257_76_3898), .ZN(n_257_76_3899));
   NAND2_X1 i_257_76_3906 (.A1(n_257_76_3600), .A2(n_257_76_3899), .ZN(
      n_257_76_3900));
   INV_X1 i_257_76_3907 (.A(n_257_76_3900), .ZN(n_257_76_3901));
   NAND2_X1 i_257_76_3908 (.A1(n_257_76_18067), .A2(n_257_76_3901), .ZN(
      n_257_76_3902));
   NAND2_X1 i_257_76_3909 (.A1(n_257_316), .A2(n_257_422), .ZN(n_257_76_3903));
   NAND3_X1 i_257_76_3910 (.A1(n_257_76_3638), .A2(n_257_76_3903), .A3(
      n_257_76_3696), .ZN(n_257_76_3904));
   INV_X1 i_257_76_3911 (.A(n_257_76_3904), .ZN(n_257_76_3905));
   NAND2_X1 i_257_76_3912 (.A1(n_257_76_3691), .A2(n_257_76_3637), .ZN(
      n_257_76_3906));
   INV_X1 i_257_76_3913 (.A(n_257_76_3906), .ZN(n_257_76_3907));
   NAND3_X1 i_257_76_3914 (.A1(n_257_76_3603), .A2(n_257_442), .A3(n_257_897), 
      .ZN(n_257_76_3908));
   INV_X1 i_257_76_3915 (.A(n_257_76_3908), .ZN(n_257_76_3909));
   NAND3_X1 i_257_76_3916 (.A1(n_257_420), .A2(n_257_76_3698), .A3(n_257_76_3909), 
      .ZN(n_257_76_3910));
   INV_X1 i_257_76_3917 (.A(n_257_76_3910), .ZN(n_257_76_3911));
   NAND4_X1 i_257_76_3918 (.A1(n_257_76_3911), .A2(n_257_76_3693), .A3(
      n_257_76_3632), .A4(n_257_76_3697), .ZN(n_257_76_3912));
   INV_X1 i_257_76_3919 (.A(n_257_76_3912), .ZN(n_257_76_3913));
   NAND3_X1 i_257_76_3920 (.A1(n_257_76_3905), .A2(n_257_76_3907), .A3(
      n_257_76_3913), .ZN(n_257_76_3914));
   NAND4_X1 i_257_76_3921 (.A1(n_257_76_3641), .A2(n_257_76_3687), .A3(
      n_257_76_3688), .A4(n_257_76_3631), .ZN(n_257_76_3915));
   NOR2_X1 i_257_76_3922 (.A1(n_257_76_3914), .A2(n_257_76_3915), .ZN(
      n_257_76_3916));
   NAND4_X1 i_257_76_3923 (.A1(n_257_76_3684), .A2(n_257_76_3602), .A3(
      n_257_76_3674), .A4(n_257_76_3623), .ZN(n_257_76_3917));
   INV_X1 i_257_76_3924 (.A(n_257_76_3917), .ZN(n_257_76_3918));
   NAND2_X1 i_257_76_3925 (.A1(n_257_76_3625), .A2(n_257_76_3626), .ZN(
      n_257_76_3919));
   NAND2_X1 i_257_76_3926 (.A1(n_257_278), .A2(n_257_423), .ZN(n_257_76_3920));
   NAND3_X1 i_257_76_3927 (.A1(n_257_76_3920), .A2(n_257_76_3627), .A3(
      n_257_76_3640), .ZN(n_257_76_3921));
   NOR2_X1 i_257_76_3928 (.A1(n_257_76_3919), .A2(n_257_76_3921), .ZN(
      n_257_76_3922));
   NAND4_X1 i_257_76_3929 (.A1(n_257_76_3916), .A2(n_257_76_3918), .A3(
      n_257_76_3922), .A4(n_257_76_3679), .ZN(n_257_76_3923));
   NAND2_X1 i_257_76_3930 (.A1(n_257_355), .A2(n_257_421), .ZN(n_257_76_3924));
   NAND3_X1 i_257_76_3931 (.A1(n_257_76_3630), .A2(n_257_76_3678), .A3(
      n_257_76_3924), .ZN(n_257_76_3925));
   NOR2_X1 i_257_76_3932 (.A1(n_257_76_3923), .A2(n_257_76_3925), .ZN(
      n_257_76_3926));
   NAND2_X1 i_257_76_3933 (.A1(n_257_76_3601), .A2(n_257_76_3681), .ZN(
      n_257_76_3927));
   INV_X1 i_257_76_3934 (.A(n_257_76_3927), .ZN(n_257_76_3928));
   NAND3_X1 i_257_76_3935 (.A1(n_257_76_3926), .A2(n_257_76_3600), .A3(
      n_257_76_3928), .ZN(n_257_76_3929));
   INV_X1 i_257_76_3936 (.A(n_257_76_3929), .ZN(n_257_76_3930));
   NAND2_X1 i_257_76_3937 (.A1(n_257_76_18073), .A2(n_257_76_3930), .ZN(
      n_257_76_3931));
   NAND2_X1 i_257_76_3938 (.A1(n_257_430), .A2(n_257_76_3616), .ZN(n_257_76_3932));
   INV_X1 i_257_76_3939 (.A(n_257_76_3932), .ZN(n_257_76_3933));
   NAND2_X1 i_257_76_3940 (.A1(n_257_76_3697), .A2(n_257_76_3933), .ZN(
      n_257_76_3934));
   INV_X1 i_257_76_3941 (.A(n_257_76_3934), .ZN(n_257_76_3935));
   NAND3_X1 i_257_76_3942 (.A1(n_257_76_3696), .A2(n_257_76_3632), .A3(
      n_257_76_3935), .ZN(n_257_76_3936));
   INV_X1 i_257_76_3943 (.A(n_257_76_3936), .ZN(n_257_76_3937));
   NAND3_X1 i_257_76_3944 (.A1(n_257_76_3816), .A2(n_257_76_3937), .A3(
      n_257_76_3631), .ZN(n_257_76_3938));
   NAND3_X1 i_257_76_3945 (.A1(n_257_76_3640), .A2(n_257_76_3641), .A3(
      n_257_76_3687), .ZN(n_257_76_3939));
   NOR2_X1 i_257_76_3946 (.A1(n_257_76_3938), .A2(n_257_76_3939), .ZN(
      n_257_76_3940));
   NAND3_X1 i_257_76_3947 (.A1(n_257_76_3602), .A2(n_257_76_3674), .A3(
      n_257_76_3623), .ZN(n_257_76_3941));
   INV_X1 i_257_76_3948 (.A(n_257_76_3941), .ZN(n_257_76_3942));
   NAND4_X1 i_257_76_3949 (.A1(n_257_76_3625), .A2(n_257_76_3626), .A3(n_257_119), 
      .A4(n_257_76_3627), .ZN(n_257_76_3943));
   INV_X1 i_257_76_3950 (.A(n_257_76_3943), .ZN(n_257_76_3944));
   NAND3_X1 i_257_76_3951 (.A1(n_257_76_3940), .A2(n_257_76_3942), .A3(
      n_257_76_3944), .ZN(n_257_76_3945));
   INV_X1 i_257_76_3952 (.A(n_257_76_3945), .ZN(n_257_76_3946));
   NAND2_X1 i_257_76_3953 (.A1(n_257_76_3630), .A2(n_257_76_3679), .ZN(
      n_257_76_3947));
   INV_X1 i_257_76_3954 (.A(n_257_76_3947), .ZN(n_257_76_3948));
   NAND3_X1 i_257_76_3955 (.A1(n_257_76_3946), .A2(n_257_76_3601), .A3(
      n_257_76_3948), .ZN(n_257_76_3949));
   NOR2_X1 i_257_76_3956 (.A1(n_257_76_3622), .A2(n_257_76_3949), .ZN(
      n_257_76_3950));
   NAND2_X1 i_257_76_3957 (.A1(n_257_76_18068), .A2(n_257_76_3950), .ZN(
      n_257_76_3951));
   NAND3_X1 i_257_76_3958 (.A1(n_257_76_3902), .A2(n_257_76_3931), .A3(
      n_257_76_3951), .ZN(n_257_76_3952));
   INV_X1 i_257_76_3959 (.A(n_257_76_3952), .ZN(n_257_76_3953));
   NAND3_X1 i_257_76_3960 (.A1(n_257_76_3602), .A2(n_257_76_3623), .A3(
      n_257_76_3626), .ZN(n_257_76_3954));
   NAND2_X1 i_257_76_3961 (.A1(n_257_76_3631), .A2(n_257_447), .ZN(n_257_76_3955));
   INV_X1 i_257_76_3962 (.A(n_257_76_3955), .ZN(n_257_76_3956));
   INV_X1 i_257_76_3963 (.A(n_257_771), .ZN(n_257_76_3957));
   NOR2_X1 i_257_76_3964 (.A1(n_257_76_3604), .A2(n_257_76_3957), .ZN(
      n_257_76_3958));
   NAND3_X1 i_257_76_3965 (.A1(n_257_76_3637), .A2(n_257_76_3638), .A3(
      n_257_76_3958), .ZN(n_257_76_3959));
   INV_X1 i_257_76_3966 (.A(n_257_76_3959), .ZN(n_257_76_3960));
   NAND3_X1 i_257_76_3967 (.A1(n_257_76_3956), .A2(n_257_76_3960), .A3(
      n_257_76_3627), .ZN(n_257_76_3961));
   NOR2_X1 i_257_76_3968 (.A1(n_257_76_3954), .A2(n_257_76_3961), .ZN(
      n_257_76_3962));
   NAND2_X1 i_257_76_3969 (.A1(n_257_76_3601), .A2(n_257_76_3962), .ZN(
      n_257_76_3963));
   INV_X1 i_257_76_3970 (.A(n_257_76_3963), .ZN(n_257_76_3964));
   NAND2_X1 i_257_76_3971 (.A1(n_257_76_3600), .A2(n_257_76_3964), .ZN(
      n_257_76_3965));
   INV_X1 i_257_76_3972 (.A(n_257_76_3965), .ZN(n_257_76_3966));
   NAND2_X1 i_257_76_3973 (.A1(n_257_81), .A2(n_257_76_3602), .ZN(n_257_76_3967));
   NAND3_X1 i_257_76_3974 (.A1(n_257_76_3674), .A2(n_257_76_3623), .A3(
      n_257_76_3625), .ZN(n_257_76_3968));
   NOR2_X1 i_257_76_3975 (.A1(n_257_76_3967), .A2(n_257_76_3968), .ZN(
      n_257_76_3969));
   NAND2_X1 i_257_76_3976 (.A1(n_257_431), .A2(n_257_76_3616), .ZN(n_257_76_3970));
   INV_X1 i_257_76_3977 (.A(n_257_76_3970), .ZN(n_257_76_3971));
   NAND2_X1 i_257_76_3978 (.A1(n_257_76_3697), .A2(n_257_76_3971), .ZN(
      n_257_76_3972));
   INV_X1 i_257_76_3979 (.A(n_257_76_3972), .ZN(n_257_76_3973));
   NAND3_X1 i_257_76_3980 (.A1(n_257_76_3696), .A2(n_257_76_3632), .A3(
      n_257_76_3973), .ZN(n_257_76_3974));
   INV_X1 i_257_76_3981 (.A(n_257_76_3974), .ZN(n_257_76_3975));
   NAND4_X1 i_257_76_3982 (.A1(n_257_76_3816), .A2(n_257_76_3975), .A3(
      n_257_76_3687), .A4(n_257_76_3631), .ZN(n_257_76_3976));
   NOR2_X1 i_257_76_3983 (.A1(n_257_76_3807), .A2(n_257_76_3976), .ZN(
      n_257_76_3977));
   NAND3_X1 i_257_76_3984 (.A1(n_257_76_3630), .A2(n_257_76_3969), .A3(
      n_257_76_3977), .ZN(n_257_76_3978));
   INV_X1 i_257_76_3985 (.A(n_257_76_3978), .ZN(n_257_76_3979));
   NAND2_X1 i_257_76_3986 (.A1(n_257_76_3979), .A2(n_257_76_3601), .ZN(
      n_257_76_3980));
   NOR2_X1 i_257_76_3987 (.A1(n_257_76_3980), .A2(n_257_76_3622), .ZN(
      n_257_76_3981));
   AOI22_X1 i_257_76_3988 (.A1(n_257_76_18085), .A2(n_257_76_3966), .B1(
      n_257_76_18080), .B2(n_257_76_3981), .ZN(n_257_76_3982));
   NAND3_X1 i_257_76_3989 (.A1(n_257_76_3889), .A2(n_257_76_3953), .A3(
      n_257_76_3982), .ZN(n_257_76_3983));
   INV_X1 i_257_76_3990 (.A(n_257_76_3723), .ZN(n_257_76_3984));
   NAND3_X1 i_257_76_3991 (.A1(n_257_76_3627), .A2(n_257_76_3641), .A3(
      n_257_76_3631), .ZN(n_257_76_3985));
   NAND4_X1 i_257_76_3992 (.A1(n_257_76_3637), .A2(n_257_76_3638), .A3(n_257_448), 
      .A4(n_257_76_3865), .ZN(n_257_76_3986));
   NOR2_X1 i_257_76_3993 (.A1(n_257_76_3985), .A2(n_257_76_3986), .ZN(
      n_257_76_3987));
   NAND3_X1 i_257_76_3994 (.A1(n_257_76_3984), .A2(n_257_675), .A3(n_257_76_3987), 
      .ZN(n_257_76_3988));
   INV_X1 i_257_76_3995 (.A(n_257_76_3988), .ZN(n_257_76_3989));
   NAND2_X1 i_257_76_3996 (.A1(n_257_76_3601), .A2(n_257_76_3989), .ZN(
      n_257_76_3990));
   INV_X1 i_257_76_3997 (.A(n_257_76_3990), .ZN(n_257_76_3991));
   NAND2_X1 i_257_76_3998 (.A1(n_257_76_3600), .A2(n_257_76_3991), .ZN(
      n_257_76_3992));
   INV_X1 i_257_76_3999 (.A(n_257_76_3992), .ZN(n_257_76_3993));
   NAND2_X1 i_257_76_4000 (.A1(n_257_76_18079), .A2(n_257_76_3993), .ZN(
      n_257_76_3994));
   NAND2_X1 i_257_76_4001 (.A1(n_257_425), .A2(n_257_76_3616), .ZN(n_257_76_3995));
   INV_X1 i_257_76_4002 (.A(n_257_76_3995), .ZN(n_257_76_3996));
   NAND3_X1 i_257_76_4003 (.A1(n_257_76_3697), .A2(n_257_76_3698), .A3(
      n_257_76_3996), .ZN(n_257_76_3997));
   NOR2_X1 i_257_76_4004 (.A1(n_257_76_3778), .A2(n_257_76_3997), .ZN(
      n_257_76_3998));
   NAND4_X1 i_257_76_4005 (.A1(n_257_76_3998), .A2(n_257_76_3637), .A3(
      n_257_76_3638), .A4(n_257_76_3696), .ZN(n_257_76_3999));
   NAND3_X1 i_257_76_4006 (.A1(n_257_76_3688), .A2(n_257_76_3631), .A3(
      n_257_76_3691), .ZN(n_257_76_4000));
   NOR2_X1 i_257_76_4007 (.A1(n_257_76_3999), .A2(n_257_76_4000), .ZN(
      n_257_76_4001));
   NAND3_X1 i_257_76_4008 (.A1(n_257_76_3623), .A2(n_257_76_3625), .A3(
      n_257_76_3626), .ZN(n_257_76_4002));
   INV_X1 i_257_76_4009 (.A(n_257_76_4002), .ZN(n_257_76_4003));
   NAND4_X1 i_257_76_4010 (.A1(n_257_76_3627), .A2(n_257_76_3640), .A3(
      n_257_76_3641), .A4(n_257_76_3687), .ZN(n_257_76_4004));
   INV_X1 i_257_76_4011 (.A(n_257_76_4004), .ZN(n_257_76_4005));
   NAND3_X1 i_257_76_4012 (.A1(n_257_76_4001), .A2(n_257_76_4003), .A3(
      n_257_76_4005), .ZN(n_257_76_4006));
   INV_X1 i_257_76_4013 (.A(n_257_76_4006), .ZN(n_257_76_4007));
   NAND3_X1 i_257_76_4014 (.A1(n_257_76_3740), .A2(n_257_76_3679), .A3(n_257_238), 
      .ZN(n_257_76_4008));
   INV_X1 i_257_76_4015 (.A(n_257_76_4008), .ZN(n_257_76_4009));
   NAND4_X1 i_257_76_4016 (.A1(n_257_76_4007), .A2(n_257_76_4009), .A3(
      n_257_76_3681), .A4(n_257_76_3630), .ZN(n_257_76_4010));
   INV_X1 i_257_76_4017 (.A(n_257_76_4010), .ZN(n_257_76_4011));
   NAND3_X1 i_257_76_4018 (.A1(n_257_76_4011), .A2(n_257_76_3600), .A3(
      n_257_76_3601), .ZN(n_257_76_4012));
   INV_X1 i_257_76_4019 (.A(n_257_76_4012), .ZN(n_257_76_4013));
   NAND2_X1 i_257_76_4020 (.A1(n_257_76_18064), .A2(n_257_76_4013), .ZN(
      n_257_76_4014));
   NAND2_X1 i_257_76_4021 (.A1(n_257_76_3600), .A2(n_257_76_3601), .ZN(
      n_257_76_4015));
   NAND2_X1 i_257_76_4022 (.A1(n_257_421), .A2(n_257_76_3616), .ZN(n_257_76_4016));
   INV_X1 i_257_76_4023 (.A(n_257_76_4016), .ZN(n_257_76_4017));
   NAND3_X1 i_257_76_4024 (.A1(n_257_76_3697), .A2(n_257_76_3698), .A3(
      n_257_76_4017), .ZN(n_257_76_4018));
   INV_X1 i_257_76_4025 (.A(n_257_76_4018), .ZN(n_257_76_4019));
   NAND3_X1 i_257_76_4026 (.A1(n_257_76_4019), .A2(n_257_76_3693), .A3(
      n_257_76_3632), .ZN(n_257_76_4020));
   INV_X1 i_257_76_4027 (.A(n_257_76_4020), .ZN(n_257_76_4021));
   NAND3_X1 i_257_76_4028 (.A1(n_257_76_3905), .A2(n_257_76_3907), .A3(
      n_257_76_4021), .ZN(n_257_76_4022));
   NOR2_X1 i_257_76_4029 (.A1(n_257_76_4022), .A2(n_257_76_3915), .ZN(
      n_257_76_4023));
   NAND3_X1 i_257_76_4030 (.A1(n_257_76_4023), .A2(n_257_76_3918), .A3(
      n_257_76_3922), .ZN(n_257_76_4024));
   INV_X1 i_257_76_4031 (.A(n_257_76_4024), .ZN(n_257_76_4025));
   INV_X1 i_257_76_4032 (.A(n_257_76_3678), .ZN(n_257_76_4026));
   NAND2_X1 i_257_76_4033 (.A1(n_257_76_3679), .A2(n_257_355), .ZN(n_257_76_4027));
   NOR2_X1 i_257_76_4034 (.A1(n_257_76_4026), .A2(n_257_76_4027), .ZN(
      n_257_76_4028));
   NAND3_X1 i_257_76_4035 (.A1(n_257_76_4025), .A2(n_257_76_3754), .A3(
      n_257_76_4028), .ZN(n_257_76_4029));
   NOR2_X1 i_257_76_4036 (.A1(n_257_76_4015), .A2(n_257_76_4029), .ZN(
      n_257_76_4030));
   NAND2_X1 i_257_76_4037 (.A1(n_257_76_18082), .A2(n_257_76_4030), .ZN(
      n_257_76_4031));
   NAND3_X1 i_257_76_4038 (.A1(n_257_76_3994), .A2(n_257_76_4014), .A3(
      n_257_76_4031), .ZN(n_257_76_4032));
   INV_X1 i_257_76_4039 (.A(n_257_76_4032), .ZN(n_257_76_4033));
   NAND4_X1 i_257_76_4040 (.A1(n_257_76_3687), .A2(n_257_76_3631), .A3(
      n_257_76_3637), .A4(n_257_76_3638), .ZN(n_257_76_4034));
   NOR2_X1 i_257_76_4041 (.A1(n_257_76_3676), .A2(n_257_76_4034), .ZN(
      n_257_76_4035));
   NAND4_X1 i_257_76_4042 (.A1(n_257_76_3674), .A2(n_257_76_3623), .A3(
      n_257_76_3625), .A4(n_257_76_3626), .ZN(n_257_76_4036));
   INV_X1 i_257_76_4043 (.A(n_257_76_4036), .ZN(n_257_76_4037));
   INV_X1 i_257_76_4044 (.A(n_257_571), .ZN(n_257_76_4038));
   NAND3_X1 i_257_76_4045 (.A1(n_257_76_3603), .A2(n_257_76_4038), .A3(n_257_442), 
      .ZN(n_257_76_4039));
   OAI21_X1 i_257_76_4046 (.A(n_257_76_4039), .B1(n_257_428), .B2(n_257_76_3604), 
      .ZN(n_257_76_4040));
   NAND3_X1 i_257_76_4047 (.A1(n_257_427), .A2(n_257_76_4040), .A3(n_257_76_3697), 
      .ZN(n_257_76_4041));
   INV_X1 i_257_76_4048 (.A(n_257_76_4041), .ZN(n_257_76_4042));
   NAND4_X1 i_257_76_4049 (.A1(n_257_76_4042), .A2(n_257_76_3696), .A3(n_257_198), 
      .A4(n_257_76_3632), .ZN(n_257_76_4043));
   INV_X1 i_257_76_4050 (.A(n_257_76_4043), .ZN(n_257_76_4044));
   NAND3_X1 i_257_76_4051 (.A1(n_257_76_3684), .A2(n_257_76_3602), .A3(
      n_257_76_4044), .ZN(n_257_76_4045));
   INV_X1 i_257_76_4052 (.A(n_257_76_4045), .ZN(n_257_76_4046));
   NAND4_X1 i_257_76_4053 (.A1(n_257_76_4035), .A2(n_257_76_4037), .A3(
      n_257_76_4046), .A4(n_257_76_3679), .ZN(n_257_76_4047));
   INV_X1 i_257_76_4054 (.A(n_257_76_4047), .ZN(n_257_76_4048));
   NAND3_X1 i_257_76_4055 (.A1(n_257_76_4048), .A2(n_257_76_3754), .A3(
      n_257_76_3601), .ZN(n_257_76_4049));
   NOR2_X1 i_257_76_4056 (.A1(n_257_76_4049), .A2(n_257_76_3622), .ZN(
      n_257_76_4050));
   NAND2_X1 i_257_76_4057 (.A1(n_257_76_18065), .A2(n_257_76_4050), .ZN(
      n_257_76_4051));
   NAND3_X1 i_257_76_4058 (.A1(n_257_76_3696), .A2(n_257_76_3865), .A3(n_257_458), 
      .ZN(n_257_76_4052));
   INV_X1 i_257_76_4059 (.A(n_257_76_4052), .ZN(n_257_76_4053));
   NAND3_X1 i_257_76_4060 (.A1(n_257_76_4053), .A2(n_257_76_3816), .A3(
      n_257_76_3631), .ZN(n_257_76_4054));
   NAND3_X1 i_257_76_4061 (.A1(n_257_76_3640), .A2(n_257_76_3641), .A3(n_257_451), 
      .ZN(n_257_76_4055));
   NOR2_X1 i_257_76_4062 (.A1(n_257_76_4054), .A2(n_257_76_4055), .ZN(
      n_257_76_4056));
   NAND3_X1 i_257_76_4063 (.A1(n_257_76_3629), .A2(n_257_76_3630), .A3(
      n_257_76_4056), .ZN(n_257_76_4057));
   INV_X1 i_257_76_4064 (.A(n_257_76_4057), .ZN(n_257_76_4058));
   NAND2_X1 i_257_76_4065 (.A1(n_257_76_4058), .A2(n_257_76_3601), .ZN(
      n_257_76_4059));
   NOR2_X1 i_257_76_4066 (.A1(n_257_76_3622), .A2(n_257_76_4059), .ZN(
      n_257_76_4060));
   NAND2_X1 i_257_76_4067 (.A1(n_257_76_18063), .A2(n_257_76_4060), .ZN(
      n_257_76_4061));
   NAND2_X1 i_257_76_4068 (.A1(n_257_76_3638), .A2(n_257_76_3696), .ZN(
      n_257_76_4062));
   INV_X1 i_257_76_4069 (.A(n_257_76_4062), .ZN(n_257_76_4063));
   NAND2_X1 i_257_76_4070 (.A1(n_257_76_3632), .A2(n_257_76_3697), .ZN(
      n_257_76_4064));
   NAND3_X1 i_257_76_4071 (.A1(n_257_507), .A2(n_257_76_4040), .A3(n_257_424), 
      .ZN(n_257_76_4065));
   NOR2_X1 i_257_76_4072 (.A1(n_257_76_4064), .A2(n_257_76_4065), .ZN(
      n_257_76_4066));
   NAND3_X1 i_257_76_4073 (.A1(n_257_76_3907), .A2(n_257_76_4063), .A3(
      n_257_76_4066), .ZN(n_257_76_4067));
   NOR2_X1 i_257_76_4074 (.A1(n_257_76_3915), .A2(n_257_76_4067), .ZN(
      n_257_76_4068));
   NAND4_X1 i_257_76_4075 (.A1(n_257_76_4068), .A2(n_257_76_3738), .A3(
      n_257_76_3740), .A4(n_257_76_3679), .ZN(n_257_76_4069));
   NAND2_X1 i_257_76_4076 (.A1(n_257_76_3630), .A2(n_257_76_3678), .ZN(
      n_257_76_4070));
   NOR2_X1 i_257_76_4077 (.A1(n_257_76_4069), .A2(n_257_76_4070), .ZN(
      n_257_76_4071));
   NAND3_X1 i_257_76_4078 (.A1(n_257_76_4071), .A2(n_257_76_3600), .A3(
      n_257_76_3928), .ZN(n_257_76_4072));
   INV_X1 i_257_76_4079 (.A(n_257_76_4072), .ZN(n_257_76_4073));
   NAND2_X1 i_257_76_4080 (.A1(n_257_76_18062), .A2(n_257_76_4073), .ZN(
      n_257_76_4074));
   NAND3_X1 i_257_76_4081 (.A1(n_257_76_4051), .A2(n_257_76_4061), .A3(
      n_257_76_4074), .ZN(n_257_76_4075));
   INV_X1 i_257_76_4082 (.A(n_257_76_4075), .ZN(n_257_76_4076));
   NAND3_X1 i_257_76_4083 (.A1(n_257_76_3697), .A2(n_257_76_4040), .A3(n_257_422), 
      .ZN(n_257_76_4077));
   INV_X1 i_257_76_4084 (.A(n_257_316), .ZN(n_257_76_4078));
   NOR2_X1 i_257_76_4085 (.A1(n_257_76_4077), .A2(n_257_76_4078), .ZN(
      n_257_76_4079));
   NAND3_X1 i_257_76_4086 (.A1(n_257_76_4079), .A2(n_257_76_3695), .A3(
      n_257_76_3696), .ZN(n_257_76_4080));
   INV_X1 i_257_76_4087 (.A(n_257_76_4080), .ZN(n_257_76_4081));
   NAND3_X1 i_257_76_4088 (.A1(n_257_76_4081), .A2(n_257_76_3684), .A3(
      n_257_76_3602), .ZN(n_257_76_4082));
   INV_X1 i_257_76_4089 (.A(n_257_76_4082), .ZN(n_257_76_4083));
   INV_X1 i_257_76_4090 (.A(n_257_76_3968), .ZN(n_257_76_4084));
   NAND4_X1 i_257_76_4091 (.A1(n_257_76_3626), .A2(n_257_76_3920), .A3(
      n_257_76_3627), .A4(n_257_76_3640), .ZN(n_257_76_4085));
   INV_X1 i_257_76_4092 (.A(n_257_76_4085), .ZN(n_257_76_4086));
   NAND3_X1 i_257_76_4093 (.A1(n_257_76_3641), .A2(n_257_76_3687), .A3(
      n_257_76_3688), .ZN(n_257_76_4087));
   NAND4_X1 i_257_76_4094 (.A1(n_257_76_3631), .A2(n_257_76_3691), .A3(
      n_257_76_3637), .A4(n_257_76_3638), .ZN(n_257_76_4088));
   NOR2_X1 i_257_76_4095 (.A1(n_257_76_4087), .A2(n_257_76_4088), .ZN(
      n_257_76_4089));
   NAND4_X1 i_257_76_4096 (.A1(n_257_76_4083), .A2(n_257_76_4084), .A3(
      n_257_76_4086), .A4(n_257_76_4089), .ZN(n_257_76_4090));
   NAND3_X1 i_257_76_4097 (.A1(n_257_76_3630), .A2(n_257_76_3678), .A3(
      n_257_76_3679), .ZN(n_257_76_4091));
   NOR2_X1 i_257_76_4098 (.A1(n_257_76_4090), .A2(n_257_76_4091), .ZN(
      n_257_76_4092));
   NAND3_X1 i_257_76_4099 (.A1(n_257_76_4092), .A2(n_257_76_3600), .A3(
      n_257_76_3928), .ZN(n_257_76_4093));
   INV_X1 i_257_76_4100 (.A(n_257_76_4093), .ZN(n_257_76_4094));
   NAND2_X1 i_257_76_4101 (.A1(n_257_342), .A2(n_257_76_4094), .ZN(n_257_76_4095));
   NAND2_X1 i_257_76_4102 (.A1(n_257_76_3924), .A2(n_257_76_3679), .ZN(
      n_257_76_4096));
   NOR2_X1 i_257_76_4103 (.A1(n_257_76_4070), .A2(n_257_76_4096), .ZN(
      n_257_76_4097));
   NAND2_X1 i_257_76_4104 (.A1(n_257_76_3631), .A2(n_257_76_3691), .ZN(
      n_257_76_4098));
   NOR2_X1 i_257_76_4105 (.A1(n_257_76_4098), .A2(n_257_76_3815), .ZN(
      n_257_76_4099));
   NAND3_X1 i_257_76_4106 (.A1(n_257_76_3616), .A2(n_257_394), .A3(n_257_484), 
      .ZN(n_257_76_4100));
   INV_X1 i_257_76_4107 (.A(n_257_76_4100), .ZN(n_257_76_4101));
   NAND2_X1 i_257_76_4108 (.A1(n_257_76_3698), .A2(n_257_76_4101), .ZN(
      n_257_76_4102));
   INV_X1 i_257_76_4109 (.A(n_257_76_4102), .ZN(n_257_76_4103));
   NAND2_X1 i_257_76_4110 (.A1(n_257_76_4103), .A2(n_257_76_3697), .ZN(
      n_257_76_4104));
   NAND2_X1 i_257_76_4111 (.A1(n_257_420), .A2(n_257_897), .ZN(n_257_76_4105));
   INV_X1 i_257_76_4112 (.A(n_257_76_4105), .ZN(n_257_76_4106));
   NOR2_X1 i_257_76_4113 (.A1(n_257_76_4104), .A2(n_257_76_4106), .ZN(
      n_257_76_4107));
   NAND2_X1 i_257_76_4114 (.A1(n_257_76_3695), .A2(n_257_76_4107), .ZN(
      n_257_76_4108));
   NAND2_X1 i_257_76_4115 (.A1(n_257_76_3903), .A2(n_257_76_3696), .ZN(
      n_257_76_4109));
   NOR2_X1 i_257_76_4116 (.A1(n_257_76_4108), .A2(n_257_76_4109), .ZN(
      n_257_76_4110));
   NAND2_X1 i_257_76_4117 (.A1(n_257_76_4099), .A2(n_257_76_4110), .ZN(
      n_257_76_4111));
   INV_X1 i_257_76_4118 (.A(n_257_76_4111), .ZN(n_257_76_4112));
   NAND2_X1 i_257_76_4119 (.A1(n_257_76_3687), .A2(n_257_76_3688), .ZN(
      n_257_76_4113));
   NOR2_X1 i_257_76_4120 (.A1(n_257_76_3642), .A2(n_257_76_4113), .ZN(
      n_257_76_4114));
   NAND2_X1 i_257_76_4121 (.A1(n_257_76_4112), .A2(n_257_76_4114), .ZN(
      n_257_76_4115));
   NAND2_X1 i_257_76_4122 (.A1(n_257_76_3684), .A2(n_257_76_3602), .ZN(
      n_257_76_4116));
   NAND2_X1 i_257_76_4123 (.A1(n_257_76_3674), .A2(n_257_76_3623), .ZN(
      n_257_76_4117));
   NOR2_X1 i_257_76_4124 (.A1(n_257_76_4116), .A2(n_257_76_4117), .ZN(
      n_257_76_4118));
   NAND2_X1 i_257_76_4125 (.A1(n_257_76_3920), .A2(n_257_76_3627), .ZN(
      n_257_76_4119));
   NOR2_X1 i_257_76_4126 (.A1(n_257_76_3919), .A2(n_257_76_4119), .ZN(
      n_257_76_4120));
   NAND2_X1 i_257_76_4127 (.A1(n_257_76_4118), .A2(n_257_76_4120), .ZN(
      n_257_76_4121));
   NOR2_X1 i_257_76_4128 (.A1(n_257_76_4115), .A2(n_257_76_4121), .ZN(
      n_257_76_4122));
   NAND2_X1 i_257_76_4129 (.A1(n_257_76_4097), .A2(n_257_76_4122), .ZN(
      n_257_76_4123));
   NAND2_X1 i_257_76_4130 (.A1(n_257_76_3600), .A2(n_257_76_3928), .ZN(
      n_257_76_4124));
   NOR2_X1 i_257_76_4131 (.A1(n_257_76_4123), .A2(n_257_76_4124), .ZN(
      n_257_76_4125));
   NAND2_X1 i_257_76_4132 (.A1(n_257_76_18060), .A2(n_257_76_4125), .ZN(
      n_257_76_4126));
   NAND2_X1 i_257_76_4133 (.A1(n_257_1033), .A2(n_257_76_17969), .ZN(
      n_257_76_4127));
   NAND2_X1 i_257_76_4134 (.A1(n_257_76_4010), .A2(n_257_76_4127), .ZN(
      n_257_76_4128));
   INV_X1 i_257_76_4135 (.A(n_257_76_4029), .ZN(n_257_76_4129));
   NOR2_X1 i_257_76_4136 (.A1(n_257_76_4128), .A2(n_257_76_4129), .ZN(
      n_257_76_4130));
   NAND2_X1 i_257_76_4137 (.A1(n_257_1001), .A2(n_257_76_17964), .ZN(
      n_257_76_4131));
   INV_X1 i_257_76_4138 (.A(n_257_76_4131), .ZN(n_257_76_4132));
   NAND2_X1 i_257_76_4139 (.A1(n_257_76_3788), .A2(n_257_76_3705), .ZN(
      n_257_76_4133));
   NOR2_X1 i_257_76_4140 (.A1(n_257_76_4132), .A2(n_257_76_4133), .ZN(
      n_257_76_4134));
   NAND2_X1 i_257_76_4141 (.A1(n_257_969), .A2(n_257_442), .ZN(n_257_76_4135));
   INV_X1 i_257_76_4142 (.A(n_257_76_4135), .ZN(n_257_76_4136));
   NAND2_X1 i_257_76_4143 (.A1(n_257_441), .A2(n_257_76_4136), .ZN(n_257_76_4137));
   NAND2_X1 i_257_76_4144 (.A1(n_257_76_4080), .A2(n_257_76_4137), .ZN(
      n_257_76_4138));
   NAND2_X1 i_257_76_4145 (.A1(n_257_119), .A2(n_257_76_17925), .ZN(
      n_257_76_4139));
   INV_X1 i_257_76_4146 (.A(n_257_76_4139), .ZN(n_257_76_4140));
   NOR2_X1 i_257_76_4147 (.A1(n_257_76_4138), .A2(n_257_76_4140), .ZN(
      n_257_76_4141));
   NAND2_X1 i_257_76_4148 (.A1(n_257_458), .A2(n_257_442), .ZN(n_257_76_4142));
   INV_X1 i_257_76_4149 (.A(n_257_76_4142), .ZN(n_257_76_4143));
   NAND2_X1 i_257_76_4150 (.A1(n_257_451), .A2(n_257_76_4143), .ZN(n_257_76_4144));
   NAND2_X1 i_257_76_4151 (.A1(n_257_803), .A2(n_257_76_17952), .ZN(
      n_257_76_4145));
   NAND2_X1 i_257_76_4152 (.A1(n_257_76_4144), .A2(n_257_76_4145), .ZN(
      n_257_76_4146));
   NAND2_X1 i_257_76_4153 (.A1(n_257_739), .A2(n_257_76_17935), .ZN(
      n_257_76_4147));
   NAND2_X1 i_257_76_4154 (.A1(n_257_76_4147), .A2(n_257_76_4043), .ZN(
      n_257_76_4148));
   NOR2_X1 i_257_76_4155 (.A1(n_257_76_4146), .A2(n_257_76_4148), .ZN(
      n_257_76_4149));
   NAND2_X1 i_257_76_4156 (.A1(n_257_76_4141), .A2(n_257_76_4149), .ZN(
      n_257_76_4150));
   INV_X1 i_257_76_4157 (.A(n_257_76_4150), .ZN(n_257_76_4151));
   NAND2_X1 i_257_76_4158 (.A1(n_257_635), .A2(n_257_76_17928), .ZN(
      n_257_76_4152));
   NAND2_X1 i_257_76_4159 (.A1(n_257_76_4152), .A2(n_257_76_4065), .ZN(
      n_257_76_4153));
   NAND2_X1 i_257_76_4160 (.A1(n_257_438), .A2(n_257_76_7160), .ZN(n_257_76_4154));
   INV_X1 i_257_76_4161 (.A(n_257_76_4154), .ZN(n_257_76_4155));
   NOR2_X1 i_257_76_4162 (.A1(n_257_76_4153), .A2(n_257_76_4155), .ZN(
      n_257_76_4156));
   NAND2_X1 i_257_76_4163 (.A1(n_257_76_15655), .A2(n_257_707), .ZN(
      n_257_76_4157));
   NAND2_X1 i_257_76_4164 (.A1(n_257_76_4157), .A2(n_257_76_3910), .ZN(
      n_257_76_4158));
   INV_X1 i_257_76_4165 (.A(Small_Packet_Data_Size[6]), .ZN(n_257_76_4159));
   NAND2_X1 i_257_76_4166 (.A1(n_257_76_4100), .A2(n_257_76_18051), .ZN(
      n_257_76_4160));
   NOR2_X1 i_257_76_4167 (.A1(n_257_76_4160), .A2(n_257_76_3745), .ZN(
      n_257_76_4161));
   NAND2_X1 i_257_76_4168 (.A1(n_257_603), .A2(n_257_442), .ZN(n_257_76_4162));
   INV_X1 i_257_76_4169 (.A(n_257_76_4162), .ZN(n_257_76_4163));
   NAND2_X1 i_257_76_4170 (.A1(n_257_432), .A2(n_257_76_4163), .ZN(n_257_76_4164));
   NAND2_X1 i_257_76_4171 (.A1(n_257_76_4161), .A2(n_257_76_4164), .ZN(
      n_257_76_4165));
   NOR2_X1 i_257_76_4172 (.A1(n_257_76_4158), .A2(n_257_76_4165), .ZN(
      n_257_76_4166));
   NAND2_X1 i_257_76_4173 (.A1(n_257_76_4156), .A2(n_257_76_4166), .ZN(
      n_257_76_4167));
   INV_X1 i_257_76_4174 (.A(n_257_76_4167), .ZN(n_257_76_4168));
   NAND3_X1 i_257_76_4175 (.A1(n_257_905), .A2(n_257_439), .A3(n_257_442), 
      .ZN(n_257_76_4169));
   NAND2_X1 i_257_76_4176 (.A1(n_257_937), .A2(n_257_442), .ZN(n_257_76_4170));
   INV_X1 i_257_76_4177 (.A(n_257_76_4170), .ZN(n_257_76_4171));
   NAND2_X1 i_257_76_4178 (.A1(n_257_440), .A2(n_257_76_4171), .ZN(n_257_76_4172));
   NAND2_X1 i_257_76_4179 (.A1(n_257_76_4169), .A2(n_257_76_4172), .ZN(
      n_257_76_4173));
   NAND2_X1 i_257_76_4180 (.A1(n_257_41), .A2(n_257_76_17918), .ZN(n_257_76_4174));
   INV_X1 i_257_76_4181 (.A(n_257_76_4174), .ZN(n_257_76_4175));
   NOR2_X1 i_257_76_4182 (.A1(n_257_76_4173), .A2(n_257_76_4175), .ZN(
      n_257_76_4176));
   NAND2_X1 i_257_76_4183 (.A1(n_257_76_4168), .A2(n_257_76_4176), .ZN(
      n_257_76_4177));
   NAND2_X1 i_257_76_4184 (.A1(n_257_835), .A2(n_257_442), .ZN(n_257_76_4178));
   INV_X1 i_257_76_4185 (.A(n_257_76_4178), .ZN(n_257_76_4179));
   AOI22_X1 i_257_76_4186 (.A1(n_257_867), .A2(n_257_76_17903), .B1(n_257_446), 
      .B2(n_257_76_4179), .ZN(n_257_76_4180));
   NAND2_X1 i_257_76_4187 (.A1(n_257_771), .A2(n_257_442), .ZN(n_257_76_4181));
   INV_X1 i_257_76_4188 (.A(n_257_76_4181), .ZN(n_257_76_4182));
   AOI22_X1 i_257_76_4189 (.A1(n_257_449), .A2(n_257_76_11546), .B1(n_257_447), 
      .B2(n_257_76_4182), .ZN(n_257_76_4183));
   NAND2_X1 i_257_76_4190 (.A1(n_257_76_4180), .A2(n_257_76_4183), .ZN(
      n_257_76_4184));
   NOR2_X1 i_257_76_4191 (.A1(n_257_76_4177), .A2(n_257_76_4184), .ZN(
      n_257_76_4185));
   NAND2_X1 i_257_76_4192 (.A1(n_257_76_4151), .A2(n_257_76_4185), .ZN(
      n_257_76_4186));
   AOI22_X1 i_257_76_4193 (.A1(n_257_675), .A2(n_257_76_17958), .B1(n_257_81), 
      .B2(n_257_76_17932), .ZN(n_257_76_4187));
   NAND2_X1 i_257_76_4194 (.A1(n_257_158), .A2(n_257_76_17331), .ZN(
      n_257_76_4188));
   NAND2_X1 i_257_76_4195 (.A1(n_257_76_4187), .A2(n_257_76_4188), .ZN(
      n_257_76_4189));
   NOR2_X1 i_257_76_4196 (.A1(n_257_76_4186), .A2(n_257_76_4189), .ZN(
      n_257_76_4190));
   NAND2_X1 i_257_76_4197 (.A1(n_257_76_4134), .A2(n_257_76_4190), .ZN(
      n_257_76_4191));
   INV_X1 i_257_76_4198 (.A(n_257_76_4191), .ZN(n_257_76_4192));
   NAND2_X1 i_257_76_4199 (.A1(n_257_76_4130), .A2(n_257_76_4192), .ZN(
      n_257_76_4193));
   NAND3_X1 i_257_76_4200 (.A1(n_257_76_4095), .A2(n_257_76_4126), .A3(
      n_257_76_4193), .ZN(n_257_76_4194));
   INV_X1 i_257_76_4201 (.A(n_257_76_4194), .ZN(n_257_76_4195));
   NAND3_X1 i_257_76_4202 (.A1(n_257_76_4033), .A2(n_257_76_4076), .A3(
      n_257_76_4195), .ZN(n_257_76_4196));
   NOR2_X1 i_257_76_4203 (.A1(n_257_76_3983), .A2(n_257_76_4196), .ZN(
      n_257_76_4197));
   NAND2_X1 i_257_76_4204 (.A1(n_257_76_3849), .A2(n_257_76_4197), .ZN(n_6));
   NAND2_X1 i_257_76_4205 (.A1(n_257_1002), .A2(n_257_444), .ZN(n_257_76_4198));
   NAND2_X1 i_257_76_4206 (.A1(n_257_441), .A2(n_257_970), .ZN(n_257_76_4199));
   INV_X1 i_257_76_4207 (.A(n_257_1066), .ZN(n_257_76_4200));
   NAND2_X1 i_257_76_4208 (.A1(n_257_76_4200), .A2(n_257_442), .ZN(n_257_76_4201));
   INV_X1 i_257_76_4209 (.A(n_257_938), .ZN(n_257_76_4202));
   NOR2_X1 i_257_76_4210 (.A1(n_257_76_4201), .A2(n_257_76_4202), .ZN(
      n_257_76_4203));
   NAND2_X1 i_257_76_4211 (.A1(n_257_440), .A2(n_257_76_4203), .ZN(n_257_76_4204));
   INV_X1 i_257_76_4212 (.A(n_257_76_4204), .ZN(n_257_76_4205));
   NAND2_X1 i_257_76_4213 (.A1(n_257_76_4199), .A2(n_257_76_4205), .ZN(
      n_257_76_4206));
   INV_X1 i_257_76_4214 (.A(n_257_76_4206), .ZN(n_257_76_4207));
   NAND2_X1 i_257_76_4215 (.A1(n_257_76_4198), .A2(n_257_76_4207), .ZN(
      n_257_76_4208));
   INV_X1 i_257_76_4216 (.A(n_257_76_4208), .ZN(n_257_76_4209));
   NAND2_X1 i_257_76_4217 (.A1(n_257_1034), .A2(n_257_443), .ZN(n_257_76_4210));
   NAND2_X1 i_257_76_4218 (.A1(n_257_76_4209), .A2(n_257_76_4210), .ZN(
      n_257_76_4211));
   INV_X1 i_257_76_4219 (.A(n_257_76_4211), .ZN(n_257_76_4212));
   NAND2_X1 i_257_76_4220 (.A1(n_257_17), .A2(n_257_76_4212), .ZN(n_257_76_4213));
   INV_X1 i_257_76_4221 (.A(n_257_76_4201), .ZN(n_257_76_4214));
   NAND2_X1 i_257_76_4222 (.A1(n_257_443), .A2(n_257_76_4214), .ZN(n_257_76_4215));
   INV_X1 i_257_76_4223 (.A(n_257_76_4215), .ZN(n_257_76_4216));
   NAND2_X1 i_257_76_4224 (.A1(n_257_1034), .A2(n_257_76_4216), .ZN(
      n_257_76_4217));
   INV_X1 i_257_76_4225 (.A(n_257_76_4217), .ZN(n_257_76_4218));
   NAND2_X1 i_257_76_4226 (.A1(n_257_76_18072), .A2(n_257_76_4218), .ZN(
      n_257_76_4219));
   NAND2_X1 i_257_76_4227 (.A1(n_257_868), .A2(n_257_445), .ZN(n_257_76_4220));
   NAND2_X1 i_257_76_4228 (.A1(n_257_76_4199), .A2(n_257_76_4220), .ZN(
      n_257_76_4221));
   NAND2_X1 i_257_76_4229 (.A1(n_257_740), .A2(n_257_436), .ZN(n_257_76_4222));
   NAND2_X1 i_257_76_4230 (.A1(n_257_804), .A2(n_257_437), .ZN(n_257_76_4223));
   NAND2_X1 i_257_76_4231 (.A1(n_257_446), .A2(n_257_836), .ZN(n_257_76_4224));
   NAND3_X1 i_257_76_4232 (.A1(n_257_76_4222), .A2(n_257_76_4223), .A3(
      n_257_76_4224), .ZN(n_257_76_4225));
   NOR2_X1 i_257_76_4233 (.A1(n_257_76_4221), .A2(n_257_76_4225), .ZN(
      n_257_76_4226));
   NAND2_X1 i_257_76_4234 (.A1(n_257_676), .A2(n_257_448), .ZN(n_257_76_4227));
   NAND2_X1 i_257_76_4235 (.A1(n_257_906), .A2(n_257_439), .ZN(n_257_76_4228));
   NAND2_X1 i_257_76_4236 (.A1(n_257_708), .A2(n_257_435), .ZN(n_257_76_4229));
   NAND2_X1 i_257_76_4237 (.A1(n_257_450), .A2(n_257_76_4214), .ZN(n_257_76_4230));
   INV_X1 i_257_76_4238 (.A(n_257_76_4230), .ZN(n_257_76_4231));
   NAND3_X1 i_257_76_4239 (.A1(n_257_76_4229), .A2(n_257_636), .A3(n_257_76_4231), 
      .ZN(n_257_76_4232));
   INV_X1 i_257_76_4240 (.A(n_257_76_4232), .ZN(n_257_76_4233));
   NAND2_X1 i_257_76_4241 (.A1(n_257_440), .A2(n_257_938), .ZN(n_257_76_4234));
   NAND2_X1 i_257_76_4242 (.A1(n_257_438), .A2(n_257_1072), .ZN(n_257_76_4235));
   NAND4_X1 i_257_76_4243 (.A1(n_257_76_4228), .A2(n_257_76_4233), .A3(
      n_257_76_4234), .A4(n_257_76_4235), .ZN(n_257_76_4236));
   NAND2_X1 i_257_76_4244 (.A1(n_257_449), .A2(n_257_1080), .ZN(n_257_76_4237));
   NAND2_X1 i_257_76_4245 (.A1(n_257_447), .A2(n_257_772), .ZN(n_257_76_4238));
   NAND2_X1 i_257_76_4246 (.A1(n_257_76_4237), .A2(n_257_76_4238), .ZN(
      n_257_76_4239));
   NOR2_X1 i_257_76_4247 (.A1(n_257_76_4236), .A2(n_257_76_4239), .ZN(
      n_257_76_4240));
   NAND3_X1 i_257_76_4248 (.A1(n_257_76_4226), .A2(n_257_76_4227), .A3(
      n_257_76_4240), .ZN(n_257_76_4241));
   INV_X1 i_257_76_4249 (.A(n_257_76_4241), .ZN(n_257_76_4242));
   NAND2_X1 i_257_76_4250 (.A1(n_257_76_4242), .A2(n_257_76_4198), .ZN(
      n_257_76_4243));
   INV_X1 i_257_76_4251 (.A(n_257_76_4210), .ZN(n_257_76_4244));
   NOR2_X1 i_257_76_4252 (.A1(n_257_76_4243), .A2(n_257_76_4244), .ZN(
      n_257_76_4245));
   NAND2_X1 i_257_76_4253 (.A1(n_257_28), .A2(n_257_76_4245), .ZN(n_257_76_4246));
   NAND3_X1 i_257_76_4254 (.A1(n_257_76_4213), .A2(n_257_76_4219), .A3(
      n_257_76_4246), .ZN(n_257_76_4247));
   NAND2_X1 i_257_76_4255 (.A1(n_257_76_4228), .A2(n_257_446), .ZN(n_257_76_4248));
   INV_X1 i_257_76_4256 (.A(n_257_76_4248), .ZN(n_257_76_4249));
   NAND2_X1 i_257_76_4257 (.A1(n_257_836), .A2(n_257_76_4214), .ZN(n_257_76_4250));
   INV_X1 i_257_76_4258 (.A(n_257_76_4250), .ZN(n_257_76_4251));
   NAND3_X1 i_257_76_4259 (.A1(n_257_76_4234), .A2(n_257_76_4235), .A3(
      n_257_76_4251), .ZN(n_257_76_4252));
   INV_X1 i_257_76_4260 (.A(n_257_76_4252), .ZN(n_257_76_4253));
   NAND4_X1 i_257_76_4261 (.A1(n_257_76_4199), .A2(n_257_76_4220), .A3(
      n_257_76_4249), .A4(n_257_76_4253), .ZN(n_257_76_4254));
   INV_X1 i_257_76_4262 (.A(n_257_76_4254), .ZN(n_257_76_4255));
   NAND2_X1 i_257_76_4263 (.A1(n_257_76_4198), .A2(n_257_76_4255), .ZN(
      n_257_76_4256));
   INV_X1 i_257_76_4264 (.A(n_257_76_4256), .ZN(n_257_76_4257));
   NAND2_X1 i_257_76_4265 (.A1(n_257_76_4257), .A2(n_257_76_4210), .ZN(
      n_257_76_4258));
   INV_X1 i_257_76_4266 (.A(n_257_76_4258), .ZN(n_257_76_4259));
   NAND2_X1 i_257_76_4267 (.A1(n_257_76_18070), .A2(n_257_76_4259), .ZN(
      n_257_76_4260));
   NAND2_X1 i_257_76_4268 (.A1(n_257_439), .A2(n_257_76_4214), .ZN(n_257_76_4261));
   INV_X1 i_257_76_4269 (.A(n_257_76_4261), .ZN(n_257_76_4262));
   NAND3_X1 i_257_76_4270 (.A1(n_257_76_4262), .A2(n_257_76_4234), .A3(n_257_906), 
      .ZN(n_257_76_4263));
   INV_X1 i_257_76_4271 (.A(n_257_76_4263), .ZN(n_257_76_4264));
   NAND2_X1 i_257_76_4272 (.A1(n_257_76_4199), .A2(n_257_76_4264), .ZN(
      n_257_76_4265));
   INV_X1 i_257_76_4273 (.A(n_257_76_4265), .ZN(n_257_76_4266));
   NAND2_X1 i_257_76_4274 (.A1(n_257_76_4198), .A2(n_257_76_4266), .ZN(
      n_257_76_4267));
   INV_X1 i_257_76_4275 (.A(n_257_76_4267), .ZN(n_257_76_4268));
   NAND2_X1 i_257_76_4276 (.A1(n_257_76_4268), .A2(n_257_76_4210), .ZN(
      n_257_76_4269));
   INV_X1 i_257_76_4277 (.A(n_257_76_4269), .ZN(n_257_76_4270));
   NAND2_X1 i_257_76_4278 (.A1(n_257_76_18084), .A2(n_257_76_4270), .ZN(
      n_257_76_4271));
   NAND2_X1 i_257_76_4279 (.A1(n_257_451), .A2(n_257_459), .ZN(n_257_76_4272));
   NAND2_X1 i_257_76_4280 (.A1(n_257_76_4199), .A2(n_257_76_4272), .ZN(
      n_257_76_4273));
   NAND3_X1 i_257_76_4281 (.A1(n_257_76_4224), .A2(n_257_76_4237), .A3(
      n_257_76_4238), .ZN(n_257_76_4274));
   NOR2_X1 i_257_76_4282 (.A1(n_257_76_4273), .A2(n_257_76_4274), .ZN(
      n_257_76_4275));
   NAND2_X1 i_257_76_4283 (.A1(n_257_159), .A2(n_257_429), .ZN(n_257_76_4276));
   NAND2_X1 i_257_76_4284 (.A1(n_257_82), .A2(n_257_431), .ZN(n_257_76_4277));
   NAND3_X1 i_257_76_4285 (.A1(n_257_76_4275), .A2(n_257_76_4276), .A3(
      n_257_76_4277), .ZN(n_257_76_4278));
   NAND2_X1 i_257_76_4286 (.A1(n_257_239), .A2(n_257_425), .ZN(n_257_76_4279));
   NAND2_X1 i_257_76_4287 (.A1(n_257_76_4227), .A2(n_257_76_4279), .ZN(
      n_257_76_4280));
   NOR2_X1 i_257_76_4288 (.A1(n_257_76_4278), .A2(n_257_76_4280), .ZN(
      n_257_76_4281));
   NAND2_X1 i_257_76_4289 (.A1(n_257_120), .A2(n_257_430), .ZN(n_257_76_4282));
   NAND2_X1 i_257_76_4290 (.A1(n_257_76_4220), .A2(n_257_76_4282), .ZN(
      n_257_76_4283));
   INV_X1 i_257_76_4291 (.A(n_257_76_4283), .ZN(n_257_76_4284));
   NAND2_X1 i_257_76_4292 (.A1(n_257_199), .A2(n_257_427), .ZN(n_257_76_4285));
   NAND3_X1 i_257_76_4293 (.A1(n_257_76_4234), .A2(n_257_76_4235), .A3(
      n_257_76_4285), .ZN(n_257_76_4286));
   NAND2_X1 i_257_76_4294 (.A1(n_257_636), .A2(n_257_450), .ZN(n_257_76_4287));
   NAND2_X1 i_257_76_4295 (.A1(n_257_432), .A2(n_257_604), .ZN(n_257_76_4288));
   NAND2_X1 i_257_76_4296 (.A1(n_257_428), .A2(n_257_572), .ZN(n_257_76_4289));
   NAND2_X1 i_257_76_4297 (.A1(n_257_423), .A2(n_257_76_4214), .ZN(n_257_76_4290));
   INV_X1 i_257_76_4298 (.A(n_257_76_4290), .ZN(n_257_76_4291));
   NAND3_X1 i_257_76_4299 (.A1(n_257_76_4288), .A2(n_257_76_4289), .A3(
      n_257_76_4291), .ZN(n_257_76_4292));
   INV_X1 i_257_76_4300 (.A(n_257_76_4292), .ZN(n_257_76_4293));
   NAND2_X1 i_257_76_4301 (.A1(n_257_508), .A2(n_257_424), .ZN(n_257_76_4294));
   NAND4_X1 i_257_76_4302 (.A1(n_257_76_4287), .A2(n_257_76_4293), .A3(
      n_257_76_4294), .A4(n_257_76_4229), .ZN(n_257_76_4295));
   NOR2_X1 i_257_76_4303 (.A1(n_257_76_4286), .A2(n_257_76_4295), .ZN(
      n_257_76_4296));
   NAND2_X1 i_257_76_4304 (.A1(n_257_540), .A2(n_257_426), .ZN(n_257_76_4297));
   NAND2_X1 i_257_76_4305 (.A1(n_257_42), .A2(n_257_433), .ZN(n_257_76_4298));
   NAND4_X1 i_257_76_4306 (.A1(n_257_76_4297), .A2(n_257_279), .A3(n_257_76_4298), 
      .A4(n_257_76_4228), .ZN(n_257_76_4299));
   INV_X1 i_257_76_4307 (.A(n_257_76_4299), .ZN(n_257_76_4300));
   NAND2_X1 i_257_76_4308 (.A1(n_257_76_4222), .A2(n_257_76_4223), .ZN(
      n_257_76_4301));
   INV_X1 i_257_76_4309 (.A(n_257_76_4301), .ZN(n_257_76_4302));
   NAND4_X1 i_257_76_4310 (.A1(n_257_76_4284), .A2(n_257_76_4296), .A3(
      n_257_76_4300), .A4(n_257_76_4302), .ZN(n_257_76_4303));
   INV_X1 i_257_76_4311 (.A(n_257_76_4303), .ZN(n_257_76_4304));
   NAND2_X1 i_257_76_4312 (.A1(n_257_76_4198), .A2(n_257_76_4304), .ZN(
      n_257_76_4305));
   INV_X1 i_257_76_4313 (.A(n_257_76_4305), .ZN(n_257_76_4306));
   NAND3_X1 i_257_76_4314 (.A1(n_257_76_4281), .A2(n_257_76_4306), .A3(
      n_257_76_4210), .ZN(n_257_76_4307));
   INV_X1 i_257_76_4315 (.A(n_257_76_4307), .ZN(n_257_76_4308));
   NAND2_X1 i_257_76_4316 (.A1(n_257_76_18066), .A2(n_257_76_4308), .ZN(
      n_257_76_4309));
   NAND3_X1 i_257_76_4317 (.A1(n_257_76_4260), .A2(n_257_76_4271), .A3(
      n_257_76_4309), .ZN(n_257_76_4310));
   NOR2_X1 i_257_76_4318 (.A1(n_257_76_4247), .A2(n_257_76_4310), .ZN(
      n_257_76_4311));
   NAND2_X1 i_257_76_4319 (.A1(n_257_970), .A2(n_257_76_4214), .ZN(n_257_76_4312));
   INV_X1 i_257_76_4320 (.A(n_257_76_4312), .ZN(n_257_76_4313));
   NAND2_X1 i_257_76_4321 (.A1(n_257_441), .A2(n_257_76_4313), .ZN(n_257_76_4314));
   INV_X1 i_257_76_4322 (.A(n_257_76_4314), .ZN(n_257_76_4315));
   NAND2_X1 i_257_76_4323 (.A1(n_257_76_4198), .A2(n_257_76_4315), .ZN(
      n_257_76_4316));
   INV_X1 i_257_76_4324 (.A(n_257_76_4316), .ZN(n_257_76_4317));
   NAND2_X1 i_257_76_4325 (.A1(n_257_76_4317), .A2(n_257_76_4210), .ZN(
      n_257_76_4318));
   INV_X1 i_257_76_4326 (.A(n_257_76_4318), .ZN(n_257_76_4319));
   NAND2_X1 i_257_76_4327 (.A1(n_257_76_18071), .A2(n_257_76_4319), .ZN(
      n_257_76_4320));
   NAND4_X1 i_257_76_4328 (.A1(n_257_76_4199), .A2(n_257_76_4220), .A3(
      n_257_76_4222), .A4(n_257_76_4223), .ZN(n_257_76_4321));
   INV_X1 i_257_76_4329 (.A(n_257_708), .ZN(n_257_76_4322));
   NAND2_X1 i_257_76_4330 (.A1(n_257_435), .A2(n_257_76_4214), .ZN(n_257_76_4323));
   NOR2_X1 i_257_76_4331 (.A1(n_257_76_4322), .A2(n_257_76_4323), .ZN(
      n_257_76_4324));
   NAND3_X1 i_257_76_4332 (.A1(n_257_76_4234), .A2(n_257_76_4235), .A3(
      n_257_76_4324), .ZN(n_257_76_4325));
   INV_X1 i_257_76_4333 (.A(n_257_76_4325), .ZN(n_257_76_4326));
   NAND4_X1 i_257_76_4334 (.A1(n_257_76_4326), .A2(n_257_76_4224), .A3(
      n_257_76_4238), .A4(n_257_76_4228), .ZN(n_257_76_4327));
   NOR2_X1 i_257_76_4335 (.A1(n_257_76_4321), .A2(n_257_76_4327), .ZN(
      n_257_76_4328));
   NAND2_X1 i_257_76_4336 (.A1(n_257_76_4198), .A2(n_257_76_4328), .ZN(
      n_257_76_4329));
   INV_X1 i_257_76_4337 (.A(n_257_76_4329), .ZN(n_257_76_4330));
   NAND2_X1 i_257_76_4338 (.A1(n_257_76_4330), .A2(n_257_76_4210), .ZN(
      n_257_76_4331));
   INV_X1 i_257_76_4339 (.A(n_257_76_4331), .ZN(n_257_76_4332));
   NAND2_X1 i_257_76_4340 (.A1(n_257_76_18078), .A2(n_257_76_4332), .ZN(
      n_257_76_4333));
   NAND2_X1 i_257_76_4341 (.A1(n_257_76_4234), .A2(n_257_76_4235), .ZN(
      n_257_76_4334));
   INV_X1 i_257_76_4342 (.A(n_257_76_4334), .ZN(n_257_76_4335));
   NAND3_X1 i_257_76_4343 (.A1(n_257_76_4200), .A2(n_257_442), .A3(n_257_572), 
      .ZN(n_257_76_4336));
   INV_X1 i_257_76_4344 (.A(n_257_76_4336), .ZN(n_257_76_4337));
   NAND2_X1 i_257_76_4345 (.A1(n_257_428), .A2(n_257_76_4337), .ZN(n_257_76_4338));
   INV_X1 i_257_76_4346 (.A(n_257_76_4338), .ZN(n_257_76_4339));
   NAND2_X1 i_257_76_4347 (.A1(n_257_76_4288), .A2(n_257_76_4339), .ZN(
      n_257_76_4340));
   INV_X1 i_257_76_4348 (.A(n_257_76_4340), .ZN(n_257_76_4341));
   NAND3_X1 i_257_76_4349 (.A1(n_257_76_4287), .A2(n_257_76_4229), .A3(
      n_257_76_4341), .ZN(n_257_76_4342));
   INV_X1 i_257_76_4350 (.A(n_257_76_4342), .ZN(n_257_76_4343));
   NAND3_X1 i_257_76_4351 (.A1(n_257_76_4335), .A2(n_257_76_4343), .A3(
      n_257_76_4228), .ZN(n_257_76_4344));
   NAND3_X1 i_257_76_4352 (.A1(n_257_76_4237), .A2(n_257_76_4238), .A3(
      n_257_76_4298), .ZN(n_257_76_4345));
   NOR2_X1 i_257_76_4353 (.A1(n_257_76_4344), .A2(n_257_76_4345), .ZN(
      n_257_76_4346));
   NAND4_X1 i_257_76_4354 (.A1(n_257_76_4282), .A2(n_257_76_4222), .A3(
      n_257_76_4223), .A4(n_257_76_4224), .ZN(n_257_76_4347));
   INV_X1 i_257_76_4355 (.A(n_257_76_4347), .ZN(n_257_76_4348));
   NAND3_X1 i_257_76_4356 (.A1(n_257_76_4199), .A2(n_257_76_4272), .A3(
      n_257_76_4220), .ZN(n_257_76_4349));
   INV_X1 i_257_76_4357 (.A(n_257_76_4349), .ZN(n_257_76_4350));
   NAND4_X1 i_257_76_4358 (.A1(n_257_76_4346), .A2(n_257_76_4348), .A3(
      n_257_76_4350), .A4(n_257_76_4277), .ZN(n_257_76_4351));
   NAND2_X1 i_257_76_4359 (.A1(n_257_76_4227), .A2(n_257_76_4276), .ZN(
      n_257_76_4352));
   NOR2_X1 i_257_76_4360 (.A1(n_257_76_4351), .A2(n_257_76_4352), .ZN(
      n_257_76_4353));
   NAND3_X1 i_257_76_4361 (.A1(n_257_76_4353), .A2(n_257_76_4210), .A3(
      n_257_76_4198), .ZN(n_257_76_4354));
   INV_X1 i_257_76_4362 (.A(n_257_76_4354), .ZN(n_257_76_4355));
   NAND2_X1 i_257_76_4363 (.A1(n_257_76_18074), .A2(n_257_76_4355), .ZN(
      n_257_76_4356));
   NAND3_X1 i_257_76_4364 (.A1(n_257_76_4320), .A2(n_257_76_4333), .A3(
      n_257_76_4356), .ZN(n_257_76_4357));
   NAND2_X1 i_257_76_4365 (.A1(n_257_1066), .A2(n_257_442), .ZN(n_257_76_4358));
   INV_X1 i_257_76_4366 (.A(n_257_76_4358), .ZN(n_257_76_4359));
   NAND2_X1 i_257_76_4367 (.A1(n_257_13), .A2(n_257_76_4359), .ZN(n_257_76_4360));
   NAND2_X1 i_257_76_4368 (.A1(n_257_868), .A2(n_257_76_4228), .ZN(n_257_76_4361));
   INV_X1 i_257_76_4369 (.A(n_257_76_4361), .ZN(n_257_76_4362));
   NAND2_X1 i_257_76_4370 (.A1(n_257_445), .A2(n_257_76_4214), .ZN(n_257_76_4363));
   INV_X1 i_257_76_4371 (.A(n_257_76_4363), .ZN(n_257_76_4364));
   NAND3_X1 i_257_76_4372 (.A1(n_257_76_4234), .A2(n_257_76_4235), .A3(
      n_257_76_4364), .ZN(n_257_76_4365));
   INV_X1 i_257_76_4373 (.A(n_257_76_4365), .ZN(n_257_76_4366));
   NAND3_X1 i_257_76_4374 (.A1(n_257_76_4362), .A2(n_257_76_4199), .A3(
      n_257_76_4366), .ZN(n_257_76_4367));
   INV_X1 i_257_76_4375 (.A(n_257_76_4367), .ZN(n_257_76_4368));
   NAND2_X1 i_257_76_4376 (.A1(n_257_76_4198), .A2(n_257_76_4368), .ZN(
      n_257_76_4369));
   INV_X1 i_257_76_4377 (.A(n_257_76_4369), .ZN(n_257_76_4370));
   NAND2_X1 i_257_76_4378 (.A1(n_257_76_4370), .A2(n_257_76_4210), .ZN(
      n_257_76_4371));
   INV_X1 i_257_76_4379 (.A(n_257_76_4371), .ZN(n_257_76_4372));
   NAND2_X1 i_257_76_4380 (.A1(n_257_76_18077), .A2(n_257_76_4372), .ZN(
      n_257_76_4373));
   NAND2_X1 i_257_76_4381 (.A1(n_257_76_4360), .A2(n_257_76_4373), .ZN(
      n_257_76_4374));
   NOR2_X1 i_257_76_4382 (.A1(n_257_76_4357), .A2(n_257_76_4374), .ZN(
      n_257_76_4375));
   INV_X1 i_257_76_4383 (.A(n_257_76_4198), .ZN(n_257_76_4376));
   INV_X1 i_257_76_4384 (.A(n_257_76_4229), .ZN(n_257_76_4377));
   NAND2_X1 i_257_76_4385 (.A1(n_257_426), .A2(n_257_76_4214), .ZN(n_257_76_4378));
   INV_X1 i_257_76_4386 (.A(n_257_76_4378), .ZN(n_257_76_4379));
   NAND3_X1 i_257_76_4387 (.A1(n_257_76_4288), .A2(n_257_76_4289), .A3(
      n_257_76_4379), .ZN(n_257_76_4380));
   NOR2_X1 i_257_76_4388 (.A1(n_257_76_4377), .A2(n_257_76_4380), .ZN(
      n_257_76_4381));
   NAND4_X1 i_257_76_4389 (.A1(n_257_76_4381), .A2(n_257_540), .A3(n_257_76_4285), 
      .A4(n_257_76_4287), .ZN(n_257_76_4382));
   NAND3_X1 i_257_76_4390 (.A1(n_257_76_4228), .A2(n_257_76_4234), .A3(
      n_257_76_4235), .ZN(n_257_76_4383));
   NOR2_X1 i_257_76_4391 (.A1(n_257_76_4382), .A2(n_257_76_4383), .ZN(
      n_257_76_4384));
   NAND3_X1 i_257_76_4392 (.A1(n_257_76_4222), .A2(n_257_76_4223), .A3(
      n_257_76_4298), .ZN(n_257_76_4385));
   INV_X1 i_257_76_4393 (.A(n_257_76_4385), .ZN(n_257_76_4386));
   NAND3_X1 i_257_76_4394 (.A1(n_257_76_4384), .A2(n_257_76_4284), .A3(
      n_257_76_4386), .ZN(n_257_76_4387));
   NOR2_X1 i_257_76_4395 (.A1(n_257_76_4376), .A2(n_257_76_4387), .ZN(
      n_257_76_4388));
   NAND4_X1 i_257_76_4396 (.A1(n_257_76_4227), .A2(n_257_76_4275), .A3(
      n_257_76_4276), .A4(n_257_76_4277), .ZN(n_257_76_4389));
   INV_X1 i_257_76_4397 (.A(n_257_76_4389), .ZN(n_257_76_4390));
   NAND3_X1 i_257_76_4398 (.A1(n_257_76_4388), .A2(n_257_76_4210), .A3(
      n_257_76_4390), .ZN(n_257_76_4391));
   INV_X1 i_257_76_4399 (.A(n_257_76_4391), .ZN(n_257_76_4392));
   NAND2_X1 i_257_76_4400 (.A1(n_257_76_18076), .A2(n_257_76_4392), .ZN(
      n_257_76_4393));
   NAND2_X1 i_257_76_4401 (.A1(n_257_740), .A2(n_257_76_4228), .ZN(n_257_76_4394));
   INV_X1 i_257_76_4402 (.A(n_257_76_4394), .ZN(n_257_76_4395));
   NAND2_X1 i_257_76_4403 (.A1(n_257_436), .A2(n_257_76_4214), .ZN(n_257_76_4396));
   INV_X1 i_257_76_4404 (.A(n_257_76_4396), .ZN(n_257_76_4397));
   NAND3_X1 i_257_76_4405 (.A1(n_257_76_4234), .A2(n_257_76_4235), .A3(
      n_257_76_4397), .ZN(n_257_76_4398));
   INV_X1 i_257_76_4406 (.A(n_257_76_4398), .ZN(n_257_76_4399));
   NAND4_X1 i_257_76_4407 (.A1(n_257_76_4395), .A2(n_257_76_4399), .A3(
      n_257_76_4224), .A4(n_257_76_4238), .ZN(n_257_76_4400));
   NAND3_X1 i_257_76_4408 (.A1(n_257_76_4199), .A2(n_257_76_4220), .A3(
      n_257_76_4223), .ZN(n_257_76_4401));
   NOR2_X1 i_257_76_4409 (.A1(n_257_76_4400), .A2(n_257_76_4401), .ZN(
      n_257_76_4402));
   NAND2_X1 i_257_76_4410 (.A1(n_257_76_4198), .A2(n_257_76_4402), .ZN(
      n_257_76_4403));
   INV_X1 i_257_76_4411 (.A(n_257_76_4403), .ZN(n_257_76_4404));
   NAND2_X1 i_257_76_4412 (.A1(n_257_76_4404), .A2(n_257_76_4210), .ZN(
      n_257_76_4405));
   INV_X1 i_257_76_4413 (.A(n_257_76_4405), .ZN(n_257_76_4406));
   NAND2_X1 i_257_76_4414 (.A1(n_257_76_18069), .A2(n_257_76_4406), .ZN(
      n_257_76_4407));
   INV_X1 i_257_76_4415 (.A(n_257_76_4287), .ZN(n_257_76_4408));
   INV_X1 i_257_76_4416 (.A(n_257_604), .ZN(n_257_76_4409));
   NOR2_X1 i_257_76_4417 (.A1(n_257_76_4201), .A2(n_257_76_4409), .ZN(
      n_257_76_4410));
   NAND2_X1 i_257_76_4418 (.A1(n_257_432), .A2(n_257_76_4410), .ZN(n_257_76_4411));
   INV_X1 i_257_76_4419 (.A(n_257_76_4411), .ZN(n_257_76_4412));
   NAND2_X1 i_257_76_4420 (.A1(n_257_76_4229), .A2(n_257_76_4412), .ZN(
      n_257_76_4413));
   NOR2_X1 i_257_76_4421 (.A1(n_257_76_4408), .A2(n_257_76_4413), .ZN(
      n_257_76_4414));
   NAND4_X1 i_257_76_4422 (.A1(n_257_76_4414), .A2(n_257_76_4335), .A3(
      n_257_76_4298), .A4(n_257_76_4228), .ZN(n_257_76_4415));
   NAND4_X1 i_257_76_4423 (.A1(n_257_76_4223), .A2(n_257_76_4224), .A3(
      n_257_76_4237), .A4(n_257_76_4238), .ZN(n_257_76_4416));
   NOR2_X1 i_257_76_4424 (.A1(n_257_76_4415), .A2(n_257_76_4416), .ZN(
      n_257_76_4417));
   NAND4_X1 i_257_76_4425 (.A1(n_257_76_4199), .A2(n_257_76_4272), .A3(
      n_257_76_4220), .A4(n_257_76_4222), .ZN(n_257_76_4418));
   INV_X1 i_257_76_4426 (.A(n_257_76_4418), .ZN(n_257_76_4419));
   NAND3_X1 i_257_76_4427 (.A1(n_257_76_4417), .A2(n_257_76_4227), .A3(
      n_257_76_4419), .ZN(n_257_76_4420));
   INV_X1 i_257_76_4428 (.A(n_257_76_4420), .ZN(n_257_76_4421));
   NAND2_X1 i_257_76_4429 (.A1(n_257_76_4421), .A2(n_257_76_4198), .ZN(
      n_257_76_4422));
   NOR2_X1 i_257_76_4430 (.A1(n_257_76_4422), .A2(n_257_76_4244), .ZN(
      n_257_76_4423));
   NAND2_X1 i_257_76_4431 (.A1(n_257_68), .A2(n_257_76_4423), .ZN(n_257_76_4424));
   NAND3_X1 i_257_76_4432 (.A1(n_257_76_4393), .A2(n_257_76_4407), .A3(
      n_257_76_4424), .ZN(n_257_76_4425));
   NAND2_X1 i_257_76_4433 (.A1(n_257_804), .A2(n_257_76_4228), .ZN(n_257_76_4426));
   INV_X1 i_257_76_4434 (.A(n_257_76_4426), .ZN(n_257_76_4427));
   NAND2_X1 i_257_76_4435 (.A1(n_257_437), .A2(n_257_76_4214), .ZN(n_257_76_4428));
   INV_X1 i_257_76_4436 (.A(n_257_76_4428), .ZN(n_257_76_4429));
   NAND3_X1 i_257_76_4437 (.A1(n_257_76_4234), .A2(n_257_76_4235), .A3(
      n_257_76_4429), .ZN(n_257_76_4430));
   INV_X1 i_257_76_4438 (.A(n_257_76_4430), .ZN(n_257_76_4431));
   NAND3_X1 i_257_76_4439 (.A1(n_257_76_4427), .A2(n_257_76_4431), .A3(
      n_257_76_4224), .ZN(n_257_76_4432));
   NOR2_X1 i_257_76_4440 (.A1(n_257_76_4432), .A2(n_257_76_4221), .ZN(
      n_257_76_4433));
   NAND2_X1 i_257_76_4441 (.A1(n_257_76_4198), .A2(n_257_76_4433), .ZN(
      n_257_76_4434));
   INV_X1 i_257_76_4442 (.A(n_257_76_4434), .ZN(n_257_76_4435));
   NAND2_X1 i_257_76_4443 (.A1(n_257_76_4435), .A2(n_257_76_4210), .ZN(
      n_257_76_4436));
   INV_X1 i_257_76_4444 (.A(n_257_76_4436), .ZN(n_257_76_4437));
   NAND2_X1 i_257_76_4445 (.A1(n_257_22), .A2(n_257_76_4437), .ZN(n_257_76_4438));
   NAND2_X1 i_257_76_4446 (.A1(n_257_444), .A2(n_257_76_4214), .ZN(n_257_76_4439));
   INV_X1 i_257_76_4447 (.A(n_257_76_4439), .ZN(n_257_76_4440));
   NAND2_X1 i_257_76_4448 (.A1(n_257_1002), .A2(n_257_76_4440), .ZN(
      n_257_76_4441));
   INV_X1 i_257_76_4449 (.A(n_257_76_4441), .ZN(n_257_76_4442));
   NAND2_X1 i_257_76_4450 (.A1(n_257_76_4210), .A2(n_257_76_4442), .ZN(
      n_257_76_4443));
   INV_X1 i_257_76_4451 (.A(n_257_76_4443), .ZN(n_257_76_4444));
   NAND2_X1 i_257_76_4452 (.A1(n_257_76_18075), .A2(n_257_76_4444), .ZN(
      n_257_76_4445));
   NAND2_X1 i_257_76_4453 (.A1(n_257_76_4438), .A2(n_257_76_4445), .ZN(
      n_257_76_4446));
   NOR2_X1 i_257_76_4454 (.A1(n_257_76_4425), .A2(n_257_76_4446), .ZN(
      n_257_76_4447));
   NAND3_X1 i_257_76_4455 (.A1(n_257_76_4311), .A2(n_257_76_4375), .A3(
      n_257_76_4447), .ZN(n_257_76_4448));
   INV_X1 i_257_76_4456 (.A(n_257_76_4448), .ZN(n_257_76_4449));
   NAND2_X1 i_257_76_4457 (.A1(n_257_42), .A2(n_257_76_4287), .ZN(n_257_76_4450));
   INV_X1 i_257_76_4458 (.A(n_257_76_4450), .ZN(n_257_76_4451));
   NAND2_X1 i_257_76_4459 (.A1(n_257_433), .A2(n_257_76_4214), .ZN(n_257_76_4452));
   INV_X1 i_257_76_4460 (.A(n_257_76_4452), .ZN(n_257_76_4453));
   NAND2_X1 i_257_76_4461 (.A1(n_257_76_4229), .A2(n_257_76_4453), .ZN(
      n_257_76_4454));
   INV_X1 i_257_76_4462 (.A(n_257_76_4454), .ZN(n_257_76_4455));
   NAND4_X1 i_257_76_4463 (.A1(n_257_76_4335), .A2(n_257_76_4451), .A3(
      n_257_76_4228), .A4(n_257_76_4455), .ZN(n_257_76_4456));
   NOR2_X1 i_257_76_4464 (.A1(n_257_76_4416), .A2(n_257_76_4456), .ZN(
      n_257_76_4457));
   NAND3_X1 i_257_76_4465 (.A1(n_257_76_4457), .A2(n_257_76_4227), .A3(
      n_257_76_4419), .ZN(n_257_76_4458));
   INV_X1 i_257_76_4466 (.A(n_257_76_4458), .ZN(n_257_76_4459));
   NAND2_X1 i_257_76_4467 (.A1(n_257_76_4459), .A2(n_257_76_4198), .ZN(
      n_257_76_4460));
   NOR2_X1 i_257_76_4468 (.A1(n_257_76_4460), .A2(n_257_76_4244), .ZN(
      n_257_76_4461));
   NAND2_X1 i_257_76_4469 (.A1(n_257_76_18081), .A2(n_257_76_4461), .ZN(
      n_257_76_4462));
   NAND3_X1 i_257_76_4470 (.A1(n_257_76_4238), .A2(n_257_76_4228), .A3(n_257_449), 
      .ZN(n_257_76_4463));
   NAND2_X1 i_257_76_4471 (.A1(n_257_76_17760), .A2(n_257_76_4214), .ZN(
      n_257_76_4464));
   OAI21_X1 i_257_76_4472 (.A(n_257_76_4464), .B1(n_257_708), .B2(n_257_76_4201), 
      .ZN(n_257_76_4465));
   NAND4_X1 i_257_76_4473 (.A1(n_257_76_4234), .A2(n_257_76_4235), .A3(
      n_257_76_4465), .A4(n_257_1080), .ZN(n_257_76_4466));
   NOR2_X1 i_257_76_4474 (.A1(n_257_76_4463), .A2(n_257_76_4466), .ZN(
      n_257_76_4467));
   NAND3_X1 i_257_76_4475 (.A1(n_257_76_4226), .A2(n_257_76_4227), .A3(
      n_257_76_4467), .ZN(n_257_76_4468));
   INV_X1 i_257_76_4476 (.A(n_257_76_4468), .ZN(n_257_76_4469));
   NAND2_X1 i_257_76_4477 (.A1(n_257_76_4469), .A2(n_257_76_4198), .ZN(
      n_257_76_4470));
   NOR2_X1 i_257_76_4478 (.A1(n_257_76_4470), .A2(n_257_76_4244), .ZN(
      n_257_76_4471));
   NAND2_X1 i_257_76_4479 (.A1(n_257_76_18083), .A2(n_257_76_4471), .ZN(
      n_257_76_4472));
   NAND2_X1 i_257_76_4480 (.A1(n_257_76_4277), .A2(n_257_159), .ZN(n_257_76_4473));
   INV_X1 i_257_76_4481 (.A(n_257_76_4473), .ZN(n_257_76_4474));
   NAND2_X1 i_257_76_4482 (.A1(n_257_429), .A2(n_257_76_4214), .ZN(n_257_76_4475));
   INV_X1 i_257_76_4483 (.A(n_257_76_4475), .ZN(n_257_76_4476));
   NAND2_X1 i_257_76_4484 (.A1(n_257_76_4288), .A2(n_257_76_4476), .ZN(
      n_257_76_4477));
   INV_X1 i_257_76_4485 (.A(n_257_76_4477), .ZN(n_257_76_4478));
   NAND3_X1 i_257_76_4486 (.A1(n_257_76_4287), .A2(n_257_76_4229), .A3(
      n_257_76_4478), .ZN(n_257_76_4479));
   INV_X1 i_257_76_4487 (.A(n_257_76_4479), .ZN(n_257_76_4480));
   NAND4_X1 i_257_76_4488 (.A1(n_257_76_4335), .A2(n_257_76_4480), .A3(
      n_257_76_4298), .A4(n_257_76_4228), .ZN(n_257_76_4481));
   NOR2_X1 i_257_76_4489 (.A1(n_257_76_4416), .A2(n_257_76_4481), .ZN(
      n_257_76_4482));
   NAND3_X1 i_257_76_4490 (.A1(n_257_76_4220), .A2(n_257_76_4282), .A3(
      n_257_76_4222), .ZN(n_257_76_4483));
   NOR2_X1 i_257_76_4491 (.A1(n_257_76_4483), .A2(n_257_76_4273), .ZN(
      n_257_76_4484));
   NAND4_X1 i_257_76_4492 (.A1(n_257_76_4474), .A2(n_257_76_4482), .A3(
      n_257_76_4227), .A4(n_257_76_4484), .ZN(n_257_76_4485));
   INV_X1 i_257_76_4493 (.A(n_257_76_4485), .ZN(n_257_76_4486));
   NAND3_X1 i_257_76_4494 (.A1(n_257_76_4486), .A2(n_257_76_4210), .A3(
      n_257_76_4198), .ZN(n_257_76_4487));
   INV_X1 i_257_76_4495 (.A(n_257_76_4487), .ZN(n_257_76_4488));
   NAND2_X1 i_257_76_4496 (.A1(n_257_76_18061), .A2(n_257_76_4488), .ZN(
      n_257_76_4489));
   NAND3_X1 i_257_76_4497 (.A1(n_257_76_4462), .A2(n_257_76_4472), .A3(
      n_257_76_4489), .ZN(n_257_76_4490));
   INV_X1 i_257_76_4498 (.A(n_257_76_4490), .ZN(n_257_76_4491));
   NAND2_X1 i_257_76_4499 (.A1(n_257_1072), .A2(n_257_76_4214), .ZN(
      n_257_76_4492));
   INV_X1 i_257_76_4500 (.A(n_257_76_4492), .ZN(n_257_76_4493));
   NAND2_X1 i_257_76_4501 (.A1(n_257_438), .A2(n_257_76_4493), .ZN(n_257_76_4494));
   INV_X1 i_257_76_4502 (.A(n_257_76_4494), .ZN(n_257_76_4495));
   NAND3_X1 i_257_76_4503 (.A1(n_257_76_4228), .A2(n_257_76_4495), .A3(
      n_257_76_4234), .ZN(n_257_76_4496));
   INV_X1 i_257_76_4504 (.A(n_257_76_4496), .ZN(n_257_76_4497));
   NAND2_X1 i_257_76_4505 (.A1(n_257_76_4497), .A2(n_257_76_4199), .ZN(
      n_257_76_4498));
   INV_X1 i_257_76_4506 (.A(n_257_76_4498), .ZN(n_257_76_4499));
   NAND2_X1 i_257_76_4507 (.A1(n_257_76_4198), .A2(n_257_76_4499), .ZN(
      n_257_76_4500));
   INV_X1 i_257_76_4508 (.A(n_257_76_4500), .ZN(n_257_76_4501));
   NAND2_X1 i_257_76_4509 (.A1(n_257_76_4501), .A2(n_257_76_4210), .ZN(
      n_257_76_4502));
   INV_X1 i_257_76_4510 (.A(n_257_76_4502), .ZN(n_257_76_4503));
   NAND2_X1 i_257_76_4511 (.A1(n_257_76_18067), .A2(n_257_76_4503), .ZN(
      n_257_76_4504));
   NAND2_X1 i_257_76_4512 (.A1(n_257_279), .A2(n_257_423), .ZN(n_257_76_4505));
   NAND3_X1 i_257_76_4513 (.A1(n_257_76_4222), .A2(n_257_76_4505), .A3(
      n_257_76_4223), .ZN(n_257_76_4506));
   INV_X1 i_257_76_4514 (.A(n_257_76_4506), .ZN(n_257_76_4507));
   NAND3_X1 i_257_76_4515 (.A1(n_257_76_4200), .A2(n_257_442), .A3(n_257_898), 
      .ZN(n_257_76_4508));
   INV_X1 i_257_76_4516 (.A(n_257_76_4508), .ZN(n_257_76_4509));
   NAND3_X1 i_257_76_4517 (.A1(n_257_420), .A2(n_257_76_4289), .A3(n_257_76_4509), 
      .ZN(n_257_76_4510));
   INV_X1 i_257_76_4518 (.A(n_257_76_4510), .ZN(n_257_76_4511));
   NAND2_X1 i_257_76_4519 (.A1(n_257_76_4294), .A2(n_257_76_4511), .ZN(
      n_257_76_4512));
   INV_X1 i_257_76_4520 (.A(n_257_76_4512), .ZN(n_257_76_4513));
   NAND2_X1 i_257_76_4521 (.A1(n_257_76_4229), .A2(n_257_76_4288), .ZN(
      n_257_76_4514));
   INV_X1 i_257_76_4522 (.A(n_257_76_4514), .ZN(n_257_76_4515));
   NAND4_X1 i_257_76_4523 (.A1(n_257_76_4513), .A2(n_257_76_4515), .A3(
      n_257_76_4285), .A4(n_257_76_4287), .ZN(n_257_76_4516));
   NAND2_X1 i_257_76_4524 (.A1(n_257_317), .A2(n_257_422), .ZN(n_257_76_4517));
   NAND4_X1 i_257_76_4525 (.A1(n_257_76_4228), .A2(n_257_76_4517), .A3(
      n_257_76_4234), .A4(n_257_76_4235), .ZN(n_257_76_4518));
   NOR2_X1 i_257_76_4526 (.A1(n_257_76_4516), .A2(n_257_76_4518), .ZN(
      n_257_76_4519));
   NAND3_X1 i_257_76_4527 (.A1(n_257_76_4238), .A2(n_257_76_4297), .A3(
      n_257_76_4298), .ZN(n_257_76_4520));
   NAND2_X1 i_257_76_4528 (.A1(n_257_76_4224), .A2(n_257_76_4237), .ZN(
      n_257_76_4521));
   NOR2_X1 i_257_76_4529 (.A1(n_257_76_4520), .A2(n_257_76_4521), .ZN(
      n_257_76_4522));
   NAND3_X1 i_257_76_4530 (.A1(n_257_76_4507), .A2(n_257_76_4519), .A3(
      n_257_76_4522), .ZN(n_257_76_4523));
   NAND2_X1 i_257_76_4531 (.A1(n_257_356), .A2(n_257_421), .ZN(n_257_76_4524));
   NAND2_X1 i_257_76_4532 (.A1(n_257_76_4524), .A2(n_257_76_4199), .ZN(
      n_257_76_4525));
   INV_X1 i_257_76_4533 (.A(n_257_76_4525), .ZN(n_257_76_4526));
   NAND3_X1 i_257_76_4534 (.A1(n_257_76_4272), .A2(n_257_76_4220), .A3(
      n_257_76_4282), .ZN(n_257_76_4527));
   INV_X1 i_257_76_4535 (.A(n_257_76_4527), .ZN(n_257_76_4528));
   NAND3_X1 i_257_76_4536 (.A1(n_257_76_4526), .A2(n_257_76_4528), .A3(
      n_257_76_4277), .ZN(n_257_76_4529));
   NOR2_X1 i_257_76_4537 (.A1(n_257_76_4523), .A2(n_257_76_4529), .ZN(
      n_257_76_4530));
   NAND3_X1 i_257_76_4538 (.A1(n_257_76_4227), .A2(n_257_76_4279), .A3(
      n_257_76_4276), .ZN(n_257_76_4531));
   INV_X1 i_257_76_4539 (.A(n_257_76_4531), .ZN(n_257_76_4532));
   NAND3_X1 i_257_76_4540 (.A1(n_257_76_4530), .A2(n_257_76_4532), .A3(
      n_257_76_4198), .ZN(n_257_76_4533));
   NOR2_X1 i_257_76_4541 (.A1(n_257_76_4533), .A2(n_257_76_4244), .ZN(
      n_257_76_4534));
   NAND2_X1 i_257_76_4542 (.A1(n_257_76_18073), .A2(n_257_76_4534), .ZN(
      n_257_76_4535));
   NAND2_X1 i_257_76_4543 (.A1(n_257_430), .A2(n_257_76_4214), .ZN(n_257_76_4536));
   INV_X1 i_257_76_4544 (.A(n_257_76_4536), .ZN(n_257_76_4537));
   NAND2_X1 i_257_76_4545 (.A1(n_257_76_4288), .A2(n_257_76_4537), .ZN(
      n_257_76_4538));
   INV_X1 i_257_76_4546 (.A(n_257_76_4538), .ZN(n_257_76_4539));
   NAND3_X1 i_257_76_4547 (.A1(n_257_76_4287), .A2(n_257_76_4229), .A3(
      n_257_76_4539), .ZN(n_257_76_4540));
   INV_X1 i_257_76_4548 (.A(n_257_76_4540), .ZN(n_257_76_4541));
   NAND4_X1 i_257_76_4549 (.A1(n_257_76_4335), .A2(n_257_76_4541), .A3(
      n_257_76_4298), .A4(n_257_76_4228), .ZN(n_257_76_4542));
   NAND4_X1 i_257_76_4550 (.A1(n_257_76_4224), .A2(n_257_76_4237), .A3(
      n_257_76_4238), .A4(n_257_120), .ZN(n_257_76_4543));
   NOR2_X1 i_257_76_4551 (.A1(n_257_76_4542), .A2(n_257_76_4543), .ZN(
      n_257_76_4544));
   NAND3_X1 i_257_76_4552 (.A1(n_257_76_4220), .A2(n_257_76_4222), .A3(
      n_257_76_4223), .ZN(n_257_76_4545));
   NOR2_X1 i_257_76_4553 (.A1(n_257_76_4545), .A2(n_257_76_4273), .ZN(
      n_257_76_4546));
   NAND4_X1 i_257_76_4554 (.A1(n_257_76_4227), .A2(n_257_76_4544), .A3(
      n_257_76_4546), .A4(n_257_76_4277), .ZN(n_257_76_4547));
   INV_X1 i_257_76_4555 (.A(n_257_76_4547), .ZN(n_257_76_4548));
   NAND3_X1 i_257_76_4556 (.A1(n_257_76_4548), .A2(n_257_76_4210), .A3(
      n_257_76_4198), .ZN(n_257_76_4549));
   INV_X1 i_257_76_4557 (.A(n_257_76_4549), .ZN(n_257_76_4550));
   NAND2_X1 i_257_76_4558 (.A1(n_257_76_18068), .A2(n_257_76_4550), .ZN(
      n_257_76_4551));
   NAND3_X1 i_257_76_4559 (.A1(n_257_76_4504), .A2(n_257_76_4535), .A3(
      n_257_76_4551), .ZN(n_257_76_4552));
   INV_X1 i_257_76_4560 (.A(n_257_76_4552), .ZN(n_257_76_4553));
   NAND2_X1 i_257_76_4561 (.A1(n_257_76_4228), .A2(n_257_447), .ZN(n_257_76_4554));
   INV_X1 i_257_76_4562 (.A(n_257_76_4554), .ZN(n_257_76_4555));
   INV_X1 i_257_76_4563 (.A(n_257_772), .ZN(n_257_76_4556));
   NOR2_X1 i_257_76_4564 (.A1(n_257_76_4201), .A2(n_257_76_4556), .ZN(
      n_257_76_4557));
   NAND3_X1 i_257_76_4565 (.A1(n_257_76_4234), .A2(n_257_76_4235), .A3(
      n_257_76_4557), .ZN(n_257_76_4558));
   INV_X1 i_257_76_4566 (.A(n_257_76_4558), .ZN(n_257_76_4559));
   NAND3_X1 i_257_76_4567 (.A1(n_257_76_4555), .A2(n_257_76_4559), .A3(
      n_257_76_4224), .ZN(n_257_76_4560));
   NOR2_X1 i_257_76_4568 (.A1(n_257_76_4401), .A2(n_257_76_4560), .ZN(
      n_257_76_4561));
   NAND2_X1 i_257_76_4569 (.A1(n_257_76_4198), .A2(n_257_76_4561), .ZN(
      n_257_76_4562));
   INV_X1 i_257_76_4570 (.A(n_257_76_4562), .ZN(n_257_76_4563));
   NAND2_X1 i_257_76_4571 (.A1(n_257_76_4563), .A2(n_257_76_4210), .ZN(
      n_257_76_4564));
   INV_X1 i_257_76_4572 (.A(n_257_76_4564), .ZN(n_257_76_4565));
   NAND2_X1 i_257_76_4573 (.A1(n_257_431), .A2(n_257_76_4214), .ZN(n_257_76_4566));
   INV_X1 i_257_76_4574 (.A(n_257_76_4566), .ZN(n_257_76_4567));
   NAND2_X1 i_257_76_4575 (.A1(n_257_76_4288), .A2(n_257_76_4567), .ZN(
      n_257_76_4568));
   INV_X1 i_257_76_4576 (.A(n_257_76_4568), .ZN(n_257_76_4569));
   NAND2_X1 i_257_76_4577 (.A1(n_257_76_4569), .A2(n_257_76_4229), .ZN(
      n_257_76_4570));
   INV_X1 i_257_76_4578 (.A(n_257_76_4570), .ZN(n_257_76_4571));
   NAND4_X1 i_257_76_4579 (.A1(n_257_76_4571), .A2(n_257_76_4234), .A3(
      n_257_76_4235), .A4(n_257_76_4287), .ZN(n_257_76_4572));
   NAND2_X1 i_257_76_4580 (.A1(n_257_76_4298), .A2(n_257_76_4228), .ZN(
      n_257_76_4573));
   NOR2_X1 i_257_76_4581 (.A1(n_257_76_4572), .A2(n_257_76_4573), .ZN(
      n_257_76_4574));
   INV_X1 i_257_76_4582 (.A(n_257_76_4274), .ZN(n_257_76_4575));
   NAND3_X1 i_257_76_4583 (.A1(n_257_76_4574), .A2(n_257_76_4302), .A3(
      n_257_76_4575), .ZN(n_257_76_4576));
   NAND4_X1 i_257_76_4584 (.A1(n_257_82), .A2(n_257_76_4199), .A3(n_257_76_4272), 
      .A4(n_257_76_4220), .ZN(n_257_76_4577));
   NOR2_X1 i_257_76_4585 (.A1(n_257_76_4576), .A2(n_257_76_4577), .ZN(
      n_257_76_4578));
   NAND3_X1 i_257_76_4586 (.A1(n_257_76_4578), .A2(n_257_76_4198), .A3(
      n_257_76_4227), .ZN(n_257_76_4579));
   NOR2_X1 i_257_76_4587 (.A1(n_257_76_4579), .A2(n_257_76_4244), .ZN(
      n_257_76_4580));
   AOI22_X1 i_257_76_4588 (.A1(n_257_76_18085), .A2(n_257_76_4565), .B1(
      n_257_76_18080), .B2(n_257_76_4580), .ZN(n_257_76_4581));
   NAND3_X1 i_257_76_4589 (.A1(n_257_76_4491), .A2(n_257_76_4553), .A3(
      n_257_76_4581), .ZN(n_257_76_4582));
   NAND3_X1 i_257_76_4590 (.A1(n_257_76_4223), .A2(n_257_76_4224), .A3(
      n_257_76_4238), .ZN(n_257_76_4583));
   NAND2_X1 i_257_76_4591 (.A1(n_257_448), .A2(n_257_76_4465), .ZN(n_257_76_4584));
   INV_X1 i_257_76_4592 (.A(n_257_76_4584), .ZN(n_257_76_4585));
   NAND3_X1 i_257_76_4593 (.A1(n_257_76_4335), .A2(n_257_76_4585), .A3(
      n_257_76_4228), .ZN(n_257_76_4586));
   NOR2_X1 i_257_76_4594 (.A1(n_257_76_4583), .A2(n_257_76_4586), .ZN(
      n_257_76_4587));
   NAND3_X1 i_257_76_4595 (.A1(n_257_76_4199), .A2(n_257_76_4220), .A3(
      n_257_76_4222), .ZN(n_257_76_4588));
   INV_X1 i_257_76_4596 (.A(n_257_76_4588), .ZN(n_257_76_4589));
   NAND3_X1 i_257_76_4597 (.A1(n_257_76_4587), .A2(n_257_676), .A3(n_257_76_4589), 
      .ZN(n_257_76_4590));
   INV_X1 i_257_76_4598 (.A(n_257_76_4590), .ZN(n_257_76_4591));
   NAND2_X1 i_257_76_4599 (.A1(n_257_76_4198), .A2(n_257_76_4591), .ZN(
      n_257_76_4592));
   NOR2_X1 i_257_76_4600 (.A1(n_257_76_4244), .A2(n_257_76_4592), .ZN(
      n_257_76_4593));
   NAND2_X1 i_257_76_4601 (.A1(n_257_76_18079), .A2(n_257_76_4593), .ZN(
      n_257_76_4594));
   NAND2_X1 i_257_76_4602 (.A1(n_257_425), .A2(n_257_76_4214), .ZN(n_257_76_4595));
   INV_X1 i_257_76_4603 (.A(n_257_76_4595), .ZN(n_257_76_4596));
   NAND3_X1 i_257_76_4604 (.A1(n_257_76_4288), .A2(n_257_76_4289), .A3(
      n_257_76_4596), .ZN(n_257_76_4597));
   INV_X1 i_257_76_4605 (.A(n_257_76_4597), .ZN(n_257_76_4598));
   NAND3_X1 i_257_76_4606 (.A1(n_257_76_4287), .A2(n_257_76_4229), .A3(
      n_257_76_4598), .ZN(n_257_76_4599));
   NOR2_X1 i_257_76_4607 (.A1(n_257_76_4286), .A2(n_257_76_4599), .ZN(
      n_257_76_4600));
   INV_X1 i_257_76_4608 (.A(n_257_76_4239), .ZN(n_257_76_4601));
   NAND3_X1 i_257_76_4609 (.A1(n_257_76_4297), .A2(n_257_76_4298), .A3(
      n_257_76_4228), .ZN(n_257_76_4602));
   INV_X1 i_257_76_4610 (.A(n_257_76_4602), .ZN(n_257_76_4603));
   NAND3_X1 i_257_76_4611 (.A1(n_257_76_4600), .A2(n_257_76_4601), .A3(
      n_257_76_4603), .ZN(n_257_76_4604));
   NOR2_X1 i_257_76_4612 (.A1(n_257_76_4604), .A2(n_257_76_4347), .ZN(
      n_257_76_4605));
   NAND3_X1 i_257_76_4613 (.A1(n_257_76_4350), .A2(n_257_76_4277), .A3(n_257_239), 
      .ZN(n_257_76_4606));
   INV_X1 i_257_76_4614 (.A(n_257_76_4606), .ZN(n_257_76_4607));
   NAND4_X1 i_257_76_4615 (.A1(n_257_76_4605), .A2(n_257_76_4607), .A3(
      n_257_76_4227), .A4(n_257_76_4276), .ZN(n_257_76_4608));
   INV_X1 i_257_76_4616 (.A(n_257_76_4608), .ZN(n_257_76_4609));
   NAND3_X1 i_257_76_4617 (.A1(n_257_76_4609), .A2(n_257_76_4210), .A3(
      n_257_76_4198), .ZN(n_257_76_4610));
   INV_X1 i_257_76_4618 (.A(n_257_76_4610), .ZN(n_257_76_4611));
   NAND2_X1 i_257_76_4619 (.A1(n_257_76_18064), .A2(n_257_76_4611), .ZN(
      n_257_76_4612));
   NAND3_X1 i_257_76_4620 (.A1(n_257_76_4282), .A2(n_257_76_4222), .A3(
      n_257_76_4505), .ZN(n_257_76_4613));
   NAND3_X1 i_257_76_4621 (.A1(n_257_356), .A2(n_257_76_4223), .A3(n_257_76_4224), 
      .ZN(n_257_76_4614));
   NOR2_X1 i_257_76_4622 (.A1(n_257_76_4613), .A2(n_257_76_4614), .ZN(
      n_257_76_4615));
   NAND2_X1 i_257_76_4623 (.A1(n_257_76_4228), .A2(n_257_76_4517), .ZN(
      n_257_76_4616));
   INV_X1 i_257_76_4624 (.A(n_257_76_4616), .ZN(n_257_76_4617));
   INV_X1 i_257_76_4625 (.A(n_257_76_4286), .ZN(n_257_76_4618));
   NAND2_X1 i_257_76_4626 (.A1(n_257_421), .A2(n_257_76_4214), .ZN(n_257_76_4619));
   INV_X1 i_257_76_4627 (.A(n_257_76_4619), .ZN(n_257_76_4620));
   NAND3_X1 i_257_76_4628 (.A1(n_257_76_4288), .A2(n_257_76_4289), .A3(
      n_257_76_4620), .ZN(n_257_76_4621));
   INV_X1 i_257_76_4629 (.A(n_257_76_4621), .ZN(n_257_76_4622));
   NAND4_X1 i_257_76_4630 (.A1(n_257_76_4287), .A2(n_257_76_4622), .A3(
      n_257_76_4294), .A4(n_257_76_4229), .ZN(n_257_76_4623));
   INV_X1 i_257_76_4631 (.A(n_257_76_4623), .ZN(n_257_76_4624));
   NAND3_X1 i_257_76_4632 (.A1(n_257_76_4617), .A2(n_257_76_4618), .A3(
      n_257_76_4624), .ZN(n_257_76_4625));
   NAND4_X1 i_257_76_4633 (.A1(n_257_76_4237), .A2(n_257_76_4238), .A3(
      n_257_76_4297), .A4(n_257_76_4298), .ZN(n_257_76_4626));
   NOR2_X1 i_257_76_4634 (.A1(n_257_76_4625), .A2(n_257_76_4626), .ZN(
      n_257_76_4627));
   NAND4_X1 i_257_76_4635 (.A1(n_257_76_4615), .A2(n_257_76_4627), .A3(
      n_257_76_4350), .A4(n_257_76_4277), .ZN(n_257_76_4628));
   INV_X1 i_257_76_4636 (.A(n_257_76_4628), .ZN(n_257_76_4629));
   NAND4_X1 i_257_76_4637 (.A1(n_257_76_4629), .A2(n_257_76_4210), .A3(
      n_257_76_4198), .A4(n_257_76_4532), .ZN(n_257_76_4630));
   INV_X1 i_257_76_4638 (.A(n_257_76_4630), .ZN(n_257_76_4631));
   NAND2_X1 i_257_76_4639 (.A1(n_257_76_18082), .A2(n_257_76_4631), .ZN(
      n_257_76_4632));
   NAND3_X1 i_257_76_4640 (.A1(n_257_76_4594), .A2(n_257_76_4612), .A3(
      n_257_76_4632), .ZN(n_257_76_4633));
   INV_X1 i_257_76_4641 (.A(n_257_76_4633), .ZN(n_257_76_4634));
   NAND4_X1 i_257_76_4642 (.A1(n_257_76_4298), .A2(n_257_76_4228), .A3(
      n_257_76_4234), .A4(n_257_76_4235), .ZN(n_257_76_4635));
   NOR2_X1 i_257_76_4643 (.A1(n_257_76_4274), .A2(n_257_76_4635), .ZN(
      n_257_76_4636));
   NAND2_X1 i_257_76_4644 (.A1(n_257_76_4229), .A2(n_257_199), .ZN(n_257_76_4637));
   INV_X1 i_257_76_4645 (.A(n_257_76_4637), .ZN(n_257_76_4638));
   INV_X1 i_257_76_4646 (.A(n_257_572), .ZN(n_257_76_4639));
   NAND3_X1 i_257_76_4647 (.A1(n_257_76_4200), .A2(n_257_76_4639), .A3(n_257_442), 
      .ZN(n_257_76_4640));
   OAI21_X1 i_257_76_4648 (.A(n_257_76_4640), .B1(n_257_428), .B2(n_257_76_4201), 
      .ZN(n_257_76_4641));
   NAND3_X1 i_257_76_4649 (.A1(n_257_427), .A2(n_257_76_4641), .A3(n_257_76_4288), 
      .ZN(n_257_76_4642));
   INV_X1 i_257_76_4650 (.A(n_257_76_4642), .ZN(n_257_76_4643));
   NAND3_X1 i_257_76_4651 (.A1(n_257_76_4638), .A2(n_257_76_4287), .A3(
      n_257_76_4643), .ZN(n_257_76_4644));
   INV_X1 i_257_76_4652 (.A(n_257_76_4644), .ZN(n_257_76_4645));
   NAND4_X1 i_257_76_4653 (.A1(n_257_76_4282), .A2(n_257_76_4645), .A3(
      n_257_76_4222), .A4(n_257_76_4223), .ZN(n_257_76_4646));
   INV_X1 i_257_76_4654 (.A(n_257_76_4646), .ZN(n_257_76_4647));
   NAND4_X1 i_257_76_4655 (.A1(n_257_76_4636), .A2(n_257_76_4647), .A3(
      n_257_76_4350), .A4(n_257_76_4277), .ZN(n_257_76_4648));
   NOR2_X1 i_257_76_4656 (.A1(n_257_76_4648), .A2(n_257_76_4352), .ZN(
      n_257_76_4649));
   NAND3_X1 i_257_76_4657 (.A1(n_257_76_4649), .A2(n_257_76_4210), .A3(
      n_257_76_4198), .ZN(n_257_76_4650));
   INV_X1 i_257_76_4658 (.A(n_257_76_4650), .ZN(n_257_76_4651));
   NAND2_X1 i_257_76_4659 (.A1(n_257_76_18065), .A2(n_257_76_4651), .ZN(
      n_257_76_4652));
   NAND3_X1 i_257_76_4660 (.A1(n_257_76_4287), .A2(n_257_76_4465), .A3(n_257_459), 
      .ZN(n_257_76_4653));
   INV_X1 i_257_76_4661 (.A(n_257_76_4653), .ZN(n_257_76_4654));
   NAND3_X1 i_257_76_4662 (.A1(n_257_76_4654), .A2(n_257_76_4335), .A3(
      n_257_76_4228), .ZN(n_257_76_4655));
   NAND3_X1 i_257_76_4663 (.A1(n_257_76_4237), .A2(n_257_76_4238), .A3(n_257_451), 
      .ZN(n_257_76_4656));
   NOR2_X1 i_257_76_4664 (.A1(n_257_76_4655), .A2(n_257_76_4656), .ZN(
      n_257_76_4657));
   NAND3_X1 i_257_76_4665 (.A1(n_257_76_4226), .A2(n_257_76_4227), .A3(
      n_257_76_4657), .ZN(n_257_76_4658));
   INV_X1 i_257_76_4666 (.A(n_257_76_4658), .ZN(n_257_76_4659));
   NAND2_X1 i_257_76_4667 (.A1(n_257_76_4659), .A2(n_257_76_4198), .ZN(
      n_257_76_4660));
   NOR2_X1 i_257_76_4668 (.A1(n_257_76_4660), .A2(n_257_76_4244), .ZN(
      n_257_76_4661));
   NAND2_X1 i_257_76_4669 (.A1(n_257_76_18063), .A2(n_257_76_4661), .ZN(
      n_257_76_4662));
   NAND4_X1 i_257_76_4670 (.A1(n_257_76_4228), .A2(n_257_76_4234), .A3(
      n_257_76_4235), .A4(n_257_76_4285), .ZN(n_257_76_4663));
   NAND2_X1 i_257_76_4671 (.A1(n_257_76_4297), .A2(n_257_76_4298), .ZN(
      n_257_76_4664));
   NOR2_X1 i_257_76_4672 (.A1(n_257_76_4663), .A2(n_257_76_4664), .ZN(
      n_257_76_4665));
   INV_X1 i_257_76_4673 (.A(n_257_76_4416), .ZN(n_257_76_4666));
   NAND2_X1 i_257_76_4674 (.A1(n_257_76_4282), .A2(n_257_76_4222), .ZN(
      n_257_76_4667));
   INV_X1 i_257_76_4675 (.A(n_257_76_4667), .ZN(n_257_76_4668));
   NAND3_X1 i_257_76_4676 (.A1(n_257_76_4665), .A2(n_257_76_4666), .A3(
      n_257_76_4668), .ZN(n_257_76_4669));
   INV_X1 i_257_76_4677 (.A(n_257_76_4273), .ZN(n_257_76_4670));
   NAND3_X1 i_257_76_4678 (.A1(n_257_76_4288), .A2(n_257_76_4641), .A3(n_257_424), 
      .ZN(n_257_76_4671));
   INV_X1 i_257_76_4679 (.A(n_257_76_4671), .ZN(n_257_76_4672));
   NAND4_X1 i_257_76_4680 (.A1(n_257_76_4287), .A2(n_257_76_4672), .A3(
      n_257_76_4229), .A4(n_257_508), .ZN(n_257_76_4673));
   INV_X1 i_257_76_4681 (.A(n_257_76_4673), .ZN(n_257_76_4674));
   NAND2_X1 i_257_76_4682 (.A1(n_257_76_4220), .A2(n_257_76_4674), .ZN(
      n_257_76_4675));
   INV_X1 i_257_76_4683 (.A(n_257_76_4675), .ZN(n_257_76_4676));
   NAND3_X1 i_257_76_4684 (.A1(n_257_76_4277), .A2(n_257_76_4670), .A3(
      n_257_76_4676), .ZN(n_257_76_4677));
   NOR2_X1 i_257_76_4685 (.A1(n_257_76_4669), .A2(n_257_76_4677), .ZN(
      n_257_76_4678));
   NAND3_X1 i_257_76_4686 (.A1(n_257_76_4678), .A2(n_257_76_4532), .A3(
      n_257_76_4198), .ZN(n_257_76_4679));
   NOR2_X1 i_257_76_4687 (.A1(n_257_76_4679), .A2(n_257_76_4244), .ZN(
      n_257_76_4680));
   NAND2_X1 i_257_76_4688 (.A1(n_257_76_18062), .A2(n_257_76_4680), .ZN(
      n_257_76_4681));
   NAND3_X1 i_257_76_4689 (.A1(n_257_76_4652), .A2(n_257_76_4662), .A3(
      n_257_76_4681), .ZN(n_257_76_4682));
   INV_X1 i_257_76_4690 (.A(n_257_76_4682), .ZN(n_257_76_4683));
   INV_X1 i_257_76_4691 (.A(n_257_76_4199), .ZN(n_257_76_4684));
   NAND3_X1 i_257_76_4692 (.A1(n_257_76_4288), .A2(n_257_76_4641), .A3(n_257_422), 
      .ZN(n_257_76_4685));
   NOR2_X1 i_257_76_4693 (.A1(n_257_76_4685), .A2(n_257_76_4377), .ZN(
      n_257_76_4686));
   NAND2_X1 i_257_76_4694 (.A1(n_257_76_4294), .A2(n_257_317), .ZN(n_257_76_4687));
   INV_X1 i_257_76_4695 (.A(n_257_76_4687), .ZN(n_257_76_4688));
   NAND3_X1 i_257_76_4696 (.A1(n_257_76_4686), .A2(n_257_76_4688), .A3(
      n_257_76_4287), .ZN(n_257_76_4689));
   NOR2_X1 i_257_76_4697 (.A1(n_257_76_4684), .A2(n_257_76_4689), .ZN(
      n_257_76_4690));
   NAND3_X1 i_257_76_4698 (.A1(n_257_76_4690), .A2(n_257_76_4528), .A3(
      n_257_76_4277), .ZN(n_257_76_4691));
   NAND2_X1 i_257_76_4699 (.A1(n_257_76_4222), .A2(n_257_76_4505), .ZN(
      n_257_76_4692));
   INV_X1 i_257_76_4700 (.A(n_257_76_4692), .ZN(n_257_76_4693));
   NAND3_X1 i_257_76_4701 (.A1(n_257_76_4665), .A2(n_257_76_4666), .A3(
      n_257_76_4693), .ZN(n_257_76_4694));
   NOR2_X1 i_257_76_4702 (.A1(n_257_76_4691), .A2(n_257_76_4694), .ZN(
      n_257_76_4695));
   NAND3_X1 i_257_76_4703 (.A1(n_257_76_4695), .A2(n_257_76_4532), .A3(
      n_257_76_4198), .ZN(n_257_76_4696));
   NOR2_X1 i_257_76_4704 (.A1(n_257_76_4696), .A2(n_257_76_4244), .ZN(
      n_257_76_4697));
   NAND2_X1 i_257_76_4705 (.A1(n_257_342), .A2(n_257_76_4697), .ZN(n_257_76_4698));
   NAND2_X1 i_257_76_4706 (.A1(n_257_76_4276), .A2(n_257_76_4277), .ZN(
      n_257_76_4699));
   NOR2_X1 i_257_76_4707 (.A1(n_257_76_4280), .A2(n_257_76_4699), .ZN(
      n_257_76_4700));
   INV_X1 i_257_76_4708 (.A(n_257_76_4664), .ZN(n_257_76_4701));
   NAND2_X1 i_257_76_4709 (.A1(n_257_76_4517), .A2(n_257_76_4234), .ZN(
      n_257_76_4702));
   INV_X1 i_257_76_4710 (.A(n_257_76_4228), .ZN(n_257_76_4703));
   NOR2_X1 i_257_76_4711 (.A1(n_257_76_4702), .A2(n_257_76_4703), .ZN(
      n_257_76_4704));
   NAND2_X1 i_257_76_4712 (.A1(n_257_76_4701), .A2(n_257_76_4704), .ZN(
      n_257_76_4705));
   NAND2_X1 i_257_76_4713 (.A1(n_257_76_4285), .A2(n_257_76_4287), .ZN(
      n_257_76_4706));
   INV_X1 i_257_76_4714 (.A(n_257_76_4235), .ZN(n_257_76_4707));
   NOR2_X1 i_257_76_4715 (.A1(n_257_76_4706), .A2(n_257_76_4707), .ZN(
      n_257_76_4708));
   INV_X1 i_257_76_4716 (.A(n_257_76_4288), .ZN(n_257_76_4709));
   NAND3_X1 i_257_76_4717 (.A1(n_257_76_4214), .A2(n_257_395), .A3(n_257_484), 
      .ZN(n_257_76_4710));
   INV_X1 i_257_76_4718 (.A(n_257_76_4710), .ZN(n_257_76_4711));
   NAND2_X1 i_257_76_4719 (.A1(n_257_76_4289), .A2(n_257_76_4711), .ZN(
      n_257_76_4712));
   NOR2_X1 i_257_76_4720 (.A1(n_257_76_4709), .A2(n_257_76_4712), .ZN(
      n_257_76_4713));
   NAND2_X1 i_257_76_4721 (.A1(n_257_420), .A2(n_257_898), .ZN(n_257_76_4714));
   NAND2_X1 i_257_76_4722 (.A1(n_257_76_4713), .A2(n_257_76_4714), .ZN(
      n_257_76_4715));
   NAND2_X1 i_257_76_4723 (.A1(n_257_76_4294), .A2(n_257_76_4229), .ZN(
      n_257_76_4716));
   NOR2_X1 i_257_76_4724 (.A1(n_257_76_4715), .A2(n_257_76_4716), .ZN(
      n_257_76_4717));
   NAND2_X1 i_257_76_4725 (.A1(n_257_76_4708), .A2(n_257_76_4717), .ZN(
      n_257_76_4718));
   NOR2_X1 i_257_76_4726 (.A1(n_257_76_4705), .A2(n_257_76_4718), .ZN(
      n_257_76_4719));
   NAND2_X1 i_257_76_4727 (.A1(n_257_76_4223), .A2(n_257_76_4224), .ZN(
      n_257_76_4720));
   NOR2_X1 i_257_76_4728 (.A1(n_257_76_4720), .A2(n_257_76_4239), .ZN(
      n_257_76_4721));
   NAND2_X1 i_257_76_4729 (.A1(n_257_76_4719), .A2(n_257_76_4721), .ZN(
      n_257_76_4722));
   INV_X1 i_257_76_4730 (.A(n_257_76_4524), .ZN(n_257_76_4723));
   NOR2_X1 i_257_76_4731 (.A1(n_257_76_4273), .A2(n_257_76_4723), .ZN(
      n_257_76_4724));
   NOR2_X1 i_257_76_4732 (.A1(n_257_76_4283), .A2(n_257_76_4692), .ZN(
      n_257_76_4725));
   NAND2_X1 i_257_76_4733 (.A1(n_257_76_4724), .A2(n_257_76_4725), .ZN(
      n_257_76_4726));
   NOR2_X1 i_257_76_4734 (.A1(n_257_76_4722), .A2(n_257_76_4726), .ZN(
      n_257_76_4727));
   NAND2_X1 i_257_76_4735 (.A1(n_257_76_4700), .A2(n_257_76_4727), .ZN(
      n_257_76_4728));
   NAND2_X1 i_257_76_4736 (.A1(n_257_76_4210), .A2(n_257_76_4198), .ZN(
      n_257_76_4729));
   NOR2_X1 i_257_76_4737 (.A1(n_257_76_4728), .A2(n_257_76_4729), .ZN(
      n_257_76_4730));
   NAND2_X1 i_257_76_4738 (.A1(n_257_76_18060), .A2(n_257_76_4730), .ZN(
      n_257_76_4731));
   INV_X1 i_257_76_4739 (.A(n_257_1034), .ZN(n_257_76_4732));
   OAI21_X1 i_257_76_4740 (.A(n_257_76_4628), .B1(n_257_76_4732), .B2(
      n_257_76_17968), .ZN(n_257_76_4733));
   NOR2_X1 i_257_76_4741 (.A1(n_257_76_4733), .A2(n_257_76_4609), .ZN(
      n_257_76_4734));
   AOI22_X1 i_257_76_4742 (.A1(n_257_159), .A2(n_257_76_17331), .B1(n_257_82), 
      .B2(n_257_76_17932), .ZN(n_257_76_4735));
   NAND2_X1 i_257_76_4743 (.A1(n_257_676), .A2(n_257_76_17958), .ZN(
      n_257_76_4736));
   NAND2_X1 i_257_76_4744 (.A1(n_257_76_4735), .A2(n_257_76_4736), .ZN(
      n_257_76_4737));
   INV_X1 i_257_76_4745 (.A(n_257_76_4737), .ZN(n_257_76_4738));
   NAND2_X1 i_257_76_4746 (.A1(n_257_970), .A2(n_257_442), .ZN(n_257_76_4739));
   INV_X1 i_257_76_4747 (.A(n_257_76_4739), .ZN(n_257_76_4740));
   NAND2_X1 i_257_76_4748 (.A1(n_257_441), .A2(n_257_76_4740), .ZN(n_257_76_4741));
   NAND2_X1 i_257_76_4749 (.A1(n_257_76_4689), .A2(n_257_76_4741), .ZN(
      n_257_76_4742));
   NAND2_X1 i_257_76_4750 (.A1(n_257_459), .A2(n_257_442), .ZN(n_257_76_4743));
   INV_X1 i_257_76_4751 (.A(n_257_76_4743), .ZN(n_257_76_4744));
   NAND2_X1 i_257_76_4752 (.A1(n_257_451), .A2(n_257_76_4744), .ZN(n_257_76_4745));
   NAND2_X1 i_257_76_4753 (.A1(n_257_868), .A2(n_257_76_17903), .ZN(
      n_257_76_4746));
   NAND2_X1 i_257_76_4754 (.A1(n_257_76_4745), .A2(n_257_76_4746), .ZN(
      n_257_76_4747));
   NOR2_X1 i_257_76_4755 (.A1(n_257_76_4742), .A2(n_257_76_4747), .ZN(
      n_257_76_4748));
   NAND2_X1 i_257_76_4756 (.A1(n_257_120), .A2(n_257_76_17925), .ZN(
      n_257_76_4749));
   NAND2_X1 i_257_76_4757 (.A1(n_257_740), .A2(n_257_76_17935), .ZN(
      n_257_76_4750));
   NAND2_X1 i_257_76_4758 (.A1(n_257_76_4749), .A2(n_257_76_4750), .ZN(
      n_257_76_4751));
   NAND2_X1 i_257_76_4759 (.A1(n_257_804), .A2(n_257_76_17952), .ZN(
      n_257_76_4752));
   NAND2_X1 i_257_76_4760 (.A1(n_257_76_4673), .A2(n_257_76_4752), .ZN(
      n_257_76_4753));
   NOR2_X1 i_257_76_4761 (.A1(n_257_76_4751), .A2(n_257_76_4753), .ZN(
      n_257_76_4754));
   NAND2_X1 i_257_76_4762 (.A1(n_257_76_4748), .A2(n_257_76_4754), .ZN(
      n_257_76_4755));
   NAND2_X1 i_257_76_4763 (.A1(n_257_836), .A2(n_257_442), .ZN(n_257_76_4756));
   INV_X1 i_257_76_4764 (.A(n_257_76_4756), .ZN(n_257_76_4757));
   NAND2_X1 i_257_76_4765 (.A1(n_257_446), .A2(n_257_76_4757), .ZN(n_257_76_4758));
   NAND2_X1 i_257_76_4766 (.A1(n_257_76_4644), .A2(n_257_76_4758), .ZN(
      n_257_76_4759));
   NAND2_X1 i_257_76_4767 (.A1(n_257_449), .A2(n_257_76_12076), .ZN(
      n_257_76_4760));
   NAND2_X1 i_257_76_4768 (.A1(n_257_772), .A2(n_257_442), .ZN(n_257_76_4761));
   INV_X1 i_257_76_4769 (.A(n_257_76_4761), .ZN(n_257_76_4762));
   NAND2_X1 i_257_76_4770 (.A1(n_257_447), .A2(n_257_76_4762), .ZN(n_257_76_4763));
   NAND2_X1 i_257_76_4771 (.A1(n_257_76_4760), .A2(n_257_76_4763), .ZN(
      n_257_76_4764));
   NOR2_X1 i_257_76_4772 (.A1(n_257_76_4759), .A2(n_257_76_4764), .ZN(
      n_257_76_4765));
   NAND2_X1 i_257_76_4773 (.A1(n_257_938), .A2(n_257_442), .ZN(n_257_76_4766));
   INV_X1 i_257_76_4774 (.A(n_257_76_4766), .ZN(n_257_76_4767));
   AOI22_X1 i_257_76_4775 (.A1(n_257_42), .A2(n_257_76_17918), .B1(n_257_440), 
      .B2(n_257_76_4767), .ZN(n_257_76_4768));
   NAND3_X1 i_257_76_4776 (.A1(n_257_906), .A2(n_257_439), .A3(n_257_442), 
      .ZN(n_257_76_4769));
   NAND2_X1 i_257_76_4777 (.A1(n_257_76_4768), .A2(n_257_76_4769), .ZN(
      n_257_76_4770));
   NAND2_X1 i_257_76_4778 (.A1(n_257_76_15655), .A2(n_257_708), .ZN(
      n_257_76_4771));
   NAND2_X1 i_257_76_4779 (.A1(n_257_76_4771), .A2(n_257_76_4510), .ZN(
      n_257_76_4772));
   NAND2_X1 i_257_76_4780 (.A1(n_257_604), .A2(n_257_442), .ZN(n_257_76_4773));
   OAI21_X1 i_257_76_4781 (.A(n_257_76_4338), .B1(n_257_76_15481), .B2(
      n_257_76_4773), .ZN(n_257_76_4774));
   INV_X1 i_257_76_4782 (.A(n_257_76_4774), .ZN(n_257_76_4775));
   INV_X1 i_257_76_4783 (.A(Small_Packet_Data_Size[7]), .ZN(n_257_76_4776));
   NAND2_X1 i_257_76_4784 (.A1(n_257_76_4710), .A2(n_257_76_18050), .ZN(
      n_257_76_4777));
   INV_X1 i_257_76_4785 (.A(n_257_76_4777), .ZN(n_257_76_4778));
   NAND2_X1 i_257_76_4786 (.A1(n_257_76_4775), .A2(n_257_76_4778), .ZN(
      n_257_76_4779));
   NOR2_X1 i_257_76_4787 (.A1(n_257_76_4772), .A2(n_257_76_4779), .ZN(
      n_257_76_4780));
   AOI22_X1 i_257_76_4788 (.A1(n_257_438), .A2(n_257_76_7724), .B1(n_257_636), 
      .B2(n_257_76_17928), .ZN(n_257_76_4781));
   NAND2_X1 i_257_76_4789 (.A1(n_257_76_4780), .A2(n_257_76_4781), .ZN(
      n_257_76_4782));
   NOR2_X1 i_257_76_4790 (.A1(n_257_76_4770), .A2(n_257_76_4782), .ZN(
      n_257_76_4783));
   NAND2_X1 i_257_76_4791 (.A1(n_257_76_4765), .A2(n_257_76_4783), .ZN(
      n_257_76_4784));
   NOR2_X1 i_257_76_4792 (.A1(n_257_76_4755), .A2(n_257_76_4784), .ZN(
      n_257_76_4785));
   NAND2_X1 i_257_76_4793 (.A1(n_257_76_4738), .A2(n_257_76_4785), .ZN(
      n_257_76_4786));
   NAND2_X1 i_257_76_4794 (.A1(n_257_76_4387), .A2(n_257_76_4303), .ZN(
      n_257_76_4787));
   INV_X1 i_257_76_4795 (.A(n_257_76_4787), .ZN(n_257_76_4788));
   NAND2_X1 i_257_76_4796 (.A1(n_257_1002), .A2(n_257_76_17964), .ZN(
      n_257_76_4789));
   NAND2_X1 i_257_76_4797 (.A1(n_257_76_4788), .A2(n_257_76_4789), .ZN(
      n_257_76_4790));
   NOR2_X1 i_257_76_4798 (.A1(n_257_76_4786), .A2(n_257_76_4790), .ZN(
      n_257_76_4791));
   NAND2_X1 i_257_76_4799 (.A1(n_257_76_4734), .A2(n_257_76_4791), .ZN(
      n_257_76_4792));
   NAND3_X1 i_257_76_4800 (.A1(n_257_76_4698), .A2(n_257_76_4731), .A3(
      n_257_76_4792), .ZN(n_257_76_4793));
   INV_X1 i_257_76_4801 (.A(n_257_76_4793), .ZN(n_257_76_4794));
   NAND3_X1 i_257_76_4802 (.A1(n_257_76_4634), .A2(n_257_76_4683), .A3(
      n_257_76_4794), .ZN(n_257_76_4795));
   NOR2_X1 i_257_76_4803 (.A1(n_257_76_4582), .A2(n_257_76_4795), .ZN(
      n_257_76_4796));
   NAND2_X1 i_257_76_4804 (.A1(n_257_76_4449), .A2(n_257_76_4796), .ZN(n_7));
   NAND2_X1 i_257_76_4805 (.A1(n_257_1003), .A2(n_257_444), .ZN(n_257_76_4797));
   NAND2_X1 i_257_76_4806 (.A1(n_257_441), .A2(n_257_971), .ZN(n_257_76_4798));
   NAND2_X1 i_257_76_4807 (.A1(n_257_939), .A2(n_257_442), .ZN(n_257_76_4799));
   NOR2_X1 i_257_76_4808 (.A1(n_257_1067), .A2(n_257_76_4799), .ZN(n_257_76_4800));
   NAND2_X1 i_257_76_4809 (.A1(n_257_440), .A2(n_257_76_4800), .ZN(n_257_76_4801));
   INV_X1 i_257_76_4810 (.A(n_257_76_4801), .ZN(n_257_76_4802));
   NAND2_X1 i_257_76_4811 (.A1(n_257_76_4798), .A2(n_257_76_4802), .ZN(
      n_257_76_4803));
   INV_X1 i_257_76_4812 (.A(n_257_76_4803), .ZN(n_257_76_4804));
   NAND2_X1 i_257_76_4813 (.A1(n_257_76_4797), .A2(n_257_76_4804), .ZN(
      n_257_76_4805));
   INV_X1 i_257_76_4814 (.A(n_257_76_4805), .ZN(n_257_76_4806));
   NAND2_X1 i_257_76_4815 (.A1(n_257_1035), .A2(n_257_443), .ZN(n_257_76_4807));
   NAND2_X1 i_257_76_4816 (.A1(n_257_76_4806), .A2(n_257_76_4807), .ZN(
      n_257_76_4808));
   INV_X1 i_257_76_4817 (.A(n_257_76_4808), .ZN(n_257_76_4809));
   NAND2_X1 i_257_76_4818 (.A1(n_257_17), .A2(n_257_76_4809), .ZN(n_257_76_4810));
   NOR2_X1 i_257_76_4819 (.A1(n_257_1067), .A2(n_257_76_17412), .ZN(
      n_257_76_4811));
   NAND2_X1 i_257_76_4820 (.A1(n_257_443), .A2(n_257_76_4811), .ZN(n_257_76_4812));
   INV_X1 i_257_76_4821 (.A(n_257_76_4812), .ZN(n_257_76_4813));
   NAND2_X1 i_257_76_4822 (.A1(n_257_1035), .A2(n_257_76_4813), .ZN(
      n_257_76_4814));
   INV_X1 i_257_76_4823 (.A(n_257_76_4814), .ZN(n_257_76_4815));
   NAND2_X1 i_257_76_4824 (.A1(n_257_76_18072), .A2(n_257_76_4815), .ZN(
      n_257_76_4816));
   NAND2_X1 i_257_76_4825 (.A1(n_257_907), .A2(n_257_439), .ZN(n_257_76_4817));
   NAND2_X1 i_257_76_4826 (.A1(n_257_446), .A2(n_257_837), .ZN(n_257_76_4818));
   NAND2_X1 i_257_76_4827 (.A1(n_257_76_4817), .A2(n_257_76_4818), .ZN(
      n_257_76_4819));
   INV_X1 i_257_76_4828 (.A(n_257_76_4819), .ZN(n_257_76_4820));
   NAND3_X1 i_257_76_4829 (.A1(n_257_76_4811), .A2(n_257_637), .A3(n_257_450), 
      .ZN(n_257_76_4821));
   INV_X1 i_257_76_4830 (.A(n_257_76_4821), .ZN(n_257_76_4822));
   NAND2_X1 i_257_76_4831 (.A1(n_257_709), .A2(n_257_435), .ZN(n_257_76_4823));
   NAND2_X1 i_257_76_4832 (.A1(n_257_440), .A2(n_257_939), .ZN(n_257_76_4824));
   NAND2_X1 i_257_76_4833 (.A1(n_257_438), .A2(n_257_1073), .ZN(n_257_76_4825));
   NAND4_X1 i_257_76_4834 (.A1(n_257_76_4822), .A2(n_257_76_4823), .A3(
      n_257_76_4824), .A4(n_257_76_4825), .ZN(n_257_76_4826));
   INV_X1 i_257_76_4835 (.A(n_257_76_4826), .ZN(n_257_76_4827));
   NAND2_X1 i_257_76_4836 (.A1(n_257_449), .A2(n_257_1081), .ZN(n_257_76_4828));
   NAND2_X1 i_257_76_4837 (.A1(n_257_447), .A2(n_257_773), .ZN(n_257_76_4829));
   NAND2_X1 i_257_76_4838 (.A1(n_257_76_4828), .A2(n_257_76_4829), .ZN(
      n_257_76_4830));
   INV_X1 i_257_76_4839 (.A(n_257_76_4830), .ZN(n_257_76_4831));
   NAND4_X1 i_257_76_4840 (.A1(n_257_76_4820), .A2(n_257_76_4827), .A3(
      n_257_76_4831), .A4(n_257_76_4798), .ZN(n_257_76_4832));
   NAND2_X1 i_257_76_4841 (.A1(n_257_741), .A2(n_257_436), .ZN(n_257_76_4833));
   NAND2_X1 i_257_76_4842 (.A1(n_257_805), .A2(n_257_437), .ZN(n_257_76_4834));
   NAND2_X1 i_257_76_4843 (.A1(n_257_869), .A2(n_257_445), .ZN(n_257_76_4835));
   NAND3_X1 i_257_76_4844 (.A1(n_257_76_4833), .A2(n_257_76_4834), .A3(
      n_257_76_4835), .ZN(n_257_76_4836));
   NOR2_X1 i_257_76_4845 (.A1(n_257_76_4832), .A2(n_257_76_4836), .ZN(
      n_257_76_4837));
   NAND2_X1 i_257_76_4846 (.A1(n_257_677), .A2(n_257_448), .ZN(n_257_76_4838));
   NAND3_X1 i_257_76_4847 (.A1(n_257_76_4837), .A2(n_257_76_4838), .A3(
      n_257_76_4797), .ZN(n_257_76_4839));
   INV_X1 i_257_76_4848 (.A(n_257_76_4807), .ZN(n_257_76_4840));
   NOR2_X1 i_257_76_4849 (.A1(n_257_76_4839), .A2(n_257_76_4840), .ZN(
      n_257_76_4841));
   NAND2_X1 i_257_76_4850 (.A1(n_257_28), .A2(n_257_76_4841), .ZN(n_257_76_4842));
   NAND3_X1 i_257_76_4851 (.A1(n_257_76_4810), .A2(n_257_76_4816), .A3(
      n_257_76_4842), .ZN(n_257_76_4843));
   INV_X1 i_257_76_4852 (.A(n_257_76_4811), .ZN(n_257_76_4844));
   INV_X1 i_257_76_4853 (.A(n_257_837), .ZN(n_257_76_4845));
   NOR2_X1 i_257_76_4854 (.A1(n_257_76_4844), .A2(n_257_76_4845), .ZN(
      n_257_76_4846));
   NAND4_X1 i_257_76_4855 (.A1(n_257_446), .A2(n_257_76_4846), .A3(n_257_76_4824), 
      .A4(n_257_76_4825), .ZN(n_257_76_4847));
   INV_X1 i_257_76_4856 (.A(n_257_76_4847), .ZN(n_257_76_4848));
   NAND4_X1 i_257_76_4857 (.A1(n_257_76_4835), .A2(n_257_76_4848), .A3(
      n_257_76_4798), .A4(n_257_76_4817), .ZN(n_257_76_4849));
   INV_X1 i_257_76_4858 (.A(n_257_76_4849), .ZN(n_257_76_4850));
   NAND2_X1 i_257_76_4859 (.A1(n_257_76_4797), .A2(n_257_76_4850), .ZN(
      n_257_76_4851));
   INV_X1 i_257_76_4860 (.A(n_257_76_4851), .ZN(n_257_76_4852));
   NAND2_X1 i_257_76_4861 (.A1(n_257_76_4852), .A2(n_257_76_4807), .ZN(
      n_257_76_4853));
   INV_X1 i_257_76_4862 (.A(n_257_76_4853), .ZN(n_257_76_4854));
   NAND2_X1 i_257_76_4863 (.A1(n_257_76_18070), .A2(n_257_76_4854), .ZN(
      n_257_76_4855));
   NAND2_X1 i_257_76_4864 (.A1(n_257_439), .A2(n_257_76_4811), .ZN(n_257_76_4856));
   INV_X1 i_257_76_4865 (.A(n_257_76_4856), .ZN(n_257_76_4857));
   NAND3_X1 i_257_76_4866 (.A1(n_257_907), .A2(n_257_76_4857), .A3(n_257_76_4824), 
      .ZN(n_257_76_4858));
   INV_X1 i_257_76_4867 (.A(n_257_76_4858), .ZN(n_257_76_4859));
   NAND2_X1 i_257_76_4868 (.A1(n_257_76_4859), .A2(n_257_76_4798), .ZN(
      n_257_76_4860));
   INV_X1 i_257_76_4869 (.A(n_257_76_4860), .ZN(n_257_76_4861));
   NAND2_X1 i_257_76_4870 (.A1(n_257_76_4797), .A2(n_257_76_4861), .ZN(
      n_257_76_4862));
   INV_X1 i_257_76_4871 (.A(n_257_76_4862), .ZN(n_257_76_4863));
   NAND2_X1 i_257_76_4872 (.A1(n_257_76_4863), .A2(n_257_76_4807), .ZN(
      n_257_76_4864));
   INV_X1 i_257_76_4873 (.A(n_257_76_4864), .ZN(n_257_76_4865));
   NAND2_X1 i_257_76_4874 (.A1(n_257_76_18084), .A2(n_257_76_4865), .ZN(
      n_257_76_4866));
   NAND2_X1 i_257_76_4875 (.A1(n_257_160), .A2(n_257_429), .ZN(n_257_76_4867));
   NAND2_X1 i_257_76_4876 (.A1(n_257_541), .A2(n_257_426), .ZN(n_257_76_4868));
   NAND2_X1 i_257_76_4877 (.A1(n_257_43), .A2(n_257_433), .ZN(n_257_76_4869));
   NAND3_X1 i_257_76_4878 (.A1(n_257_76_4868), .A2(n_257_280), .A3(n_257_76_4869), 
      .ZN(n_257_76_4870));
   INV_X1 i_257_76_4879 (.A(n_257_76_4870), .ZN(n_257_76_4871));
   NAND2_X1 i_257_76_4880 (.A1(n_257_432), .A2(n_257_605), .ZN(n_257_76_4872));
   INV_X1 i_257_76_4881 (.A(n_257_1067), .ZN(n_257_76_4873));
   INV_X1 i_257_76_4882 (.A(n_257_573), .ZN(n_257_76_4874));
   NAND2_X1 i_257_76_4883 (.A1(n_257_76_4874), .A2(n_257_442), .ZN(n_257_76_4875));
   OAI21_X1 i_257_76_4884 (.A(n_257_76_4875), .B1(n_257_428), .B2(n_257_76_17412), 
      .ZN(n_257_76_4876));
   NAND4_X1 i_257_76_4885 (.A1(n_257_76_4872), .A2(n_257_76_4873), .A3(
      n_257_76_4876), .A4(n_257_423), .ZN(n_257_76_4877));
   INV_X1 i_257_76_4886 (.A(n_257_76_4877), .ZN(n_257_76_4878));
   NAND2_X1 i_257_76_4887 (.A1(n_257_637), .A2(n_257_450), .ZN(n_257_76_4879));
   NAND2_X1 i_257_76_4888 (.A1(n_257_200), .A2(n_257_427), .ZN(n_257_76_4880));
   NAND2_X1 i_257_76_4889 (.A1(n_257_509), .A2(n_257_424), .ZN(n_257_76_4881));
   NAND4_X1 i_257_76_4890 (.A1(n_257_76_4878), .A2(n_257_76_4879), .A3(
      n_257_76_4880), .A4(n_257_76_4881), .ZN(n_257_76_4882));
   INV_X1 i_257_76_4891 (.A(n_257_76_4882), .ZN(n_257_76_4883));
   NAND3_X1 i_257_76_4892 (.A1(n_257_76_4823), .A2(n_257_76_4824), .A3(
      n_257_76_4825), .ZN(n_257_76_4884));
   INV_X1 i_257_76_4893 (.A(n_257_76_4884), .ZN(n_257_76_4885));
   NAND4_X1 i_257_76_4894 (.A1(n_257_76_4871), .A2(n_257_76_4883), .A3(
      n_257_76_4817), .A4(n_257_76_4885), .ZN(n_257_76_4886));
   INV_X1 i_257_76_4895 (.A(n_257_76_4886), .ZN(n_257_76_4887));
   NAND2_X1 i_257_76_4896 (.A1(n_257_83), .A2(n_257_431), .ZN(n_257_76_4888));
   NAND3_X1 i_257_76_4897 (.A1(n_257_76_4867), .A2(n_257_76_4887), .A3(
      n_257_76_4888), .ZN(n_257_76_4889));
   INV_X1 i_257_76_4898 (.A(n_257_76_4889), .ZN(n_257_76_4890));
   NAND3_X1 i_257_76_4899 (.A1(n_257_76_4818), .A2(n_257_76_4828), .A3(
      n_257_76_4829), .ZN(n_257_76_4891));
   INV_X1 i_257_76_4900 (.A(n_257_76_4891), .ZN(n_257_76_4892));
   NAND2_X1 i_257_76_4901 (.A1(n_257_121), .A2(n_257_430), .ZN(n_257_76_4893));
   NAND2_X1 i_257_76_4902 (.A1(n_257_451), .A2(n_257_460), .ZN(n_257_76_4894));
   NAND4_X1 i_257_76_4903 (.A1(n_257_76_4892), .A2(n_257_76_4893), .A3(
      n_257_76_4798), .A4(n_257_76_4894), .ZN(n_257_76_4895));
   NOR2_X1 i_257_76_4904 (.A1(n_257_76_4895), .A2(n_257_76_4836), .ZN(
      n_257_76_4896));
   NAND4_X1 i_257_76_4905 (.A1(n_257_76_4890), .A2(n_257_76_4896), .A3(
      n_257_76_4838), .A4(n_257_76_4797), .ZN(n_257_76_4897));
   NAND2_X1 i_257_76_4906 (.A1(n_257_240), .A2(n_257_425), .ZN(n_257_76_4898));
   NAND2_X1 i_257_76_4907 (.A1(n_257_76_4807), .A2(n_257_76_4898), .ZN(
      n_257_76_4899));
   NOR2_X1 i_257_76_4908 (.A1(n_257_76_4897), .A2(n_257_76_4899), .ZN(
      n_257_76_4900));
   NAND2_X1 i_257_76_4909 (.A1(n_257_76_18066), .A2(n_257_76_4900), .ZN(
      n_257_76_4901));
   NAND3_X1 i_257_76_4910 (.A1(n_257_76_4855), .A2(n_257_76_4866), .A3(
      n_257_76_4901), .ZN(n_257_76_4902));
   NOR2_X1 i_257_76_4911 (.A1(n_257_76_4843), .A2(n_257_76_4902), .ZN(
      n_257_76_4903));
   INV_X1 i_257_76_4912 (.A(n_257_971), .ZN(n_257_76_4904));
   NOR2_X1 i_257_76_4913 (.A1(n_257_76_4844), .A2(n_257_76_4904), .ZN(
      n_257_76_4905));
   NAND2_X1 i_257_76_4914 (.A1(n_257_441), .A2(n_257_76_4905), .ZN(n_257_76_4906));
   INV_X1 i_257_76_4915 (.A(n_257_76_4906), .ZN(n_257_76_4907));
   NAND2_X1 i_257_76_4916 (.A1(n_257_76_4797), .A2(n_257_76_4907), .ZN(
      n_257_76_4908));
   INV_X1 i_257_76_4917 (.A(n_257_76_4908), .ZN(n_257_76_4909));
   NAND2_X1 i_257_76_4918 (.A1(n_257_76_4909), .A2(n_257_76_4807), .ZN(
      n_257_76_4910));
   INV_X1 i_257_76_4919 (.A(n_257_76_4910), .ZN(n_257_76_4911));
   NAND2_X1 i_257_76_4920 (.A1(n_257_76_18071), .A2(n_257_76_4911), .ZN(
      n_257_76_4912));
   NAND2_X1 i_257_76_4921 (.A1(n_257_76_4818), .A2(n_257_76_4829), .ZN(
      n_257_76_4913));
   INV_X1 i_257_76_4922 (.A(n_257_76_4913), .ZN(n_257_76_4914));
   NOR2_X1 i_257_76_4923 (.A1(n_257_76_4844), .A2(n_257_76_17760), .ZN(
      n_257_76_4915));
   NAND4_X1 i_257_76_4924 (.A1(n_257_76_4915), .A2(n_257_76_4824), .A3(
      n_257_76_4825), .A4(n_257_709), .ZN(n_257_76_4916));
   INV_X1 i_257_76_4925 (.A(n_257_76_4916), .ZN(n_257_76_4917));
   NAND4_X1 i_257_76_4926 (.A1(n_257_76_4914), .A2(n_257_76_4917), .A3(
      n_257_76_4798), .A4(n_257_76_4817), .ZN(n_257_76_4918));
   NOR2_X1 i_257_76_4927 (.A1(n_257_76_4836), .A2(n_257_76_4918), .ZN(
      n_257_76_4919));
   NAND2_X1 i_257_76_4928 (.A1(n_257_76_4797), .A2(n_257_76_4919), .ZN(
      n_257_76_4920));
   NOR2_X1 i_257_76_4929 (.A1(n_257_76_4840), .A2(n_257_76_4920), .ZN(
      n_257_76_4921));
   NAND2_X1 i_257_76_4930 (.A1(n_257_76_18078), .A2(n_257_76_4921), .ZN(
      n_257_76_4922));
   NAND4_X1 i_257_76_4931 (.A1(n_257_76_4894), .A2(n_257_76_4817), .A3(
      n_257_76_4818), .A4(n_257_76_4828), .ZN(n_257_76_4923));
   NAND2_X1 i_257_76_4932 (.A1(n_257_442), .A2(n_257_573), .ZN(n_257_76_4924));
   INV_X1 i_257_76_4933 (.A(n_257_76_4924), .ZN(n_257_76_4925));
   NAND2_X1 i_257_76_4934 (.A1(n_257_428), .A2(n_257_76_4925), .ZN(n_257_76_4926));
   INV_X1 i_257_76_4935 (.A(n_257_76_4926), .ZN(n_257_76_4927));
   NAND3_X1 i_257_76_4936 (.A1(n_257_76_4872), .A2(n_257_76_4873), .A3(
      n_257_76_4927), .ZN(n_257_76_4928));
   INV_X1 i_257_76_4937 (.A(n_257_76_4928), .ZN(n_257_76_4929));
   NAND3_X1 i_257_76_4938 (.A1(n_257_76_4825), .A2(n_257_76_4879), .A3(
      n_257_76_4929), .ZN(n_257_76_4930));
   INV_X1 i_257_76_4939 (.A(n_257_76_4930), .ZN(n_257_76_4931));
   NAND2_X1 i_257_76_4940 (.A1(n_257_76_4823), .A2(n_257_76_4824), .ZN(
      n_257_76_4932));
   INV_X1 i_257_76_4941 (.A(n_257_76_4932), .ZN(n_257_76_4933));
   NAND4_X1 i_257_76_4942 (.A1(n_257_76_4931), .A2(n_257_76_4933), .A3(
      n_257_76_4829), .A4(n_257_76_4869), .ZN(n_257_76_4934));
   NOR2_X1 i_257_76_4943 (.A1(n_257_76_4923), .A2(n_257_76_4934), .ZN(
      n_257_76_4935));
   NAND2_X1 i_257_76_4944 (.A1(n_257_76_4888), .A2(n_257_76_4833), .ZN(
      n_257_76_4936));
   INV_X1 i_257_76_4945 (.A(n_257_76_4936), .ZN(n_257_76_4937));
   NAND4_X1 i_257_76_4946 (.A1(n_257_76_4834), .A2(n_257_76_4835), .A3(
      n_257_76_4893), .A4(n_257_76_4798), .ZN(n_257_76_4938));
   INV_X1 i_257_76_4947 (.A(n_257_76_4938), .ZN(n_257_76_4939));
   NAND4_X1 i_257_76_4948 (.A1(n_257_76_4935), .A2(n_257_76_4937), .A3(
      n_257_76_4939), .A4(n_257_76_4867), .ZN(n_257_76_4940));
   INV_X1 i_257_76_4949 (.A(n_257_76_4940), .ZN(n_257_76_4941));
   NAND2_X1 i_257_76_4950 (.A1(n_257_76_4838), .A2(n_257_76_4797), .ZN(
      n_257_76_4942));
   INV_X1 i_257_76_4951 (.A(n_257_76_4942), .ZN(n_257_76_4943));
   NAND3_X1 i_257_76_4952 (.A1(n_257_76_4941), .A2(n_257_76_4943), .A3(
      n_257_76_4807), .ZN(n_257_76_4944));
   INV_X1 i_257_76_4953 (.A(n_257_76_4944), .ZN(n_257_76_4945));
   NAND2_X1 i_257_76_4954 (.A1(n_257_76_18074), .A2(n_257_76_4945), .ZN(
      n_257_76_4946));
   NAND3_X1 i_257_76_4955 (.A1(n_257_76_4912), .A2(n_257_76_4922), .A3(
      n_257_76_4946), .ZN(n_257_76_4947));
   NAND2_X1 i_257_76_4956 (.A1(n_257_1067), .A2(n_257_442), .ZN(n_257_76_4948));
   INV_X1 i_257_76_4957 (.A(n_257_76_4948), .ZN(n_257_76_4949));
   NAND2_X1 i_257_76_4958 (.A1(n_257_13), .A2(n_257_76_4949), .ZN(n_257_76_4950));
   NOR2_X1 i_257_76_4959 (.A1(n_257_76_4844), .A2(n_257_76_11918), .ZN(
      n_257_76_4951));
   NAND3_X1 i_257_76_4960 (.A1(n_257_76_4951), .A2(n_257_76_4824), .A3(
      n_257_76_4825), .ZN(n_257_76_4952));
   INV_X1 i_257_76_4961 (.A(n_257_76_4952), .ZN(n_257_76_4953));
   NAND4_X1 i_257_76_4962 (.A1(n_257_76_4798), .A2(n_257_76_4953), .A3(n_257_869), 
      .A4(n_257_76_4817), .ZN(n_257_76_4954));
   INV_X1 i_257_76_4963 (.A(n_257_76_4954), .ZN(n_257_76_4955));
   NAND2_X1 i_257_76_4964 (.A1(n_257_76_4797), .A2(n_257_76_4955), .ZN(
      n_257_76_4956));
   INV_X1 i_257_76_4965 (.A(n_257_76_4956), .ZN(n_257_76_4957));
   NAND2_X1 i_257_76_4966 (.A1(n_257_76_4957), .A2(n_257_76_4807), .ZN(
      n_257_76_4958));
   INV_X1 i_257_76_4967 (.A(n_257_76_4958), .ZN(n_257_76_4959));
   NAND2_X1 i_257_76_4968 (.A1(n_257_76_18077), .A2(n_257_76_4959), .ZN(
      n_257_76_4960));
   NAND2_X1 i_257_76_4969 (.A1(n_257_76_4950), .A2(n_257_76_4960), .ZN(
      n_257_76_4961));
   NOR2_X1 i_257_76_4970 (.A1(n_257_76_4947), .A2(n_257_76_4961), .ZN(
      n_257_76_4962));
   NAND2_X1 i_257_76_4971 (.A1(n_257_76_4869), .A2(n_257_76_4823), .ZN(
      n_257_76_4963));
   INV_X1 i_257_76_4972 (.A(n_257_76_4963), .ZN(n_257_76_4964));
   NAND3_X1 i_257_76_4973 (.A1(n_257_76_4824), .A2(n_257_76_4825), .A3(n_257_541), 
      .ZN(n_257_76_4965));
   INV_X1 i_257_76_4974 (.A(n_257_76_4965), .ZN(n_257_76_4966));
   NAND4_X1 i_257_76_4975 (.A1(n_257_76_4872), .A2(n_257_76_4873), .A3(
      n_257_76_4876), .A4(n_257_426), .ZN(n_257_76_4967));
   INV_X1 i_257_76_4976 (.A(n_257_76_4967), .ZN(n_257_76_4968));
   NAND3_X1 i_257_76_4977 (.A1(n_257_76_4968), .A2(n_257_76_4879), .A3(
      n_257_76_4880), .ZN(n_257_76_4969));
   INV_X1 i_257_76_4978 (.A(n_257_76_4969), .ZN(n_257_76_4970));
   NAND4_X1 i_257_76_4979 (.A1(n_257_76_4964), .A2(n_257_76_4966), .A3(
      n_257_76_4970), .A4(n_257_76_4817), .ZN(n_257_76_4971));
   INV_X1 i_257_76_4980 (.A(n_257_76_4971), .ZN(n_257_76_4972));
   NAND3_X1 i_257_76_4981 (.A1(n_257_76_4867), .A2(n_257_76_4972), .A3(
      n_257_76_4888), .ZN(n_257_76_4973));
   NAND2_X1 i_257_76_4982 (.A1(n_257_76_4833), .A2(n_257_76_4834), .ZN(
      n_257_76_4974));
   INV_X1 i_257_76_4983 (.A(n_257_76_4974), .ZN(n_257_76_4975));
   NAND3_X1 i_257_76_4984 (.A1(n_257_76_4835), .A2(n_257_76_4893), .A3(
      n_257_76_4798), .ZN(n_257_76_4976));
   INV_X1 i_257_76_4985 (.A(n_257_76_4976), .ZN(n_257_76_4977));
   INV_X1 i_257_76_4986 (.A(n_257_76_4894), .ZN(n_257_76_4978));
   NOR2_X1 i_257_76_4987 (.A1(n_257_76_4891), .A2(n_257_76_4978), .ZN(
      n_257_76_4979));
   NAND3_X1 i_257_76_4988 (.A1(n_257_76_4975), .A2(n_257_76_4977), .A3(
      n_257_76_4979), .ZN(n_257_76_4980));
   NOR2_X1 i_257_76_4989 (.A1(n_257_76_4973), .A2(n_257_76_4980), .ZN(
      n_257_76_4981));
   NAND3_X1 i_257_76_4990 (.A1(n_257_76_4981), .A2(n_257_76_4943), .A3(
      n_257_76_4807), .ZN(n_257_76_4982));
   INV_X1 i_257_76_4991 (.A(n_257_76_4982), .ZN(n_257_76_4983));
   NAND2_X1 i_257_76_4992 (.A1(n_257_76_18076), .A2(n_257_76_4983), .ZN(
      n_257_76_4984));
   NAND3_X1 i_257_76_4993 (.A1(n_257_76_4834), .A2(n_257_76_4835), .A3(n_257_741), 
      .ZN(n_257_76_4985));
   NOR2_X1 i_257_76_4994 (.A1(n_257_76_4844), .A2(n_257_76_8311), .ZN(
      n_257_76_4986));
   NAND3_X1 i_257_76_4995 (.A1(n_257_76_4986), .A2(n_257_76_4824), .A3(
      n_257_76_4825), .ZN(n_257_76_4987));
   INV_X1 i_257_76_4996 (.A(n_257_76_4987), .ZN(n_257_76_4988));
   NAND4_X1 i_257_76_4997 (.A1(n_257_76_4914), .A2(n_257_76_4798), .A3(
      n_257_76_4817), .A4(n_257_76_4988), .ZN(n_257_76_4989));
   NOR2_X1 i_257_76_4998 (.A1(n_257_76_4985), .A2(n_257_76_4989), .ZN(
      n_257_76_4990));
   NAND2_X1 i_257_76_4999 (.A1(n_257_76_4797), .A2(n_257_76_4990), .ZN(
      n_257_76_4991));
   NOR2_X1 i_257_76_5000 (.A1(n_257_76_4840), .A2(n_257_76_4991), .ZN(
      n_257_76_4992));
   NAND2_X1 i_257_76_5001 (.A1(n_257_76_18069), .A2(n_257_76_4992), .ZN(
      n_257_76_4993));
   NAND4_X1 i_257_76_5002 (.A1(n_257_76_4833), .A2(n_257_76_4834), .A3(
      n_257_76_4835), .A4(n_257_76_4798), .ZN(n_257_76_4994));
   NAND2_X1 i_257_76_5003 (.A1(n_257_605), .A2(n_257_442), .ZN(n_257_76_4995));
   INV_X1 i_257_76_5004 (.A(n_257_76_4995), .ZN(n_257_76_4996));
   NAND2_X1 i_257_76_5005 (.A1(n_257_432), .A2(n_257_76_4996), .ZN(n_257_76_4997));
   NOR2_X1 i_257_76_5006 (.A1(n_257_76_4997), .A2(n_257_1067), .ZN(n_257_76_4998));
   NAND4_X1 i_257_76_5007 (.A1(n_257_76_4824), .A2(n_257_76_4825), .A3(
      n_257_76_4879), .A4(n_257_76_4998), .ZN(n_257_76_4999));
   NOR2_X1 i_257_76_5008 (.A1(n_257_76_4999), .A2(n_257_76_4963), .ZN(
      n_257_76_5000));
   NAND2_X1 i_257_76_5009 (.A1(n_257_76_4894), .A2(n_257_76_4817), .ZN(
      n_257_76_5001));
   INV_X1 i_257_76_5010 (.A(n_257_76_5001), .ZN(n_257_76_5002));
   NAND3_X1 i_257_76_5011 (.A1(n_257_76_5000), .A2(n_257_76_5002), .A3(
      n_257_76_4892), .ZN(n_257_76_5003));
   NOR2_X1 i_257_76_5012 (.A1(n_257_76_4994), .A2(n_257_76_5003), .ZN(
      n_257_76_5004));
   NAND3_X1 i_257_76_5013 (.A1(n_257_76_5004), .A2(n_257_76_4838), .A3(
      n_257_76_4797), .ZN(n_257_76_5005));
   NOR2_X1 i_257_76_5014 (.A1(n_257_76_5005), .A2(n_257_76_4840), .ZN(
      n_257_76_5006));
   NAND2_X1 i_257_76_5015 (.A1(n_257_68), .A2(n_257_76_5006), .ZN(n_257_76_5007));
   NAND3_X1 i_257_76_5016 (.A1(n_257_76_4984), .A2(n_257_76_4993), .A3(
      n_257_76_5007), .ZN(n_257_76_5008));
   NOR2_X1 i_257_76_5017 (.A1(n_257_76_4844), .A2(n_257_76_15924), .ZN(
      n_257_76_5009));
   NAND3_X1 i_257_76_5018 (.A1(n_257_76_5009), .A2(n_257_76_4824), .A3(
      n_257_76_4825), .ZN(n_257_76_5010));
   INV_X1 i_257_76_5019 (.A(n_257_76_5010), .ZN(n_257_76_5011));
   NAND4_X1 i_257_76_5020 (.A1(n_257_805), .A2(n_257_76_5011), .A3(n_257_76_4817), 
      .A4(n_257_76_4818), .ZN(n_257_76_5012));
   NAND2_X1 i_257_76_5021 (.A1(n_257_76_4835), .A2(n_257_76_4798), .ZN(
      n_257_76_5013));
   NOR2_X1 i_257_76_5022 (.A1(n_257_76_5012), .A2(n_257_76_5013), .ZN(
      n_257_76_5014));
   NAND2_X1 i_257_76_5023 (.A1(n_257_76_4797), .A2(n_257_76_5014), .ZN(
      n_257_76_5015));
   INV_X1 i_257_76_5024 (.A(n_257_76_5015), .ZN(n_257_76_5016));
   NAND2_X1 i_257_76_5025 (.A1(n_257_76_5016), .A2(n_257_76_4807), .ZN(
      n_257_76_5017));
   INV_X1 i_257_76_5026 (.A(n_257_76_5017), .ZN(n_257_76_5018));
   NAND2_X1 i_257_76_5027 (.A1(n_257_22), .A2(n_257_76_5018), .ZN(n_257_76_5019));
   NAND2_X1 i_257_76_5028 (.A1(n_257_444), .A2(n_257_76_4811), .ZN(n_257_76_5020));
   INV_X1 i_257_76_5029 (.A(n_257_76_5020), .ZN(n_257_76_5021));
   NAND2_X1 i_257_76_5030 (.A1(n_257_1003), .A2(n_257_76_5021), .ZN(
      n_257_76_5022));
   INV_X1 i_257_76_5031 (.A(n_257_76_5022), .ZN(n_257_76_5023));
   NAND2_X1 i_257_76_5032 (.A1(n_257_76_4807), .A2(n_257_76_5023), .ZN(
      n_257_76_5024));
   INV_X1 i_257_76_5033 (.A(n_257_76_5024), .ZN(n_257_76_5025));
   NAND2_X1 i_257_76_5034 (.A1(n_257_76_18075), .A2(n_257_76_5025), .ZN(
      n_257_76_5026));
   NAND2_X1 i_257_76_5035 (.A1(n_257_76_5019), .A2(n_257_76_5026), .ZN(
      n_257_76_5027));
   NOR2_X1 i_257_76_5036 (.A1(n_257_76_5008), .A2(n_257_76_5027), .ZN(
      n_257_76_5028));
   NAND3_X1 i_257_76_5037 (.A1(n_257_76_4903), .A2(n_257_76_4962), .A3(
      n_257_76_5028), .ZN(n_257_76_5029));
   INV_X1 i_257_76_5038 (.A(n_257_76_5029), .ZN(n_257_76_5030));
   NOR2_X1 i_257_76_5039 (.A1(n_257_1067), .A2(n_257_76_17633), .ZN(
      n_257_76_5031));
   NAND3_X1 i_257_76_5040 (.A1(n_257_76_4879), .A2(n_257_43), .A3(n_257_76_5031), 
      .ZN(n_257_76_5032));
   NOR2_X1 i_257_76_5041 (.A1(n_257_76_4884), .A2(n_257_76_5032), .ZN(
      n_257_76_5033));
   NAND3_X1 i_257_76_5042 (.A1(n_257_76_5002), .A2(n_257_76_5033), .A3(
      n_257_76_4892), .ZN(n_257_76_5034));
   NOR2_X1 i_257_76_5043 (.A1(n_257_76_4994), .A2(n_257_76_5034), .ZN(
      n_257_76_5035));
   NAND3_X1 i_257_76_5044 (.A1(n_257_76_5035), .A2(n_257_76_4838), .A3(
      n_257_76_4797), .ZN(n_257_76_5036));
   NOR2_X1 i_257_76_5045 (.A1(n_257_76_5036), .A2(n_257_76_4840), .ZN(
      n_257_76_5037));
   NAND2_X1 i_257_76_5046 (.A1(n_257_76_18081), .A2(n_257_76_5037), .ZN(
      n_257_76_5038));
   NAND2_X1 i_257_76_5047 (.A1(n_257_1081), .A2(n_257_76_4811), .ZN(
      n_257_76_5039));
   INV_X1 i_257_76_5048 (.A(n_257_76_5039), .ZN(n_257_76_5040));
   NAND3_X1 i_257_76_5049 (.A1(n_257_76_5040), .A2(n_257_76_4824), .A3(
      n_257_76_4825), .ZN(n_257_76_5041));
   NAND2_X1 i_257_76_5050 (.A1(n_257_76_4823), .A2(n_257_449), .ZN(n_257_76_5042));
   NOR2_X1 i_257_76_5051 (.A1(n_257_76_5041), .A2(n_257_76_5042), .ZN(
      n_257_76_5043));
   NAND4_X1 i_257_76_5052 (.A1(n_257_76_5043), .A2(n_257_76_4914), .A3(
      n_257_76_4798), .A4(n_257_76_4817), .ZN(n_257_76_5044));
   NOR2_X1 i_257_76_5053 (.A1(n_257_76_5044), .A2(n_257_76_4836), .ZN(
      n_257_76_5045));
   NAND3_X1 i_257_76_5054 (.A1(n_257_76_5045), .A2(n_257_76_4838), .A3(
      n_257_76_4797), .ZN(n_257_76_5046));
   NOR2_X1 i_257_76_5055 (.A1(n_257_76_5046), .A2(n_257_76_4840), .ZN(
      n_257_76_5047));
   NAND2_X1 i_257_76_5056 (.A1(n_257_76_18083), .A2(n_257_76_5047), .ZN(
      n_257_76_5048));
   NAND3_X1 i_257_76_5057 (.A1(n_257_76_4828), .A2(n_257_76_4829), .A3(
      n_257_76_4869), .ZN(n_257_76_5049));
   INV_X1 i_257_76_5058 (.A(n_257_76_5049), .ZN(n_257_76_5050));
   NAND3_X1 i_257_76_5059 (.A1(n_257_76_4872), .A2(n_257_76_4873), .A3(
      n_257_76_17331), .ZN(n_257_76_5051));
   INV_X1 i_257_76_5060 (.A(n_257_76_5051), .ZN(n_257_76_5052));
   NAND3_X1 i_257_76_5061 (.A1(n_257_76_4825), .A2(n_257_76_4879), .A3(
      n_257_76_5052), .ZN(n_257_76_5053));
   NOR2_X1 i_257_76_5062 (.A1(n_257_76_5053), .A2(n_257_76_4932), .ZN(
      n_257_76_5054));
   NAND3_X1 i_257_76_5063 (.A1(n_257_76_5050), .A2(n_257_76_4820), .A3(
      n_257_76_5054), .ZN(n_257_76_5055));
   NAND4_X1 i_257_76_5064 (.A1(n_257_76_4835), .A2(n_257_76_4893), .A3(
      n_257_76_4798), .A4(n_257_76_4894), .ZN(n_257_76_5056));
   NOR2_X1 i_257_76_5065 (.A1(n_257_76_5055), .A2(n_257_76_5056), .ZN(
      n_257_76_5057));
   NAND4_X1 i_257_76_5066 (.A1(n_257_76_4888), .A2(n_257_160), .A3(n_257_76_4833), 
      .A4(n_257_76_4834), .ZN(n_257_76_5058));
   INV_X1 i_257_76_5067 (.A(n_257_76_5058), .ZN(n_257_76_5059));
   NAND4_X1 i_257_76_5068 (.A1(n_257_76_5057), .A2(n_257_76_4838), .A3(
      n_257_76_5059), .A4(n_257_76_4797), .ZN(n_257_76_5060));
   NOR2_X1 i_257_76_5069 (.A1(n_257_76_5060), .A2(n_257_76_4840), .ZN(
      n_257_76_5061));
   NAND2_X1 i_257_76_5070 (.A1(n_257_76_18061), .A2(n_257_76_5061), .ZN(
      n_257_76_5062));
   NAND3_X1 i_257_76_5071 (.A1(n_257_76_5038), .A2(n_257_76_5048), .A3(
      n_257_76_5062), .ZN(n_257_76_5063));
   INV_X1 i_257_76_5072 (.A(n_257_76_5063), .ZN(n_257_76_5064));
   NOR2_X1 i_257_76_5073 (.A1(n_257_76_4844), .A2(n_257_76_8215), .ZN(
      n_257_76_5065));
   NAND3_X1 i_257_76_5074 (.A1(n_257_76_5065), .A2(n_257_76_4824), .A3(n_257_438), 
      .ZN(n_257_76_5066));
   INV_X1 i_257_76_5075 (.A(n_257_76_5066), .ZN(n_257_76_5067));
   NAND3_X1 i_257_76_5076 (.A1(n_257_76_4798), .A2(n_257_76_5067), .A3(
      n_257_76_4817), .ZN(n_257_76_5068));
   INV_X1 i_257_76_5077 (.A(n_257_76_5068), .ZN(n_257_76_5069));
   NAND2_X1 i_257_76_5078 (.A1(n_257_76_4797), .A2(n_257_76_5069), .ZN(
      n_257_76_5070));
   INV_X1 i_257_76_5079 (.A(n_257_76_5070), .ZN(n_257_76_5071));
   NAND2_X1 i_257_76_5080 (.A1(n_257_76_5071), .A2(n_257_76_4807), .ZN(
      n_257_76_5072));
   INV_X1 i_257_76_5081 (.A(n_257_76_5072), .ZN(n_257_76_5073));
   NAND2_X1 i_257_76_5082 (.A1(n_257_76_18067), .A2(n_257_76_5073), .ZN(
      n_257_76_5074));
   NAND2_X1 i_257_76_5083 (.A1(n_257_76_4867), .A2(n_257_76_4888), .ZN(
      n_257_76_5075));
   INV_X1 i_257_76_5084 (.A(n_257_76_5075), .ZN(n_257_76_5076));
   NAND2_X1 i_257_76_5085 (.A1(n_257_76_5076), .A2(n_257_76_4797), .ZN(
      n_257_76_5077));
   INV_X1 i_257_76_5086 (.A(n_257_76_5077), .ZN(n_257_76_5078));
   NAND2_X1 i_257_76_5087 (.A1(n_257_280), .A2(n_257_423), .ZN(n_257_76_5079));
   NAND2_X1 i_257_76_5088 (.A1(n_257_76_4820), .A2(n_257_76_5079), .ZN(
      n_257_76_5080));
   NAND2_X1 i_257_76_5089 (.A1(n_257_76_4798), .A2(n_257_76_4894), .ZN(
      n_257_76_5081));
   NOR2_X1 i_257_76_5090 (.A1(n_257_76_5080), .A2(n_257_76_5081), .ZN(
      n_257_76_5082));
   NAND2_X1 i_257_76_5091 (.A1(n_257_318), .A2(n_257_422), .ZN(n_257_76_5083));
   NAND2_X1 i_257_76_5092 (.A1(n_257_76_5083), .A2(n_257_76_4825), .ZN(
      n_257_76_5084));
   NOR2_X1 i_257_76_5093 (.A1(n_257_76_4932), .A2(n_257_76_5084), .ZN(
      n_257_76_5085));
   NAND2_X1 i_257_76_5094 (.A1(n_257_76_4872), .A2(n_257_76_4873), .ZN(
      n_257_76_5086));
   NAND2_X1 i_257_76_5095 (.A1(n_257_76_14086), .A2(n_257_76_4874), .ZN(
      n_257_76_5087));
   OAI21_X1 i_257_76_5096 (.A(n_257_76_5087), .B1(n_257_428), .B2(n_257_76_13825), 
      .ZN(n_257_76_5088));
   NAND2_X1 i_257_76_5097 (.A1(n_257_420), .A2(n_257_76_5088), .ZN(n_257_76_5089));
   NOR2_X1 i_257_76_5098 (.A1(n_257_76_5086), .A2(n_257_76_5089), .ZN(
      n_257_76_5090));
   NAND2_X1 i_257_76_5099 (.A1(n_257_76_5090), .A2(n_257_76_4881), .ZN(
      n_257_76_5091));
   NAND2_X1 i_257_76_5100 (.A1(n_257_76_4879), .A2(n_257_76_4880), .ZN(
      n_257_76_5092));
   NOR2_X1 i_257_76_5101 (.A1(n_257_76_5091), .A2(n_257_76_5092), .ZN(
      n_257_76_5093));
   NAND2_X1 i_257_76_5102 (.A1(n_257_76_5085), .A2(n_257_76_5093), .ZN(
      n_257_76_5094));
   NAND2_X1 i_257_76_5103 (.A1(n_257_76_4868), .A2(n_257_76_4869), .ZN(
      n_257_76_5095));
   INV_X1 i_257_76_5104 (.A(n_257_76_5095), .ZN(n_257_76_5096));
   NAND2_X1 i_257_76_5105 (.A1(n_257_76_4831), .A2(n_257_76_5096), .ZN(
      n_257_76_5097));
   NOR2_X1 i_257_76_5106 (.A1(n_257_76_5094), .A2(n_257_76_5097), .ZN(
      n_257_76_5098));
   NAND2_X1 i_257_76_5107 (.A1(n_257_76_5082), .A2(n_257_76_5098), .ZN(
      n_257_76_5099));
   NAND2_X1 i_257_76_5108 (.A1(n_257_357), .A2(n_257_421), .ZN(n_257_76_5100));
   NAND2_X1 i_257_76_5109 (.A1(n_257_76_5100), .A2(n_257_76_4893), .ZN(
      n_257_76_5101));
   INV_X1 i_257_76_5110 (.A(n_257_76_4835), .ZN(n_257_76_5102));
   NOR2_X1 i_257_76_5111 (.A1(n_257_76_5101), .A2(n_257_76_5102), .ZN(
      n_257_76_5103));
   NAND2_X1 i_257_76_5112 (.A1(n_257_76_4975), .A2(n_257_76_5103), .ZN(
      n_257_76_5104));
   NOR2_X1 i_257_76_5113 (.A1(n_257_76_5099), .A2(n_257_76_5104), .ZN(
      n_257_76_5105));
   NAND2_X1 i_257_76_5114 (.A1(n_257_76_5078), .A2(n_257_76_5105), .ZN(
      n_257_76_5106));
   NAND2_X1 i_257_76_5115 (.A1(n_257_76_4898), .A2(n_257_76_4838), .ZN(
      n_257_76_5107));
   INV_X1 i_257_76_5116 (.A(n_257_76_5107), .ZN(n_257_76_5108));
   NAND2_X1 i_257_76_5117 (.A1(n_257_76_5108), .A2(n_257_76_4807), .ZN(
      n_257_76_5109));
   NOR2_X1 i_257_76_5118 (.A1(n_257_76_5106), .A2(n_257_76_5109), .ZN(
      n_257_76_5110));
   NAND2_X1 i_257_76_5119 (.A1(n_257_76_18073), .A2(n_257_76_5110), .ZN(
      n_257_76_5111));
   INV_X1 i_257_76_5120 (.A(n_257_76_4888), .ZN(n_257_76_5112));
   NOR2_X1 i_257_76_5121 (.A1(n_257_76_4836), .A2(n_257_76_5112), .ZN(
      n_257_76_5113));
   NAND3_X1 i_257_76_5122 (.A1(n_257_76_4872), .A2(n_257_76_4873), .A3(
      n_257_76_17925), .ZN(n_257_76_5114));
   INV_X1 i_257_76_5123 (.A(n_257_76_5114), .ZN(n_257_76_5115));
   NAND3_X1 i_257_76_5124 (.A1(n_257_76_4825), .A2(n_257_76_4879), .A3(
      n_257_76_5115), .ZN(n_257_76_5116));
   NOR2_X1 i_257_76_5125 (.A1(n_257_76_5116), .A2(n_257_76_4932), .ZN(
      n_257_76_5117));
   NAND2_X1 i_257_76_5126 (.A1(n_257_76_4818), .A2(n_257_76_4828), .ZN(
      n_257_76_5118));
   INV_X1 i_257_76_5127 (.A(n_257_76_5118), .ZN(n_257_76_5119));
   NAND2_X1 i_257_76_5128 (.A1(n_257_76_4829), .A2(n_257_76_4869), .ZN(
      n_257_76_5120));
   INV_X1 i_257_76_5129 (.A(n_257_76_5120), .ZN(n_257_76_5121));
   NAND3_X1 i_257_76_5130 (.A1(n_257_76_5117), .A2(n_257_76_5119), .A3(
      n_257_76_5121), .ZN(n_257_76_5122));
   NAND4_X1 i_257_76_5131 (.A1(n_257_76_4798), .A2(n_257_76_4894), .A3(
      n_257_76_4817), .A4(n_257_121), .ZN(n_257_76_5123));
   NOR2_X1 i_257_76_5132 (.A1(n_257_76_5122), .A2(n_257_76_5123), .ZN(
      n_257_76_5124));
   NAND4_X1 i_257_76_5133 (.A1(n_257_76_4838), .A2(n_257_76_4797), .A3(
      n_257_76_5113), .A4(n_257_76_5124), .ZN(n_257_76_5125));
   NOR2_X1 i_257_76_5134 (.A1(n_257_76_5125), .A2(n_257_76_4840), .ZN(
      n_257_76_5126));
   NAND2_X1 i_257_76_5135 (.A1(n_257_76_18068), .A2(n_257_76_5126), .ZN(
      n_257_76_5127));
   NAND3_X1 i_257_76_5136 (.A1(n_257_76_5074), .A2(n_257_76_5111), .A3(
      n_257_76_5127), .ZN(n_257_76_5128));
   INV_X1 i_257_76_5137 (.A(n_257_76_5128), .ZN(n_257_76_5129));
   NAND2_X1 i_257_76_5138 (.A1(n_257_773), .A2(n_257_442), .ZN(n_257_76_5130));
   NOR2_X1 i_257_76_5139 (.A1(n_257_1067), .A2(n_257_76_5130), .ZN(n_257_76_5131));
   NAND4_X1 i_257_76_5140 (.A1(n_257_447), .A2(n_257_76_4824), .A3(n_257_76_4825), 
      .A4(n_257_76_5131), .ZN(n_257_76_5132));
   INV_X1 i_257_76_5141 (.A(n_257_76_5132), .ZN(n_257_76_5133));
   NAND4_X1 i_257_76_5142 (.A1(n_257_76_5133), .A2(n_257_76_4798), .A3(
      n_257_76_4817), .A4(n_257_76_4818), .ZN(n_257_76_5134));
   NAND2_X1 i_257_76_5143 (.A1(n_257_76_4834), .A2(n_257_76_4835), .ZN(
      n_257_76_5135));
   NOR2_X1 i_257_76_5144 (.A1(n_257_76_5134), .A2(n_257_76_5135), .ZN(
      n_257_76_5136));
   NAND2_X1 i_257_76_5145 (.A1(n_257_76_4797), .A2(n_257_76_5136), .ZN(
      n_257_76_5137));
   INV_X1 i_257_76_5146 (.A(n_257_76_5137), .ZN(n_257_76_5138));
   NAND2_X1 i_257_76_5147 (.A1(n_257_76_5138), .A2(n_257_76_4807), .ZN(
      n_257_76_5139));
   INV_X1 i_257_76_5148 (.A(n_257_76_5139), .ZN(n_257_76_5140));
   NAND4_X1 i_257_76_5149 (.A1(n_257_76_4817), .A2(n_257_76_4818), .A3(
      n_257_76_4828), .A4(n_257_76_4829), .ZN(n_257_76_5141));
   INV_X1 i_257_76_5150 (.A(n_257_76_5141), .ZN(n_257_76_5142));
   INV_X1 i_257_76_5151 (.A(n_257_76_5081), .ZN(n_257_76_5143));
   NAND3_X1 i_257_76_5152 (.A1(n_257_76_4872), .A2(n_257_76_4873), .A3(
      n_257_76_17932), .ZN(n_257_76_5144));
   INV_X1 i_257_76_5153 (.A(n_257_76_5144), .ZN(n_257_76_5145));
   NAND4_X1 i_257_76_5154 (.A1(n_257_76_4824), .A2(n_257_76_4825), .A3(
      n_257_76_4879), .A4(n_257_76_5145), .ZN(n_257_76_5146));
   NOR2_X1 i_257_76_5155 (.A1(n_257_76_5146), .A2(n_257_76_4963), .ZN(
      n_257_76_5147));
   NAND3_X1 i_257_76_5156 (.A1(n_257_76_5142), .A2(n_257_76_5143), .A3(
      n_257_76_5147), .ZN(n_257_76_5148));
   NAND4_X1 i_257_76_5157 (.A1(n_257_76_4833), .A2(n_257_76_4834), .A3(n_257_83), 
      .A4(n_257_76_4835), .ZN(n_257_76_5149));
   NOR2_X1 i_257_76_5158 (.A1(n_257_76_5148), .A2(n_257_76_5149), .ZN(
      n_257_76_5150));
   NAND3_X1 i_257_76_5159 (.A1(n_257_76_5150), .A2(n_257_76_4838), .A3(
      n_257_76_4797), .ZN(n_257_76_5151));
   NOR2_X1 i_257_76_5160 (.A1(n_257_76_5151), .A2(n_257_76_4840), .ZN(
      n_257_76_5152));
   AOI22_X1 i_257_76_5161 (.A1(n_257_76_18085), .A2(n_257_76_5140), .B1(
      n_257_76_18080), .B2(n_257_76_5152), .ZN(n_257_76_5153));
   NAND3_X1 i_257_76_5162 (.A1(n_257_76_5064), .A2(n_257_76_5129), .A3(
      n_257_76_5153), .ZN(n_257_76_5154));
   INV_X1 i_257_76_5163 (.A(n_257_76_4829), .ZN(n_257_76_5155));
   NAND3_X1 i_257_76_5164 (.A1(n_257_76_4824), .A2(n_257_76_4825), .A3(n_257_448), 
      .ZN(n_257_76_5156));
   NOR2_X1 i_257_76_5165 (.A1(n_257_76_5155), .A2(n_257_76_5156), .ZN(
      n_257_76_5157));
   NAND2_X1 i_257_76_5166 (.A1(n_257_76_4811), .A2(n_257_76_17760), .ZN(
      n_257_76_5158));
   OAI21_X1 i_257_76_5167 (.A(n_257_76_5158), .B1(n_257_709), .B2(n_257_76_4844), 
      .ZN(n_257_76_5159));
   NAND2_X1 i_257_76_5168 (.A1(n_257_76_4818), .A2(n_257_76_5159), .ZN(
      n_257_76_5160));
   INV_X1 i_257_76_5169 (.A(n_257_76_5160), .ZN(n_257_76_5161));
   NAND4_X1 i_257_76_5170 (.A1(n_257_76_5157), .A2(n_257_76_5161), .A3(
      n_257_76_4798), .A4(n_257_76_4817), .ZN(n_257_76_5162));
   NOR2_X1 i_257_76_5171 (.A1(n_257_76_5162), .A2(n_257_76_4836), .ZN(
      n_257_76_5163));
   NAND3_X1 i_257_76_5172 (.A1(n_257_76_5163), .A2(n_257_76_4797), .A3(n_257_677), 
      .ZN(n_257_76_5164));
   NOR2_X1 i_257_76_5173 (.A1(n_257_76_5164), .A2(n_257_76_4840), .ZN(
      n_257_76_5165));
   NAND2_X1 i_257_76_5174 (.A1(n_257_76_18079), .A2(n_257_76_5165), .ZN(
      n_257_76_5166));
   NAND4_X1 i_257_76_5175 (.A1(n_257_76_4872), .A2(n_257_76_4873), .A3(
      n_257_76_4876), .A4(n_257_425), .ZN(n_257_76_5167));
   INV_X1 i_257_76_5176 (.A(n_257_76_5167), .ZN(n_257_76_5168));
   NAND4_X1 i_257_76_5177 (.A1(n_257_76_5168), .A2(n_257_76_4825), .A3(
      n_257_76_4879), .A4(n_257_76_4880), .ZN(n_257_76_5169));
   NAND3_X1 i_257_76_5178 (.A1(n_257_76_4869), .A2(n_257_76_4823), .A3(
      n_257_76_4824), .ZN(n_257_76_5170));
   NOR2_X1 i_257_76_5179 (.A1(n_257_76_5169), .A2(n_257_76_5170), .ZN(
      n_257_76_5171));
   NAND3_X1 i_257_76_5180 (.A1(n_257_76_4828), .A2(n_257_76_4829), .A3(
      n_257_76_4868), .ZN(n_257_76_5172));
   INV_X1 i_257_76_5181 (.A(n_257_76_5172), .ZN(n_257_76_5173));
   NAND3_X1 i_257_76_5182 (.A1(n_257_76_5171), .A2(n_257_76_5173), .A3(
      n_257_76_4820), .ZN(n_257_76_5174));
   NOR2_X1 i_257_76_5183 (.A1(n_257_76_5174), .A2(n_257_76_5056), .ZN(
      n_257_76_5175));
   NAND3_X1 i_257_76_5184 (.A1(n_257_76_4867), .A2(n_257_76_4975), .A3(
      n_257_76_4888), .ZN(n_257_76_5176));
   INV_X1 i_257_76_5185 (.A(n_257_76_5176), .ZN(n_257_76_5177));
   NAND4_X1 i_257_76_5186 (.A1(n_257_76_5175), .A2(n_257_76_5177), .A3(
      n_257_76_4838), .A4(n_257_240), .ZN(n_257_76_5178));
   NAND2_X1 i_257_76_5187 (.A1(n_257_76_4807), .A2(n_257_76_4797), .ZN(
      n_257_76_5179));
   NOR2_X1 i_257_76_5188 (.A1(n_257_76_5178), .A2(n_257_76_5179), .ZN(
      n_257_76_5180));
   NAND2_X1 i_257_76_5189 (.A1(n_257_76_18064), .A2(n_257_76_5180), .ZN(
      n_257_76_5181));
   INV_X1 i_257_76_5190 (.A(n_257_76_4836), .ZN(n_257_76_5182));
   NAND4_X1 i_257_76_5191 (.A1(n_257_76_4894), .A2(n_257_76_5079), .A3(
      n_257_76_4817), .A4(n_257_357), .ZN(n_257_76_5183));
   NAND2_X1 i_257_76_5192 (.A1(n_257_76_4893), .A2(n_257_76_4798), .ZN(
      n_257_76_5184));
   NOR2_X1 i_257_76_5193 (.A1(n_257_76_5183), .A2(n_257_76_5184), .ZN(
      n_257_76_5185));
   NAND4_X1 i_257_76_5194 (.A1(n_257_76_4872), .A2(n_257_76_4873), .A3(
      n_257_76_4876), .A4(n_257_421), .ZN(n_257_76_5186));
   INV_X1 i_257_76_5195 (.A(n_257_76_5186), .ZN(n_257_76_5187));
   NAND4_X1 i_257_76_5196 (.A1(n_257_76_5187), .A2(n_257_76_4879), .A3(
      n_257_76_4880), .A4(n_257_76_4881), .ZN(n_257_76_5188));
   INV_X1 i_257_76_5197 (.A(n_257_76_5188), .ZN(n_257_76_5189));
   NAND3_X1 i_257_76_5198 (.A1(n_257_76_4824), .A2(n_257_76_5083), .A3(
      n_257_76_4825), .ZN(n_257_76_5190));
   INV_X1 i_257_76_5199 (.A(n_257_76_5190), .ZN(n_257_76_5191));
   NAND3_X1 i_257_76_5200 (.A1(n_257_76_5189), .A2(n_257_76_4964), .A3(
      n_257_76_5191), .ZN(n_257_76_5192));
   NAND4_X1 i_257_76_5201 (.A1(n_257_76_4818), .A2(n_257_76_4828), .A3(
      n_257_76_4829), .A4(n_257_76_4868), .ZN(n_257_76_5193));
   NOR2_X1 i_257_76_5202 (.A1(n_257_76_5192), .A2(n_257_76_5193), .ZN(
      n_257_76_5194));
   NAND4_X1 i_257_76_5203 (.A1(n_257_76_5182), .A2(n_257_76_5185), .A3(
      n_257_76_5194), .A4(n_257_76_4888), .ZN(n_257_76_5195));
   INV_X1 i_257_76_5204 (.A(n_257_76_5195), .ZN(n_257_76_5196));
   NAND2_X1 i_257_76_5205 (.A1(n_257_76_4807), .A2(n_257_76_5196), .ZN(
      n_257_76_5197));
   NAND4_X1 i_257_76_5206 (.A1(n_257_76_4898), .A2(n_257_76_4838), .A3(
      n_257_76_4797), .A4(n_257_76_4867), .ZN(n_257_76_5198));
   NOR2_X1 i_257_76_5207 (.A1(n_257_76_5197), .A2(n_257_76_5198), .ZN(
      n_257_76_5199));
   NAND2_X1 i_257_76_5208 (.A1(n_257_76_18082), .A2(n_257_76_5199), .ZN(
      n_257_76_5200));
   NAND3_X1 i_257_76_5209 (.A1(n_257_76_5166), .A2(n_257_76_5181), .A3(
      n_257_76_5200), .ZN(n_257_76_5201));
   INV_X1 i_257_76_5210 (.A(n_257_76_5201), .ZN(n_257_76_5202));
   NAND3_X1 i_257_76_5211 (.A1(n_257_76_4824), .A2(n_257_76_4825), .A3(
      n_257_76_4879), .ZN(n_257_76_5203));
   INV_X1 i_257_76_5212 (.A(n_257_76_5203), .ZN(n_257_76_5204));
   NAND2_X1 i_257_76_5213 (.A1(n_257_76_4964), .A2(n_257_76_5204), .ZN(
      n_257_76_5205));
   NOR2_X1 i_257_76_5214 (.A1(n_257_76_5205), .A2(n_257_76_4891), .ZN(
      n_257_76_5206));
   NAND2_X1 i_257_76_5215 (.A1(n_257_76_4835), .A2(n_257_76_4893), .ZN(
      n_257_76_5207));
   INV_X1 i_257_76_5216 (.A(n_257_76_5207), .ZN(n_257_76_5208));
   INV_X1 i_257_76_5217 (.A(n_257_76_4876), .ZN(n_257_76_5209));
   NOR2_X1 i_257_76_5218 (.A1(n_257_76_5209), .A2(n_257_1067), .ZN(n_257_76_5210));
   NAND4_X1 i_257_76_5219 (.A1(n_257_76_5210), .A2(n_257_200), .A3(n_257_427), 
      .A4(n_257_76_4872), .ZN(n_257_76_5211));
   INV_X1 i_257_76_5220 (.A(n_257_76_5211), .ZN(n_257_76_5212));
   NAND4_X1 i_257_76_5221 (.A1(n_257_76_4798), .A2(n_257_76_4894), .A3(
      n_257_76_4817), .A4(n_257_76_5212), .ZN(n_257_76_5213));
   INV_X1 i_257_76_5222 (.A(n_257_76_5213), .ZN(n_257_76_5214));
   NAND3_X1 i_257_76_5223 (.A1(n_257_76_5206), .A2(n_257_76_5208), .A3(
      n_257_76_5214), .ZN(n_257_76_5215));
   NOR2_X1 i_257_76_5224 (.A1(n_257_76_5176), .A2(n_257_76_5215), .ZN(
      n_257_76_5216));
   NAND3_X1 i_257_76_5225 (.A1(n_257_76_5216), .A2(n_257_76_4943), .A3(
      n_257_76_4807), .ZN(n_257_76_5217));
   INV_X1 i_257_76_5226 (.A(n_257_76_5217), .ZN(n_257_76_5218));
   NAND2_X1 i_257_76_5227 (.A1(n_257_76_18065), .A2(n_257_76_5218), .ZN(
      n_257_76_5219));
   INV_X1 i_257_76_5228 (.A(n_257_460), .ZN(n_257_76_5220));
   NOR2_X1 i_257_76_5229 (.A1(n_257_76_4844), .A2(n_257_76_5220), .ZN(
      n_257_76_5221));
   NAND3_X1 i_257_76_5230 (.A1(n_257_76_5221), .A2(n_257_76_4825), .A3(
      n_257_76_4879), .ZN(n_257_76_5222));
   NOR2_X1 i_257_76_5231 (.A1(n_257_76_5222), .A2(n_257_76_4932), .ZN(
      n_257_76_5223));
   NAND3_X1 i_257_76_5232 (.A1(n_257_76_4828), .A2(n_257_76_4829), .A3(n_257_451), 
      .ZN(n_257_76_5224));
   INV_X1 i_257_76_5233 (.A(n_257_76_5224), .ZN(n_257_76_5225));
   NAND4_X1 i_257_76_5234 (.A1(n_257_76_5223), .A2(n_257_76_5225), .A3(
      n_257_76_4820), .A4(n_257_76_4798), .ZN(n_257_76_5226));
   NOR2_X1 i_257_76_5235 (.A1(n_257_76_5226), .A2(n_257_76_4836), .ZN(
      n_257_76_5227));
   NAND3_X1 i_257_76_5236 (.A1(n_257_76_5227), .A2(n_257_76_4838), .A3(
      n_257_76_4797), .ZN(n_257_76_5228));
   NOR2_X1 i_257_76_5237 (.A1(n_257_76_5228), .A2(n_257_76_4840), .ZN(
      n_257_76_5229));
   NAND2_X1 i_257_76_5238 (.A1(n_257_76_18063), .A2(n_257_76_5229), .ZN(
      n_257_76_5230));
   NAND4_X1 i_257_76_5239 (.A1(n_257_76_4824), .A2(n_257_76_4825), .A3(
      n_257_76_4879), .A4(n_257_76_4880), .ZN(n_257_76_5231));
   NOR2_X1 i_257_76_5240 (.A1(n_257_76_5231), .A2(n_257_76_4963), .ZN(
      n_257_76_5232));
   NAND3_X1 i_257_76_5241 (.A1(n_257_76_4817), .A2(n_257_76_4818), .A3(
      n_257_76_4828), .ZN(n_257_76_5233));
   INV_X1 i_257_76_5242 (.A(n_257_76_5233), .ZN(n_257_76_5234));
   NAND2_X1 i_257_76_5243 (.A1(n_257_76_4876), .A2(n_257_424), .ZN(n_257_76_5235));
   INV_X1 i_257_76_5244 (.A(n_257_76_5235), .ZN(n_257_76_5236));
   NAND4_X1 i_257_76_5245 (.A1(n_257_76_5236), .A2(n_257_509), .A3(n_257_76_4872), 
      .A4(n_257_76_4873), .ZN(n_257_76_5237));
   INV_X1 i_257_76_5246 (.A(n_257_76_5237), .ZN(n_257_76_5238));
   NAND3_X1 i_257_76_5247 (.A1(n_257_76_4829), .A2(n_257_76_5238), .A3(
      n_257_76_4868), .ZN(n_257_76_5239));
   INV_X1 i_257_76_5248 (.A(n_257_76_5239), .ZN(n_257_76_5240));
   NAND3_X1 i_257_76_5249 (.A1(n_257_76_5232), .A2(n_257_76_5234), .A3(
      n_257_76_5240), .ZN(n_257_76_5241));
   NOR2_X1 i_257_76_5250 (.A1(n_257_76_5241), .A2(n_257_76_5056), .ZN(
      n_257_76_5242));
   NAND4_X1 i_257_76_5251 (.A1(n_257_76_5242), .A2(n_257_76_5177), .A3(
      n_257_76_4838), .A4(n_257_76_4797), .ZN(n_257_76_5243));
   NOR2_X1 i_257_76_5252 (.A1(n_257_76_5243), .A2(n_257_76_4899), .ZN(
      n_257_76_5244));
   NAND2_X1 i_257_76_5253 (.A1(n_257_76_18062), .A2(n_257_76_5244), .ZN(
      n_257_76_5245));
   NAND3_X1 i_257_76_5254 (.A1(n_257_76_5219), .A2(n_257_76_5230), .A3(
      n_257_76_5245), .ZN(n_257_76_5246));
   INV_X1 i_257_76_5255 (.A(n_257_76_5246), .ZN(n_257_76_5247));
   NAND3_X1 i_257_76_5256 (.A1(n_257_76_4868), .A2(n_257_76_4869), .A3(
      n_257_76_4823), .ZN(n_257_76_5248));
   NOR2_X1 i_257_76_5257 (.A1(n_257_76_5248), .A2(n_257_76_5231), .ZN(
      n_257_76_5249));
   INV_X1 i_257_76_5258 (.A(n_257_76_5086), .ZN(n_257_76_5250));
   NAND2_X1 i_257_76_5259 (.A1(n_257_76_4876), .A2(n_257_422), .ZN(n_257_76_5251));
   INV_X1 i_257_76_5260 (.A(n_257_76_5251), .ZN(n_257_76_5252));
   NAND4_X1 i_257_76_5261 (.A1(n_257_76_4881), .A2(n_257_76_5250), .A3(n_257_318), 
      .A4(n_257_76_5252), .ZN(n_257_76_5253));
   INV_X1 i_257_76_5262 (.A(n_257_76_5253), .ZN(n_257_76_5254));
   NAND3_X1 i_257_76_5263 (.A1(n_257_76_5079), .A2(n_257_76_4817), .A3(
      n_257_76_5254), .ZN(n_257_76_5255));
   INV_X1 i_257_76_5264 (.A(n_257_76_5255), .ZN(n_257_76_5256));
   NAND3_X1 i_257_76_5265 (.A1(n_257_76_5249), .A2(n_257_76_5256), .A3(
      n_257_76_4892), .ZN(n_257_76_5257));
   NOR2_X1 i_257_76_5266 (.A1(n_257_76_5257), .A2(n_257_76_5056), .ZN(
      n_257_76_5258));
   NAND4_X1 i_257_76_5267 (.A1(n_257_76_5258), .A2(n_257_76_5177), .A3(
      n_257_76_4838), .A4(n_257_76_4797), .ZN(n_257_76_5259));
   NOR2_X1 i_257_76_5268 (.A1(n_257_76_5259), .A2(n_257_76_4899), .ZN(
      n_257_76_5260));
   NAND2_X1 i_257_76_5269 (.A1(n_257_342), .A2(n_257_76_5260), .ZN(n_257_76_5261));
   NAND3_X1 i_257_76_5270 (.A1(n_257_76_4823), .A2(n_257_76_4824), .A3(
      n_257_76_5083), .ZN(n_257_76_5262));
   INV_X1 i_257_76_5271 (.A(n_257_76_5262), .ZN(n_257_76_5263));
   NAND3_X1 i_257_76_5272 (.A1(n_257_76_4825), .A2(n_257_76_4879), .A3(
      n_257_76_4880), .ZN(n_257_76_5264));
   INV_X1 i_257_76_5273 (.A(n_257_76_5264), .ZN(n_257_76_5265));
   NAND2_X1 i_257_76_5274 (.A1(n_257_428), .A2(n_257_573), .ZN(n_257_76_5266));
   NAND3_X1 i_257_76_5275 (.A1(n_257_396), .A2(n_257_484), .A3(n_257_442), 
      .ZN(n_257_76_5267));
   INV_X1 i_257_76_5276 (.A(n_257_76_5267), .ZN(n_257_76_5268));
   NAND2_X1 i_257_76_5277 (.A1(n_257_76_5266), .A2(n_257_76_5268), .ZN(
      n_257_76_5269));
   NOR2_X1 i_257_76_5278 (.A1(n_257_76_5269), .A2(n_257_1067), .ZN(n_257_76_5270));
   NAND2_X1 i_257_76_5279 (.A1(n_257_420), .A2(n_257_661), .ZN(n_257_76_5271));
   NAND4_X1 i_257_76_5280 (.A1(n_257_76_5270), .A2(n_257_76_4881), .A3(
      n_257_76_5271), .A4(n_257_76_4872), .ZN(n_257_76_5272));
   INV_X1 i_257_76_5281 (.A(n_257_76_5272), .ZN(n_257_76_5273));
   NAND3_X1 i_257_76_5282 (.A1(n_257_76_5263), .A2(n_257_76_5265), .A3(
      n_257_76_5273), .ZN(n_257_76_5274));
   NAND4_X1 i_257_76_5283 (.A1(n_257_76_4828), .A2(n_257_76_4829), .A3(
      n_257_76_4868), .A4(n_257_76_4869), .ZN(n_257_76_5275));
   NOR2_X1 i_257_76_5284 (.A1(n_257_76_5274), .A2(n_257_76_5275), .ZN(
      n_257_76_5276));
   NAND3_X1 i_257_76_5285 (.A1(n_257_76_5276), .A2(n_257_76_4867), .A3(
      n_257_76_4888), .ZN(n_257_76_5277));
   NAND3_X1 i_257_76_5286 (.A1(n_257_76_5079), .A2(n_257_76_4817), .A3(
      n_257_76_4818), .ZN(n_257_76_5278));
   NOR2_X1 i_257_76_5287 (.A1(n_257_76_5081), .A2(n_257_76_5278), .ZN(
      n_257_76_5279));
   NAND3_X1 i_257_76_5288 (.A1(n_257_76_4835), .A2(n_257_76_5100), .A3(
      n_257_76_4893), .ZN(n_257_76_5280));
   INV_X1 i_257_76_5289 (.A(n_257_76_5280), .ZN(n_257_76_5281));
   NAND3_X1 i_257_76_5290 (.A1(n_257_76_5279), .A2(n_257_76_4975), .A3(
      n_257_76_5281), .ZN(n_257_76_5282));
   NOR2_X1 i_257_76_5291 (.A1(n_257_76_5277), .A2(n_257_76_5282), .ZN(
      n_257_76_5283));
   NAND4_X1 i_257_76_5292 (.A1(n_257_76_5283), .A2(n_257_76_4943), .A3(
      n_257_76_4807), .A4(n_257_76_4898), .ZN(n_257_76_5284));
   INV_X1 i_257_76_5293 (.A(n_257_76_5284), .ZN(n_257_76_5285));
   NAND2_X1 i_257_76_5294 (.A1(n_257_76_18060), .A2(n_257_76_5285), .ZN(
      n_257_76_5286));
   INV_X1 i_257_76_5295 (.A(n_257_76_5130), .ZN(n_257_76_5287));
   NAND2_X1 i_257_76_5296 (.A1(n_257_447), .A2(n_257_76_5287), .ZN(n_257_76_5288));
   INV_X1 i_257_76_5297 (.A(Small_Packet_Data_Size[8]), .ZN(n_257_76_5289));
   NAND2_X1 i_257_76_5298 (.A1(n_257_76_5266), .A2(n_257_76_18049), .ZN(
      n_257_76_5290));
   INV_X1 i_257_76_5299 (.A(n_257_76_5290), .ZN(n_257_76_5291));
   NAND3_X1 i_257_76_5300 (.A1(n_257_76_5291), .A2(n_257_76_5271), .A3(
      n_257_76_4873), .ZN(n_257_76_5292));
   NAND2_X1 i_257_76_5301 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[8]), 
      .ZN(n_257_76_5293));
   NAND2_X1 i_257_76_5302 (.A1(n_257_76_5292), .A2(n_257_76_5293), .ZN(
      n_257_76_5294));
   NAND3_X1 i_257_76_5303 (.A1(n_257_76_5253), .A2(n_257_76_5288), .A3(
      n_257_76_5294), .ZN(n_257_76_5295));
   NAND2_X1 i_257_76_5304 (.A1(n_257_837), .A2(n_257_442), .ZN(n_257_76_5296));
   INV_X1 i_257_76_5305 (.A(n_257_76_5296), .ZN(n_257_76_5297));
   NAND2_X1 i_257_76_5306 (.A1(n_257_446), .A2(n_257_76_5297), .ZN(n_257_76_5298));
   NAND2_X1 i_257_76_5307 (.A1(n_257_449), .A2(n_257_76_12626), .ZN(
      n_257_76_5299));
   NAND2_X1 i_257_76_5308 (.A1(n_257_76_5298), .A2(n_257_76_5299), .ZN(
      n_257_76_5300));
   NOR2_X1 i_257_76_5309 (.A1(n_257_76_5295), .A2(n_257_76_5300), .ZN(
      n_257_76_5301));
   NAND2_X1 i_257_76_5310 (.A1(n_257_971), .A2(n_257_442), .ZN(n_257_76_5302));
   INV_X1 i_257_76_5311 (.A(n_257_76_5302), .ZN(n_257_76_5303));
   NAND2_X1 i_257_76_5312 (.A1(n_257_441), .A2(n_257_76_5303), .ZN(n_257_76_5304));
   NAND2_X1 i_257_76_5313 (.A1(n_257_460), .A2(n_257_442), .ZN(n_257_76_5305));
   INV_X1 i_257_76_5314 (.A(n_257_76_5305), .ZN(n_257_76_5306));
   NAND2_X1 i_257_76_5315 (.A1(n_257_451), .A2(n_257_76_5306), .ZN(n_257_76_5307));
   NAND2_X1 i_257_76_5316 (.A1(n_257_907), .A2(n_257_76_17940), .ZN(
      n_257_76_5308));
   NAND3_X1 i_257_76_5317 (.A1(n_257_76_5304), .A2(n_257_76_5307), .A3(
      n_257_76_5308), .ZN(n_257_76_5309));
   INV_X1 i_257_76_5318 (.A(n_257_76_5309), .ZN(n_257_76_5310));
   NAND2_X1 i_257_76_5319 (.A1(n_257_43), .A2(n_257_76_17918), .ZN(n_257_76_5311));
   NAND2_X1 i_257_76_5320 (.A1(n_257_709), .A2(n_257_76_15655), .ZN(
      n_257_76_5312));
   NAND4_X1 i_257_76_5321 (.A1(n_257_76_5311), .A2(n_257_76_5211), .A3(
      n_257_76_5312), .A4(n_257_76_5237), .ZN(n_257_76_5313));
   INV_X1 i_257_76_5322 (.A(n_257_76_4799), .ZN(n_257_76_5314));
   NAND2_X1 i_257_76_5323 (.A1(n_257_440), .A2(n_257_76_5314), .ZN(n_257_76_5315));
   NAND2_X1 i_257_76_5324 (.A1(n_257_438), .A2(n_257_76_8280), .ZN(n_257_76_5316));
   NAND2_X1 i_257_76_5325 (.A1(n_257_637), .A2(n_257_76_17928), .ZN(
      n_257_76_5317));
   NAND4_X1 i_257_76_5326 (.A1(n_257_76_5315), .A2(n_257_76_5316), .A3(
      n_257_76_5317), .A4(n_257_76_4997), .ZN(n_257_76_5318));
   NOR2_X1 i_257_76_5327 (.A1(n_257_76_5313), .A2(n_257_76_5318), .ZN(
      n_257_76_5319));
   NAND3_X1 i_257_76_5328 (.A1(n_257_76_5301), .A2(n_257_76_5310), .A3(
      n_257_76_5319), .ZN(n_257_76_5320));
   NAND2_X1 i_257_76_5329 (.A1(n_257_741), .A2(n_257_76_17935), .ZN(
      n_257_76_5321));
   NAND2_X1 i_257_76_5330 (.A1(n_257_805), .A2(n_257_76_17952), .ZN(
      n_257_76_5322));
   NAND2_X1 i_257_76_5331 (.A1(n_257_869), .A2(n_257_76_17903), .ZN(
      n_257_76_5323));
   NAND2_X1 i_257_76_5332 (.A1(n_257_121), .A2(n_257_76_17925), .ZN(
      n_257_76_5324));
   NAND4_X1 i_257_76_5333 (.A1(n_257_76_5321), .A2(n_257_76_5322), .A3(
      n_257_76_5323), .A4(n_257_76_5324), .ZN(n_257_76_5325));
   NOR2_X1 i_257_76_5334 (.A1(n_257_76_5320), .A2(n_257_76_5325), .ZN(
      n_257_76_5326));
   NAND2_X1 i_257_76_5335 (.A1(n_257_83), .A2(n_257_76_17932), .ZN(n_257_76_5327));
   NAND3_X1 i_257_76_5336 (.A1(n_257_76_4886), .A2(n_257_76_5327), .A3(
      n_257_76_4971), .ZN(n_257_76_5328));
   NAND2_X1 i_257_76_5337 (.A1(n_257_160), .A2(n_257_76_17331), .ZN(
      n_257_76_5329));
   INV_X1 i_257_76_5338 (.A(n_257_76_5329), .ZN(n_257_76_5330));
   NOR2_X1 i_257_76_5339 (.A1(n_257_76_5328), .A2(n_257_76_5330), .ZN(
      n_257_76_5331));
   NAND2_X1 i_257_76_5340 (.A1(n_257_677), .A2(n_257_76_17958), .ZN(
      n_257_76_5332));
   NAND2_X1 i_257_76_5341 (.A1(n_257_1003), .A2(n_257_76_17964), .ZN(
      n_257_76_5333));
   NAND4_X1 i_257_76_5342 (.A1(n_257_76_5326), .A2(n_257_76_5331), .A3(
      n_257_76_5332), .A4(n_257_76_5333), .ZN(n_257_76_5334));
   INV_X1 i_257_76_5343 (.A(n_257_76_5334), .ZN(n_257_76_5335));
   INV_X1 i_257_76_5344 (.A(n_257_1035), .ZN(n_257_76_5336));
   OAI21_X1 i_257_76_5345 (.A(n_257_76_5195), .B1(n_257_76_5336), .B2(
      n_257_76_17968), .ZN(n_257_76_5337));
   INV_X1 i_257_76_5346 (.A(n_257_76_5337), .ZN(n_257_76_5338));
   NAND3_X1 i_257_76_5347 (.A1(n_257_76_5335), .A2(n_257_76_5338), .A3(
      n_257_76_5178), .ZN(n_257_76_5339));
   NAND3_X1 i_257_76_5348 (.A1(n_257_76_5261), .A2(n_257_76_5286), .A3(
      n_257_76_5339), .ZN(n_257_76_5340));
   INV_X1 i_257_76_5349 (.A(n_257_76_5340), .ZN(n_257_76_5341));
   NAND3_X1 i_257_76_5350 (.A1(n_257_76_5202), .A2(n_257_76_5247), .A3(
      n_257_76_5341), .ZN(n_257_76_5342));
   NOR2_X1 i_257_76_5351 (.A1(n_257_76_5154), .A2(n_257_76_5342), .ZN(
      n_257_76_5343));
   NAND2_X1 i_257_76_5352 (.A1(n_257_76_5030), .A2(n_257_76_5343), .ZN(n_8));
   NAND2_X1 i_257_76_5353 (.A1(n_257_1036), .A2(n_257_443), .ZN(n_257_76_5344));
   NAND2_X1 i_257_76_5354 (.A1(n_257_1004), .A2(n_257_444), .ZN(n_257_76_5345));
   NAND2_X1 i_257_76_5355 (.A1(n_257_441), .A2(n_257_972), .ZN(n_257_76_5346));
   INV_X1 i_257_76_5356 (.A(n_257_1068), .ZN(n_257_76_5347));
   NAND2_X1 i_257_76_5357 (.A1(n_257_940), .A2(n_257_442), .ZN(n_257_76_5348));
   INV_X1 i_257_76_5358 (.A(n_257_76_5348), .ZN(n_257_76_5349));
   NAND3_X1 i_257_76_5359 (.A1(n_257_76_5347), .A2(n_257_440), .A3(n_257_76_5349), 
      .ZN(n_257_76_5350));
   INV_X1 i_257_76_5360 (.A(n_257_76_5350), .ZN(n_257_76_5351));
   NAND2_X1 i_257_76_5361 (.A1(n_257_76_5346), .A2(n_257_76_5351), .ZN(
      n_257_76_5352));
   INV_X1 i_257_76_5362 (.A(n_257_76_5352), .ZN(n_257_76_5353));
   NAND2_X1 i_257_76_5363 (.A1(n_257_76_5345), .A2(n_257_76_5353), .ZN(
      n_257_76_5354));
   INV_X1 i_257_76_5364 (.A(n_257_76_5354), .ZN(n_257_76_5355));
   NAND2_X1 i_257_76_5365 (.A1(n_257_76_5344), .A2(n_257_76_5355), .ZN(
      n_257_76_5356));
   INV_X1 i_257_76_5366 (.A(n_257_76_5356), .ZN(n_257_76_5357));
   NAND2_X1 i_257_76_5367 (.A1(n_257_17), .A2(n_257_76_5357), .ZN(n_257_76_5358));
   NOR2_X1 i_257_76_5368 (.A1(n_257_1068), .A2(n_257_76_17412), .ZN(
      n_257_76_5359));
   INV_X1 i_257_76_5369 (.A(n_257_76_5359), .ZN(n_257_76_5360));
   NOR2_X1 i_257_76_5370 (.A1(n_257_76_5360), .A2(n_257_76_15197), .ZN(
      n_257_76_5361));
   NAND2_X1 i_257_76_5371 (.A1(n_257_1036), .A2(n_257_76_5361), .ZN(
      n_257_76_5362));
   INV_X1 i_257_76_5372 (.A(n_257_76_5362), .ZN(n_257_76_5363));
   NAND2_X1 i_257_76_5373 (.A1(n_257_76_18072), .A2(n_257_76_5363), .ZN(
      n_257_76_5364));
   NAND2_X1 i_257_76_5374 (.A1(n_257_710), .A2(n_257_435), .ZN(n_257_76_5365));
   NAND2_X1 i_257_76_5375 (.A1(n_257_446), .A2(n_257_838), .ZN(n_257_76_5366));
   NAND2_X1 i_257_76_5376 (.A1(n_257_449), .A2(n_257_1082), .ZN(n_257_76_5367));
   NAND3_X1 i_257_76_5377 (.A1(n_257_76_5365), .A2(n_257_76_5366), .A3(
      n_257_76_5367), .ZN(n_257_76_5368));
   NAND3_X1 i_257_76_5378 (.A1(n_257_638), .A2(n_257_76_5347), .A3(
      n_257_76_17928), .ZN(n_257_76_5369));
   INV_X1 i_257_76_5379 (.A(n_257_76_5369), .ZN(n_257_76_5370));
   NAND2_X1 i_257_76_5380 (.A1(n_257_447), .A2(n_257_774), .ZN(n_257_76_5371));
   NAND2_X1 i_257_76_5381 (.A1(n_257_438), .A2(n_257_1074), .ZN(n_257_76_5372));
   NAND2_X1 i_257_76_5382 (.A1(n_257_440), .A2(n_257_940), .ZN(n_257_76_5373));
   NAND2_X1 i_257_76_5383 (.A1(n_257_76_5372), .A2(n_257_76_5373), .ZN(
      n_257_76_5374));
   INV_X1 i_257_76_5384 (.A(n_257_76_5374), .ZN(n_257_76_5375));
   NAND3_X1 i_257_76_5385 (.A1(n_257_76_5370), .A2(n_257_76_5371), .A3(
      n_257_76_5375), .ZN(n_257_76_5376));
   NOR2_X1 i_257_76_5386 (.A1(n_257_76_5368), .A2(n_257_76_5376), .ZN(
      n_257_76_5377));
   NAND2_X1 i_257_76_5387 (.A1(n_257_908), .A2(n_257_439), .ZN(n_257_76_5378));
   NAND2_X1 i_257_76_5388 (.A1(n_257_76_5378), .A2(n_257_76_5346), .ZN(
      n_257_76_5379));
   INV_X1 i_257_76_5389 (.A(n_257_76_5379), .ZN(n_257_76_5380));
   NAND2_X1 i_257_76_5390 (.A1(n_257_870), .A2(n_257_445), .ZN(n_257_76_5381));
   NAND3_X1 i_257_76_5391 (.A1(n_257_76_5377), .A2(n_257_76_5380), .A3(
      n_257_76_5381), .ZN(n_257_76_5382));
   NAND2_X1 i_257_76_5392 (.A1(n_257_806), .A2(n_257_437), .ZN(n_257_76_5383));
   NAND2_X1 i_257_76_5393 (.A1(n_257_742), .A2(n_257_436), .ZN(n_257_76_5384));
   NAND2_X1 i_257_76_5394 (.A1(n_257_76_5383), .A2(n_257_76_5384), .ZN(
      n_257_76_5385));
   NOR2_X1 i_257_76_5395 (.A1(n_257_76_5382), .A2(n_257_76_5385), .ZN(
      n_257_76_5386));
   NAND2_X1 i_257_76_5396 (.A1(n_257_76_5345), .A2(n_257_76_5386), .ZN(
      n_257_76_5387));
   INV_X1 i_257_76_5397 (.A(n_257_76_5387), .ZN(n_257_76_5388));
   NAND2_X1 i_257_76_5398 (.A1(n_257_678), .A2(n_257_448), .ZN(n_257_76_5389));
   NAND3_X1 i_257_76_5399 (.A1(n_257_76_5388), .A2(n_257_76_5344), .A3(
      n_257_76_5389), .ZN(n_257_76_5390));
   INV_X1 i_257_76_5400 (.A(n_257_76_5390), .ZN(n_257_76_5391));
   NAND2_X1 i_257_76_5401 (.A1(n_257_28), .A2(n_257_76_5391), .ZN(n_257_76_5392));
   NAND3_X1 i_257_76_5402 (.A1(n_257_76_5358), .A2(n_257_76_5364), .A3(
      n_257_76_5392), .ZN(n_257_76_5393));
   NAND2_X1 i_257_76_5403 (.A1(n_257_446), .A2(n_257_76_5359), .ZN(n_257_76_5394));
   NAND3_X1 i_257_76_5404 (.A1(n_257_76_5372), .A2(n_257_76_5373), .A3(n_257_838), 
      .ZN(n_257_76_5395));
   NOR2_X1 i_257_76_5405 (.A1(n_257_76_5394), .A2(n_257_76_5395), .ZN(
      n_257_76_5396));
   NAND3_X1 i_257_76_5406 (.A1(n_257_76_5396), .A2(n_257_76_5378), .A3(
      n_257_76_5346), .ZN(n_257_76_5397));
   INV_X1 i_257_76_5407 (.A(n_257_76_5381), .ZN(n_257_76_5398));
   NOR2_X1 i_257_76_5408 (.A1(n_257_76_5397), .A2(n_257_76_5398), .ZN(
      n_257_76_5399));
   NAND2_X1 i_257_76_5409 (.A1(n_257_76_5345), .A2(n_257_76_5399), .ZN(
      n_257_76_5400));
   INV_X1 i_257_76_5410 (.A(n_257_76_5400), .ZN(n_257_76_5401));
   NAND2_X1 i_257_76_5411 (.A1(n_257_76_5344), .A2(n_257_76_5401), .ZN(
      n_257_76_5402));
   INV_X1 i_257_76_5412 (.A(n_257_76_5402), .ZN(n_257_76_5403));
   NAND2_X1 i_257_76_5413 (.A1(n_257_76_18070), .A2(n_257_76_5403), .ZN(
      n_257_76_5404));
   NAND3_X1 i_257_76_5414 (.A1(n_257_76_5359), .A2(n_257_76_5373), .A3(n_257_439), 
      .ZN(n_257_76_5405));
   INV_X1 i_257_76_5415 (.A(n_257_76_5405), .ZN(n_257_76_5406));
   NAND3_X1 i_257_76_5416 (.A1(n_257_76_5406), .A2(n_257_76_5346), .A3(n_257_908), 
      .ZN(n_257_76_5407));
   INV_X1 i_257_76_5417 (.A(n_257_76_5407), .ZN(n_257_76_5408));
   NAND2_X1 i_257_76_5418 (.A1(n_257_76_5345), .A2(n_257_76_5408), .ZN(
      n_257_76_5409));
   INV_X1 i_257_76_5419 (.A(n_257_76_5409), .ZN(n_257_76_5410));
   NAND2_X1 i_257_76_5420 (.A1(n_257_76_5344), .A2(n_257_76_5410), .ZN(
      n_257_76_5411));
   INV_X1 i_257_76_5421 (.A(n_257_76_5411), .ZN(n_257_76_5412));
   NAND2_X1 i_257_76_5422 (.A1(n_257_76_18084), .A2(n_257_76_5412), .ZN(
      n_257_76_5413));
   NAND2_X1 i_257_76_5423 (.A1(n_257_201), .A2(n_257_427), .ZN(n_257_76_5414));
   NAND2_X1 i_257_76_5424 (.A1(n_257_638), .A2(n_257_450), .ZN(n_257_76_5415));
   NAND2_X1 i_257_76_5425 (.A1(n_257_510), .A2(n_257_424), .ZN(n_257_76_5416));
   NAND3_X1 i_257_76_5426 (.A1(n_257_76_5414), .A2(n_257_76_5415), .A3(
      n_257_76_5416), .ZN(n_257_76_5417));
   INV_X1 i_257_76_5427 (.A(n_257_574), .ZN(n_257_76_5418));
   NAND2_X1 i_257_76_5428 (.A1(n_257_76_5418), .A2(n_257_442), .ZN(n_257_76_5419));
   OAI21_X1 i_257_76_5429 (.A(n_257_76_5419), .B1(n_257_428), .B2(n_257_76_17412), 
      .ZN(n_257_76_5420));
   INV_X1 i_257_76_5430 (.A(n_257_76_5420), .ZN(n_257_76_5421));
   NOR2_X1 i_257_76_5431 (.A1(n_257_1068), .A2(n_257_76_5421), .ZN(n_257_76_5422));
   NAND2_X1 i_257_76_5432 (.A1(n_257_432), .A2(n_257_606), .ZN(n_257_76_5423));
   NAND2_X1 i_257_76_5433 (.A1(n_257_76_5423), .A2(n_257_423), .ZN(n_257_76_5424));
   INV_X1 i_257_76_5434 (.A(n_257_76_5424), .ZN(n_257_76_5425));
   NAND4_X1 i_257_76_5435 (.A1(n_257_76_5422), .A2(n_257_76_5372), .A3(
      n_257_76_5373), .A4(n_257_76_5425), .ZN(n_257_76_5426));
   NOR2_X1 i_257_76_5436 (.A1(n_257_76_5417), .A2(n_257_76_5426), .ZN(
      n_257_76_5427));
   NAND3_X1 i_257_76_5437 (.A1(n_257_76_5366), .A2(n_257_76_5367), .A3(
      n_257_76_5371), .ZN(n_257_76_5428));
   INV_X1 i_257_76_5438 (.A(n_257_76_5428), .ZN(n_257_76_5429));
   NAND2_X1 i_257_76_5439 (.A1(n_257_44), .A2(n_257_433), .ZN(n_257_76_5430));
   NAND2_X1 i_257_76_5440 (.A1(n_257_76_5430), .A2(n_257_76_5365), .ZN(
      n_257_76_5431));
   INV_X1 i_257_76_5441 (.A(n_257_76_5431), .ZN(n_257_76_5432));
   NAND3_X1 i_257_76_5442 (.A1(n_257_76_5427), .A2(n_257_76_5429), .A3(
      n_257_76_5432), .ZN(n_257_76_5433));
   NAND2_X1 i_257_76_5443 (.A1(n_257_542), .A2(n_257_426), .ZN(n_257_76_5434));
   NAND2_X1 i_257_76_5444 (.A1(n_257_76_5434), .A2(n_257_76_5346), .ZN(
      n_257_76_5435));
   INV_X1 i_257_76_5445 (.A(n_257_76_5435), .ZN(n_257_76_5436));
   NAND2_X1 i_257_76_5446 (.A1(n_257_122), .A2(n_257_430), .ZN(n_257_76_5437));
   NAND3_X1 i_257_76_5447 (.A1(n_257_76_5436), .A2(n_257_76_5437), .A3(
      n_257_76_5378), .ZN(n_257_76_5438));
   NOR2_X1 i_257_76_5448 (.A1(n_257_76_5433), .A2(n_257_76_5438), .ZN(
      n_257_76_5439));
   NAND2_X1 i_257_76_5449 (.A1(n_257_451), .A2(n_257_461), .ZN(n_257_76_5440));
   NAND2_X1 i_257_76_5450 (.A1(n_257_281), .A2(n_257_76_5440), .ZN(n_257_76_5441));
   INV_X1 i_257_76_5451 (.A(n_257_76_5441), .ZN(n_257_76_5442));
   NAND3_X1 i_257_76_5452 (.A1(n_257_76_5442), .A2(n_257_76_5384), .A3(
      n_257_76_5381), .ZN(n_257_76_5443));
   INV_X1 i_257_76_5453 (.A(n_257_76_5443), .ZN(n_257_76_5444));
   NAND2_X1 i_257_76_5454 (.A1(n_257_84), .A2(n_257_431), .ZN(n_257_76_5445));
   NAND2_X1 i_257_76_5455 (.A1(n_257_76_5383), .A2(n_257_76_5445), .ZN(
      n_257_76_5446));
   INV_X1 i_257_76_5456 (.A(n_257_76_5446), .ZN(n_257_76_5447));
   NAND2_X1 i_257_76_5457 (.A1(n_257_161), .A2(n_257_429), .ZN(n_257_76_5448));
   NAND4_X1 i_257_76_5458 (.A1(n_257_76_5439), .A2(n_257_76_5444), .A3(
      n_257_76_5447), .A4(n_257_76_5448), .ZN(n_257_76_5449));
   INV_X1 i_257_76_5459 (.A(n_257_76_5449), .ZN(n_257_76_5450));
   NAND2_X1 i_257_76_5460 (.A1(n_257_76_5344), .A2(n_257_76_5450), .ZN(
      n_257_76_5451));
   NAND2_X1 i_257_76_5461 (.A1(n_257_241), .A2(n_257_425), .ZN(n_257_76_5452));
   NAND3_X1 i_257_76_5462 (.A1(n_257_76_5389), .A2(n_257_76_5452), .A3(
      n_257_76_5345), .ZN(n_257_76_5453));
   NOR2_X1 i_257_76_5463 (.A1(n_257_76_5451), .A2(n_257_76_5453), .ZN(
      n_257_76_5454));
   NAND2_X1 i_257_76_5464 (.A1(n_257_76_18066), .A2(n_257_76_5454), .ZN(
      n_257_76_5455));
   NAND3_X1 i_257_76_5465 (.A1(n_257_76_5404), .A2(n_257_76_5413), .A3(
      n_257_76_5455), .ZN(n_257_76_5456));
   NOR2_X1 i_257_76_5466 (.A1(n_257_76_5393), .A2(n_257_76_5456), .ZN(
      n_257_76_5457));
   NAND2_X1 i_257_76_5467 (.A1(n_257_76_5359), .A2(n_257_972), .ZN(n_257_76_5458));
   NOR2_X1 i_257_76_5468 (.A1(n_257_76_13147), .A2(n_257_76_5458), .ZN(
      n_257_76_5459));
   NAND2_X1 i_257_76_5469 (.A1(n_257_76_5345), .A2(n_257_76_5459), .ZN(
      n_257_76_5460));
   INV_X1 i_257_76_5470 (.A(n_257_76_5460), .ZN(n_257_76_5461));
   NAND2_X1 i_257_76_5471 (.A1(n_257_76_5344), .A2(n_257_76_5461), .ZN(
      n_257_76_5462));
   INV_X1 i_257_76_5472 (.A(n_257_76_5462), .ZN(n_257_76_5463));
   NAND2_X1 i_257_76_5473 (.A1(n_257_76_18071), .A2(n_257_76_5463), .ZN(
      n_257_76_5464));
   NAND2_X1 i_257_76_5474 (.A1(n_257_76_5366), .A2(n_257_76_5371), .ZN(
      n_257_76_5465));
   INV_X1 i_257_76_5475 (.A(n_257_76_5465), .ZN(n_257_76_5466));
   NOR2_X1 i_257_76_5476 (.A1(n_257_1068), .A2(n_257_76_15289), .ZN(
      n_257_76_5467));
   NAND4_X1 i_257_76_5477 (.A1(n_257_710), .A2(n_257_76_5467), .A3(n_257_76_5372), 
      .A4(n_257_76_5373), .ZN(n_257_76_5468));
   INV_X1 i_257_76_5478 (.A(n_257_76_5468), .ZN(n_257_76_5469));
   NAND4_X1 i_257_76_5479 (.A1(n_257_76_5466), .A2(n_257_76_5378), .A3(
      n_257_76_5469), .A4(n_257_76_5346), .ZN(n_257_76_5470));
   INV_X1 i_257_76_5480 (.A(n_257_76_5470), .ZN(n_257_76_5471));
   NAND4_X1 i_257_76_5481 (.A1(n_257_76_5471), .A2(n_257_76_5383), .A3(
      n_257_76_5384), .A4(n_257_76_5381), .ZN(n_257_76_5472));
   INV_X1 i_257_76_5482 (.A(n_257_76_5472), .ZN(n_257_76_5473));
   NAND2_X1 i_257_76_5483 (.A1(n_257_76_5345), .A2(n_257_76_5473), .ZN(
      n_257_76_5474));
   INV_X1 i_257_76_5484 (.A(n_257_76_5474), .ZN(n_257_76_5475));
   NAND2_X1 i_257_76_5485 (.A1(n_257_76_5344), .A2(n_257_76_5475), .ZN(
      n_257_76_5476));
   INV_X1 i_257_76_5486 (.A(n_257_76_5476), .ZN(n_257_76_5477));
   NAND2_X1 i_257_76_5487 (.A1(n_257_76_18078), .A2(n_257_76_5477), .ZN(
      n_257_76_5478));
   NAND3_X1 i_257_76_5488 (.A1(n_257_76_5383), .A2(n_257_76_5445), .A3(
      n_257_76_5384), .ZN(n_257_76_5479));
   INV_X1 i_257_76_5489 (.A(n_257_76_5448), .ZN(n_257_76_5480));
   NOR2_X1 i_257_76_5490 (.A1(n_257_76_5479), .A2(n_257_76_5480), .ZN(
      n_257_76_5481));
   NAND2_X1 i_257_76_5491 (.A1(n_257_442), .A2(n_257_574), .ZN(n_257_76_5482));
   INV_X1 i_257_76_5492 (.A(n_257_76_5482), .ZN(n_257_76_5483));
   NAND2_X1 i_257_76_5493 (.A1(n_257_428), .A2(n_257_76_5483), .ZN(n_257_76_5484));
   INV_X1 i_257_76_5494 (.A(n_257_76_5484), .ZN(n_257_76_5485));
   NAND2_X1 i_257_76_5495 (.A1(n_257_76_5485), .A2(n_257_76_5423), .ZN(
      n_257_76_5486));
   NOR2_X1 i_257_76_5496 (.A1(n_257_76_5486), .A2(n_257_1068), .ZN(n_257_76_5487));
   NAND4_X1 i_257_76_5497 (.A1(n_257_76_5371), .A2(n_257_76_5375), .A3(
      n_257_76_5415), .A4(n_257_76_5487), .ZN(n_257_76_5488));
   INV_X1 i_257_76_5498 (.A(n_257_76_5488), .ZN(n_257_76_5489));
   NAND2_X1 i_257_76_5499 (.A1(n_257_76_5346), .A2(n_257_76_5430), .ZN(
      n_257_76_5490));
   INV_X1 i_257_76_5500 (.A(n_257_76_5490), .ZN(n_257_76_5491));
   INV_X1 i_257_76_5501 (.A(n_257_76_5368), .ZN(n_257_76_5492));
   NAND4_X1 i_257_76_5502 (.A1(n_257_76_5489), .A2(n_257_76_5491), .A3(
      n_257_76_5492), .A4(n_257_76_5378), .ZN(n_257_76_5493));
   NAND3_X1 i_257_76_5503 (.A1(n_257_76_5381), .A2(n_257_76_5440), .A3(
      n_257_76_5437), .ZN(n_257_76_5494));
   NOR2_X1 i_257_76_5504 (.A1(n_257_76_5493), .A2(n_257_76_5494), .ZN(
      n_257_76_5495));
   NAND4_X1 i_257_76_5505 (.A1(n_257_76_5481), .A2(n_257_76_5389), .A3(
      n_257_76_5345), .A4(n_257_76_5495), .ZN(n_257_76_5496));
   INV_X1 i_257_76_5506 (.A(n_257_76_5344), .ZN(n_257_76_5497));
   NOR2_X1 i_257_76_5507 (.A1(n_257_76_5496), .A2(n_257_76_5497), .ZN(
      n_257_76_5498));
   NAND2_X1 i_257_76_5508 (.A1(n_257_76_18074), .A2(n_257_76_5498), .ZN(
      n_257_76_5499));
   NAND3_X1 i_257_76_5509 (.A1(n_257_76_5464), .A2(n_257_76_5478), .A3(
      n_257_76_5499), .ZN(n_257_76_5500));
   NAND2_X1 i_257_76_5510 (.A1(n_257_1068), .A2(n_257_442), .ZN(n_257_76_5501));
   INV_X1 i_257_76_5511 (.A(n_257_76_5501), .ZN(n_257_76_5502));
   NAND2_X1 i_257_76_5512 (.A1(n_257_13), .A2(n_257_76_5502), .ZN(n_257_76_5503));
   INV_X1 i_257_76_5513 (.A(n_257_76_5346), .ZN(n_257_76_5504));
   NOR2_X1 i_257_76_5514 (.A1(n_257_76_17902), .A2(n_257_1068), .ZN(
      n_257_76_5505));
   NAND3_X1 i_257_76_5515 (.A1(n_257_76_5505), .A2(n_257_76_5372), .A3(
      n_257_76_5373), .ZN(n_257_76_5506));
   NOR2_X1 i_257_76_5516 (.A1(n_257_76_5504), .A2(n_257_76_5506), .ZN(
      n_257_76_5507));
   NAND3_X1 i_257_76_5517 (.A1(n_257_76_5507), .A2(n_257_870), .A3(n_257_76_5378), 
      .ZN(n_257_76_5508));
   INV_X1 i_257_76_5518 (.A(n_257_76_5508), .ZN(n_257_76_5509));
   NAND2_X1 i_257_76_5519 (.A1(n_257_76_5345), .A2(n_257_76_5509), .ZN(
      n_257_76_5510));
   INV_X1 i_257_76_5520 (.A(n_257_76_5510), .ZN(n_257_76_5511));
   NAND2_X1 i_257_76_5521 (.A1(n_257_76_5344), .A2(n_257_76_5511), .ZN(
      n_257_76_5512));
   INV_X1 i_257_76_5522 (.A(n_257_76_5512), .ZN(n_257_76_5513));
   NAND2_X1 i_257_76_5523 (.A1(n_257_76_18077), .A2(n_257_76_5513), .ZN(
      n_257_76_5514));
   NAND2_X1 i_257_76_5524 (.A1(n_257_76_5503), .A2(n_257_76_5514), .ZN(
      n_257_76_5515));
   NOR2_X1 i_257_76_5525 (.A1(n_257_76_5500), .A2(n_257_76_5515), .ZN(
      n_257_76_5516));
   NAND2_X1 i_257_76_5526 (.A1(n_257_76_5437), .A2(n_257_76_5378), .ZN(
      n_257_76_5517));
   INV_X1 i_257_76_5527 (.A(n_257_76_5517), .ZN(n_257_76_5518));
   NAND4_X1 i_257_76_5528 (.A1(n_257_76_5346), .A2(n_257_76_5366), .A3(
      n_257_76_5367), .A4(n_257_76_5371), .ZN(n_257_76_5519));
   INV_X1 i_257_76_5529 (.A(n_257_76_5519), .ZN(n_257_76_5520));
   NAND4_X1 i_257_76_5530 (.A1(n_257_76_5518), .A2(n_257_76_5520), .A3(
      n_257_76_5381), .A4(n_257_76_5440), .ZN(n_257_76_5521));
   NAND2_X1 i_257_76_5531 (.A1(n_257_76_5445), .A2(n_257_76_5384), .ZN(
      n_257_76_5522));
   NOR2_X1 i_257_76_5532 (.A1(n_257_76_5521), .A2(n_257_76_5522), .ZN(
      n_257_76_5523));
   NAND3_X1 i_257_76_5533 (.A1(n_257_542), .A2(n_257_76_5414), .A3(n_257_76_5415), 
      .ZN(n_257_76_5524));
   INV_X1 i_257_76_5534 (.A(n_257_76_5524), .ZN(n_257_76_5525));
   NAND2_X1 i_257_76_5535 (.A1(n_257_76_5423), .A2(n_257_426), .ZN(n_257_76_5526));
   INV_X1 i_257_76_5536 (.A(n_257_76_5526), .ZN(n_257_76_5527));
   NAND3_X1 i_257_76_5537 (.A1(n_257_76_5527), .A2(n_257_76_5347), .A3(
      n_257_76_5420), .ZN(n_257_76_5528));
   NOR2_X1 i_257_76_5538 (.A1(n_257_76_5374), .A2(n_257_76_5528), .ZN(
      n_257_76_5529));
   NAND4_X1 i_257_76_5539 (.A1(n_257_76_5525), .A2(n_257_76_5529), .A3(
      n_257_76_5430), .A4(n_257_76_5365), .ZN(n_257_76_5530));
   INV_X1 i_257_76_5540 (.A(n_257_76_5530), .ZN(n_257_76_5531));
   NAND3_X1 i_257_76_5541 (.A1(n_257_76_5448), .A2(n_257_76_5531), .A3(
      n_257_76_5383), .ZN(n_257_76_5532));
   INV_X1 i_257_76_5542 (.A(n_257_76_5532), .ZN(n_257_76_5533));
   NAND4_X1 i_257_76_5543 (.A1(n_257_76_5389), .A2(n_257_76_5523), .A3(
      n_257_76_5345), .A4(n_257_76_5533), .ZN(n_257_76_5534));
   NOR2_X1 i_257_76_5544 (.A1(n_257_76_5534), .A2(n_257_76_5497), .ZN(
      n_257_76_5535));
   NAND2_X1 i_257_76_5545 (.A1(n_257_76_18076), .A2(n_257_76_5535), .ZN(
      n_257_76_5536));
   NOR2_X1 i_257_76_5546 (.A1(n_257_1068), .A2(n_257_76_17934), .ZN(
      n_257_76_5537));
   NAND3_X1 i_257_76_5547 (.A1(n_257_76_5537), .A2(n_257_76_5372), .A3(
      n_257_76_5373), .ZN(n_257_76_5538));
   INV_X1 i_257_76_5548 (.A(n_257_76_5538), .ZN(n_257_76_5539));
   NAND4_X1 i_257_76_5549 (.A1(n_257_76_5346), .A2(n_257_76_5539), .A3(
      n_257_76_5366), .A4(n_257_76_5371), .ZN(n_257_76_5540));
   INV_X1 i_257_76_5550 (.A(n_257_76_5378), .ZN(n_257_76_5541));
   NOR2_X1 i_257_76_5551 (.A1(n_257_76_5540), .A2(n_257_76_5541), .ZN(
      n_257_76_5542));
   NAND2_X1 i_257_76_5552 (.A1(n_257_76_5381), .A2(n_257_742), .ZN(n_257_76_5543));
   INV_X1 i_257_76_5553 (.A(n_257_76_5543), .ZN(n_257_76_5544));
   NAND3_X1 i_257_76_5554 (.A1(n_257_76_5542), .A2(n_257_76_5544), .A3(
      n_257_76_5383), .ZN(n_257_76_5545));
   INV_X1 i_257_76_5555 (.A(n_257_76_5545), .ZN(n_257_76_5546));
   NAND2_X1 i_257_76_5556 (.A1(n_257_76_5345), .A2(n_257_76_5546), .ZN(
      n_257_76_5547));
   INV_X1 i_257_76_5557 (.A(n_257_76_5547), .ZN(n_257_76_5548));
   NAND2_X1 i_257_76_5558 (.A1(n_257_76_5344), .A2(n_257_76_5548), .ZN(
      n_257_76_5549));
   INV_X1 i_257_76_5559 (.A(n_257_76_5549), .ZN(n_257_76_5550));
   NAND2_X1 i_257_76_5560 (.A1(n_257_76_18069), .A2(n_257_76_5550), .ZN(
      n_257_76_5551));
   NAND2_X1 i_257_76_5561 (.A1(n_257_606), .A2(n_257_442), .ZN(n_257_76_5552));
   INV_X1 i_257_76_5562 (.A(n_257_76_5552), .ZN(n_257_76_5553));
   NAND2_X1 i_257_76_5563 (.A1(n_257_432), .A2(n_257_76_5553), .ZN(n_257_76_5554));
   NOR2_X1 i_257_76_5564 (.A1(n_257_1068), .A2(n_257_76_5554), .ZN(n_257_76_5555));
   NAND3_X1 i_257_76_5565 (.A1(n_257_76_5555), .A2(n_257_76_5372), .A3(
      n_257_76_5373), .ZN(n_257_76_5556));
   INV_X1 i_257_76_5566 (.A(n_257_76_5556), .ZN(n_257_76_5557));
   NAND4_X1 i_257_76_5567 (.A1(n_257_76_5557), .A2(n_257_76_5367), .A3(
      n_257_76_5371), .A4(n_257_76_5415), .ZN(n_257_76_5558));
   NAND3_X1 i_257_76_5568 (.A1(n_257_76_5430), .A2(n_257_76_5365), .A3(
      n_257_76_5366), .ZN(n_257_76_5559));
   NOR2_X1 i_257_76_5569 (.A1(n_257_76_5558), .A2(n_257_76_5559), .ZN(
      n_257_76_5560));
   NAND4_X1 i_257_76_5570 (.A1(n_257_76_5560), .A2(n_257_76_5380), .A3(
      n_257_76_5381), .A4(n_257_76_5440), .ZN(n_257_76_5561));
   NOR2_X1 i_257_76_5571 (.A1(n_257_76_5561), .A2(n_257_76_5385), .ZN(
      n_257_76_5562));
   NAND3_X1 i_257_76_5572 (.A1(n_257_76_5562), .A2(n_257_76_5389), .A3(
      n_257_76_5345), .ZN(n_257_76_5563));
   NOR2_X1 i_257_76_5573 (.A1(n_257_76_5563), .A2(n_257_76_5497), .ZN(
      n_257_76_5564));
   NAND2_X1 i_257_76_5574 (.A1(n_257_68), .A2(n_257_76_5564), .ZN(n_257_76_5565));
   NAND3_X1 i_257_76_5575 (.A1(n_257_76_5536), .A2(n_257_76_5551), .A3(
      n_257_76_5565), .ZN(n_257_76_5566));
   NOR2_X1 i_257_76_5576 (.A1(n_257_1068), .A2(n_257_76_17951), .ZN(
      n_257_76_5567));
   NAND3_X1 i_257_76_5577 (.A1(n_257_76_5567), .A2(n_257_76_5372), .A3(
      n_257_76_5373), .ZN(n_257_76_5568));
   INV_X1 i_257_76_5578 (.A(n_257_76_5568), .ZN(n_257_76_5569));
   NAND3_X1 i_257_76_5579 (.A1(n_257_76_5569), .A2(n_257_76_5346), .A3(
      n_257_76_5366), .ZN(n_257_76_5570));
   INV_X1 i_257_76_5580 (.A(n_257_76_5570), .ZN(n_257_76_5571));
   NAND4_X1 i_257_76_5581 (.A1(n_257_806), .A2(n_257_76_5381), .A3(n_257_76_5571), 
      .A4(n_257_76_5378), .ZN(n_257_76_5572));
   INV_X1 i_257_76_5582 (.A(n_257_76_5572), .ZN(n_257_76_5573));
   NAND2_X1 i_257_76_5583 (.A1(n_257_76_5345), .A2(n_257_76_5573), .ZN(
      n_257_76_5574));
   INV_X1 i_257_76_5584 (.A(n_257_76_5574), .ZN(n_257_76_5575));
   NAND2_X1 i_257_76_5585 (.A1(n_257_76_5344), .A2(n_257_76_5575), .ZN(
      n_257_76_5576));
   INV_X1 i_257_76_5586 (.A(n_257_76_5576), .ZN(n_257_76_5577));
   NAND2_X1 i_257_76_5587 (.A1(n_257_22), .A2(n_257_76_5577), .ZN(n_257_76_5578));
   NAND2_X1 i_257_76_5588 (.A1(n_257_444), .A2(n_257_76_5359), .ZN(n_257_76_5579));
   INV_X1 i_257_76_5589 (.A(n_257_76_5579), .ZN(n_257_76_5580));
   NAND2_X1 i_257_76_5590 (.A1(n_257_1004), .A2(n_257_76_5580), .ZN(
      n_257_76_5581));
   INV_X1 i_257_76_5591 (.A(n_257_76_5581), .ZN(n_257_76_5582));
   NAND2_X1 i_257_76_5592 (.A1(n_257_76_5344), .A2(n_257_76_5582), .ZN(
      n_257_76_5583));
   INV_X1 i_257_76_5593 (.A(n_257_76_5583), .ZN(n_257_76_5584));
   NAND2_X1 i_257_76_5594 (.A1(n_257_76_18075), .A2(n_257_76_5584), .ZN(
      n_257_76_5585));
   NAND2_X1 i_257_76_5595 (.A1(n_257_76_5578), .A2(n_257_76_5585), .ZN(
      n_257_76_5586));
   NOR2_X1 i_257_76_5596 (.A1(n_257_76_5566), .A2(n_257_76_5586), .ZN(
      n_257_76_5587));
   NAND3_X1 i_257_76_5597 (.A1(n_257_76_5457), .A2(n_257_76_5516), .A3(
      n_257_76_5587), .ZN(n_257_76_5588));
   INV_X1 i_257_76_5598 (.A(n_257_76_5588), .ZN(n_257_76_5589));
   NOR2_X1 i_257_76_5599 (.A1(n_257_1068), .A2(n_257_76_17633), .ZN(
      n_257_76_5590));
   NAND3_X1 i_257_76_5600 (.A1(n_257_76_5590), .A2(n_257_76_5372), .A3(
      n_257_76_5373), .ZN(n_257_76_5591));
   INV_X1 i_257_76_5601 (.A(n_257_76_5591), .ZN(n_257_76_5592));
   NAND4_X1 i_257_76_5602 (.A1(n_257_76_5592), .A2(n_257_76_5371), .A3(n_257_44), 
      .A4(n_257_76_5415), .ZN(n_257_76_5593));
   NAND4_X1 i_257_76_5603 (.A1(n_257_76_5346), .A2(n_257_76_5365), .A3(
      n_257_76_5366), .A4(n_257_76_5367), .ZN(n_257_76_5594));
   NOR2_X1 i_257_76_5604 (.A1(n_257_76_5593), .A2(n_257_76_5594), .ZN(
      n_257_76_5595));
   NAND2_X1 i_257_76_5605 (.A1(n_257_76_5440), .A2(n_257_76_5378), .ZN(
      n_257_76_5596));
   INV_X1 i_257_76_5606 (.A(n_257_76_5596), .ZN(n_257_76_5597));
   NAND3_X1 i_257_76_5607 (.A1(n_257_76_5595), .A2(n_257_76_5597), .A3(
      n_257_76_5381), .ZN(n_257_76_5598));
   NOR2_X1 i_257_76_5608 (.A1(n_257_76_5598), .A2(n_257_76_5385), .ZN(
      n_257_76_5599));
   NAND2_X1 i_257_76_5609 (.A1(n_257_76_5345), .A2(n_257_76_5599), .ZN(
      n_257_76_5600));
   INV_X1 i_257_76_5610 (.A(n_257_76_5600), .ZN(n_257_76_5601));
   NAND3_X1 i_257_76_5611 (.A1(n_257_76_5601), .A2(n_257_76_5344), .A3(
      n_257_76_5389), .ZN(n_257_76_5602));
   INV_X1 i_257_76_5612 (.A(n_257_76_5602), .ZN(n_257_76_5603));
   NAND2_X1 i_257_76_5613 (.A1(n_257_76_18081), .A2(n_257_76_5603), .ZN(
      n_257_76_5604));
   NAND2_X1 i_257_76_5614 (.A1(n_257_76_5373), .A2(n_257_76_5347), .ZN(
      n_257_76_5605));
   INV_X1 i_257_76_5615 (.A(n_257_76_5605), .ZN(n_257_76_5606));
   NAND3_X1 i_257_76_5616 (.A1(n_257_76_5365), .A2(n_257_76_18047), .A3(
      n_257_76_5606), .ZN(n_257_76_5607));
   NOR2_X1 i_257_76_5617 (.A1(n_257_76_5541), .A2(n_257_76_5607), .ZN(
      n_257_76_5608));
   INV_X1 i_257_76_5618 (.A(n_257_76_5367), .ZN(n_257_76_5609));
   NAND4_X1 i_257_76_5619 (.A1(n_257_76_5346), .A2(n_257_76_5609), .A3(
      n_257_76_5366), .A4(n_257_76_5371), .ZN(n_257_76_5610));
   INV_X1 i_257_76_5620 (.A(n_257_76_5610), .ZN(n_257_76_5611));
   NAND3_X1 i_257_76_5621 (.A1(n_257_76_5608), .A2(n_257_76_5381), .A3(
      n_257_76_5611), .ZN(n_257_76_5612));
   NOR2_X1 i_257_76_5622 (.A1(n_257_76_5612), .A2(n_257_76_5385), .ZN(
      n_257_76_5613));
   NAND2_X1 i_257_76_5623 (.A1(n_257_76_5345), .A2(n_257_76_5613), .ZN(
      n_257_76_5614));
   INV_X1 i_257_76_5624 (.A(n_257_76_5614), .ZN(n_257_76_5615));
   NAND3_X1 i_257_76_5625 (.A1(n_257_76_5615), .A2(n_257_76_5344), .A3(
      n_257_76_5389), .ZN(n_257_76_5616));
   INV_X1 i_257_76_5626 (.A(n_257_76_5616), .ZN(n_257_76_5617));
   NAND2_X1 i_257_76_5627 (.A1(n_257_76_18083), .A2(n_257_76_5617), .ZN(
      n_257_76_5618));
   NAND2_X1 i_257_76_5628 (.A1(n_257_76_5440), .A2(n_257_76_5437), .ZN(
      n_257_76_5619));
   INV_X1 i_257_76_5629 (.A(n_257_76_5619), .ZN(n_257_76_5620));
   INV_X1 i_257_76_5630 (.A(n_257_606), .ZN(n_257_76_5621));
   NAND2_X1 i_257_76_5631 (.A1(n_257_76_5621), .A2(n_257_442), .ZN(n_257_76_5622));
   OAI21_X1 i_257_76_5632 (.A(n_257_76_5622), .B1(n_257_432), .B2(n_257_76_17412), 
      .ZN(n_257_76_5623));
   NAND3_X1 i_257_76_5633 (.A1(n_257_76_5347), .A2(n_257_76_5623), .A3(n_257_429), 
      .ZN(n_257_76_5624));
   INV_X1 i_257_76_5634 (.A(n_257_76_5624), .ZN(n_257_76_5625));
   NAND4_X1 i_257_76_5635 (.A1(n_257_76_5371), .A2(n_257_76_5375), .A3(
      n_257_76_5415), .A4(n_257_76_5625), .ZN(n_257_76_5626));
   NOR2_X1 i_257_76_5636 (.A1(n_257_76_5626), .A2(n_257_76_5368), .ZN(
      n_257_76_5627));
   NOR2_X1 i_257_76_5637 (.A1(n_257_76_5541), .A2(n_257_76_5490), .ZN(
      n_257_76_5628));
   NAND4_X1 i_257_76_5638 (.A1(n_257_76_5620), .A2(n_257_76_5627), .A3(
      n_257_76_5628), .A4(n_257_76_5381), .ZN(n_257_76_5629));
   NAND4_X1 i_257_76_5639 (.A1(n_257_76_5383), .A2(n_257_76_5445), .A3(n_257_161), 
      .A4(n_257_76_5384), .ZN(n_257_76_5630));
   NOR2_X1 i_257_76_5640 (.A1(n_257_76_5629), .A2(n_257_76_5630), .ZN(
      n_257_76_5631));
   NAND3_X1 i_257_76_5641 (.A1(n_257_76_5631), .A2(n_257_76_5389), .A3(
      n_257_76_5345), .ZN(n_257_76_5632));
   NOR2_X1 i_257_76_5642 (.A1(n_257_76_5632), .A2(n_257_76_5497), .ZN(
      n_257_76_5633));
   NAND2_X1 i_257_76_5643 (.A1(n_257_76_18061), .A2(n_257_76_5633), .ZN(
      n_257_76_5634));
   NAND3_X1 i_257_76_5644 (.A1(n_257_76_5604), .A2(n_257_76_5618), .A3(
      n_257_76_5634), .ZN(n_257_76_5635));
   INV_X1 i_257_76_5645 (.A(n_257_76_5635), .ZN(n_257_76_5636));
   INV_X1 i_257_76_5646 (.A(n_257_76_5372), .ZN(n_257_76_5637));
   NAND3_X1 i_257_76_5647 (.A1(n_257_76_5359), .A2(n_257_76_5637), .A3(
      n_257_76_5373), .ZN(n_257_76_5638));
   INV_X1 i_257_76_5648 (.A(n_257_76_5638), .ZN(n_257_76_5639));
   NAND2_X1 i_257_76_5649 (.A1(n_257_76_5639), .A2(n_257_76_5346), .ZN(
      n_257_76_5640));
   NOR2_X1 i_257_76_5650 (.A1(n_257_76_5541), .A2(n_257_76_5640), .ZN(
      n_257_76_5641));
   NAND2_X1 i_257_76_5651 (.A1(n_257_76_5345), .A2(n_257_76_5641), .ZN(
      n_257_76_5642));
   INV_X1 i_257_76_5652 (.A(n_257_76_5642), .ZN(n_257_76_5643));
   NAND2_X1 i_257_76_5653 (.A1(n_257_76_5344), .A2(n_257_76_5643), .ZN(
      n_257_76_5644));
   INV_X1 i_257_76_5654 (.A(n_257_76_5644), .ZN(n_257_76_5645));
   NAND2_X1 i_257_76_5655 (.A1(n_257_76_18067), .A2(n_257_76_5645), .ZN(
      n_257_76_5646));
   NAND3_X1 i_257_76_5656 (.A1(n_257_76_5346), .A2(n_257_76_5430), .A3(
      n_257_76_5365), .ZN(n_257_76_5647));
   NOR2_X1 i_257_76_5657 (.A1(n_257_76_14354), .A2(n_257_574), .ZN(n_257_76_5648));
   AOI21_X1 i_257_76_5658 (.A(n_257_76_5648), .B1(n_257_76_16810), .B2(
      n_257_76_14600), .ZN(n_257_76_5649));
   NOR2_X1 i_257_76_5659 (.A1(n_257_1068), .A2(n_257_76_5649), .ZN(n_257_76_5650));
   NAND2_X1 i_257_76_5660 (.A1(n_257_420), .A2(n_257_76_5423), .ZN(n_257_76_5651));
   INV_X1 i_257_76_5661 (.A(n_257_76_5651), .ZN(n_257_76_5652));
   NAND3_X1 i_257_76_5662 (.A1(n_257_76_5650), .A2(n_257_76_5416), .A3(
      n_257_76_5652), .ZN(n_257_76_5653));
   INV_X1 i_257_76_5663 (.A(n_257_76_5653), .ZN(n_257_76_5654));
   NAND2_X1 i_257_76_5664 (.A1(n_257_76_5434), .A2(n_257_76_5654), .ZN(
      n_257_76_5655));
   NOR2_X1 i_257_76_5665 (.A1(n_257_76_5647), .A2(n_257_76_5655), .ZN(
      n_257_76_5656));
   NAND2_X1 i_257_76_5666 (.A1(n_257_319), .A2(n_257_422), .ZN(n_257_76_5657));
   NAND4_X1 i_257_76_5667 (.A1(n_257_76_5375), .A2(n_257_76_5657), .A3(
      n_257_76_5414), .A4(n_257_76_5415), .ZN(n_257_76_5658));
   NOR2_X1 i_257_76_5668 (.A1(n_257_76_5658), .A2(n_257_76_5428), .ZN(
      n_257_76_5659));
   NAND3_X1 i_257_76_5669 (.A1(n_257_76_5656), .A2(n_257_76_5518), .A3(
      n_257_76_5659), .ZN(n_257_76_5660));
   NAND2_X1 i_257_76_5670 (.A1(n_257_281), .A2(n_257_423), .ZN(n_257_76_5661));
   NAND2_X1 i_257_76_5671 (.A1(n_257_358), .A2(n_257_421), .ZN(n_257_76_5662));
   NAND4_X1 i_257_76_5672 (.A1(n_257_76_5661), .A2(n_257_76_5381), .A3(
      n_257_76_5662), .A4(n_257_76_5440), .ZN(n_257_76_5663));
   NOR2_X1 i_257_76_5673 (.A1(n_257_76_5660), .A2(n_257_76_5663), .ZN(
      n_257_76_5664));
   NAND3_X1 i_257_76_5674 (.A1(n_257_76_5664), .A2(n_257_76_5345), .A3(
      n_257_76_5481), .ZN(n_257_76_5665));
   INV_X1 i_257_76_5675 (.A(n_257_76_5665), .ZN(n_257_76_5666));
   NAND2_X1 i_257_76_5676 (.A1(n_257_76_5389), .A2(n_257_76_5452), .ZN(
      n_257_76_5667));
   INV_X1 i_257_76_5677 (.A(n_257_76_5667), .ZN(n_257_76_5668));
   NAND3_X1 i_257_76_5678 (.A1(n_257_76_5666), .A2(n_257_76_5668), .A3(
      n_257_76_5344), .ZN(n_257_76_5669));
   INV_X1 i_257_76_5679 (.A(n_257_76_5669), .ZN(n_257_76_5670));
   NAND2_X1 i_257_76_5680 (.A1(n_257_76_18073), .A2(n_257_76_5670), .ZN(
      n_257_76_5671));
   NAND3_X1 i_257_76_5681 (.A1(n_257_76_5347), .A2(n_257_76_5623), .A3(n_257_430), 
      .ZN(n_257_76_5672));
   INV_X1 i_257_76_5682 (.A(n_257_76_5672), .ZN(n_257_76_5673));
   NAND4_X1 i_257_76_5683 (.A1(n_257_76_5673), .A2(n_257_76_5415), .A3(
      n_257_76_5372), .A4(n_257_76_5373), .ZN(n_257_76_5674));
   NOR2_X1 i_257_76_5684 (.A1(n_257_76_5428), .A2(n_257_76_5674), .ZN(
      n_257_76_5675));
   NAND4_X1 i_257_76_5685 (.A1(n_257_122), .A2(n_257_76_5346), .A3(n_257_76_5430), 
      .A4(n_257_76_5365), .ZN(n_257_76_5676));
   INV_X1 i_257_76_5686 (.A(n_257_76_5676), .ZN(n_257_76_5677));
   NAND4_X1 i_257_76_5687 (.A1(n_257_76_5597), .A2(n_257_76_5675), .A3(
      n_257_76_5381), .A4(n_257_76_5677), .ZN(n_257_76_5678));
   NOR2_X1 i_257_76_5688 (.A1(n_257_76_5678), .A2(n_257_76_5479), .ZN(
      n_257_76_5679));
   NAND3_X1 i_257_76_5689 (.A1(n_257_76_5679), .A2(n_257_76_5389), .A3(
      n_257_76_5345), .ZN(n_257_76_5680));
   NOR2_X1 i_257_76_5690 (.A1(n_257_76_5680), .A2(n_257_76_5497), .ZN(
      n_257_76_5681));
   NAND2_X1 i_257_76_5691 (.A1(n_257_76_18068), .A2(n_257_76_5681), .ZN(
      n_257_76_5682));
   NAND3_X1 i_257_76_5692 (.A1(n_257_76_5646), .A2(n_257_76_5671), .A3(
      n_257_76_5682), .ZN(n_257_76_5683));
   INV_X1 i_257_76_5693 (.A(n_257_76_5683), .ZN(n_257_76_5684));
   NAND2_X1 i_257_76_5694 (.A1(n_257_774), .A2(n_257_442), .ZN(n_257_76_5685));
   NOR2_X1 i_257_76_5695 (.A1(n_257_1068), .A2(n_257_76_5685), .ZN(n_257_76_5686));
   NAND4_X1 i_257_76_5696 (.A1(n_257_447), .A2(n_257_76_5686), .A3(n_257_76_5372), 
      .A4(n_257_76_5373), .ZN(n_257_76_5687));
   INV_X1 i_257_76_5697 (.A(n_257_76_5687), .ZN(n_257_76_5688));
   NAND4_X1 i_257_76_5698 (.A1(n_257_76_5378), .A2(n_257_76_5688), .A3(
      n_257_76_5346), .A4(n_257_76_5366), .ZN(n_257_76_5689));
   INV_X1 i_257_76_5699 (.A(n_257_76_5689), .ZN(n_257_76_5690));
   NAND3_X1 i_257_76_5700 (.A1(n_257_76_5690), .A2(n_257_76_5383), .A3(
      n_257_76_5381), .ZN(n_257_76_5691));
   INV_X1 i_257_76_5701 (.A(n_257_76_5691), .ZN(n_257_76_5692));
   NAND2_X1 i_257_76_5702 (.A1(n_257_76_5345), .A2(n_257_76_5692), .ZN(
      n_257_76_5693));
   INV_X1 i_257_76_5703 (.A(n_257_76_5693), .ZN(n_257_76_5694));
   NAND2_X1 i_257_76_5704 (.A1(n_257_76_5344), .A2(n_257_76_5694), .ZN(
      n_257_76_5695));
   INV_X1 i_257_76_5705 (.A(n_257_76_5695), .ZN(n_257_76_5696));
   NOR2_X1 i_257_76_5706 (.A1(n_257_76_5490), .A2(n_257_76_5368), .ZN(
      n_257_76_5697));
   NAND3_X1 i_257_76_5707 (.A1(n_257_76_5347), .A2(n_257_76_5623), .A3(n_257_431), 
      .ZN(n_257_76_5698));
   INV_X1 i_257_76_5708 (.A(n_257_76_5698), .ZN(n_257_76_5699));
   NAND4_X1 i_257_76_5709 (.A1(n_257_76_5371), .A2(n_257_76_5375), .A3(
      n_257_76_5415), .A4(n_257_76_5699), .ZN(n_257_76_5700));
   INV_X1 i_257_76_5710 (.A(n_257_76_5700), .ZN(n_257_76_5701));
   NAND4_X1 i_257_76_5711 (.A1(n_257_76_5697), .A2(n_257_76_5597), .A3(n_257_84), 
      .A4(n_257_76_5701), .ZN(n_257_76_5702));
   NAND3_X1 i_257_76_5712 (.A1(n_257_76_5383), .A2(n_257_76_5384), .A3(
      n_257_76_5381), .ZN(n_257_76_5703));
   NOR2_X1 i_257_76_5713 (.A1(n_257_76_5702), .A2(n_257_76_5703), .ZN(
      n_257_76_5704));
   NAND3_X1 i_257_76_5714 (.A1(n_257_76_5704), .A2(n_257_76_5389), .A3(
      n_257_76_5345), .ZN(n_257_76_5705));
   NOR2_X1 i_257_76_5715 (.A1(n_257_76_5705), .A2(n_257_76_5497), .ZN(
      n_257_76_5706));
   AOI22_X1 i_257_76_5716 (.A1(n_257_76_18085), .A2(n_257_76_5696), .B1(
      n_257_76_18080), .B2(n_257_76_5706), .ZN(n_257_76_5707));
   NAND3_X1 i_257_76_5717 (.A1(n_257_76_5636), .A2(n_257_76_5684), .A3(
      n_257_76_5707), .ZN(n_257_76_5708));
   NAND2_X1 i_257_76_5718 (.A1(n_257_76_5448), .A2(n_257_76_5383), .ZN(
      n_257_76_5709));
   NAND4_X1 i_257_76_5719 (.A1(n_257_76_5445), .A2(n_257_76_5384), .A3(
      n_257_76_5661), .A4(n_257_76_5440), .ZN(n_257_76_5710));
   NOR2_X1 i_257_76_5720 (.A1(n_257_76_5709), .A2(n_257_76_5710), .ZN(
      n_257_76_5711));
   NAND3_X1 i_257_76_5721 (.A1(n_257_76_5437), .A2(n_257_76_5378), .A3(n_257_358), 
      .ZN(n_257_76_5712));
   INV_X1 i_257_76_5722 (.A(n_257_76_5712), .ZN(n_257_76_5713));
   NAND4_X1 i_257_76_5723 (.A1(n_257_76_5367), .A2(n_257_76_5371), .A3(
      n_257_76_5657), .A4(n_257_76_5414), .ZN(n_257_76_5714));
   NAND2_X1 i_257_76_5724 (.A1(n_257_76_5423), .A2(n_257_421), .ZN(n_257_76_5715));
   INV_X1 i_257_76_5725 (.A(n_257_76_5715), .ZN(n_257_76_5716));
   NAND3_X1 i_257_76_5726 (.A1(n_257_76_5716), .A2(n_257_76_5347), .A3(
      n_257_76_5420), .ZN(n_257_76_5717));
   INV_X1 i_257_76_5727 (.A(n_257_76_5717), .ZN(n_257_76_5718));
   NAND4_X1 i_257_76_5728 (.A1(n_257_76_5375), .A2(n_257_76_5718), .A3(
      n_257_76_5415), .A4(n_257_76_5416), .ZN(n_257_76_5719));
   NOR2_X1 i_257_76_5729 (.A1(n_257_76_5714), .A2(n_257_76_5719), .ZN(
      n_257_76_5720));
   NOR2_X1 i_257_76_5730 (.A1(n_257_76_5559), .A2(n_257_76_5435), .ZN(
      n_257_76_5721));
   NAND4_X1 i_257_76_5731 (.A1(n_257_76_5713), .A2(n_257_76_5720), .A3(
      n_257_76_5721), .A4(n_257_76_5381), .ZN(n_257_76_5722));
   INV_X1 i_257_76_5732 (.A(n_257_76_5722), .ZN(n_257_76_5723));
   NAND4_X1 i_257_76_5733 (.A1(n_257_76_5711), .A2(n_257_76_5452), .A3(
      n_257_76_5723), .A4(n_257_76_5345), .ZN(n_257_76_5724));
   NAND2_X1 i_257_76_5734 (.A1(n_257_76_5344), .A2(n_257_76_5389), .ZN(
      n_257_76_5725));
   NOR2_X1 i_257_76_5735 (.A1(n_257_76_5724), .A2(n_257_76_5725), .ZN(
      n_257_76_5726));
   NAND2_X1 i_257_76_5736 (.A1(n_257_76_18082), .A2(n_257_76_5726), .ZN(
      n_257_76_5727));
   NAND2_X1 i_257_76_5737 (.A1(n_257_201), .A2(n_257_76_5373), .ZN(n_257_76_5728));
   NAND4_X1 i_257_76_5738 (.A1(n_257_76_5347), .A2(n_257_76_5420), .A3(n_257_427), 
      .A4(n_257_76_5423), .ZN(n_257_76_5729));
   NOR2_X1 i_257_76_5739 (.A1(n_257_76_5728), .A2(n_257_76_5729), .ZN(
      n_257_76_5730));
   NAND2_X1 i_257_76_5740 (.A1(n_257_76_5415), .A2(n_257_76_5372), .ZN(
      n_257_76_5731));
   INV_X1 i_257_76_5741 (.A(n_257_76_5731), .ZN(n_257_76_5732));
   NAND4_X1 i_257_76_5742 (.A1(n_257_76_5730), .A2(n_257_76_5732), .A3(
      n_257_76_5430), .A4(n_257_76_5365), .ZN(n_257_76_5733));
   INV_X1 i_257_76_5743 (.A(n_257_76_5733), .ZN(n_257_76_5734));
   NAND3_X1 i_257_76_5744 (.A1(n_257_76_5383), .A2(n_257_76_5445), .A3(
      n_257_76_5734), .ZN(n_257_76_5735));
   NOR2_X1 i_257_76_5745 (.A1(n_257_76_5735), .A2(n_257_76_5480), .ZN(
      n_257_76_5736));
   NOR2_X1 i_257_76_5746 (.A1(n_257_76_5519), .A2(n_257_76_5541), .ZN(
      n_257_76_5737));
   NAND4_X1 i_257_76_5747 (.A1(n_257_76_5737), .A2(n_257_76_5620), .A3(
      n_257_76_5384), .A4(n_257_76_5381), .ZN(n_257_76_5738));
   INV_X1 i_257_76_5748 (.A(n_257_76_5738), .ZN(n_257_76_5739));
   NAND4_X1 i_257_76_5749 (.A1(n_257_76_5736), .A2(n_257_76_5389), .A3(
      n_257_76_5345), .A4(n_257_76_5739), .ZN(n_257_76_5740));
   NOR2_X1 i_257_76_5750 (.A1(n_257_76_5740), .A2(n_257_76_5497), .ZN(
      n_257_76_5741));
   NAND2_X1 i_257_76_5751 (.A1(n_257_76_18065), .A2(n_257_76_5741), .ZN(
      n_257_76_5742));
   INV_X1 i_257_76_5752 (.A(n_257_76_5385), .ZN(n_257_76_5743));
   NAND2_X1 i_257_76_5753 (.A1(n_257_76_5372), .A2(n_257_76_5359), .ZN(
      n_257_76_5744));
   INV_X1 i_257_76_5754 (.A(n_257_76_5744), .ZN(n_257_76_5745));
   NAND2_X1 i_257_76_5755 (.A1(n_257_76_5373), .A2(n_257_461), .ZN(n_257_76_5746));
   INV_X1 i_257_76_5756 (.A(n_257_76_5746), .ZN(n_257_76_5747));
   NAND4_X1 i_257_76_5757 (.A1(n_257_76_5745), .A2(n_257_76_5371), .A3(
      n_257_76_5747), .A4(n_257_76_5415), .ZN(n_257_76_5748));
   NOR2_X1 i_257_76_5758 (.A1(n_257_76_5748), .A2(n_257_76_5368), .ZN(
      n_257_76_5749));
   NAND3_X1 i_257_76_5759 (.A1(n_257_76_5378), .A2(n_257_451), .A3(n_257_76_5346), 
      .ZN(n_257_76_5750));
   INV_X1 i_257_76_5760 (.A(n_257_76_5750), .ZN(n_257_76_5751));
   NAND3_X1 i_257_76_5761 (.A1(n_257_76_5749), .A2(n_257_76_5751), .A3(
      n_257_76_5381), .ZN(n_257_76_5752));
   INV_X1 i_257_76_5762 (.A(n_257_76_5752), .ZN(n_257_76_5753));
   NAND2_X1 i_257_76_5763 (.A1(n_257_76_5743), .A2(n_257_76_5753), .ZN(
      n_257_76_5754));
   INV_X1 i_257_76_5764 (.A(n_257_76_5345), .ZN(n_257_76_5755));
   NOR2_X1 i_257_76_5765 (.A1(n_257_76_5754), .A2(n_257_76_5755), .ZN(
      n_257_76_5756));
   NAND3_X1 i_257_76_5766 (.A1(n_257_76_5756), .A2(n_257_76_5344), .A3(
      n_257_76_5389), .ZN(n_257_76_5757));
   INV_X1 i_257_76_5767 (.A(n_257_76_5757), .ZN(n_257_76_5758));
   NAND2_X1 i_257_76_5768 (.A1(n_257_76_18063), .A2(n_257_76_5758), .ZN(
      n_257_76_5759));
   NAND3_X1 i_257_76_5769 (.A1(n_257_76_5727), .A2(n_257_76_5742), .A3(
      n_257_76_5759), .ZN(n_257_76_5760));
   INV_X1 i_257_76_5770 (.A(n_257_76_5760), .ZN(n_257_76_5761));
   NAND3_X1 i_257_76_5771 (.A1(n_257_76_5620), .A2(n_257_76_5384), .A3(
      n_257_76_5381), .ZN(n_257_76_5762));
   NAND4_X1 i_257_76_5772 (.A1(n_257_76_5414), .A2(n_257_76_5415), .A3(
      n_257_76_5372), .A4(n_257_76_5373), .ZN(n_257_76_5763));
   NOR2_X1 i_257_76_5773 (.A1(n_257_76_5428), .A2(n_257_76_5763), .ZN(
      n_257_76_5764));
   NAND2_X1 i_257_76_5774 (.A1(n_257_76_5378), .A2(n_257_76_5434), .ZN(
      n_257_76_5765));
   INV_X1 i_257_76_5775 (.A(n_257_76_5765), .ZN(n_257_76_5766));
   NAND2_X1 i_257_76_5776 (.A1(n_257_76_5423), .A2(n_257_424), .ZN(n_257_76_5767));
   INV_X1 i_257_76_5777 (.A(n_257_76_5767), .ZN(n_257_76_5768));
   NAND4_X1 i_257_76_5778 (.A1(n_257_76_5768), .A2(n_257_76_5347), .A3(n_257_510), 
      .A4(n_257_76_5420), .ZN(n_257_76_5769));
   INV_X1 i_257_76_5779 (.A(n_257_76_5769), .ZN(n_257_76_5770));
   NAND4_X1 i_257_76_5780 (.A1(n_257_76_5346), .A2(n_257_76_5430), .A3(
      n_257_76_5770), .A4(n_257_76_5365), .ZN(n_257_76_5771));
   INV_X1 i_257_76_5781 (.A(n_257_76_5771), .ZN(n_257_76_5772));
   NAND3_X1 i_257_76_5782 (.A1(n_257_76_5764), .A2(n_257_76_5766), .A3(
      n_257_76_5772), .ZN(n_257_76_5773));
   NOR2_X1 i_257_76_5783 (.A1(n_257_76_5762), .A2(n_257_76_5773), .ZN(
      n_257_76_5774));
   NAND3_X1 i_257_76_5784 (.A1(n_257_76_5448), .A2(n_257_76_5383), .A3(
      n_257_76_5445), .ZN(n_257_76_5775));
   INV_X1 i_257_76_5785 (.A(n_257_76_5775), .ZN(n_257_76_5776));
   NAND3_X1 i_257_76_5786 (.A1(n_257_76_5774), .A2(n_257_76_5776), .A3(
      n_257_76_5345), .ZN(n_257_76_5777));
   INV_X1 i_257_76_5787 (.A(n_257_76_5777), .ZN(n_257_76_5778));
   NAND3_X1 i_257_76_5788 (.A1(n_257_76_5778), .A2(n_257_76_5668), .A3(
      n_257_76_5344), .ZN(n_257_76_5779));
   INV_X1 i_257_76_5789 (.A(n_257_76_5779), .ZN(n_257_76_5780));
   NAND2_X1 i_257_76_5790 (.A1(n_257_76_18062), .A2(n_257_76_5780), .ZN(
      n_257_76_5781));
   NAND3_X1 i_257_76_5791 (.A1(n_257_76_5445), .A2(n_257_76_5384), .A3(
      n_257_76_5661), .ZN(n_257_76_5782));
   NOR2_X1 i_257_76_5792 (.A1(n_257_76_5782), .A2(n_257_76_5521), .ZN(
      n_257_76_5783));
   NAND2_X1 i_257_76_5793 (.A1(n_257_76_5434), .A2(n_257_76_5430), .ZN(
      n_257_76_5784));
   INV_X1 i_257_76_5794 (.A(n_257_76_5784), .ZN(n_257_76_5785));
   NAND2_X1 i_257_76_5795 (.A1(n_257_422), .A2(n_257_76_5423), .ZN(n_257_76_5786));
   INV_X1 i_257_76_5796 (.A(n_257_76_5786), .ZN(n_257_76_5787));
   NAND4_X1 i_257_76_5797 (.A1(n_257_76_5373), .A2(n_257_76_5787), .A3(
      n_257_76_5347), .A4(n_257_76_5420), .ZN(n_257_76_5788));
   NAND3_X1 i_257_76_5798 (.A1(n_257_76_5416), .A2(n_257_319), .A3(n_257_76_5372), 
      .ZN(n_257_76_5789));
   NOR2_X1 i_257_76_5799 (.A1(n_257_76_5788), .A2(n_257_76_5789), .ZN(
      n_257_76_5790));
   NAND3_X1 i_257_76_5800 (.A1(n_257_76_5365), .A2(n_257_76_5414), .A3(
      n_257_76_5415), .ZN(n_257_76_5791));
   INV_X1 i_257_76_5801 (.A(n_257_76_5791), .ZN(n_257_76_5792));
   NAND3_X1 i_257_76_5802 (.A1(n_257_76_5785), .A2(n_257_76_5790), .A3(
      n_257_76_5792), .ZN(n_257_76_5793));
   INV_X1 i_257_76_5803 (.A(n_257_76_5793), .ZN(n_257_76_5794));
   NAND3_X1 i_257_76_5804 (.A1(n_257_76_5448), .A2(n_257_76_5794), .A3(
      n_257_76_5383), .ZN(n_257_76_5795));
   INV_X1 i_257_76_5805 (.A(n_257_76_5795), .ZN(n_257_76_5796));
   NAND3_X1 i_257_76_5806 (.A1(n_257_76_5783), .A2(n_257_76_5345), .A3(
      n_257_76_5796), .ZN(n_257_76_5797));
   INV_X1 i_257_76_5807 (.A(n_257_76_5797), .ZN(n_257_76_5798));
   NAND3_X1 i_257_76_5808 (.A1(n_257_76_5798), .A2(n_257_76_5668), .A3(
      n_257_76_5344), .ZN(n_257_76_5799));
   INV_X1 i_257_76_5809 (.A(n_257_76_5799), .ZN(n_257_76_5800));
   NAND2_X1 i_257_76_5810 (.A1(n_257_342), .A2(n_257_76_5800), .ZN(n_257_76_5801));
   NAND2_X1 i_257_76_5811 (.A1(n_257_742), .A2(n_257_76_17935), .ZN(
      n_257_76_5802));
   NAND3_X1 i_257_76_5812 (.A1(n_257_76_5802), .A2(n_257_76_5530), .A3(
      n_257_76_5733), .ZN(n_257_76_5803));
   NAND2_X1 i_257_76_5813 (.A1(n_257_84), .A2(n_257_76_17932), .ZN(n_257_76_5804));
   NAND2_X1 i_257_76_5814 (.A1(n_257_76_5793), .A2(n_257_76_5804), .ZN(
      n_257_76_5805));
   NOR2_X1 i_257_76_5815 (.A1(n_257_76_5803), .A2(n_257_76_5805), .ZN(
      n_257_76_5806));
   NAND3_X1 i_257_76_5816 (.A1(n_257_76_18047), .A2(n_257_449), .A3(n_257_1082), 
      .ZN(n_257_76_5807));
   NAND2_X1 i_257_76_5817 (.A1(n_257_972), .A2(n_257_442), .ZN(n_257_76_5808));
   INV_X1 i_257_76_5818 (.A(n_257_76_5808), .ZN(n_257_76_5809));
   NAND2_X1 i_257_76_5819 (.A1(n_257_441), .A2(n_257_76_5809), .ZN(n_257_76_5810));
   NAND2_X1 i_257_76_5820 (.A1(n_257_76_5807), .A2(n_257_76_5810), .ZN(
      n_257_76_5811));
   INV_X1 i_257_76_5821 (.A(n_257_76_5811), .ZN(n_257_76_5812));
   NAND2_X1 i_257_76_5822 (.A1(n_257_44), .A2(n_257_76_17918), .ZN(n_257_76_5813));
   NAND2_X1 i_257_76_5823 (.A1(n_257_428), .A2(n_257_574), .ZN(n_257_76_5814));
   NAND2_X1 i_257_76_5824 (.A1(n_257_76_5423), .A2(n_257_76_5814), .ZN(
      n_257_76_5815));
   INV_X1 i_257_76_5825 (.A(n_257_76_5815), .ZN(n_257_76_5816));
   INV_X1 i_257_76_5826 (.A(Small_Packet_Data_Size[9]), .ZN(n_257_76_5817));
   NAND3_X1 i_257_76_5827 (.A1(n_257_76_5816), .A2(n_257_76_5347), .A3(
      n_257_76_18048), .ZN(n_257_76_5818));
   NAND2_X1 i_257_76_5828 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[9]), 
      .ZN(n_257_76_5819));
   NAND2_X1 i_257_76_5829 (.A1(n_257_76_5818), .A2(n_257_76_5819), .ZN(
      n_257_76_5820));
   NAND3_X1 i_257_76_5830 (.A1(n_257_76_5653), .A2(n_257_76_5813), .A3(
      n_257_76_5820), .ZN(n_257_76_5821));
   INV_X1 i_257_76_5831 (.A(n_257_76_5821), .ZN(n_257_76_5822));
   NAND2_X1 i_257_76_5832 (.A1(n_257_838), .A2(n_257_442), .ZN(n_257_76_5823));
   INV_X1 i_257_76_5833 (.A(n_257_76_5823), .ZN(n_257_76_5824));
   NAND2_X1 i_257_76_5834 (.A1(n_257_446), .A2(n_257_76_5824), .ZN(n_257_76_5825));
   NAND2_X1 i_257_76_5835 (.A1(n_257_710), .A2(n_257_76_15655), .ZN(
      n_257_76_5826));
   INV_X1 i_257_76_5836 (.A(n_257_76_5685), .ZN(n_257_76_5827));
   NAND2_X1 i_257_76_5837 (.A1(n_257_447), .A2(n_257_76_5827), .ZN(n_257_76_5828));
   NAND3_X1 i_257_76_5838 (.A1(n_257_76_5825), .A2(n_257_76_5826), .A3(
      n_257_76_5828), .ZN(n_257_76_5829));
   INV_X1 i_257_76_5839 (.A(n_257_76_5829), .ZN(n_257_76_5830));
   NAND2_X1 i_257_76_5840 (.A1(n_257_638), .A2(n_257_76_17928), .ZN(
      n_257_76_5831));
   NAND3_X1 i_257_76_5841 (.A1(n_257_438), .A2(n_257_1074), .A3(n_257_442), 
      .ZN(n_257_76_5832));
   NAND2_X1 i_257_76_5842 (.A1(n_257_440), .A2(n_257_76_5349), .ZN(n_257_76_5833));
   NAND4_X1 i_257_76_5843 (.A1(n_257_76_5769), .A2(n_257_76_5831), .A3(
      n_257_76_5832), .A4(n_257_76_5833), .ZN(n_257_76_5834));
   INV_X1 i_257_76_5844 (.A(n_257_76_5834), .ZN(n_257_76_5835));
   NAND4_X1 i_257_76_5845 (.A1(n_257_76_5812), .A2(n_257_76_5822), .A3(
      n_257_76_5830), .A4(n_257_76_5835), .ZN(n_257_76_5836));
   NAND2_X1 i_257_76_5846 (.A1(n_257_870), .A2(n_257_76_17903), .ZN(
      n_257_76_5837));
   NAND2_X1 i_257_76_5847 (.A1(n_257_461), .A2(n_257_442), .ZN(n_257_76_5838));
   INV_X1 i_257_76_5848 (.A(n_257_76_5838), .ZN(n_257_76_5839));
   NAND2_X1 i_257_76_5849 (.A1(n_257_451), .A2(n_257_76_5839), .ZN(n_257_76_5840));
   NAND2_X1 i_257_76_5850 (.A1(n_257_122), .A2(n_257_76_17925), .ZN(
      n_257_76_5841));
   NAND2_X1 i_257_76_5851 (.A1(n_257_908), .A2(n_257_76_17940), .ZN(
      n_257_76_5842));
   NAND4_X1 i_257_76_5852 (.A1(n_257_76_5837), .A2(n_257_76_5840), .A3(
      n_257_76_5841), .A4(n_257_76_5842), .ZN(n_257_76_5843));
   NOR2_X1 i_257_76_5853 (.A1(n_257_76_5836), .A2(n_257_76_5843), .ZN(
      n_257_76_5844));
   AOI22_X1 i_257_76_5854 (.A1(n_257_161), .A2(n_257_76_17331), .B1(n_257_806), 
      .B2(n_257_76_17952), .ZN(n_257_76_5845));
   NAND4_X1 i_257_76_5855 (.A1(n_257_76_5722), .A2(n_257_76_5806), .A3(
      n_257_76_5844), .A4(n_257_76_5845), .ZN(n_257_76_5846));
   NAND2_X1 i_257_76_5856 (.A1(n_257_678), .A2(n_257_76_17958), .ZN(
      n_257_76_5847));
   NAND2_X1 i_257_76_5857 (.A1(n_257_1004), .A2(n_257_76_17964), .ZN(
      n_257_76_5848));
   NAND2_X1 i_257_76_5858 (.A1(n_257_76_5847), .A2(n_257_76_5848), .ZN(
      n_257_76_5849));
   NOR2_X1 i_257_76_5859 (.A1(n_257_76_5846), .A2(n_257_76_5849), .ZN(
      n_257_76_5850));
   INV_X1 i_257_76_5860 (.A(n_257_1036), .ZN(n_257_76_5851));
   OAI21_X1 i_257_76_5861 (.A(n_257_76_5449), .B1(n_257_76_5851), .B2(
      n_257_76_17968), .ZN(n_257_76_5852));
   INV_X1 i_257_76_5862 (.A(n_257_76_5852), .ZN(n_257_76_5853));
   NAND2_X1 i_257_76_5863 (.A1(n_257_76_5423), .A2(n_257_425), .ZN(n_257_76_5854));
   INV_X1 i_257_76_5864 (.A(n_257_76_5854), .ZN(n_257_76_5855));
   NAND3_X1 i_257_76_5865 (.A1(n_257_76_5855), .A2(n_257_76_5347), .A3(
      n_257_76_5420), .ZN(n_257_76_5856));
   NOR2_X1 i_257_76_5866 (.A1(n_257_76_5374), .A2(n_257_76_5856), .ZN(
      n_257_76_5857));
   NAND2_X1 i_257_76_5867 (.A1(n_257_76_5414), .A2(n_257_76_5415), .ZN(
      n_257_76_5858));
   INV_X1 i_257_76_5868 (.A(n_257_76_5858), .ZN(n_257_76_5859));
   NAND3_X1 i_257_76_5869 (.A1(n_257_76_5857), .A2(n_257_76_5859), .A3(
      n_257_76_5371), .ZN(n_257_76_5860));
   NAND4_X1 i_257_76_5870 (.A1(n_257_76_5430), .A2(n_257_76_5365), .A3(
      n_257_76_5366), .A4(n_257_76_5367), .ZN(n_257_76_5861));
   NOR2_X1 i_257_76_5871 (.A1(n_257_76_5860), .A2(n_257_76_5861), .ZN(
      n_257_76_5862));
   NAND3_X1 i_257_76_5872 (.A1(n_257_76_5378), .A2(n_257_76_5434), .A3(
      n_257_76_5346), .ZN(n_257_76_5863));
   INV_X1 i_257_76_5873 (.A(n_257_76_5863), .ZN(n_257_76_5864));
   NAND4_X1 i_257_76_5874 (.A1(n_257_76_5862), .A2(n_257_76_5620), .A3(
      n_257_76_5381), .A4(n_257_76_5864), .ZN(n_257_76_5865));
   NOR2_X1 i_257_76_5875 (.A1(n_257_76_5865), .A2(n_257_76_5479), .ZN(
      n_257_76_5866));
   NAND2_X1 i_257_76_5876 (.A1(n_257_241), .A2(n_257_76_5448), .ZN(n_257_76_5867));
   INV_X1 i_257_76_5877 (.A(n_257_76_5867), .ZN(n_257_76_5868));
   NAND3_X1 i_257_76_5878 (.A1(n_257_76_5866), .A2(n_257_76_5868), .A3(
      n_257_76_5389), .ZN(n_257_76_5869));
   NAND3_X1 i_257_76_5879 (.A1(n_257_76_5850), .A2(n_257_76_5853), .A3(
      n_257_76_5869), .ZN(n_257_76_5870));
   INV_X1 i_257_76_5880 (.A(n_257_76_5870), .ZN(n_257_76_5871));
   NAND4_X1 i_257_76_5881 (.A1(n_257_76_5371), .A2(n_257_76_5657), .A3(
      n_257_76_5414), .A4(n_257_76_5415), .ZN(n_257_76_5872));
   NAND2_X1 i_257_76_5882 (.A1(n_257_76_5416), .A2(n_257_76_5372), .ZN(
      n_257_76_5873));
   INV_X1 i_257_76_5883 (.A(n_257_76_5873), .ZN(n_257_76_5874));
   NAND2_X1 i_257_76_5884 (.A1(n_257_420), .A2(n_257_662), .ZN(n_257_76_5875));
   NAND2_X1 i_257_76_5885 (.A1(n_257_76_5373), .A2(n_257_76_5875), .ZN(
      n_257_76_5876));
   INV_X1 i_257_76_5886 (.A(n_257_76_5876), .ZN(n_257_76_5877));
   NAND3_X1 i_257_76_5887 (.A1(n_257_397), .A2(n_257_484), .A3(n_257_442), 
      .ZN(n_257_76_5878));
   INV_X1 i_257_76_5888 (.A(n_257_76_5878), .ZN(n_257_76_5879));
   NAND3_X1 i_257_76_5889 (.A1(n_257_76_5423), .A2(n_257_76_5814), .A3(
      n_257_76_5879), .ZN(n_257_76_5880));
   NOR2_X1 i_257_76_5890 (.A1(n_257_76_5880), .A2(n_257_1068), .ZN(n_257_76_5881));
   NAND3_X1 i_257_76_5891 (.A1(n_257_76_5874), .A2(n_257_76_5877), .A3(
      n_257_76_5881), .ZN(n_257_76_5882));
   NOR3_X1 i_257_76_5892 (.A1(n_257_76_5861), .A2(n_257_76_5872), .A3(
      n_257_76_5882), .ZN(n_257_76_5883));
   NAND3_X1 i_257_76_5893 (.A1(n_257_76_5883), .A2(n_257_76_5448), .A3(
      n_257_76_5383), .ZN(n_257_76_5884));
   INV_X1 i_257_76_5894 (.A(n_257_76_5884), .ZN(n_257_76_5885));
   NAND4_X1 i_257_76_5895 (.A1(n_257_76_5620), .A2(n_257_76_5864), .A3(
      n_257_76_5381), .A4(n_257_76_5662), .ZN(n_257_76_5886));
   NOR2_X1 i_257_76_5896 (.A1(n_257_76_5886), .A2(n_257_76_5782), .ZN(
      n_257_76_5887));
   NAND3_X1 i_257_76_5897 (.A1(n_257_76_5885), .A2(n_257_76_5345), .A3(
      n_257_76_5887), .ZN(n_257_76_5888));
   NOR3_X1 i_257_76_5898 (.A1(n_257_76_5888), .A2(n_257_76_5497), .A3(
      n_257_76_5667), .ZN(n_257_76_5889));
   AOI21_X1 i_257_76_5899 (.A(n_257_76_5871), .B1(n_257_76_18060), .B2(
      n_257_76_5889), .ZN(n_257_76_5890));
   NAND3_X1 i_257_76_5900 (.A1(n_257_76_5781), .A2(n_257_76_5801), .A3(
      n_257_76_5890), .ZN(n_257_76_5891));
   INV_X1 i_257_76_5901 (.A(n_257_76_5891), .ZN(n_257_76_5892));
   NAND4_X1 i_257_76_5902 (.A1(n_257_76_5346), .A2(n_257_76_5366), .A3(
      n_257_76_5371), .A4(n_257_448), .ZN(n_257_76_5893));
   INV_X1 i_257_76_5903 (.A(n_257_76_5893), .ZN(n_257_76_5894));
   NAND3_X1 i_257_76_5904 (.A1(n_257_76_5608), .A2(n_257_76_5381), .A3(
      n_257_76_5894), .ZN(n_257_76_5895));
   NOR2_X1 i_257_76_5905 (.A1(n_257_76_5895), .A2(n_257_76_5385), .ZN(
      n_257_76_5896));
   NAND3_X1 i_257_76_5906 (.A1(n_257_76_5896), .A2(n_257_76_5345), .A3(n_257_678), 
      .ZN(n_257_76_5897));
   NOR2_X1 i_257_76_5907 (.A1(n_257_76_5897), .A2(n_257_76_5497), .ZN(
      n_257_76_5898));
   NAND2_X1 i_257_76_5908 (.A1(n_257_76_5344), .A2(n_257_76_5345), .ZN(
      n_257_76_5899));
   NOR2_X1 i_257_76_5909 (.A1(n_257_76_5869), .A2(n_257_76_5899), .ZN(
      n_257_76_5900));
   AOI22_X1 i_257_76_5910 (.A1(n_257_76_18079), .A2(n_257_76_5898), .B1(
      n_257_76_18064), .B2(n_257_76_5900), .ZN(n_257_76_5901));
   NAND3_X1 i_257_76_5911 (.A1(n_257_76_5761), .A2(n_257_76_5892), .A3(
      n_257_76_5901), .ZN(n_257_76_5902));
   NOR2_X1 i_257_76_5912 (.A1(n_257_76_5708), .A2(n_257_76_5902), .ZN(
      n_257_76_5903));
   NAND2_X1 i_257_76_5913 (.A1(n_257_76_5589), .A2(n_257_76_5903), .ZN(n_9));
   NAND2_X1 i_257_76_5914 (.A1(n_257_1037), .A2(n_257_443), .ZN(n_257_76_5904));
   NAND2_X1 i_257_76_5915 (.A1(n_257_1005), .A2(n_257_444), .ZN(n_257_76_5905));
   NAND2_X1 i_257_76_5916 (.A1(n_257_441), .A2(n_257_973), .ZN(n_257_76_5906));
   INV_X1 i_257_76_5917 (.A(n_257_1069), .ZN(n_257_76_5907));
   NAND2_X1 i_257_76_5918 (.A1(n_257_941), .A2(n_257_442), .ZN(n_257_76_5908));
   INV_X1 i_257_76_5919 (.A(n_257_76_5908), .ZN(n_257_76_5909));
   NAND3_X1 i_257_76_5920 (.A1(n_257_76_5907), .A2(n_257_440), .A3(n_257_76_5909), 
      .ZN(n_257_76_5910));
   INV_X1 i_257_76_5921 (.A(n_257_76_5910), .ZN(n_257_76_5911));
   NAND2_X1 i_257_76_5922 (.A1(n_257_76_5906), .A2(n_257_76_5911), .ZN(
      n_257_76_5912));
   INV_X1 i_257_76_5923 (.A(n_257_76_5912), .ZN(n_257_76_5913));
   NAND2_X1 i_257_76_5924 (.A1(n_257_76_5905), .A2(n_257_76_5913), .ZN(
      n_257_76_5914));
   INV_X1 i_257_76_5925 (.A(n_257_76_5914), .ZN(n_257_76_5915));
   NAND2_X1 i_257_76_5926 (.A1(n_257_76_5904), .A2(n_257_76_5915), .ZN(
      n_257_76_5916));
   INV_X1 i_257_76_5927 (.A(n_257_76_5916), .ZN(n_257_76_5917));
   NAND2_X1 i_257_76_5928 (.A1(n_257_17), .A2(n_257_76_5917), .ZN(n_257_76_5918));
   NOR2_X1 i_257_76_5929 (.A1(n_257_1069), .A2(n_257_76_17412), .ZN(
      n_257_76_5919));
   INV_X1 i_257_76_5930 (.A(n_257_76_5919), .ZN(n_257_76_5920));
   NOR2_X1 i_257_76_5931 (.A1(n_257_76_5920), .A2(n_257_76_15197), .ZN(
      n_257_76_5921));
   NAND2_X1 i_257_76_5932 (.A1(n_257_1037), .A2(n_257_76_5921), .ZN(
      n_257_76_5922));
   INV_X1 i_257_76_5933 (.A(n_257_76_5922), .ZN(n_257_76_5923));
   NAND2_X1 i_257_76_5934 (.A1(n_257_76_18072), .A2(n_257_76_5923), .ZN(
      n_257_76_5924));
   INV_X1 i_257_76_5935 (.A(n_257_76_5905), .ZN(n_257_76_5925));
   NOR2_X1 i_257_76_5936 (.A1(n_257_1069), .A2(n_257_76_17927), .ZN(
      n_257_76_5926));
   NAND2_X1 i_257_76_5937 (.A1(n_257_440), .A2(n_257_941), .ZN(n_257_76_5927));
   NAND3_X1 i_257_76_5938 (.A1(n_257_76_5926), .A2(n_257_76_5927), .A3(n_257_639), 
      .ZN(n_257_76_5928));
   INV_X1 i_257_76_5939 (.A(n_257_76_5928), .ZN(n_257_76_5929));
   NAND2_X1 i_257_76_5940 (.A1(n_257_449), .A2(n_257_1083), .ZN(n_257_76_5930));
   NAND2_X1 i_257_76_5941 (.A1(n_257_447), .A2(n_257_775), .ZN(n_257_76_5931));
   NAND2_X1 i_257_76_5942 (.A1(n_257_1075), .A2(n_257_438), .ZN(n_257_76_5932));
   NAND4_X1 i_257_76_5943 (.A1(n_257_76_5929), .A2(n_257_76_5930), .A3(
      n_257_76_5931), .A4(n_257_76_5932), .ZN(n_257_76_5933));
   NAND2_X1 i_257_76_5944 (.A1(n_257_711), .A2(n_257_435), .ZN(n_257_76_5934));
   NAND2_X1 i_257_76_5945 (.A1(n_257_446), .A2(n_257_839), .ZN(n_257_76_5935));
   NAND3_X1 i_257_76_5946 (.A1(n_257_76_5906), .A2(n_257_76_5934), .A3(
      n_257_76_5935), .ZN(n_257_76_5936));
   NOR2_X1 i_257_76_5947 (.A1(n_257_76_5933), .A2(n_257_76_5936), .ZN(
      n_257_76_5937));
   NAND2_X1 i_257_76_5948 (.A1(n_257_871), .A2(n_257_445), .ZN(n_257_76_5938));
   NAND2_X1 i_257_76_5949 (.A1(n_257_909), .A2(n_257_439), .ZN(n_257_76_5939));
   NAND2_X1 i_257_76_5950 (.A1(n_257_76_5938), .A2(n_257_76_5939), .ZN(
      n_257_76_5940));
   INV_X1 i_257_76_5951 (.A(n_257_76_5940), .ZN(n_257_76_5941));
   NAND2_X1 i_257_76_5952 (.A1(n_257_743), .A2(n_257_436), .ZN(n_257_76_5942));
   NAND2_X1 i_257_76_5953 (.A1(n_257_807), .A2(n_257_437), .ZN(n_257_76_5943));
   NAND4_X1 i_257_76_5954 (.A1(n_257_76_5937), .A2(n_257_76_5941), .A3(
      n_257_76_5942), .A4(n_257_76_5943), .ZN(n_257_76_5944));
   NOR2_X1 i_257_76_5955 (.A1(n_257_76_5925), .A2(n_257_76_5944), .ZN(
      n_257_76_5945));
   NAND2_X1 i_257_76_5956 (.A1(n_257_679), .A2(n_257_448), .ZN(n_257_76_5946));
   NAND3_X1 i_257_76_5957 (.A1(n_257_76_5945), .A2(n_257_76_5904), .A3(
      n_257_76_5946), .ZN(n_257_76_5947));
   INV_X1 i_257_76_5958 (.A(n_257_76_5947), .ZN(n_257_76_5948));
   NAND2_X1 i_257_76_5959 (.A1(n_257_28), .A2(n_257_76_5948), .ZN(n_257_76_5949));
   NAND3_X1 i_257_76_5960 (.A1(n_257_76_5918), .A2(n_257_76_5924), .A3(
      n_257_76_5949), .ZN(n_257_76_5950));
   NAND2_X1 i_257_76_5961 (.A1(n_257_76_5932), .A2(n_257_446), .ZN(n_257_76_5951));
   INV_X1 i_257_76_5962 (.A(n_257_76_5951), .ZN(n_257_76_5952));
   NAND3_X1 i_257_76_5963 (.A1(n_257_76_5919), .A2(n_257_76_5927), .A3(n_257_839), 
      .ZN(n_257_76_5953));
   INV_X1 i_257_76_5964 (.A(n_257_76_5953), .ZN(n_257_76_5954));
   NAND3_X1 i_257_76_5965 (.A1(n_257_76_5906), .A2(n_257_76_5952), .A3(
      n_257_76_5954), .ZN(n_257_76_5955));
   INV_X1 i_257_76_5966 (.A(n_257_76_5955), .ZN(n_257_76_5956));
   NAND3_X1 i_257_76_5967 (.A1(n_257_76_5938), .A2(n_257_76_5956), .A3(
      n_257_76_5939), .ZN(n_257_76_5957));
   INV_X1 i_257_76_5968 (.A(n_257_76_5957), .ZN(n_257_76_5958));
   NAND2_X1 i_257_76_5969 (.A1(n_257_76_5905), .A2(n_257_76_5958), .ZN(
      n_257_76_5959));
   INV_X1 i_257_76_5970 (.A(n_257_76_5959), .ZN(n_257_76_5960));
   NAND2_X1 i_257_76_5971 (.A1(n_257_76_5904), .A2(n_257_76_5960), .ZN(
      n_257_76_5961));
   INV_X1 i_257_76_5972 (.A(n_257_76_5961), .ZN(n_257_76_5962));
   NAND2_X1 i_257_76_5973 (.A1(n_257_76_18070), .A2(n_257_76_5962), .ZN(
      n_257_76_5963));
   NAND3_X1 i_257_76_5974 (.A1(n_257_76_5919), .A2(n_257_76_5927), .A3(n_257_439), 
      .ZN(n_257_76_5964));
   INV_X1 i_257_76_5975 (.A(n_257_76_5964), .ZN(n_257_76_5965));
   NAND3_X1 i_257_76_5976 (.A1(n_257_76_5906), .A2(n_257_76_5965), .A3(n_257_909), 
      .ZN(n_257_76_5966));
   INV_X1 i_257_76_5977 (.A(n_257_76_5966), .ZN(n_257_76_5967));
   NAND2_X1 i_257_76_5978 (.A1(n_257_76_5905), .A2(n_257_76_5967), .ZN(
      n_257_76_5968));
   INV_X1 i_257_76_5979 (.A(n_257_76_5968), .ZN(n_257_76_5969));
   NAND2_X1 i_257_76_5980 (.A1(n_257_76_5904), .A2(n_257_76_5969), .ZN(
      n_257_76_5970));
   INV_X1 i_257_76_5981 (.A(n_257_76_5970), .ZN(n_257_76_5971));
   NAND2_X1 i_257_76_5982 (.A1(n_257_76_18084), .A2(n_257_76_5971), .ZN(
      n_257_76_5972));
   NAND2_X1 i_257_76_5983 (.A1(n_257_45), .A2(n_257_433), .ZN(n_257_76_5973));
   NAND2_X1 i_257_76_5984 (.A1(n_257_543), .A2(n_257_426), .ZN(n_257_76_5974));
   NAND3_X1 i_257_76_5985 (.A1(n_257_76_5973), .A2(n_257_76_5974), .A3(
      n_257_76_5906), .ZN(n_257_76_5975));
   NAND3_X1 i_257_76_5986 (.A1(n_257_282), .A2(n_257_76_5934), .A3(n_257_76_5935), 
      .ZN(n_257_76_5976));
   NOR2_X1 i_257_76_5987 (.A1(n_257_76_5975), .A2(n_257_76_5976), .ZN(
      n_257_76_5977));
   NAND2_X1 i_257_76_5988 (.A1(n_257_202), .A2(n_257_427), .ZN(n_257_76_5978));
   NAND2_X1 i_257_76_5989 (.A1(n_257_639), .A2(n_257_450), .ZN(n_257_76_5979));
   NAND4_X1 i_257_76_5990 (.A1(n_257_76_5930), .A2(n_257_76_5931), .A3(
      n_257_76_5978), .A4(n_257_76_5979), .ZN(n_257_76_5980));
   NAND2_X1 i_257_76_5991 (.A1(n_257_432), .A2(n_257_607), .ZN(n_257_76_5981));
   NAND2_X1 i_257_76_5992 (.A1(n_257_76_5981), .A2(n_257_423), .ZN(n_257_76_5982));
   INV_X1 i_257_76_5993 (.A(n_257_76_5982), .ZN(n_257_76_5983));
   INV_X1 i_257_76_5994 (.A(n_257_575), .ZN(n_257_76_5984));
   NAND2_X1 i_257_76_5995 (.A1(n_257_76_5984), .A2(n_257_442), .ZN(n_257_76_5985));
   OAI21_X1 i_257_76_5996 (.A(n_257_76_5985), .B1(n_257_428), .B2(n_257_76_17412), 
      .ZN(n_257_76_5986));
   NAND3_X1 i_257_76_5997 (.A1(n_257_76_5983), .A2(n_257_76_5907), .A3(
      n_257_76_5986), .ZN(n_257_76_5987));
   INV_X1 i_257_76_5998 (.A(n_257_76_5987), .ZN(n_257_76_5988));
   NAND2_X1 i_257_76_5999 (.A1(n_257_511), .A2(n_257_424), .ZN(n_257_76_5989));
   NAND4_X1 i_257_76_6000 (.A1(n_257_76_5988), .A2(n_257_76_5932), .A3(
      n_257_76_5989), .A4(n_257_76_5927), .ZN(n_257_76_5990));
   NOR2_X1 i_257_76_6001 (.A1(n_257_76_5980), .A2(n_257_76_5990), .ZN(
      n_257_76_5991));
   NAND2_X1 i_257_76_6002 (.A1(n_257_123), .A2(n_257_430), .ZN(n_257_76_5992));
   NAND2_X1 i_257_76_6003 (.A1(n_257_76_5992), .A2(n_257_76_5939), .ZN(
      n_257_76_5993));
   INV_X1 i_257_76_6004 (.A(n_257_76_5993), .ZN(n_257_76_5994));
   NAND4_X1 i_257_76_6005 (.A1(n_257_76_5977), .A2(n_257_76_5991), .A3(
      n_257_76_5994), .A4(n_257_76_5938), .ZN(n_257_76_5995));
   INV_X1 i_257_76_6006 (.A(n_257_76_5995), .ZN(n_257_76_5996));
   NAND2_X1 i_257_76_6007 (.A1(n_257_76_5946), .A2(n_257_76_5996), .ZN(
      n_257_76_5997));
   INV_X1 i_257_76_6008 (.A(n_257_76_5997), .ZN(n_257_76_5998));
   NAND2_X1 i_257_76_6009 (.A1(n_257_242), .A2(n_257_425), .ZN(n_257_76_5999));
   NAND2_X1 i_257_76_6010 (.A1(n_257_162), .A2(n_257_429), .ZN(n_257_76_6000));
   NAND2_X1 i_257_76_6011 (.A1(n_257_76_5999), .A2(n_257_76_6000), .ZN(
      n_257_76_6001));
   INV_X1 i_257_76_6012 (.A(n_257_76_6001), .ZN(n_257_76_6002));
   NAND2_X1 i_257_76_6013 (.A1(n_257_85), .A2(n_257_431), .ZN(n_257_76_6003));
   NAND2_X1 i_257_76_6014 (.A1(n_257_451), .A2(n_257_462), .ZN(n_257_76_6004));
   NAND4_X1 i_257_76_6015 (.A1(n_257_76_5942), .A2(n_257_76_6003), .A3(
      n_257_76_5943), .A4(n_257_76_6004), .ZN(n_257_76_6005));
   INV_X1 i_257_76_6016 (.A(n_257_76_6005), .ZN(n_257_76_6006));
   NAND3_X1 i_257_76_6017 (.A1(n_257_76_5905), .A2(n_257_76_6002), .A3(
      n_257_76_6006), .ZN(n_257_76_6007));
   INV_X1 i_257_76_6018 (.A(n_257_76_6007), .ZN(n_257_76_6008));
   NAND3_X1 i_257_76_6019 (.A1(n_257_76_5998), .A2(n_257_76_6008), .A3(
      n_257_76_5904), .ZN(n_257_76_6009));
   INV_X1 i_257_76_6020 (.A(n_257_76_6009), .ZN(n_257_76_6010));
   NAND2_X1 i_257_76_6021 (.A1(n_257_76_18066), .A2(n_257_76_6010), .ZN(
      n_257_76_6011));
   NAND3_X1 i_257_76_6022 (.A1(n_257_76_5963), .A2(n_257_76_5972), .A3(
      n_257_76_6011), .ZN(n_257_76_6012));
   NOR2_X1 i_257_76_6023 (.A1(n_257_76_5950), .A2(n_257_76_6012), .ZN(
      n_257_76_6013));
   NAND2_X1 i_257_76_6024 (.A1(n_257_76_5919), .A2(n_257_973), .ZN(n_257_76_6014));
   NOR2_X1 i_257_76_6025 (.A1(n_257_76_13147), .A2(n_257_76_6014), .ZN(
      n_257_76_6015));
   NAND2_X1 i_257_76_6026 (.A1(n_257_76_5905), .A2(n_257_76_6015), .ZN(
      n_257_76_6016));
   INV_X1 i_257_76_6027 (.A(n_257_76_6016), .ZN(n_257_76_6017));
   NAND2_X1 i_257_76_6028 (.A1(n_257_76_5904), .A2(n_257_76_6017), .ZN(
      n_257_76_6018));
   INV_X1 i_257_76_6029 (.A(n_257_76_6018), .ZN(n_257_76_6019));
   NAND2_X1 i_257_76_6030 (.A1(n_257_76_18071), .A2(n_257_76_6019), .ZN(
      n_257_76_6020));
   INV_X1 i_257_76_6031 (.A(n_257_76_5904), .ZN(n_257_76_6021));
   NOR2_X1 i_257_76_6032 (.A1(n_257_1069), .A2(n_257_76_15289), .ZN(
      n_257_76_6022));
   NAND2_X1 i_257_76_6033 (.A1(n_257_76_5927), .A2(n_257_76_6022), .ZN(
      n_257_76_6023));
   INV_X1 i_257_76_6034 (.A(n_257_76_6023), .ZN(n_257_76_6024));
   NAND4_X1 i_257_76_6035 (.A1(n_257_76_6024), .A2(n_257_76_5931), .A3(n_257_711), 
      .A4(n_257_76_5932), .ZN(n_257_76_6025));
   NAND2_X1 i_257_76_6036 (.A1(n_257_76_5906), .A2(n_257_76_5935), .ZN(
      n_257_76_6026));
   NOR2_X1 i_257_76_6037 (.A1(n_257_76_6025), .A2(n_257_76_6026), .ZN(
      n_257_76_6027));
   NAND4_X1 i_257_76_6038 (.A1(n_257_76_5941), .A2(n_257_76_5942), .A3(
      n_257_76_6027), .A4(n_257_76_5943), .ZN(n_257_76_6028));
   INV_X1 i_257_76_6039 (.A(n_257_76_6028), .ZN(n_257_76_6029));
   NAND2_X1 i_257_76_6040 (.A1(n_257_76_5905), .A2(n_257_76_6029), .ZN(
      n_257_76_6030));
   NOR2_X1 i_257_76_6041 (.A1(n_257_76_6021), .A2(n_257_76_6030), .ZN(
      n_257_76_6031));
   NAND2_X1 i_257_76_6042 (.A1(n_257_76_18078), .A2(n_257_76_6031), .ZN(
      n_257_76_6032));
   NAND3_X1 i_257_76_6043 (.A1(n_257_76_5935), .A2(n_257_76_5930), .A3(
      n_257_76_5931), .ZN(n_257_76_6033));
   NAND2_X1 i_257_76_6044 (.A1(n_257_575), .A2(n_257_442), .ZN(n_257_76_6034));
   INV_X1 i_257_76_6045 (.A(n_257_76_6034), .ZN(n_257_76_6035));
   NAND2_X1 i_257_76_6046 (.A1(n_257_428), .A2(n_257_76_6035), .ZN(n_257_76_6036));
   INV_X1 i_257_76_6047 (.A(n_257_76_6036), .ZN(n_257_76_6037));
   NAND2_X1 i_257_76_6048 (.A1(n_257_76_6037), .A2(n_257_76_5981), .ZN(
      n_257_76_6038));
   NOR2_X1 i_257_76_6049 (.A1(n_257_76_6038), .A2(n_257_1069), .ZN(n_257_76_6039));
   NAND4_X1 i_257_76_6050 (.A1(n_257_76_6039), .A2(n_257_76_5979), .A3(
      n_257_76_5932), .A4(n_257_76_5927), .ZN(n_257_76_6040));
   NOR2_X1 i_257_76_6051 (.A1(n_257_76_6033), .A2(n_257_76_6040), .ZN(
      n_257_76_6041));
   NAND3_X1 i_257_76_6052 (.A1(n_257_76_5973), .A2(n_257_76_5906), .A3(
      n_257_76_5934), .ZN(n_257_76_6042));
   INV_X1 i_257_76_6053 (.A(n_257_76_6042), .ZN(n_257_76_6043));
   NAND4_X1 i_257_76_6054 (.A1(n_257_76_6041), .A2(n_257_76_6043), .A3(
      n_257_76_5992), .A4(n_257_76_5939), .ZN(n_257_76_6044));
   NAND3_X1 i_257_76_6055 (.A1(n_257_76_5943), .A2(n_257_76_5938), .A3(
      n_257_76_6004), .ZN(n_257_76_6045));
   NOR2_X1 i_257_76_6056 (.A1(n_257_76_6044), .A2(n_257_76_6045), .ZN(
      n_257_76_6046));
   NAND3_X1 i_257_76_6057 (.A1(n_257_76_6000), .A2(n_257_76_5942), .A3(
      n_257_76_6003), .ZN(n_257_76_6047));
   INV_X1 i_257_76_6058 (.A(n_257_76_6047), .ZN(n_257_76_6048));
   NAND4_X1 i_257_76_6059 (.A1(n_257_76_6046), .A2(n_257_76_5946), .A3(
      n_257_76_5905), .A4(n_257_76_6048), .ZN(n_257_76_6049));
   NOR2_X1 i_257_76_6060 (.A1(n_257_76_6049), .A2(n_257_76_6021), .ZN(
      n_257_76_6050));
   NAND2_X1 i_257_76_6061 (.A1(n_257_76_18074), .A2(n_257_76_6050), .ZN(
      n_257_76_6051));
   NAND3_X1 i_257_76_6062 (.A1(n_257_76_6020), .A2(n_257_76_6032), .A3(
      n_257_76_6051), .ZN(n_257_76_6052));
   NAND2_X1 i_257_76_6063 (.A1(n_257_1069), .A2(n_257_442), .ZN(n_257_76_6053));
   INV_X1 i_257_76_6064 (.A(n_257_76_6053), .ZN(n_257_76_6054));
   NAND2_X1 i_257_76_6065 (.A1(n_257_13), .A2(n_257_76_6054), .ZN(n_257_76_6055));
   NOR2_X1 i_257_76_6066 (.A1(n_257_76_17902), .A2(n_257_1069), .ZN(
      n_257_76_6056));
   NAND3_X1 i_257_76_6067 (.A1(n_257_76_5932), .A2(n_257_76_6056), .A3(
      n_257_76_5927), .ZN(n_257_76_6057));
   INV_X1 i_257_76_6068 (.A(n_257_76_6057), .ZN(n_257_76_6058));
   NAND4_X1 i_257_76_6069 (.A1(n_257_871), .A2(n_257_76_5939), .A3(n_257_76_6058), 
      .A4(n_257_76_5906), .ZN(n_257_76_6059));
   INV_X1 i_257_76_6070 (.A(n_257_76_6059), .ZN(n_257_76_6060));
   NAND2_X1 i_257_76_6071 (.A1(n_257_76_5905), .A2(n_257_76_6060), .ZN(
      n_257_76_6061));
   INV_X1 i_257_76_6072 (.A(n_257_76_6061), .ZN(n_257_76_6062));
   NAND2_X1 i_257_76_6073 (.A1(n_257_76_5904), .A2(n_257_76_6062), .ZN(
      n_257_76_6063));
   INV_X1 i_257_76_6074 (.A(n_257_76_6063), .ZN(n_257_76_6064));
   NAND2_X1 i_257_76_6075 (.A1(n_257_76_18077), .A2(n_257_76_6064), .ZN(
      n_257_76_6065));
   NAND2_X1 i_257_76_6076 (.A1(n_257_76_6055), .A2(n_257_76_6065), .ZN(
      n_257_76_6066));
   NOR2_X1 i_257_76_6077 (.A1(n_257_76_6052), .A2(n_257_76_6066), .ZN(
      n_257_76_6067));
   NAND4_X1 i_257_76_6078 (.A1(n_257_76_5906), .A2(n_257_76_5935), .A3(
      n_257_76_5930), .A4(n_257_76_5931), .ZN(n_257_76_6068));
   INV_X1 i_257_76_6079 (.A(n_257_76_6068), .ZN(n_257_76_6069));
   NAND4_X1 i_257_76_6080 (.A1(n_257_76_5994), .A2(n_257_76_6069), .A3(
      n_257_76_5938), .A4(n_257_76_6004), .ZN(n_257_76_6070));
   NAND2_X1 i_257_76_6081 (.A1(n_257_76_6003), .A2(n_257_76_5943), .ZN(
      n_257_76_6071));
   NOR2_X1 i_257_76_6082 (.A1(n_257_76_6070), .A2(n_257_76_6071), .ZN(
      n_257_76_6072));
   INV_X1 i_257_76_6083 (.A(n_257_76_5986), .ZN(n_257_76_6073));
   NOR2_X1 i_257_76_6084 (.A1(n_257_1069), .A2(n_257_76_6073), .ZN(n_257_76_6074));
   NAND2_X1 i_257_76_6085 (.A1(n_257_76_5981), .A2(n_257_426), .ZN(n_257_76_6075));
   INV_X1 i_257_76_6086 (.A(n_257_76_6075), .ZN(n_257_76_6076));
   NAND4_X1 i_257_76_6087 (.A1(n_257_76_5932), .A2(n_257_76_6074), .A3(
      n_257_76_5927), .A4(n_257_76_6076), .ZN(n_257_76_6077));
   INV_X1 i_257_76_6088 (.A(n_257_76_6077), .ZN(n_257_76_6078));
   NAND3_X1 i_257_76_6089 (.A1(n_257_543), .A2(n_257_76_5978), .A3(n_257_76_5979), 
      .ZN(n_257_76_6079));
   INV_X1 i_257_76_6090 (.A(n_257_76_6079), .ZN(n_257_76_6080));
   NAND4_X1 i_257_76_6091 (.A1(n_257_76_6078), .A2(n_257_76_6080), .A3(
      n_257_76_5973), .A4(n_257_76_5934), .ZN(n_257_76_6081));
   INV_X1 i_257_76_6092 (.A(n_257_76_6081), .ZN(n_257_76_6082));
   NAND3_X1 i_257_76_6093 (.A1(n_257_76_6000), .A2(n_257_76_6082), .A3(
      n_257_76_5942), .ZN(n_257_76_6083));
   INV_X1 i_257_76_6094 (.A(n_257_76_6083), .ZN(n_257_76_6084));
   NAND4_X1 i_257_76_6095 (.A1(n_257_76_5946), .A2(n_257_76_6072), .A3(
      n_257_76_5905), .A4(n_257_76_6084), .ZN(n_257_76_6085));
   NOR2_X1 i_257_76_6096 (.A1(n_257_76_6085), .A2(n_257_76_6021), .ZN(
      n_257_76_6086));
   NAND2_X1 i_257_76_6097 (.A1(n_257_76_18076), .A2(n_257_76_6086), .ZN(
      n_257_76_6087));
   NAND2_X1 i_257_76_6098 (.A1(n_257_76_5943), .A2(n_257_743), .ZN(n_257_76_6088));
   NAND2_X1 i_257_76_6099 (.A1(n_257_76_5939), .A2(n_257_76_5906), .ZN(
      n_257_76_6089));
   INV_X1 i_257_76_6100 (.A(n_257_76_6089), .ZN(n_257_76_6090));
   NAND2_X1 i_257_76_6101 (.A1(n_257_76_5935), .A2(n_257_76_5931), .ZN(
      n_257_76_6091));
   NOR2_X1 i_257_76_6102 (.A1(n_257_1069), .A2(n_257_76_17934), .ZN(
      n_257_76_6092));
   NAND3_X1 i_257_76_6103 (.A1(n_257_76_5932), .A2(n_257_76_5927), .A3(
      n_257_76_6092), .ZN(n_257_76_6093));
   NOR2_X1 i_257_76_6104 (.A1(n_257_76_6091), .A2(n_257_76_6093), .ZN(
      n_257_76_6094));
   NAND3_X1 i_257_76_6105 (.A1(n_257_76_6090), .A2(n_257_76_5938), .A3(
      n_257_76_6094), .ZN(n_257_76_6095));
   NOR2_X1 i_257_76_6106 (.A1(n_257_76_6088), .A2(n_257_76_6095), .ZN(
      n_257_76_6096));
   NAND2_X1 i_257_76_6107 (.A1(n_257_76_5905), .A2(n_257_76_6096), .ZN(
      n_257_76_6097));
   INV_X1 i_257_76_6108 (.A(n_257_76_6097), .ZN(n_257_76_6098));
   NAND2_X1 i_257_76_6109 (.A1(n_257_76_5904), .A2(n_257_76_6098), .ZN(
      n_257_76_6099));
   INV_X1 i_257_76_6110 (.A(n_257_76_6099), .ZN(n_257_76_6100));
   NAND2_X1 i_257_76_6111 (.A1(n_257_76_18069), .A2(n_257_76_6100), .ZN(
      n_257_76_6101));
   NAND2_X1 i_257_76_6112 (.A1(n_257_76_6004), .A2(n_257_76_5939), .ZN(
      n_257_76_6102));
   INV_X1 i_257_76_6113 (.A(n_257_76_6102), .ZN(n_257_76_6103));
   NAND4_X1 i_257_76_6114 (.A1(n_257_76_5973), .A2(n_257_76_5906), .A3(
      n_257_76_5934), .A4(n_257_76_5935), .ZN(n_257_76_6104));
   INV_X1 i_257_76_6115 (.A(n_257_76_6104), .ZN(n_257_76_6105));
   NAND2_X1 i_257_76_6116 (.A1(n_257_607), .A2(n_257_442), .ZN(n_257_76_6106));
   INV_X1 i_257_76_6117 (.A(n_257_76_6106), .ZN(n_257_76_6107));
   NAND2_X1 i_257_76_6118 (.A1(n_257_432), .A2(n_257_76_6107), .ZN(n_257_76_6108));
   NOR2_X1 i_257_76_6119 (.A1(n_257_1069), .A2(n_257_76_6108), .ZN(n_257_76_6109));
   NAND4_X1 i_257_76_6120 (.A1(n_257_76_5979), .A2(n_257_76_5932), .A3(
      n_257_76_5927), .A4(n_257_76_6109), .ZN(n_257_76_6110));
   NAND2_X1 i_257_76_6121 (.A1(n_257_76_5930), .A2(n_257_76_5931), .ZN(
      n_257_76_6111));
   NOR2_X1 i_257_76_6122 (.A1(n_257_76_6110), .A2(n_257_76_6111), .ZN(
      n_257_76_6112));
   NAND4_X1 i_257_76_6123 (.A1(n_257_76_6103), .A2(n_257_76_6105), .A3(
      n_257_76_6112), .A4(n_257_76_5938), .ZN(n_257_76_6113));
   NAND2_X1 i_257_76_6124 (.A1(n_257_76_5942), .A2(n_257_76_5943), .ZN(
      n_257_76_6114));
   NOR2_X1 i_257_76_6125 (.A1(n_257_76_6113), .A2(n_257_76_6114), .ZN(
      n_257_76_6115));
   NAND3_X1 i_257_76_6126 (.A1(n_257_76_6115), .A2(n_257_76_5946), .A3(
      n_257_76_5905), .ZN(n_257_76_6116));
   NOR2_X1 i_257_76_6127 (.A1(n_257_76_6116), .A2(n_257_76_6021), .ZN(
      n_257_76_6117));
   NAND2_X1 i_257_76_6128 (.A1(n_257_68), .A2(n_257_76_6117), .ZN(n_257_76_6118));
   NAND3_X1 i_257_76_6129 (.A1(n_257_76_6087), .A2(n_257_76_6101), .A3(
      n_257_76_6118), .ZN(n_257_76_6119));
   NOR2_X1 i_257_76_6130 (.A1(n_257_1069), .A2(n_257_76_17951), .ZN(
      n_257_76_6120));
   NAND2_X1 i_257_76_6131 (.A1(n_257_76_5927), .A2(n_257_76_6120), .ZN(
      n_257_76_6121));
   INV_X1 i_257_76_6132 (.A(n_257_76_6121), .ZN(n_257_76_6122));
   NAND3_X1 i_257_76_6133 (.A1(n_257_76_6122), .A2(n_257_76_5935), .A3(
      n_257_76_5932), .ZN(n_257_76_6123));
   INV_X1 i_257_76_6134 (.A(n_257_76_6123), .ZN(n_257_76_6124));
   NAND4_X1 i_257_76_6135 (.A1(n_257_76_6090), .A2(n_257_76_5938), .A3(n_257_807), 
      .A4(n_257_76_6124), .ZN(n_257_76_6125));
   INV_X1 i_257_76_6136 (.A(n_257_76_6125), .ZN(n_257_76_6126));
   NAND2_X1 i_257_76_6137 (.A1(n_257_76_5905), .A2(n_257_76_6126), .ZN(
      n_257_76_6127));
   INV_X1 i_257_76_6138 (.A(n_257_76_6127), .ZN(n_257_76_6128));
   NAND2_X1 i_257_76_6139 (.A1(n_257_76_5904), .A2(n_257_76_6128), .ZN(
      n_257_76_6129));
   INV_X1 i_257_76_6140 (.A(n_257_76_6129), .ZN(n_257_76_6130));
   NAND2_X1 i_257_76_6141 (.A1(n_257_22), .A2(n_257_76_6130), .ZN(n_257_76_6131));
   NAND2_X1 i_257_76_6142 (.A1(n_257_444), .A2(n_257_76_5919), .ZN(n_257_76_6132));
   INV_X1 i_257_76_6143 (.A(n_257_76_6132), .ZN(n_257_76_6133));
   NAND2_X1 i_257_76_6144 (.A1(n_257_1005), .A2(n_257_76_6133), .ZN(
      n_257_76_6134));
   INV_X1 i_257_76_6145 (.A(n_257_76_6134), .ZN(n_257_76_6135));
   NAND2_X1 i_257_76_6146 (.A1(n_257_76_5904), .A2(n_257_76_6135), .ZN(
      n_257_76_6136));
   INV_X1 i_257_76_6147 (.A(n_257_76_6136), .ZN(n_257_76_6137));
   NAND2_X1 i_257_76_6148 (.A1(n_257_76_18075), .A2(n_257_76_6137), .ZN(
      n_257_76_6138));
   NAND2_X1 i_257_76_6149 (.A1(n_257_76_6131), .A2(n_257_76_6138), .ZN(
      n_257_76_6139));
   NOR2_X1 i_257_76_6150 (.A1(n_257_76_6119), .A2(n_257_76_6139), .ZN(
      n_257_76_6140));
   NAND3_X1 i_257_76_6151 (.A1(n_257_76_6013), .A2(n_257_76_6067), .A3(
      n_257_76_6140), .ZN(n_257_76_6141));
   INV_X1 i_257_76_6152 (.A(n_257_76_6141), .ZN(n_257_76_6142));
   NOR2_X1 i_257_76_6153 (.A1(n_257_1069), .A2(n_257_76_17633), .ZN(
      n_257_76_6143));
   NAND4_X1 i_257_76_6154 (.A1(n_257_76_5979), .A2(n_257_76_5932), .A3(
      n_257_76_5927), .A4(n_257_76_6143), .ZN(n_257_76_6144));
   INV_X1 i_257_76_6155 (.A(n_257_76_6144), .ZN(n_257_76_6145));
   NAND2_X1 i_257_76_6156 (.A1(n_257_76_5935), .A2(n_257_76_5930), .ZN(
      n_257_76_6146));
   INV_X1 i_257_76_6157 (.A(n_257_76_6146), .ZN(n_257_76_6147));
   NAND2_X1 i_257_76_6158 (.A1(n_257_76_5931), .A2(n_257_45), .ZN(n_257_76_6148));
   INV_X1 i_257_76_6159 (.A(n_257_76_6148), .ZN(n_257_76_6149));
   NAND3_X1 i_257_76_6160 (.A1(n_257_76_6145), .A2(n_257_76_6147), .A3(
      n_257_76_6149), .ZN(n_257_76_6150));
   NAND3_X1 i_257_76_6161 (.A1(n_257_76_5939), .A2(n_257_76_5906), .A3(
      n_257_76_5934), .ZN(n_257_76_6151));
   NOR2_X1 i_257_76_6162 (.A1(n_257_76_6150), .A2(n_257_76_6151), .ZN(
      n_257_76_6152));
   NAND2_X1 i_257_76_6163 (.A1(n_257_76_5938), .A2(n_257_76_6004), .ZN(
      n_257_76_6153));
   INV_X1 i_257_76_6164 (.A(n_257_76_6153), .ZN(n_257_76_6154));
   NAND4_X1 i_257_76_6165 (.A1(n_257_76_6152), .A2(n_257_76_6154), .A3(
      n_257_76_5942), .A4(n_257_76_5943), .ZN(n_257_76_6155));
   INV_X1 i_257_76_6166 (.A(n_257_76_6155), .ZN(n_257_76_6156));
   NAND3_X1 i_257_76_6167 (.A1(n_257_76_6156), .A2(n_257_76_5946), .A3(
      n_257_76_5905), .ZN(n_257_76_6157));
   NOR2_X1 i_257_76_6168 (.A1(n_257_76_6157), .A2(n_257_76_6021), .ZN(
      n_257_76_6158));
   NAND2_X1 i_257_76_6169 (.A1(n_257_76_18081), .A2(n_257_76_6158), .ZN(
      n_257_76_6159));
   NAND2_X1 i_257_76_6170 (.A1(n_257_449), .A2(n_257_76_5919), .ZN(n_257_76_6160));
   INV_X1 i_257_76_6171 (.A(n_257_76_6160), .ZN(n_257_76_6161));
   NAND2_X1 i_257_76_6172 (.A1(n_257_76_5927), .A2(n_257_1083), .ZN(
      n_257_76_6162));
   INV_X1 i_257_76_6173 (.A(n_257_76_6162), .ZN(n_257_76_6163));
   NAND4_X1 i_257_76_6174 (.A1(n_257_76_6161), .A2(n_257_76_5931), .A3(
      n_257_76_5932), .A4(n_257_76_6163), .ZN(n_257_76_6164));
   NOR2_X1 i_257_76_6175 (.A1(n_257_76_6164), .A2(n_257_76_5936), .ZN(
      n_257_76_6165));
   NAND4_X1 i_257_76_6176 (.A1(n_257_76_6165), .A2(n_257_76_5941), .A3(
      n_257_76_5942), .A4(n_257_76_5943), .ZN(n_257_76_6166));
   NOR2_X1 i_257_76_6177 (.A1(n_257_76_5925), .A2(n_257_76_6166), .ZN(
      n_257_76_6167));
   NAND3_X1 i_257_76_6178 (.A1(n_257_76_6167), .A2(n_257_76_5904), .A3(
      n_257_76_5946), .ZN(n_257_76_6168));
   INV_X1 i_257_76_6179 (.A(n_257_76_6168), .ZN(n_257_76_6169));
   NAND2_X1 i_257_76_6180 (.A1(n_257_76_18083), .A2(n_257_76_6169), .ZN(
      n_257_76_6170));
   INV_X1 i_257_76_6181 (.A(n_257_607), .ZN(n_257_76_6171));
   NAND2_X1 i_257_76_6182 (.A1(n_257_76_6171), .A2(n_257_442), .ZN(n_257_76_6172));
   OAI21_X1 i_257_76_6183 (.A(n_257_76_6172), .B1(n_257_432), .B2(n_257_76_17412), 
      .ZN(n_257_76_6173));
   NAND3_X1 i_257_76_6184 (.A1(n_257_76_5907), .A2(n_257_76_6173), .A3(n_257_429), 
      .ZN(n_257_76_6174));
   INV_X1 i_257_76_6185 (.A(n_257_76_5927), .ZN(n_257_76_6175));
   NOR2_X1 i_257_76_6186 (.A1(n_257_76_6174), .A2(n_257_76_6175), .ZN(
      n_257_76_6176));
   NAND4_X1 i_257_76_6187 (.A1(n_257_76_6176), .A2(n_257_76_5931), .A3(
      n_257_76_5979), .A4(n_257_76_5932), .ZN(n_257_76_6177));
   NAND3_X1 i_257_76_6188 (.A1(n_257_76_5934), .A2(n_257_76_5935), .A3(
      n_257_76_5930), .ZN(n_257_76_6178));
   NOR2_X1 i_257_76_6189 (.A1(n_257_76_6177), .A2(n_257_76_6178), .ZN(
      n_257_76_6179));
   NAND2_X1 i_257_76_6190 (.A1(n_257_76_6004), .A2(n_257_76_5992), .ZN(
      n_257_76_6180));
   INV_X1 i_257_76_6191 (.A(n_257_76_6180), .ZN(n_257_76_6181));
   NAND3_X1 i_257_76_6192 (.A1(n_257_76_5939), .A2(n_257_76_5973), .A3(
      n_257_76_5906), .ZN(n_257_76_6182));
   INV_X1 i_257_76_6193 (.A(n_257_76_6182), .ZN(n_257_76_6183));
   NAND4_X1 i_257_76_6194 (.A1(n_257_76_6179), .A2(n_257_76_6181), .A3(
      n_257_76_5938), .A4(n_257_76_6183), .ZN(n_257_76_6184));
   NAND4_X1 i_257_76_6195 (.A1(n_257_76_5942), .A2(n_257_76_6003), .A3(n_257_162), 
      .A4(n_257_76_5943), .ZN(n_257_76_6185));
   NOR2_X1 i_257_76_6196 (.A1(n_257_76_6184), .A2(n_257_76_6185), .ZN(
      n_257_76_6186));
   NAND3_X1 i_257_76_6197 (.A1(n_257_76_6186), .A2(n_257_76_5946), .A3(
      n_257_76_5905), .ZN(n_257_76_6187));
   NOR2_X1 i_257_76_6198 (.A1(n_257_76_6187), .A2(n_257_76_6021), .ZN(
      n_257_76_6188));
   NAND2_X1 i_257_76_6199 (.A1(n_257_76_18061), .A2(n_257_76_6188), .ZN(
      n_257_76_6189));
   NAND3_X1 i_257_76_6200 (.A1(n_257_76_6159), .A2(n_257_76_6170), .A3(
      n_257_76_6189), .ZN(n_257_76_6190));
   INV_X1 i_257_76_6201 (.A(n_257_76_6190), .ZN(n_257_76_6191));
   NAND4_X1 i_257_76_6202 (.A1(n_257_76_5919), .A2(n_257_76_5927), .A3(
      n_257_1075), .A4(n_257_438), .ZN(n_257_76_6192));
   INV_X1 i_257_76_6203 (.A(n_257_76_6192), .ZN(n_257_76_6193));
   NAND3_X1 i_257_76_6204 (.A1(n_257_76_5939), .A2(n_257_76_5906), .A3(
      n_257_76_6193), .ZN(n_257_76_6194));
   INV_X1 i_257_76_6205 (.A(n_257_76_6194), .ZN(n_257_76_6195));
   NAND2_X1 i_257_76_6206 (.A1(n_257_76_5905), .A2(n_257_76_6195), .ZN(
      n_257_76_6196));
   INV_X1 i_257_76_6207 (.A(n_257_76_6196), .ZN(n_257_76_6197));
   NAND2_X1 i_257_76_6208 (.A1(n_257_76_5904), .A2(n_257_76_6197), .ZN(
      n_257_76_6198));
   INV_X1 i_257_76_6209 (.A(n_257_76_6198), .ZN(n_257_76_6199));
   NAND2_X1 i_257_76_6210 (.A1(n_257_76_18067), .A2(n_257_76_6199), .ZN(
      n_257_76_6200));
   NAND2_X1 i_257_76_6211 (.A1(n_257_359), .A2(n_257_421), .ZN(n_257_76_6201));
   NAND3_X1 i_257_76_6212 (.A1(n_257_76_5999), .A2(n_257_76_6000), .A3(
      n_257_76_6201), .ZN(n_257_76_6202));
   INV_X1 i_257_76_6213 (.A(n_257_76_6202), .ZN(n_257_76_6203));
   NAND4_X1 i_257_76_6214 (.A1(n_257_76_5942), .A2(n_257_76_6003), .A3(
      n_257_76_5943), .A4(n_257_76_5938), .ZN(n_257_76_6204));
   INV_X1 i_257_76_6215 (.A(n_257_76_6204), .ZN(n_257_76_6205));
   NAND2_X1 i_257_76_6216 (.A1(n_257_282), .A2(n_257_423), .ZN(n_257_76_6206));
   NAND2_X1 i_257_76_6217 (.A1(n_257_76_6206), .A2(n_257_76_5939), .ZN(
      n_257_76_6207));
   NOR2_X1 i_257_76_6218 (.A1(n_257_76_6207), .A2(n_257_76_5975), .ZN(
      n_257_76_6208));
   NAND2_X1 i_257_76_6219 (.A1(n_257_76_15125), .A2(n_257_76_5984), .ZN(
      n_257_76_6209));
   OAI21_X1 i_257_76_6220 (.A(n_257_76_6209), .B1(n_257_428), .B2(n_257_76_14977), 
      .ZN(n_257_76_6210));
   NAND4_X1 i_257_76_6221 (.A1(n_257_76_5907), .A2(n_257_76_6210), .A3(n_257_420), 
      .A4(n_257_76_5981), .ZN(n_257_76_6211));
   INV_X1 i_257_76_6222 (.A(n_257_76_6211), .ZN(n_257_76_6212));
   NAND3_X1 i_257_76_6223 (.A1(n_257_76_6212), .A2(n_257_76_5978), .A3(
      n_257_76_5989), .ZN(n_257_76_6213));
   INV_X1 i_257_76_6224 (.A(n_257_76_6213), .ZN(n_257_76_6214));
   NAND3_X1 i_257_76_6225 (.A1(n_257_76_6004), .A2(n_257_76_5992), .A3(
      n_257_76_6214), .ZN(n_257_76_6215));
   INV_X1 i_257_76_6226 (.A(n_257_76_6215), .ZN(n_257_76_6216));
   NAND4_X1 i_257_76_6227 (.A1(n_257_76_5934), .A2(n_257_76_5935), .A3(
      n_257_76_5930), .A4(n_257_76_5931), .ZN(n_257_76_6217));
   NAND2_X1 i_257_76_6228 (.A1(n_257_320), .A2(n_257_422), .ZN(n_257_76_6218));
   NAND4_X1 i_257_76_6229 (.A1(n_257_76_6218), .A2(n_257_76_5979), .A3(
      n_257_76_5932), .A4(n_257_76_5927), .ZN(n_257_76_6219));
   NOR2_X1 i_257_76_6230 (.A1(n_257_76_6217), .A2(n_257_76_6219), .ZN(
      n_257_76_6220));
   NAND3_X1 i_257_76_6231 (.A1(n_257_76_6208), .A2(n_257_76_6216), .A3(
      n_257_76_6220), .ZN(n_257_76_6221));
   INV_X1 i_257_76_6232 (.A(n_257_76_6221), .ZN(n_257_76_6222));
   NAND3_X1 i_257_76_6233 (.A1(n_257_76_6203), .A2(n_257_76_6205), .A3(
      n_257_76_6222), .ZN(n_257_76_6223));
   INV_X1 i_257_76_6234 (.A(n_257_76_6223), .ZN(n_257_76_6224));
   NAND2_X1 i_257_76_6235 (.A1(n_257_76_5946), .A2(n_257_76_5905), .ZN(
      n_257_76_6225));
   INV_X1 i_257_76_6236 (.A(n_257_76_6225), .ZN(n_257_76_6226));
   NAND3_X1 i_257_76_6237 (.A1(n_257_76_6224), .A2(n_257_76_6226), .A3(
      n_257_76_5904), .ZN(n_257_76_6227));
   INV_X1 i_257_76_6238 (.A(n_257_76_6227), .ZN(n_257_76_6228));
   NAND2_X1 i_257_76_6239 (.A1(n_257_76_18073), .A2(n_257_76_6228), .ZN(
      n_257_76_6229));
   NAND3_X1 i_257_76_6240 (.A1(n_257_76_5907), .A2(n_257_76_6173), .A3(n_257_430), 
      .ZN(n_257_76_6230));
   INV_X1 i_257_76_6241 (.A(n_257_76_6230), .ZN(n_257_76_6231));
   NAND4_X1 i_257_76_6242 (.A1(n_257_76_6231), .A2(n_257_76_5979), .A3(
      n_257_76_5932), .A4(n_257_76_5927), .ZN(n_257_76_6232));
   NOR2_X1 i_257_76_6243 (.A1(n_257_76_6033), .A2(n_257_76_6232), .ZN(
      n_257_76_6233));
   NAND4_X1 i_257_76_6244 (.A1(n_257_123), .A2(n_257_76_5973), .A3(n_257_76_5906), 
      .A4(n_257_76_5934), .ZN(n_257_76_6234));
   INV_X1 i_257_76_6245 (.A(n_257_76_6234), .ZN(n_257_76_6235));
   NAND4_X1 i_257_76_6246 (.A1(n_257_76_6103), .A2(n_257_76_6233), .A3(
      n_257_76_6235), .A4(n_257_76_5938), .ZN(n_257_76_6236));
   NAND3_X1 i_257_76_6247 (.A1(n_257_76_5942), .A2(n_257_76_6003), .A3(
      n_257_76_5943), .ZN(n_257_76_6237));
   NOR2_X1 i_257_76_6248 (.A1(n_257_76_6236), .A2(n_257_76_6237), .ZN(
      n_257_76_6238));
   NAND3_X1 i_257_76_6249 (.A1(n_257_76_6238), .A2(n_257_76_5946), .A3(
      n_257_76_5905), .ZN(n_257_76_6239));
   NOR2_X1 i_257_76_6250 (.A1(n_257_76_6239), .A2(n_257_76_6021), .ZN(
      n_257_76_6240));
   NAND2_X1 i_257_76_6251 (.A1(n_257_76_18068), .A2(n_257_76_6240), .ZN(
      n_257_76_6241));
   NAND3_X1 i_257_76_6252 (.A1(n_257_76_6200), .A2(n_257_76_6229), .A3(
      n_257_76_6241), .ZN(n_257_76_6242));
   INV_X1 i_257_76_6253 (.A(n_257_76_6242), .ZN(n_257_76_6243));
   NAND2_X1 i_257_76_6254 (.A1(n_257_775), .A2(n_257_442), .ZN(n_257_76_6244));
   NOR2_X1 i_257_76_6255 (.A1(n_257_1069), .A2(n_257_76_6244), .ZN(n_257_76_6245));
   NAND4_X1 i_257_76_6256 (.A1(n_257_76_5932), .A2(n_257_76_6245), .A3(n_257_447), 
      .A4(n_257_76_5927), .ZN(n_257_76_6246));
   INV_X1 i_257_76_6257 (.A(n_257_76_6246), .ZN(n_257_76_6247));
   NAND4_X1 i_257_76_6258 (.A1(n_257_76_5939), .A2(n_257_76_6247), .A3(
      n_257_76_5906), .A4(n_257_76_5935), .ZN(n_257_76_6248));
   INV_X1 i_257_76_6259 (.A(n_257_76_6248), .ZN(n_257_76_6249));
   NAND3_X1 i_257_76_6260 (.A1(n_257_76_6249), .A2(n_257_76_5943), .A3(
      n_257_76_5938), .ZN(n_257_76_6250));
   INV_X1 i_257_76_6261 (.A(n_257_76_6250), .ZN(n_257_76_6251));
   NAND2_X1 i_257_76_6262 (.A1(n_257_76_5905), .A2(n_257_76_6251), .ZN(
      n_257_76_6252));
   INV_X1 i_257_76_6263 (.A(n_257_76_6252), .ZN(n_257_76_6253));
   NAND2_X1 i_257_76_6264 (.A1(n_257_76_5904), .A2(n_257_76_6253), .ZN(
      n_257_76_6254));
   INV_X1 i_257_76_6265 (.A(n_257_76_6254), .ZN(n_257_76_6255));
   NAND3_X1 i_257_76_6266 (.A1(n_257_76_5907), .A2(n_257_76_6173), .A3(n_257_431), 
      .ZN(n_257_76_6256));
   INV_X1 i_257_76_6267 (.A(n_257_76_6256), .ZN(n_257_76_6257));
   NAND4_X1 i_257_76_6268 (.A1(n_257_76_6257), .A2(n_257_76_5979), .A3(
      n_257_76_5932), .A4(n_257_76_5927), .ZN(n_257_76_6258));
   NOR2_X1 i_257_76_6269 (.A1(n_257_76_6258), .A2(n_257_76_6111), .ZN(
      n_257_76_6259));
   NAND4_X1 i_257_76_6270 (.A1(n_257_76_6103), .A2(n_257_76_6105), .A3(
      n_257_76_6259), .A4(n_257_85), .ZN(n_257_76_6260));
   NAND3_X1 i_257_76_6271 (.A1(n_257_76_5942), .A2(n_257_76_5943), .A3(
      n_257_76_5938), .ZN(n_257_76_6261));
   NOR2_X1 i_257_76_6272 (.A1(n_257_76_6260), .A2(n_257_76_6261), .ZN(
      n_257_76_6262));
   NAND3_X1 i_257_76_6273 (.A1(n_257_76_6262), .A2(n_257_76_5946), .A3(
      n_257_76_5905), .ZN(n_257_76_6263));
   NOR2_X1 i_257_76_6274 (.A1(n_257_76_6263), .A2(n_257_76_6021), .ZN(
      n_257_76_6264));
   AOI22_X1 i_257_76_6275 (.A1(n_257_76_18085), .A2(n_257_76_6255), .B1(
      n_257_76_18080), .B2(n_257_76_6264), .ZN(n_257_76_6265));
   NAND3_X1 i_257_76_6276 (.A1(n_257_76_6191), .A2(n_257_76_6243), .A3(
      n_257_76_6265), .ZN(n_257_76_6266));
   NAND2_X1 i_257_76_6277 (.A1(n_257_76_5939), .A2(n_257_76_5973), .ZN(
      n_257_76_6267));
   INV_X1 i_257_76_6278 (.A(n_257_76_6267), .ZN(n_257_76_6268));
   NAND2_X1 i_257_76_6279 (.A1(n_257_76_5981), .A2(n_257_421), .ZN(n_257_76_6269));
   INV_X1 i_257_76_6280 (.A(n_257_76_6269), .ZN(n_257_76_6270));
   NAND4_X1 i_257_76_6281 (.A1(n_257_76_5989), .A2(n_257_76_6074), .A3(
      n_257_76_5927), .A4(n_257_76_6270), .ZN(n_257_76_6271));
   NAND3_X1 i_257_76_6282 (.A1(n_257_76_5978), .A2(n_257_76_5979), .A3(
      n_257_76_5932), .ZN(n_257_76_6272));
   NOR2_X1 i_257_76_6283 (.A1(n_257_76_6271), .A2(n_257_76_6272), .ZN(
      n_257_76_6273));
   NAND3_X1 i_257_76_6284 (.A1(n_257_76_5974), .A2(n_257_76_5906), .A3(
      n_257_76_5934), .ZN(n_257_76_6274));
   INV_X1 i_257_76_6285 (.A(n_257_76_6274), .ZN(n_257_76_6275));
   NAND4_X1 i_257_76_6286 (.A1(n_257_76_5935), .A2(n_257_76_5930), .A3(
      n_257_76_5931), .A4(n_257_76_6218), .ZN(n_257_76_6276));
   INV_X1 i_257_76_6287 (.A(n_257_76_6276), .ZN(n_257_76_6277));
   NAND4_X1 i_257_76_6288 (.A1(n_257_76_6268), .A2(n_257_76_6273), .A3(
      n_257_76_6275), .A4(n_257_76_6277), .ZN(n_257_76_6278));
   NAND4_X1 i_257_76_6289 (.A1(n_257_76_5938), .A2(n_257_76_6004), .A3(
      n_257_76_5992), .A4(n_257_76_6206), .ZN(n_257_76_6279));
   NOR2_X1 i_257_76_6290 (.A1(n_257_76_6278), .A2(n_257_76_6279), .ZN(
      n_257_76_6280));
   NAND4_X1 i_257_76_6291 (.A1(n_257_76_5942), .A2(n_257_76_6003), .A3(
      n_257_76_5943), .A4(n_257_359), .ZN(n_257_76_6281));
   INV_X1 i_257_76_6292 (.A(n_257_76_6281), .ZN(n_257_76_6282));
   NAND3_X1 i_257_76_6293 (.A1(n_257_76_6280), .A2(n_257_76_6002), .A3(
      n_257_76_6282), .ZN(n_257_76_6283));
   NOR3_X1 i_257_76_6294 (.A1(n_257_76_6021), .A2(n_257_76_6283), .A3(
      n_257_76_6225), .ZN(n_257_76_6284));
   NAND2_X1 i_257_76_6295 (.A1(n_257_76_18082), .A2(n_257_76_6284), .ZN(
      n_257_76_6285));
   NAND3_X1 i_257_76_6296 (.A1(n_257_76_5979), .A2(n_257_76_5932), .A3(
      n_257_76_5927), .ZN(n_257_76_6286));
   NOR2_X1 i_257_76_6297 (.A1(n_257_76_6033), .A2(n_257_76_6286), .ZN(
      n_257_76_6287));
   NAND2_X1 i_257_76_6298 (.A1(n_257_427), .A2(n_257_76_5981), .ZN(n_257_76_6288));
   INV_X1 i_257_76_6299 (.A(n_257_76_6288), .ZN(n_257_76_6289));
   NAND4_X1 i_257_76_6300 (.A1(n_257_202), .A2(n_257_76_6289), .A3(n_257_76_5907), 
      .A4(n_257_76_5986), .ZN(n_257_76_6290));
   INV_X1 i_257_76_6301 (.A(n_257_76_6290), .ZN(n_257_76_6291));
   NAND4_X1 i_257_76_6302 (.A1(n_257_76_5973), .A2(n_257_76_5906), .A3(
      n_257_76_6291), .A4(n_257_76_5934), .ZN(n_257_76_6292));
   INV_X1 i_257_76_6303 (.A(n_257_76_6292), .ZN(n_257_76_6293));
   NAND3_X1 i_257_76_6304 (.A1(n_257_76_5994), .A2(n_257_76_6287), .A3(
      n_257_76_6293), .ZN(n_257_76_6294));
   NOR2_X1 i_257_76_6305 (.A1(n_257_76_6045), .A2(n_257_76_6294), .ZN(
      n_257_76_6295));
   NAND4_X1 i_257_76_6306 (.A1(n_257_76_6295), .A2(n_257_76_5946), .A3(
      n_257_76_5905), .A4(n_257_76_6048), .ZN(n_257_76_6296));
   NOR2_X1 i_257_76_6307 (.A1(n_257_76_6296), .A2(n_257_76_6021), .ZN(
      n_257_76_6297));
   NAND2_X1 i_257_76_6308 (.A1(n_257_76_18065), .A2(n_257_76_6297), .ZN(
      n_257_76_6298));
   NAND3_X1 i_257_76_6309 (.A1(n_257_76_5919), .A2(n_257_76_5927), .A3(n_257_462), 
      .ZN(n_257_76_6299));
   INV_X1 i_257_76_6310 (.A(n_257_76_6299), .ZN(n_257_76_6300));
   NAND4_X1 i_257_76_6311 (.A1(n_257_76_6300), .A2(n_257_76_5931), .A3(
      n_257_76_5979), .A4(n_257_76_5932), .ZN(n_257_76_6301));
   NOR2_X1 i_257_76_6312 (.A1(n_257_76_6301), .A2(n_257_76_6178), .ZN(
      n_257_76_6302));
   NAND3_X1 i_257_76_6313 (.A1(n_257_76_5939), .A2(n_257_451), .A3(n_257_76_5906), 
      .ZN(n_257_76_6303));
   INV_X1 i_257_76_6314 (.A(n_257_76_6303), .ZN(n_257_76_6304));
   NAND3_X1 i_257_76_6315 (.A1(n_257_76_6302), .A2(n_257_76_6304), .A3(
      n_257_76_5938), .ZN(n_257_76_6305));
   NOR2_X1 i_257_76_6316 (.A1(n_257_76_6305), .A2(n_257_76_6114), .ZN(
      n_257_76_6306));
   NAND2_X1 i_257_76_6317 (.A1(n_257_76_5905), .A2(n_257_76_6306), .ZN(
      n_257_76_6307));
   INV_X1 i_257_76_6318 (.A(n_257_76_6307), .ZN(n_257_76_6308));
   NAND3_X1 i_257_76_6319 (.A1(n_257_76_6308), .A2(n_257_76_5904), .A3(
      n_257_76_5946), .ZN(n_257_76_6309));
   INV_X1 i_257_76_6320 (.A(n_257_76_6309), .ZN(n_257_76_6310));
   NAND2_X1 i_257_76_6321 (.A1(n_257_76_18063), .A2(n_257_76_6310), .ZN(
      n_257_76_6311));
   NAND3_X1 i_257_76_6322 (.A1(n_257_76_6285), .A2(n_257_76_6298), .A3(
      n_257_76_6311), .ZN(n_257_76_6312));
   INV_X1 i_257_76_6323 (.A(n_257_76_6312), .ZN(n_257_76_6313));
   NAND2_X1 i_257_76_6324 (.A1(n_257_76_5932), .A2(n_257_76_5927), .ZN(
      n_257_76_6314));
   INV_X1 i_257_76_6325 (.A(n_257_76_6314), .ZN(n_257_76_6315));
   NAND4_X1 i_257_76_6326 (.A1(n_257_76_6315), .A2(n_257_76_5930), .A3(
      n_257_76_5931), .A4(n_257_76_5979), .ZN(n_257_76_6316));
   NOR2_X1 i_257_76_6327 (.A1(n_257_76_6316), .A2(n_257_76_5936), .ZN(
      n_257_76_6317));
   NAND2_X1 i_257_76_6328 (.A1(n_257_511), .A2(n_257_76_5907), .ZN(n_257_76_6318));
   INV_X1 i_257_76_6329 (.A(n_257_76_6318), .ZN(n_257_76_6319));
   NAND3_X1 i_257_76_6330 (.A1(n_257_76_5986), .A2(n_257_76_5981), .A3(n_257_424), 
      .ZN(n_257_76_6320));
   INV_X1 i_257_76_6331 (.A(n_257_76_6320), .ZN(n_257_76_6321));
   NAND3_X1 i_257_76_6332 (.A1(n_257_76_5978), .A2(n_257_76_6319), .A3(
      n_257_76_6321), .ZN(n_257_76_6322));
   INV_X1 i_257_76_6333 (.A(n_257_76_6322), .ZN(n_257_76_6323));
   NAND4_X1 i_257_76_6334 (.A1(n_257_76_5939), .A2(n_257_76_6323), .A3(
      n_257_76_5973), .A4(n_257_76_5974), .ZN(n_257_76_6324));
   INV_X1 i_257_76_6335 (.A(n_257_76_6324), .ZN(n_257_76_6325));
   NAND3_X1 i_257_76_6336 (.A1(n_257_76_6317), .A2(n_257_76_6181), .A3(
      n_257_76_6325), .ZN(n_257_76_6326));
   NAND3_X1 i_257_76_6337 (.A1(n_257_76_6003), .A2(n_257_76_5943), .A3(
      n_257_76_5938), .ZN(n_257_76_6327));
   NOR2_X1 i_257_76_6338 (.A1(n_257_76_6326), .A2(n_257_76_6327), .ZN(
      n_257_76_6328));
   NAND3_X1 i_257_76_6339 (.A1(n_257_76_5999), .A2(n_257_76_6000), .A3(
      n_257_76_5942), .ZN(n_257_76_6329));
   INV_X1 i_257_76_6340 (.A(n_257_76_6329), .ZN(n_257_76_6330));
   NAND4_X1 i_257_76_6341 (.A1(n_257_76_6328), .A2(n_257_76_5946), .A3(
      n_257_76_5905), .A4(n_257_76_6330), .ZN(n_257_76_6331));
   NOR2_X1 i_257_76_6342 (.A1(n_257_76_6331), .A2(n_257_76_6021), .ZN(
      n_257_76_6332));
   NAND2_X1 i_257_76_6343 (.A1(n_257_76_18062), .A2(n_257_76_6332), .ZN(
      n_257_76_6333));
   INV_X1 i_257_76_6344 (.A(n_257_76_6207), .ZN(n_257_76_6334));
   NAND4_X1 i_257_76_6345 (.A1(n_257_76_6181), .A2(n_257_76_6334), .A3(
      n_257_76_6069), .A4(n_257_76_5938), .ZN(n_257_76_6335));
   NOR2_X1 i_257_76_6346 (.A1(n_257_76_6237), .A2(n_257_76_6335), .ZN(
      n_257_76_6336));
   NAND3_X1 i_257_76_6347 (.A1(n_257_76_5979), .A2(n_257_76_5932), .A3(
      n_257_76_5989), .ZN(n_257_76_6337));
   NAND2_X1 i_257_76_6348 (.A1(n_257_422), .A2(n_257_76_5981), .ZN(n_257_76_6338));
   INV_X1 i_257_76_6349 (.A(n_257_76_6338), .ZN(n_257_76_6339));
   NAND4_X1 i_257_76_6350 (.A1(n_257_76_6074), .A2(n_257_320), .A3(n_257_76_5927), 
      .A4(n_257_76_6339), .ZN(n_257_76_6340));
   NOR2_X1 i_257_76_6351 (.A1(n_257_76_6337), .A2(n_257_76_6340), .ZN(
      n_257_76_6341));
   NAND2_X1 i_257_76_6352 (.A1(n_257_76_5973), .A2(n_257_76_5974), .ZN(
      n_257_76_6342));
   INV_X1 i_257_76_6353 (.A(n_257_76_6342), .ZN(n_257_76_6343));
   NAND2_X1 i_257_76_6354 (.A1(n_257_76_5934), .A2(n_257_76_5978), .ZN(
      n_257_76_6344));
   INV_X1 i_257_76_6355 (.A(n_257_76_6344), .ZN(n_257_76_6345));
   NAND3_X1 i_257_76_6356 (.A1(n_257_76_6341), .A2(n_257_76_6343), .A3(
      n_257_76_6345), .ZN(n_257_76_6346));
   INV_X1 i_257_76_6357 (.A(n_257_76_6346), .ZN(n_257_76_6347));
   NAND3_X1 i_257_76_6358 (.A1(n_257_76_6347), .A2(n_257_76_5999), .A3(
      n_257_76_6000), .ZN(n_257_76_6348));
   INV_X1 i_257_76_6359 (.A(n_257_76_6348), .ZN(n_257_76_6349));
   NAND4_X1 i_257_76_6360 (.A1(n_257_76_5946), .A2(n_257_76_6336), .A3(
      n_257_76_6349), .A4(n_257_76_5905), .ZN(n_257_76_6350));
   NOR2_X1 i_257_76_6361 (.A1(n_257_76_6350), .A2(n_257_76_6021), .ZN(
      n_257_76_6351));
   NAND2_X1 i_257_76_6362 (.A1(n_257_342), .A2(n_257_76_6351), .ZN(n_257_76_6352));
   NAND2_X1 i_257_76_6363 (.A1(n_257_462), .A2(n_257_442), .ZN(n_257_76_6353));
   INV_X1 i_257_76_6364 (.A(n_257_76_6353), .ZN(n_257_76_6354));
   NAND2_X1 i_257_76_6365 (.A1(n_257_451), .A2(n_257_76_6354), .ZN(n_257_76_6355));
   NAND2_X1 i_257_76_6366 (.A1(n_257_123), .A2(n_257_76_17925), .ZN(
      n_257_76_6356));
   NAND2_X1 i_257_76_6367 (.A1(n_257_909), .A2(n_257_76_17940), .ZN(
      n_257_76_6357));
   NAND3_X1 i_257_76_6368 (.A1(n_257_76_6355), .A2(n_257_76_6356), .A3(
      n_257_76_6357), .ZN(n_257_76_6358));
   INV_X1 i_257_76_6369 (.A(n_257_76_6358), .ZN(n_257_76_6359));
   NAND2_X1 i_257_76_6370 (.A1(n_257_45), .A2(n_257_76_17918), .ZN(n_257_76_6360));
   NAND2_X1 i_257_76_6371 (.A1(n_257_973), .A2(n_257_442), .ZN(n_257_76_6361));
   INV_X1 i_257_76_6372 (.A(n_257_76_6361), .ZN(n_257_76_6362));
   NAND2_X1 i_257_76_6373 (.A1(n_257_441), .A2(n_257_76_6362), .ZN(n_257_76_6363));
   NAND2_X1 i_257_76_6374 (.A1(n_257_711), .A2(n_257_76_15655), .ZN(
      n_257_76_6364));
   NAND3_X1 i_257_76_6375 (.A1(n_257_76_6360), .A2(n_257_76_6363), .A3(
      n_257_76_6364), .ZN(n_257_76_6365));
   NAND2_X1 i_257_76_6376 (.A1(n_257_76_6213), .A2(n_257_76_6322), .ZN(
      n_257_76_6366));
   NOR2_X1 i_257_76_6377 (.A1(n_257_76_6365), .A2(n_257_76_6366), .ZN(
      n_257_76_6367));
   NAND2_X1 i_257_76_6378 (.A1(n_257_428), .A2(n_257_575), .ZN(n_257_76_6368));
   NAND2_X1 i_257_76_6379 (.A1(n_257_76_5981), .A2(n_257_76_6368), .ZN(
      n_257_76_6369));
   INV_X1 i_257_76_6380 (.A(n_257_76_6369), .ZN(n_257_76_6370));
   INV_X1 i_257_76_6381 (.A(Small_Packet_Data_Size[10]), .ZN(n_257_76_6371));
   NAND3_X1 i_257_76_6382 (.A1(n_257_76_6370), .A2(n_257_76_5907), .A3(
      n_257_76_18045), .ZN(n_257_76_6372));
   NAND2_X1 i_257_76_6383 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[10]), 
      .ZN(n_257_76_6373));
   NAND2_X1 i_257_76_6384 (.A1(n_257_76_6372), .A2(n_257_76_6373), .ZN(
      n_257_76_6374));
   NAND2_X1 i_257_76_6385 (.A1(n_257_76_13741), .A2(n_257_449), .ZN(
      n_257_76_6375));
   NAND2_X1 i_257_76_6386 (.A1(n_257_839), .A2(n_257_442), .ZN(n_257_76_6376));
   INV_X1 i_257_76_6387 (.A(n_257_76_6376), .ZN(n_257_76_6377));
   NAND2_X1 i_257_76_6388 (.A1(n_257_446), .A2(n_257_76_6377), .ZN(n_257_76_6378));
   NAND4_X1 i_257_76_6389 (.A1(n_257_76_6374), .A2(n_257_76_6375), .A3(
      n_257_76_6290), .A4(n_257_76_6378), .ZN(n_257_76_6379));
   INV_X1 i_257_76_6390 (.A(n_257_76_6244), .ZN(n_257_76_6380));
   NAND2_X1 i_257_76_6391 (.A1(n_257_447), .A2(n_257_76_6380), .ZN(n_257_76_6381));
   NAND3_X1 i_257_76_6392 (.A1(n_257_1075), .A2(n_257_438), .A3(n_257_442), 
      .ZN(n_257_76_6382));
   NAND2_X1 i_257_76_6393 (.A1(n_257_639), .A2(n_257_76_17928), .ZN(
      n_257_76_6383));
   NAND2_X1 i_257_76_6394 (.A1(n_257_440), .A2(n_257_76_5909), .ZN(n_257_76_6384));
   NAND4_X1 i_257_76_6395 (.A1(n_257_76_6381), .A2(n_257_76_6382), .A3(
      n_257_76_6383), .A4(n_257_76_6384), .ZN(n_257_76_6385));
   NOR2_X1 i_257_76_6396 (.A1(n_257_76_6379), .A2(n_257_76_6385), .ZN(
      n_257_76_6386));
   NAND3_X1 i_257_76_6397 (.A1(n_257_76_6359), .A2(n_257_76_6367), .A3(
      n_257_76_6386), .ZN(n_257_76_6387));
   NAND2_X1 i_257_76_6398 (.A1(n_257_807), .A2(n_257_76_17952), .ZN(
      n_257_76_6388));
   NAND2_X1 i_257_76_6399 (.A1(n_257_871), .A2(n_257_76_17903), .ZN(
      n_257_76_6389));
   NAND3_X1 i_257_76_6400 (.A1(n_257_76_6388), .A2(n_257_76_6081), .A3(
      n_257_76_6389), .ZN(n_257_76_6390));
   NOR2_X1 i_257_76_6401 (.A1(n_257_76_6387), .A2(n_257_76_6390), .ZN(
      n_257_76_6391));
   NAND2_X1 i_257_76_6402 (.A1(n_257_162), .A2(n_257_76_17331), .ZN(
      n_257_76_6392));
   NAND2_X1 i_257_76_6403 (.A1(n_257_743), .A2(n_257_76_17935), .ZN(
      n_257_76_6393));
   NAND2_X1 i_257_76_6404 (.A1(n_257_85), .A2(n_257_76_17932), .ZN(n_257_76_6394));
   NAND4_X1 i_257_76_6405 (.A1(n_257_76_6392), .A2(n_257_76_6346), .A3(
      n_257_76_6393), .A4(n_257_76_6394), .ZN(n_257_76_6395));
   INV_X1 i_257_76_6406 (.A(n_257_76_6395), .ZN(n_257_76_6396));
   NAND2_X1 i_257_76_6407 (.A1(n_257_1005), .A2(n_257_76_17964), .ZN(
      n_257_76_6397));
   NAND4_X1 i_257_76_6408 (.A1(n_257_76_6391), .A2(n_257_76_6396), .A3(
      n_257_76_6397), .A4(n_257_76_5995), .ZN(n_257_76_6398));
   NAND2_X1 i_257_76_6409 (.A1(n_257_1037), .A2(n_257_76_17969), .ZN(
      n_257_76_6399));
   NAND2_X1 i_257_76_6410 (.A1(n_257_76_6283), .A2(n_257_76_6399), .ZN(
      n_257_76_6400));
   NAND4_X1 i_257_76_6411 (.A1(n_257_76_5938), .A2(n_257_76_6004), .A3(
      n_257_76_5992), .A4(n_257_76_5939), .ZN(n_257_76_6401));
   INV_X1 i_257_76_6412 (.A(n_257_76_5975), .ZN(n_257_76_6402));
   INV_X1 i_257_76_6413 (.A(n_257_76_6217), .ZN(n_257_76_6403));
   NAND2_X1 i_257_76_6414 (.A1(n_257_76_5981), .A2(n_257_425), .ZN(n_257_76_6404));
   INV_X1 i_257_76_6415 (.A(n_257_76_6404), .ZN(n_257_76_6405));
   NAND3_X1 i_257_76_6416 (.A1(n_257_76_6074), .A2(n_257_76_5927), .A3(
      n_257_76_6405), .ZN(n_257_76_6406));
   NOR2_X1 i_257_76_6417 (.A1(n_257_76_6272), .A2(n_257_76_6406), .ZN(
      n_257_76_6407));
   NAND3_X1 i_257_76_6418 (.A1(n_257_76_6402), .A2(n_257_76_6403), .A3(
      n_257_76_6407), .ZN(n_257_76_6408));
   NOR2_X1 i_257_76_6419 (.A1(n_257_76_6401), .A2(n_257_76_6408), .ZN(
      n_257_76_6409));
   NAND2_X1 i_257_76_6420 (.A1(n_257_76_6000), .A2(n_257_76_5942), .ZN(
      n_257_76_6410));
   INV_X1 i_257_76_6421 (.A(n_257_76_6410), .ZN(n_257_76_6411));
   NAND3_X1 i_257_76_6422 (.A1(n_257_76_6003), .A2(n_257_242), .A3(n_257_76_5943), 
      .ZN(n_257_76_6412));
   INV_X1 i_257_76_6423 (.A(n_257_76_6412), .ZN(n_257_76_6413));
   NAND3_X1 i_257_76_6424 (.A1(n_257_76_6409), .A2(n_257_76_6411), .A3(
      n_257_76_6413), .ZN(n_257_76_6414));
   NAND2_X1 i_257_76_6425 (.A1(n_257_679), .A2(n_257_76_17958), .ZN(
      n_257_76_6415));
   NAND2_X1 i_257_76_6426 (.A1(n_257_76_6414), .A2(n_257_76_6415), .ZN(
      n_257_76_6416));
   NOR3_X1 i_257_76_6427 (.A1(n_257_76_6398), .A2(n_257_76_6400), .A3(
      n_257_76_6416), .ZN(n_257_76_6417));
   NAND3_X1 i_257_76_6428 (.A1(n_257_398), .A2(n_257_484), .A3(n_257_442), 
      .ZN(n_257_76_6418));
   INV_X1 i_257_76_6429 (.A(n_257_76_6418), .ZN(n_257_76_6419));
   NAND3_X1 i_257_76_6430 (.A1(n_257_76_5981), .A2(n_257_76_6368), .A3(
      n_257_76_6419), .ZN(n_257_76_6420));
   NOR2_X1 i_257_76_6431 (.A1(n_257_76_6420), .A2(n_257_1069), .ZN(n_257_76_6421));
   NAND2_X1 i_257_76_6432 (.A1(n_257_420), .A2(n_257_663), .ZN(n_257_76_6422));
   NAND4_X1 i_257_76_6433 (.A1(n_257_76_6421), .A2(n_257_76_5989), .A3(
      n_257_76_5927), .A4(n_257_76_6422), .ZN(n_257_76_6423));
   INV_X1 i_257_76_6434 (.A(n_257_76_6423), .ZN(n_257_76_6424));
   NAND2_X1 i_257_76_6435 (.A1(n_257_76_5931), .A2(n_257_76_6218), .ZN(
      n_257_76_6425));
   INV_X1 i_257_76_6436 (.A(n_257_76_6425), .ZN(n_257_76_6426));
   INV_X1 i_257_76_6437 (.A(n_257_76_6272), .ZN(n_257_76_6427));
   NAND3_X1 i_257_76_6438 (.A1(n_257_76_6424), .A2(n_257_76_6426), .A3(
      n_257_76_6427), .ZN(n_257_76_6428));
   NAND4_X1 i_257_76_6439 (.A1(n_257_76_5906), .A2(n_257_76_5934), .A3(
      n_257_76_5935), .A4(n_257_76_5930), .ZN(n_257_76_6429));
   NOR2_X1 i_257_76_6440 (.A1(n_257_76_6428), .A2(n_257_76_6429), .ZN(
      n_257_76_6430));
   NAND3_X1 i_257_76_6441 (.A1(n_257_76_6430), .A2(n_257_76_5999), .A3(
      n_257_76_6000), .ZN(n_257_76_6431));
   INV_X1 i_257_76_6442 (.A(n_257_76_6431), .ZN(n_257_76_6432));
   NAND3_X1 i_257_76_6443 (.A1(n_257_76_6201), .A2(n_257_76_5942), .A3(
      n_257_76_6003), .ZN(n_257_76_6433));
   INV_X1 i_257_76_6444 (.A(n_257_76_6433), .ZN(n_257_76_6434));
   NAND3_X1 i_257_76_6445 (.A1(n_257_76_6004), .A2(n_257_76_5992), .A3(
      n_257_76_6206), .ZN(n_257_76_6435));
   INV_X1 i_257_76_6446 (.A(n_257_76_6435), .ZN(n_257_76_6436));
   NAND3_X1 i_257_76_6447 (.A1(n_257_76_5939), .A2(n_257_76_5973), .A3(
      n_257_76_5974), .ZN(n_257_76_6437));
   INV_X1 i_257_76_6448 (.A(n_257_76_6437), .ZN(n_257_76_6438));
   NAND4_X1 i_257_76_6449 (.A1(n_257_76_6436), .A2(n_257_76_5943), .A3(
      n_257_76_5938), .A4(n_257_76_6438), .ZN(n_257_76_6439));
   INV_X1 i_257_76_6450 (.A(n_257_76_6439), .ZN(n_257_76_6440));
   NAND3_X1 i_257_76_6451 (.A1(n_257_76_6432), .A2(n_257_76_6434), .A3(
      n_257_76_6440), .ZN(n_257_76_6441));
   NOR3_X1 i_257_76_6452 (.A1(n_257_76_6441), .A2(n_257_76_6021), .A3(
      n_257_76_6225), .ZN(n_257_76_6442));
   AOI21_X1 i_257_76_6453 (.A(n_257_76_6417), .B1(n_257_76_18060), .B2(
      n_257_76_6442), .ZN(n_257_76_6443));
   NAND3_X1 i_257_76_6454 (.A1(n_257_76_6333), .A2(n_257_76_6352), .A3(
      n_257_76_6443), .ZN(n_257_76_6444));
   INV_X1 i_257_76_6455 (.A(n_257_76_6444), .ZN(n_257_76_6445));
   NAND3_X1 i_257_76_6456 (.A1(n_257_76_5906), .A2(n_257_76_5934), .A3(
      n_257_76_18046), .ZN(n_257_76_6446));
   NAND3_X1 i_257_76_6457 (.A1(n_257_448), .A2(n_257_76_5927), .A3(n_257_76_5907), 
      .ZN(n_257_76_6447));
   INV_X1 i_257_76_6458 (.A(n_257_76_6447), .ZN(n_257_76_6448));
   NAND3_X1 i_257_76_6459 (.A1(n_257_76_6448), .A2(n_257_76_5935), .A3(
      n_257_76_5931), .ZN(n_257_76_6449));
   NOR2_X1 i_257_76_6460 (.A1(n_257_76_6446), .A2(n_257_76_6449), .ZN(
      n_257_76_6450));
   NAND4_X1 i_257_76_6461 (.A1(n_257_76_5941), .A2(n_257_76_5942), .A3(
      n_257_76_6450), .A4(n_257_76_5943), .ZN(n_257_76_6451));
   INV_X1 i_257_76_6462 (.A(n_257_76_6451), .ZN(n_257_76_6452));
   NAND3_X1 i_257_76_6463 (.A1(n_257_76_6452), .A2(n_257_76_5905), .A3(n_257_679), 
      .ZN(n_257_76_6453));
   NOR2_X1 i_257_76_6464 (.A1(n_257_76_6021), .A2(n_257_76_6453), .ZN(
      n_257_76_6454));
   NOR3_X1 i_257_76_6465 (.A1(n_257_76_6021), .A2(n_257_76_6414), .A3(
      n_257_76_6225), .ZN(n_257_76_6455));
   AOI22_X1 i_257_76_6466 (.A1(n_257_76_18079), .A2(n_257_76_6454), .B1(
      n_257_76_18064), .B2(n_257_76_6455), .ZN(n_257_76_6456));
   NAND3_X1 i_257_76_6467 (.A1(n_257_76_6313), .A2(n_257_76_6445), .A3(
      n_257_76_6456), .ZN(n_257_76_6457));
   NOR2_X1 i_257_76_6468 (.A1(n_257_76_6266), .A2(n_257_76_6457), .ZN(
      n_257_76_6458));
   NAND2_X1 i_257_76_6469 (.A1(n_257_76_6142), .A2(n_257_76_6458), .ZN(n_10));
   NAND2_X1 i_257_76_6470 (.A1(n_257_1006), .A2(n_257_444), .ZN(n_257_76_6459));
   NAND2_X1 i_257_76_6471 (.A1(n_257_441), .A2(n_257_974), .ZN(n_257_76_6460));
   NAND2_X1 i_257_76_6472 (.A1(n_257_942), .A2(n_257_442), .ZN(n_257_76_6461));
   NOR2_X1 i_257_76_6473 (.A1(n_257_1070), .A2(n_257_76_6461), .ZN(n_257_76_6462));
   NAND2_X1 i_257_76_6474 (.A1(n_257_440), .A2(n_257_76_6462), .ZN(n_257_76_6463));
   INV_X1 i_257_76_6475 (.A(n_257_76_6463), .ZN(n_257_76_6464));
   NAND2_X1 i_257_76_6476 (.A1(n_257_76_6460), .A2(n_257_76_6464), .ZN(
      n_257_76_6465));
   INV_X1 i_257_76_6477 (.A(n_257_76_6465), .ZN(n_257_76_6466));
   NAND2_X1 i_257_76_6478 (.A1(n_257_76_6459), .A2(n_257_76_6466), .ZN(
      n_257_76_6467));
   INV_X1 i_257_76_6479 (.A(n_257_76_6467), .ZN(n_257_76_6468));
   NAND2_X1 i_257_76_6480 (.A1(n_257_1038), .A2(n_257_443), .ZN(n_257_76_6469));
   NAND2_X1 i_257_76_6481 (.A1(n_257_76_6468), .A2(n_257_76_6469), .ZN(
      n_257_76_6470));
   INV_X1 i_257_76_6482 (.A(n_257_76_6470), .ZN(n_257_76_6471));
   NAND2_X1 i_257_76_6483 (.A1(n_257_17), .A2(n_257_76_6471), .ZN(n_257_76_6472));
   NOR2_X1 i_257_76_6484 (.A1(n_257_1070), .A2(n_257_76_17412), .ZN(
      n_257_76_6473));
   NAND2_X1 i_257_76_6485 (.A1(n_257_443), .A2(n_257_76_6473), .ZN(n_257_76_6474));
   INV_X1 i_257_76_6486 (.A(n_257_76_6474), .ZN(n_257_76_6475));
   NAND2_X1 i_257_76_6487 (.A1(n_257_1038), .A2(n_257_76_6475), .ZN(
      n_257_76_6476));
   INV_X1 i_257_76_6488 (.A(n_257_76_6476), .ZN(n_257_76_6477));
   NAND2_X1 i_257_76_6489 (.A1(n_257_76_18072), .A2(n_257_76_6477), .ZN(
      n_257_76_6478));
   NAND2_X1 i_257_76_6490 (.A1(n_257_446), .A2(n_257_840), .ZN(n_257_76_6479));
   NAND2_X1 i_257_76_6491 (.A1(n_257_449), .A2(n_257_1084), .ZN(n_257_76_6480));
   NAND2_X1 i_257_76_6492 (.A1(n_257_447), .A2(n_257_776), .ZN(n_257_76_6481));
   NAND3_X1 i_257_76_6493 (.A1(n_257_76_6479), .A2(n_257_76_6480), .A3(
      n_257_76_6481), .ZN(n_257_76_6482));
   INV_X1 i_257_76_6494 (.A(n_257_76_6482), .ZN(n_257_76_6483));
   NAND2_X1 i_257_76_6495 (.A1(n_257_712), .A2(n_257_435), .ZN(n_257_76_6484));
   NAND3_X1 i_257_76_6496 (.A1(n_257_76_6473), .A2(n_257_640), .A3(n_257_450), 
      .ZN(n_257_76_6485));
   INV_X1 i_257_76_6497 (.A(n_257_76_6485), .ZN(n_257_76_6486));
   NAND2_X1 i_257_76_6498 (.A1(n_257_440), .A2(n_257_942), .ZN(n_257_76_6487));
   NAND2_X1 i_257_76_6499 (.A1(n_257_438), .A2(n_257_1076), .ZN(n_257_76_6488));
   NAND4_X1 i_257_76_6500 (.A1(n_257_76_6484), .A2(n_257_76_6486), .A3(
      n_257_76_6487), .A4(n_257_76_6488), .ZN(n_257_76_6489));
   INV_X1 i_257_76_6501 (.A(n_257_76_6489), .ZN(n_257_76_6490));
   NAND2_X1 i_257_76_6502 (.A1(n_257_910), .A2(n_257_439), .ZN(n_257_76_6491));
   NAND4_X1 i_257_76_6503 (.A1(n_257_76_6483), .A2(n_257_76_6490), .A3(
      n_257_76_6460), .A4(n_257_76_6491), .ZN(n_257_76_6492));
   NAND2_X1 i_257_76_6504 (.A1(n_257_744), .A2(n_257_436), .ZN(n_257_76_6493));
   NAND2_X1 i_257_76_6505 (.A1(n_257_872), .A2(n_257_445), .ZN(n_257_76_6494));
   NAND2_X1 i_257_76_6506 (.A1(n_257_808), .A2(n_257_437), .ZN(n_257_76_6495));
   NAND3_X1 i_257_76_6507 (.A1(n_257_76_6493), .A2(n_257_76_6494), .A3(
      n_257_76_6495), .ZN(n_257_76_6496));
   NOR2_X1 i_257_76_6508 (.A1(n_257_76_6492), .A2(n_257_76_6496), .ZN(
      n_257_76_6497));
   NAND2_X1 i_257_76_6509 (.A1(n_257_680), .A2(n_257_448), .ZN(n_257_76_6498));
   NAND3_X1 i_257_76_6510 (.A1(n_257_76_6497), .A2(n_257_76_6459), .A3(
      n_257_76_6498), .ZN(n_257_76_6499));
   INV_X1 i_257_76_6511 (.A(n_257_76_6469), .ZN(n_257_76_6500));
   NOR2_X1 i_257_76_6512 (.A1(n_257_76_6499), .A2(n_257_76_6500), .ZN(
      n_257_76_6501));
   NAND2_X1 i_257_76_6513 (.A1(n_257_28), .A2(n_257_76_6501), .ZN(n_257_76_6502));
   NAND3_X1 i_257_76_6514 (.A1(n_257_76_6472), .A2(n_257_76_6478), .A3(
      n_257_76_6502), .ZN(n_257_76_6503));
   INV_X1 i_257_76_6515 (.A(n_257_76_6473), .ZN(n_257_76_6504));
   INV_X1 i_257_76_6516 (.A(n_257_840), .ZN(n_257_76_6505));
   NOR2_X1 i_257_76_6517 (.A1(n_257_76_6504), .A2(n_257_76_6505), .ZN(
      n_257_76_6506));
   NAND4_X1 i_257_76_6518 (.A1(n_257_446), .A2(n_257_76_6506), .A3(n_257_76_6487), 
      .A4(n_257_76_6488), .ZN(n_257_76_6507));
   INV_X1 i_257_76_6519 (.A(n_257_76_6507), .ZN(n_257_76_6508));
   NAND3_X1 i_257_76_6520 (.A1(n_257_76_6508), .A2(n_257_76_6460), .A3(
      n_257_76_6491), .ZN(n_257_76_6509));
   INV_X1 i_257_76_6521 (.A(n_257_76_6494), .ZN(n_257_76_6510));
   NOR2_X1 i_257_76_6522 (.A1(n_257_76_6509), .A2(n_257_76_6510), .ZN(
      n_257_76_6511));
   NAND2_X1 i_257_76_6523 (.A1(n_257_76_6459), .A2(n_257_76_6511), .ZN(
      n_257_76_6512));
   INV_X1 i_257_76_6524 (.A(n_257_76_6512), .ZN(n_257_76_6513));
   NAND2_X1 i_257_76_6525 (.A1(n_257_76_6513), .A2(n_257_76_6469), .ZN(
      n_257_76_6514));
   INV_X1 i_257_76_6526 (.A(n_257_76_6514), .ZN(n_257_76_6515));
   NAND2_X1 i_257_76_6527 (.A1(n_257_76_18070), .A2(n_257_76_6515), .ZN(
      n_257_76_6516));
   INV_X1 i_257_76_6528 (.A(n_257_76_6460), .ZN(n_257_76_6517));
   NAND2_X1 i_257_76_6529 (.A1(n_257_439), .A2(n_257_76_6473), .ZN(n_257_76_6518));
   INV_X1 i_257_76_6530 (.A(n_257_76_6518), .ZN(n_257_76_6519));
   NAND3_X1 i_257_76_6531 (.A1(n_257_910), .A2(n_257_76_6487), .A3(n_257_76_6519), 
      .ZN(n_257_76_6520));
   NOR2_X1 i_257_76_6532 (.A1(n_257_76_6517), .A2(n_257_76_6520), .ZN(
      n_257_76_6521));
   NAND2_X1 i_257_76_6533 (.A1(n_257_76_6459), .A2(n_257_76_6521), .ZN(
      n_257_76_6522));
   INV_X1 i_257_76_6534 (.A(n_257_76_6522), .ZN(n_257_76_6523));
   NAND2_X1 i_257_76_6535 (.A1(n_257_76_6523), .A2(n_257_76_6469), .ZN(
      n_257_76_6524));
   INV_X1 i_257_76_6536 (.A(n_257_76_6524), .ZN(n_257_76_6525));
   NAND2_X1 i_257_76_6537 (.A1(n_257_76_18084), .A2(n_257_76_6525), .ZN(
      n_257_76_6526));
   NAND2_X1 i_257_76_6538 (.A1(n_257_124), .A2(n_257_430), .ZN(n_257_76_6527));
   NAND2_X1 i_257_76_6539 (.A1(n_257_451), .A2(n_257_463), .ZN(n_257_76_6528));
   NAND4_X1 i_257_76_6540 (.A1(n_257_76_6483), .A2(n_257_76_6527), .A3(
      n_257_76_6528), .A4(n_257_76_6460), .ZN(n_257_76_6529));
   NOR2_X1 i_257_76_6541 (.A1(n_257_76_6496), .A2(n_257_76_6529), .ZN(
      n_257_76_6530));
   NAND2_X1 i_257_76_6542 (.A1(n_257_544), .A2(n_257_426), .ZN(n_257_76_6531));
   NAND2_X1 i_257_76_6543 (.A1(n_257_46), .A2(n_257_433), .ZN(n_257_76_6532));
   NAND3_X1 i_257_76_6544 (.A1(n_257_76_6531), .A2(n_257_76_6484), .A3(
      n_257_76_6532), .ZN(n_257_76_6533));
   INV_X1 i_257_76_6545 (.A(n_257_76_6533), .ZN(n_257_76_6534));
   INV_X1 i_257_76_6546 (.A(n_257_576), .ZN(n_257_76_6535));
   NAND2_X1 i_257_76_6547 (.A1(n_257_76_6535), .A2(n_257_442), .ZN(n_257_76_6536));
   OAI21_X1 i_257_76_6548 (.A(n_257_76_6536), .B1(n_257_428), .B2(n_257_76_17412), 
      .ZN(n_257_76_6537));
   INV_X1 i_257_76_6549 (.A(n_257_1070), .ZN(n_257_76_6538));
   NAND2_X1 i_257_76_6550 (.A1(n_257_432), .A2(n_257_608), .ZN(n_257_76_6539));
   NAND4_X1 i_257_76_6551 (.A1(n_257_76_6537), .A2(n_257_76_6538), .A3(
      n_257_76_6539), .A4(n_257_423), .ZN(n_257_76_6540));
   INV_X1 i_257_76_6552 (.A(n_257_76_6540), .ZN(n_257_76_6541));
   NAND2_X1 i_257_76_6553 (.A1(n_257_640), .A2(n_257_450), .ZN(n_257_76_6542));
   NAND2_X1 i_257_76_6554 (.A1(n_257_512), .A2(n_257_424), .ZN(n_257_76_6543));
   NAND4_X1 i_257_76_6555 (.A1(n_257_76_6541), .A2(n_257_76_6488), .A3(
      n_257_76_6542), .A4(n_257_76_6543), .ZN(n_257_76_6544));
   INV_X1 i_257_76_6556 (.A(n_257_76_6544), .ZN(n_257_76_6545));
   NAND2_X1 i_257_76_6557 (.A1(n_257_203), .A2(n_257_427), .ZN(n_257_76_6546));
   NAND3_X1 i_257_76_6558 (.A1(n_257_283), .A2(n_257_76_6546), .A3(n_257_76_6487), 
      .ZN(n_257_76_6547));
   INV_X1 i_257_76_6559 (.A(n_257_76_6547), .ZN(n_257_76_6548));
   NAND4_X1 i_257_76_6560 (.A1(n_257_76_6534), .A2(n_257_76_6545), .A3(
      n_257_76_6491), .A4(n_257_76_6548), .ZN(n_257_76_6549));
   INV_X1 i_257_76_6561 (.A(n_257_76_6549), .ZN(n_257_76_6550));
   NAND2_X1 i_257_76_6562 (.A1(n_257_243), .A2(n_257_425), .ZN(n_257_76_6551));
   NAND2_X1 i_257_76_6563 (.A1(n_257_86), .A2(n_257_431), .ZN(n_257_76_6552));
   NAND3_X1 i_257_76_6564 (.A1(n_257_76_6550), .A2(n_257_76_6551), .A3(
      n_257_76_6552), .ZN(n_257_76_6553));
   INV_X1 i_257_76_6565 (.A(n_257_76_6553), .ZN(n_257_76_6554));
   NAND3_X1 i_257_76_6566 (.A1(n_257_76_6530), .A2(n_257_76_6498), .A3(
      n_257_76_6554), .ZN(n_257_76_6555));
   INV_X1 i_257_76_6567 (.A(n_257_76_6555), .ZN(n_257_76_6556));
   NAND2_X1 i_257_76_6568 (.A1(n_257_163), .A2(n_257_429), .ZN(n_257_76_6557));
   NAND2_X1 i_257_76_6569 (.A1(n_257_76_6557), .A2(n_257_76_6459), .ZN(
      n_257_76_6558));
   INV_X1 i_257_76_6570 (.A(n_257_76_6558), .ZN(n_257_76_6559));
   NAND3_X1 i_257_76_6571 (.A1(n_257_76_6556), .A2(n_257_76_6559), .A3(
      n_257_76_6469), .ZN(n_257_76_6560));
   INV_X1 i_257_76_6572 (.A(n_257_76_6560), .ZN(n_257_76_6561));
   NAND2_X1 i_257_76_6573 (.A1(n_257_76_18066), .A2(n_257_76_6561), .ZN(
      n_257_76_6562));
   NAND3_X1 i_257_76_6574 (.A1(n_257_76_6516), .A2(n_257_76_6526), .A3(
      n_257_76_6562), .ZN(n_257_76_6563));
   NOR2_X1 i_257_76_6575 (.A1(n_257_76_6503), .A2(n_257_76_6563), .ZN(
      n_257_76_6564));
   INV_X1 i_257_76_6576 (.A(n_257_974), .ZN(n_257_76_6565));
   NOR2_X1 i_257_76_6577 (.A1(n_257_76_6504), .A2(n_257_76_6565), .ZN(
      n_257_76_6566));
   NAND2_X1 i_257_76_6578 (.A1(n_257_441), .A2(n_257_76_6566), .ZN(n_257_76_6567));
   INV_X1 i_257_76_6579 (.A(n_257_76_6567), .ZN(n_257_76_6568));
   NAND2_X1 i_257_76_6580 (.A1(n_257_76_6459), .A2(n_257_76_6568), .ZN(
      n_257_76_6569));
   INV_X1 i_257_76_6581 (.A(n_257_76_6569), .ZN(n_257_76_6570));
   NAND2_X1 i_257_76_6582 (.A1(n_257_76_6570), .A2(n_257_76_6469), .ZN(
      n_257_76_6571));
   INV_X1 i_257_76_6583 (.A(n_257_76_6571), .ZN(n_257_76_6572));
   NAND2_X1 i_257_76_6584 (.A1(n_257_76_18071), .A2(n_257_76_6572), .ZN(
      n_257_76_6573));
   NAND2_X1 i_257_76_6585 (.A1(n_257_76_6479), .A2(n_257_76_6481), .ZN(
      n_257_76_6574));
   INV_X1 i_257_76_6586 (.A(n_257_76_6574), .ZN(n_257_76_6575));
   NOR2_X1 i_257_76_6587 (.A1(n_257_76_6504), .A2(n_257_76_17760), .ZN(
      n_257_76_6576));
   NAND4_X1 i_257_76_6588 (.A1(n_257_76_6576), .A2(n_257_76_6487), .A3(
      n_257_76_6488), .A4(n_257_712), .ZN(n_257_76_6577));
   INV_X1 i_257_76_6589 (.A(n_257_76_6577), .ZN(n_257_76_6578));
   NAND4_X1 i_257_76_6590 (.A1(n_257_76_6575), .A2(n_257_76_6578), .A3(
      n_257_76_6460), .A4(n_257_76_6491), .ZN(n_257_76_6579));
   NOR2_X1 i_257_76_6591 (.A1(n_257_76_6496), .A2(n_257_76_6579), .ZN(
      n_257_76_6580));
   NAND2_X1 i_257_76_6592 (.A1(n_257_76_6459), .A2(n_257_76_6580), .ZN(
      n_257_76_6581));
   INV_X1 i_257_76_6593 (.A(n_257_76_6581), .ZN(n_257_76_6582));
   NAND2_X1 i_257_76_6594 (.A1(n_257_76_6582), .A2(n_257_76_6469), .ZN(
      n_257_76_6583));
   INV_X1 i_257_76_6595 (.A(n_257_76_6583), .ZN(n_257_76_6584));
   NAND2_X1 i_257_76_6596 (.A1(n_257_76_18078), .A2(n_257_76_6584), .ZN(
      n_257_76_6585));
   NAND3_X1 i_257_76_6597 (.A1(n_257_76_6527), .A2(n_257_76_6528), .A3(
      n_257_76_6460), .ZN(n_257_76_6586));
   INV_X1 i_257_76_6598 (.A(n_257_76_6586), .ZN(n_257_76_6587));
   NAND4_X1 i_257_76_6599 (.A1(n_257_76_6491), .A2(n_257_76_6479), .A3(
      n_257_76_6480), .A4(n_257_76_6481), .ZN(n_257_76_6588));
   INV_X1 i_257_76_6600 (.A(n_257_76_6588), .ZN(n_257_76_6589));
   NAND2_X1 i_257_76_6601 (.A1(n_257_442), .A2(n_257_576), .ZN(n_257_76_6590));
   INV_X1 i_257_76_6602 (.A(n_257_76_6590), .ZN(n_257_76_6591));
   NAND2_X1 i_257_76_6603 (.A1(n_257_428), .A2(n_257_76_6591), .ZN(n_257_76_6592));
   INV_X1 i_257_76_6604 (.A(n_257_76_6592), .ZN(n_257_76_6593));
   NAND3_X1 i_257_76_6605 (.A1(n_257_76_6538), .A2(n_257_76_6539), .A3(
      n_257_76_6593), .ZN(n_257_76_6594));
   INV_X1 i_257_76_6606 (.A(n_257_76_6594), .ZN(n_257_76_6595));
   NAND4_X1 i_257_76_6607 (.A1(n_257_76_6487), .A2(n_257_76_6488), .A3(
      n_257_76_6542), .A4(n_257_76_6595), .ZN(n_257_76_6596));
   NAND2_X1 i_257_76_6608 (.A1(n_257_76_6484), .A2(n_257_76_6532), .ZN(
      n_257_76_6597));
   NOR2_X1 i_257_76_6609 (.A1(n_257_76_6596), .A2(n_257_76_6597), .ZN(
      n_257_76_6598));
   NAND4_X1 i_257_76_6610 (.A1(n_257_76_6587), .A2(n_257_76_6589), .A3(
      n_257_76_6598), .A4(n_257_76_6495), .ZN(n_257_76_6599));
   NAND3_X1 i_257_76_6611 (.A1(n_257_76_6552), .A2(n_257_76_6493), .A3(
      n_257_76_6494), .ZN(n_257_76_6600));
   NOR2_X1 i_257_76_6612 (.A1(n_257_76_6599), .A2(n_257_76_6600), .ZN(
      n_257_76_6601));
   NAND4_X1 i_257_76_6613 (.A1(n_257_76_6601), .A2(n_257_76_6557), .A3(
      n_257_76_6459), .A4(n_257_76_6498), .ZN(n_257_76_6602));
   NOR2_X1 i_257_76_6614 (.A1(n_257_76_6602), .A2(n_257_76_6500), .ZN(
      n_257_76_6603));
   NAND2_X1 i_257_76_6615 (.A1(n_257_76_18074), .A2(n_257_76_6603), .ZN(
      n_257_76_6604));
   NAND3_X1 i_257_76_6616 (.A1(n_257_76_6573), .A2(n_257_76_6585), .A3(
      n_257_76_6604), .ZN(n_257_76_6605));
   NAND2_X1 i_257_76_6617 (.A1(n_257_1070), .A2(n_257_442), .ZN(n_257_76_6606));
   INV_X1 i_257_76_6618 (.A(n_257_76_6606), .ZN(n_257_76_6607));
   NAND2_X1 i_257_76_6619 (.A1(n_257_13), .A2(n_257_76_6607), .ZN(n_257_76_6608));
   NOR2_X1 i_257_76_6620 (.A1(n_257_76_6504), .A2(n_257_76_11918), .ZN(
      n_257_76_6609));
   NAND3_X1 i_257_76_6621 (.A1(n_257_76_6609), .A2(n_257_76_6487), .A3(
      n_257_76_6488), .ZN(n_257_76_6610));
   INV_X1 i_257_76_6622 (.A(n_257_76_6610), .ZN(n_257_76_6611));
   NAND4_X1 i_257_76_6623 (.A1(n_257_872), .A2(n_257_76_6460), .A3(n_257_76_6611), 
      .A4(n_257_76_6491), .ZN(n_257_76_6612));
   INV_X1 i_257_76_6624 (.A(n_257_76_6612), .ZN(n_257_76_6613));
   NAND2_X1 i_257_76_6625 (.A1(n_257_76_6459), .A2(n_257_76_6613), .ZN(
      n_257_76_6614));
   INV_X1 i_257_76_6626 (.A(n_257_76_6614), .ZN(n_257_76_6615));
   NAND2_X1 i_257_76_6627 (.A1(n_257_76_6615), .A2(n_257_76_6469), .ZN(
      n_257_76_6616));
   INV_X1 i_257_76_6628 (.A(n_257_76_6616), .ZN(n_257_76_6617));
   NAND2_X1 i_257_76_6629 (.A1(n_257_76_18077), .A2(n_257_76_6617), .ZN(
      n_257_76_6618));
   NAND2_X1 i_257_76_6630 (.A1(n_257_76_6608), .A2(n_257_76_6618), .ZN(
      n_257_76_6619));
   NOR2_X1 i_257_76_6631 (.A1(n_257_76_6605), .A2(n_257_76_6619), .ZN(
      n_257_76_6620));
   NAND2_X1 i_257_76_6632 (.A1(n_257_76_6494), .A2(n_257_76_6495), .ZN(
      n_257_76_6621));
   NOR2_X1 i_257_76_6633 (.A1(n_257_76_6529), .A2(n_257_76_6621), .ZN(
      n_257_76_6622));
   INV_X1 i_257_76_6634 (.A(n_257_76_6597), .ZN(n_257_76_6623));
   NAND4_X1 i_257_76_6635 (.A1(n_257_76_6537), .A2(n_257_76_6538), .A3(
      n_257_76_6539), .A4(n_257_426), .ZN(n_257_76_6624));
   INV_X1 i_257_76_6636 (.A(n_257_76_6624), .ZN(n_257_76_6625));
   NAND3_X1 i_257_76_6637 (.A1(n_257_76_6625), .A2(n_257_76_6488), .A3(
      n_257_76_6542), .ZN(n_257_76_6626));
   INV_X1 i_257_76_6638 (.A(n_257_76_6626), .ZN(n_257_76_6627));
   NAND3_X1 i_257_76_6639 (.A1(n_257_76_6546), .A2(n_257_544), .A3(n_257_76_6487), 
      .ZN(n_257_76_6628));
   INV_X1 i_257_76_6640 (.A(n_257_76_6628), .ZN(n_257_76_6629));
   NAND4_X1 i_257_76_6641 (.A1(n_257_76_6623), .A2(n_257_76_6627), .A3(
      n_257_76_6629), .A4(n_257_76_6491), .ZN(n_257_76_6630));
   INV_X1 i_257_76_6642 (.A(n_257_76_6630), .ZN(n_257_76_6631));
   NAND3_X1 i_257_76_6643 (.A1(n_257_76_6631), .A2(n_257_76_6552), .A3(
      n_257_76_6493), .ZN(n_257_76_6632));
   INV_X1 i_257_76_6644 (.A(n_257_76_6632), .ZN(n_257_76_6633));
   NAND3_X1 i_257_76_6645 (.A1(n_257_76_6498), .A2(n_257_76_6622), .A3(
      n_257_76_6633), .ZN(n_257_76_6634));
   INV_X1 i_257_76_6646 (.A(n_257_76_6634), .ZN(n_257_76_6635));
   NAND3_X1 i_257_76_6647 (.A1(n_257_76_6635), .A2(n_257_76_6559), .A3(
      n_257_76_6469), .ZN(n_257_76_6636));
   INV_X1 i_257_76_6648 (.A(n_257_76_6636), .ZN(n_257_76_6637));
   NAND2_X1 i_257_76_6649 (.A1(n_257_76_18076), .A2(n_257_76_6637), .ZN(
      n_257_76_6638));
   NAND3_X1 i_257_76_6650 (.A1(n_257_76_6494), .A2(n_257_76_6495), .A3(n_257_744), 
      .ZN(n_257_76_6639));
   NOR2_X1 i_257_76_6651 (.A1(n_257_76_6504), .A2(n_257_76_8311), .ZN(
      n_257_76_6640));
   NAND3_X1 i_257_76_6652 (.A1(n_257_76_6640), .A2(n_257_76_6487), .A3(
      n_257_76_6488), .ZN(n_257_76_6641));
   INV_X1 i_257_76_6653 (.A(n_257_76_6641), .ZN(n_257_76_6642));
   NAND4_X1 i_257_76_6654 (.A1(n_257_76_6575), .A2(n_257_76_6460), .A3(
      n_257_76_6491), .A4(n_257_76_6642), .ZN(n_257_76_6643));
   NOR2_X1 i_257_76_6655 (.A1(n_257_76_6639), .A2(n_257_76_6643), .ZN(
      n_257_76_6644));
   NAND2_X1 i_257_76_6656 (.A1(n_257_76_6459), .A2(n_257_76_6644), .ZN(
      n_257_76_6645));
   INV_X1 i_257_76_6657 (.A(n_257_76_6645), .ZN(n_257_76_6646));
   NAND2_X1 i_257_76_6658 (.A1(n_257_76_6646), .A2(n_257_76_6469), .ZN(
      n_257_76_6647));
   INV_X1 i_257_76_6659 (.A(n_257_76_6647), .ZN(n_257_76_6648));
   NAND2_X1 i_257_76_6660 (.A1(n_257_76_18069), .A2(n_257_76_6648), .ZN(
      n_257_76_6649));
   NAND2_X1 i_257_76_6661 (.A1(n_257_76_6528), .A2(n_257_76_6460), .ZN(
      n_257_76_6650));
   INV_X1 i_257_76_6662 (.A(n_257_76_6650), .ZN(n_257_76_6651));
   NAND2_X1 i_257_76_6663 (.A1(n_257_608), .A2(n_257_442), .ZN(n_257_76_6652));
   INV_X1 i_257_76_6664 (.A(n_257_76_6652), .ZN(n_257_76_6653));
   NAND2_X1 i_257_76_6665 (.A1(n_257_432), .A2(n_257_76_6653), .ZN(n_257_76_6654));
   NOR2_X1 i_257_76_6666 (.A1(n_257_76_6654), .A2(n_257_1070), .ZN(n_257_76_6655));
   NAND4_X1 i_257_76_6667 (.A1(n_257_76_6487), .A2(n_257_76_6488), .A3(
      n_257_76_6542), .A4(n_257_76_6655), .ZN(n_257_76_6656));
   NOR2_X1 i_257_76_6668 (.A1(n_257_76_6656), .A2(n_257_76_6597), .ZN(
      n_257_76_6657));
   NAND3_X1 i_257_76_6669 (.A1(n_257_76_6589), .A2(n_257_76_6651), .A3(
      n_257_76_6657), .ZN(n_257_76_6658));
   NOR2_X1 i_257_76_6670 (.A1(n_257_76_6658), .A2(n_257_76_6496), .ZN(
      n_257_76_6659));
   NAND3_X1 i_257_76_6671 (.A1(n_257_76_6659), .A2(n_257_76_6459), .A3(
      n_257_76_6498), .ZN(n_257_76_6660));
   NOR2_X1 i_257_76_6672 (.A1(n_257_76_6660), .A2(n_257_76_6500), .ZN(
      n_257_76_6661));
   NAND2_X1 i_257_76_6673 (.A1(n_257_68), .A2(n_257_76_6661), .ZN(n_257_76_6662));
   NAND3_X1 i_257_76_6674 (.A1(n_257_76_6638), .A2(n_257_76_6649), .A3(
      n_257_76_6662), .ZN(n_257_76_6663));
   NOR2_X1 i_257_76_6675 (.A1(n_257_76_6504), .A2(n_257_76_15924), .ZN(
      n_257_76_6664));
   NAND3_X1 i_257_76_6676 (.A1(n_257_76_6664), .A2(n_257_76_6487), .A3(
      n_257_76_6488), .ZN(n_257_76_6665));
   INV_X1 i_257_76_6677 (.A(n_257_76_6665), .ZN(n_257_76_6666));
   NAND3_X1 i_257_76_6678 (.A1(n_257_76_6666), .A2(n_257_76_6491), .A3(
      n_257_76_6479), .ZN(n_257_76_6667));
   INV_X1 i_257_76_6679 (.A(n_257_76_6667), .ZN(n_257_76_6668));
   NAND2_X1 i_257_76_6680 (.A1(n_257_808), .A2(n_257_76_6460), .ZN(n_257_76_6669));
   INV_X1 i_257_76_6681 (.A(n_257_76_6669), .ZN(n_257_76_6670));
   NAND3_X1 i_257_76_6682 (.A1(n_257_76_6668), .A2(n_257_76_6670), .A3(
      n_257_76_6494), .ZN(n_257_76_6671));
   INV_X1 i_257_76_6683 (.A(n_257_76_6671), .ZN(n_257_76_6672));
   NAND2_X1 i_257_76_6684 (.A1(n_257_76_6459), .A2(n_257_76_6672), .ZN(
      n_257_76_6673));
   INV_X1 i_257_76_6685 (.A(n_257_76_6673), .ZN(n_257_76_6674));
   NAND2_X1 i_257_76_6686 (.A1(n_257_76_6674), .A2(n_257_76_6469), .ZN(
      n_257_76_6675));
   INV_X1 i_257_76_6687 (.A(n_257_76_6675), .ZN(n_257_76_6676));
   NAND2_X1 i_257_76_6688 (.A1(n_257_22), .A2(n_257_76_6676), .ZN(n_257_76_6677));
   NAND2_X1 i_257_76_6689 (.A1(n_257_444), .A2(n_257_76_6473), .ZN(n_257_76_6678));
   INV_X1 i_257_76_6690 (.A(n_257_76_6678), .ZN(n_257_76_6679));
   NAND2_X1 i_257_76_6691 (.A1(n_257_1006), .A2(n_257_76_6679), .ZN(
      n_257_76_6680));
   INV_X1 i_257_76_6692 (.A(n_257_76_6680), .ZN(n_257_76_6681));
   NAND2_X1 i_257_76_6693 (.A1(n_257_76_6469), .A2(n_257_76_6681), .ZN(
      n_257_76_6682));
   INV_X1 i_257_76_6694 (.A(n_257_76_6682), .ZN(n_257_76_6683));
   NAND2_X1 i_257_76_6695 (.A1(n_257_76_18075), .A2(n_257_76_6683), .ZN(
      n_257_76_6684));
   NAND2_X1 i_257_76_6696 (.A1(n_257_76_6677), .A2(n_257_76_6684), .ZN(
      n_257_76_6685));
   NOR2_X1 i_257_76_6697 (.A1(n_257_76_6663), .A2(n_257_76_6685), .ZN(
      n_257_76_6686));
   NAND3_X1 i_257_76_6698 (.A1(n_257_76_6564), .A2(n_257_76_6620), .A3(
      n_257_76_6686), .ZN(n_257_76_6687));
   INV_X1 i_257_76_6699 (.A(n_257_76_6687), .ZN(n_257_76_6688));
   NOR2_X1 i_257_76_6700 (.A1(n_257_1070), .A2(n_257_76_17633), .ZN(
      n_257_76_6689));
   NAND3_X1 i_257_76_6701 (.A1(n_257_46), .A2(n_257_76_6542), .A3(n_257_76_6689), 
      .ZN(n_257_76_6690));
   INV_X1 i_257_76_6702 (.A(n_257_76_6690), .ZN(n_257_76_6691));
   NAND2_X1 i_257_76_6703 (.A1(n_257_76_6487), .A2(n_257_76_6488), .ZN(
      n_257_76_6692));
   INV_X1 i_257_76_6704 (.A(n_257_76_6692), .ZN(n_257_76_6693));
   NAND4_X1 i_257_76_6705 (.A1(n_257_76_6691), .A2(n_257_76_6693), .A3(
      n_257_76_6481), .A4(n_257_76_6484), .ZN(n_257_76_6694));
   INV_X1 i_257_76_6706 (.A(n_257_76_6694), .ZN(n_257_76_6695));
   NAND3_X1 i_257_76_6707 (.A1(n_257_76_6491), .A2(n_257_76_6479), .A3(
      n_257_76_6480), .ZN(n_257_76_6696));
   INV_X1 i_257_76_6708 (.A(n_257_76_6696), .ZN(n_257_76_6697));
   NAND3_X1 i_257_76_6709 (.A1(n_257_76_6695), .A2(n_257_76_6651), .A3(
      n_257_76_6697), .ZN(n_257_76_6698));
   NOR2_X1 i_257_76_6710 (.A1(n_257_76_6698), .A2(n_257_76_6496), .ZN(
      n_257_76_6699));
   NAND3_X1 i_257_76_6711 (.A1(n_257_76_6699), .A2(n_257_76_6459), .A3(
      n_257_76_6498), .ZN(n_257_76_6700));
   NOR2_X1 i_257_76_6712 (.A1(n_257_76_6700), .A2(n_257_76_6500), .ZN(
      n_257_76_6701));
   NAND2_X1 i_257_76_6713 (.A1(n_257_76_18081), .A2(n_257_76_6701), .ZN(
      n_257_76_6702));
   NAND3_X1 i_257_76_6714 (.A1(n_257_76_6479), .A2(n_257_76_6481), .A3(
      n_257_76_6484), .ZN(n_257_76_6703));
   INV_X1 i_257_76_6715 (.A(n_257_76_6703), .ZN(n_257_76_6704));
   NAND2_X1 i_257_76_6716 (.A1(n_257_1084), .A2(n_257_76_6473), .ZN(
      n_257_76_6705));
   INV_X1 i_257_76_6717 (.A(n_257_76_6705), .ZN(n_257_76_6706));
   NAND4_X1 i_257_76_6718 (.A1(n_257_76_6706), .A2(n_257_449), .A3(n_257_76_6487), 
      .A4(n_257_76_6488), .ZN(n_257_76_6707));
   INV_X1 i_257_76_6719 (.A(n_257_76_6707), .ZN(n_257_76_6708));
   NAND4_X1 i_257_76_6720 (.A1(n_257_76_6704), .A2(n_257_76_6460), .A3(
      n_257_76_6708), .A4(n_257_76_6491), .ZN(n_257_76_6709));
   NOR2_X1 i_257_76_6721 (.A1(n_257_76_6496), .A2(n_257_76_6709), .ZN(
      n_257_76_6710));
   NAND3_X1 i_257_76_6722 (.A1(n_257_76_6710), .A2(n_257_76_6459), .A3(
      n_257_76_6498), .ZN(n_257_76_6711));
   NOR2_X1 i_257_76_6723 (.A1(n_257_76_6500), .A2(n_257_76_6711), .ZN(
      n_257_76_6712));
   NAND2_X1 i_257_76_6724 (.A1(n_257_76_18083), .A2(n_257_76_6712), .ZN(
      n_257_76_6713));
   NAND4_X1 i_257_76_6725 (.A1(n_257_76_6460), .A2(n_257_76_6491), .A3(
      n_257_76_6479), .A4(n_257_76_6480), .ZN(n_257_76_6714));
   NAND3_X1 i_257_76_6726 (.A1(n_257_76_6538), .A2(n_257_76_6539), .A3(
      n_257_76_17331), .ZN(n_257_76_6715));
   INV_X1 i_257_76_6727 (.A(n_257_76_6715), .ZN(n_257_76_6716));
   NAND4_X1 i_257_76_6728 (.A1(n_257_76_6487), .A2(n_257_76_6488), .A3(
      n_257_76_6542), .A4(n_257_76_6716), .ZN(n_257_76_6717));
   INV_X1 i_257_76_6729 (.A(n_257_76_6717), .ZN(n_257_76_6718));
   NAND3_X1 i_257_76_6730 (.A1(n_257_76_6718), .A2(n_257_76_6623), .A3(
      n_257_76_6481), .ZN(n_257_76_6719));
   NOR2_X1 i_257_76_6731 (.A1(n_257_76_6714), .A2(n_257_76_6719), .ZN(
      n_257_76_6720));
   NAND2_X1 i_257_76_6732 (.A1(n_257_76_6552), .A2(n_257_76_6493), .ZN(
      n_257_76_6721));
   INV_X1 i_257_76_6733 (.A(n_257_76_6721), .ZN(n_257_76_6722));
   NAND2_X1 i_257_76_6734 (.A1(n_257_76_6527), .A2(n_257_76_6528), .ZN(
      n_257_76_6723));
   INV_X1 i_257_76_6735 (.A(n_257_76_6723), .ZN(n_257_76_6724));
   NAND3_X1 i_257_76_6736 (.A1(n_257_76_6724), .A2(n_257_76_6494), .A3(
      n_257_76_6495), .ZN(n_257_76_6725));
   INV_X1 i_257_76_6737 (.A(n_257_76_6725), .ZN(n_257_76_6726));
   NAND4_X1 i_257_76_6738 (.A1(n_257_163), .A2(n_257_76_6720), .A3(n_257_76_6722), 
      .A4(n_257_76_6726), .ZN(n_257_76_6727));
   INV_X1 i_257_76_6739 (.A(n_257_76_6727), .ZN(n_257_76_6728));
   NAND2_X1 i_257_76_6740 (.A1(n_257_76_6459), .A2(n_257_76_6498), .ZN(
      n_257_76_6729));
   INV_X1 i_257_76_6741 (.A(n_257_76_6729), .ZN(n_257_76_6730));
   NAND3_X1 i_257_76_6742 (.A1(n_257_76_6728), .A2(n_257_76_6730), .A3(
      n_257_76_6469), .ZN(n_257_76_6731));
   INV_X1 i_257_76_6743 (.A(n_257_76_6731), .ZN(n_257_76_6732));
   NAND2_X1 i_257_76_6744 (.A1(n_257_76_18061), .A2(n_257_76_6732), .ZN(
      n_257_76_6733));
   NAND3_X1 i_257_76_6745 (.A1(n_257_76_6702), .A2(n_257_76_6713), .A3(
      n_257_76_6733), .ZN(n_257_76_6734));
   INV_X1 i_257_76_6746 (.A(n_257_76_6734), .ZN(n_257_76_6735));
   NAND3_X1 i_257_76_6747 (.A1(n_257_438), .A2(n_257_76_6473), .A3(n_257_1076), 
      .ZN(n_257_76_6736));
   INV_X1 i_257_76_6748 (.A(n_257_76_6487), .ZN(n_257_76_6737));
   NOR2_X1 i_257_76_6749 (.A1(n_257_76_6736), .A2(n_257_76_6737), .ZN(
      n_257_76_6738));
   NAND3_X1 i_257_76_6750 (.A1(n_257_76_6460), .A2(n_257_76_6738), .A3(
      n_257_76_6491), .ZN(n_257_76_6739));
   INV_X1 i_257_76_6751 (.A(n_257_76_6739), .ZN(n_257_76_6740));
   NAND2_X1 i_257_76_6752 (.A1(n_257_76_6459), .A2(n_257_76_6740), .ZN(
      n_257_76_6741));
   INV_X1 i_257_76_6753 (.A(n_257_76_6741), .ZN(n_257_76_6742));
   NAND2_X1 i_257_76_6754 (.A1(n_257_76_6742), .A2(n_257_76_6469), .ZN(
      n_257_76_6743));
   INV_X1 i_257_76_6755 (.A(n_257_76_6743), .ZN(n_257_76_6744));
   NAND2_X1 i_257_76_6756 (.A1(n_257_76_18067), .A2(n_257_76_6744), .ZN(
      n_257_76_6745));
   NAND2_X1 i_257_76_6757 (.A1(n_257_76_6551), .A2(n_257_76_6552), .ZN(
      n_257_76_6746));
   INV_X1 i_257_76_6758 (.A(n_257_76_6746), .ZN(n_257_76_6747));
   NAND2_X1 i_257_76_6759 (.A1(n_257_76_6498), .A2(n_257_76_6747), .ZN(
      n_257_76_6748));
   INV_X1 i_257_76_6760 (.A(n_257_76_6748), .ZN(n_257_76_6749));
   NAND2_X1 i_257_76_6761 (.A1(n_257_283), .A2(n_257_423), .ZN(n_257_76_6750));
   NAND2_X1 i_257_76_6762 (.A1(n_257_76_6750), .A2(n_257_76_6479), .ZN(
      n_257_76_6751));
   INV_X1 i_257_76_6763 (.A(n_257_76_6751), .ZN(n_257_76_6752));
   NAND2_X1 i_257_76_6764 (.A1(n_257_76_6752), .A2(n_257_76_6491), .ZN(
      n_257_76_6753));
   NOR2_X1 i_257_76_6765 (.A1(n_257_76_6753), .A2(n_257_76_6650), .ZN(
      n_257_76_6754));
   NAND2_X1 i_257_76_6766 (.A1(n_257_321), .A2(n_257_422), .ZN(n_257_76_6755));
   NAND2_X1 i_257_76_6767 (.A1(n_257_76_6532), .A2(n_257_76_6755), .ZN(
      n_257_76_6756));
   NAND2_X1 i_257_76_6768 (.A1(n_257_76_6546), .A2(n_257_76_6487), .ZN(
      n_257_76_6757));
   NOR2_X1 i_257_76_6769 (.A1(n_257_76_6756), .A2(n_257_76_6757), .ZN(
      n_257_76_6758));
   NAND2_X1 i_257_76_6770 (.A1(n_257_76_15674), .A2(n_257_76_6535), .ZN(
      n_257_76_6759));
   OAI21_X1 i_257_76_6771 (.A(n_257_76_6759), .B1(n_257_428), .B2(n_257_76_15412), 
      .ZN(n_257_76_6760));
   NAND2_X1 i_257_76_6772 (.A1(n_257_76_6538), .A2(n_257_76_6760), .ZN(
      n_257_76_6761));
   NAND2_X1 i_257_76_6773 (.A1(n_257_76_6539), .A2(n_257_420), .ZN(n_257_76_6762));
   NOR2_X1 i_257_76_6774 (.A1(n_257_76_6761), .A2(n_257_76_6762), .ZN(
      n_257_76_6763));
   NAND2_X1 i_257_76_6775 (.A1(n_257_76_6763), .A2(n_257_76_6543), .ZN(
      n_257_76_6764));
   NAND2_X1 i_257_76_6776 (.A1(n_257_76_6488), .A2(n_257_76_6542), .ZN(
      n_257_76_6765));
   NOR2_X1 i_257_76_6777 (.A1(n_257_76_6764), .A2(n_257_76_6765), .ZN(
      n_257_76_6766));
   NAND2_X1 i_257_76_6778 (.A1(n_257_76_6758), .A2(n_257_76_6766), .ZN(
      n_257_76_6767));
   NAND2_X1 i_257_76_6779 (.A1(n_257_76_6480), .A2(n_257_76_6481), .ZN(
      n_257_76_6768));
   INV_X1 i_257_76_6780 (.A(n_257_76_6768), .ZN(n_257_76_6769));
   NAND2_X1 i_257_76_6781 (.A1(n_257_76_6531), .A2(n_257_76_6484), .ZN(
      n_257_76_6770));
   INV_X1 i_257_76_6782 (.A(n_257_76_6770), .ZN(n_257_76_6771));
   NAND2_X1 i_257_76_6783 (.A1(n_257_76_6769), .A2(n_257_76_6771), .ZN(
      n_257_76_6772));
   NOR2_X1 i_257_76_6784 (.A1(n_257_76_6767), .A2(n_257_76_6772), .ZN(
      n_257_76_6773));
   NAND2_X1 i_257_76_6785 (.A1(n_257_76_6754), .A2(n_257_76_6773), .ZN(
      n_257_76_6774));
   NAND2_X1 i_257_76_6786 (.A1(n_257_360), .A2(n_257_421), .ZN(n_257_76_6775));
   NAND2_X1 i_257_76_6787 (.A1(n_257_76_6775), .A2(n_257_76_6527), .ZN(
      n_257_76_6776));
   INV_X1 i_257_76_6788 (.A(n_257_76_6495), .ZN(n_257_76_6777));
   NOR2_X1 i_257_76_6789 (.A1(n_257_76_6776), .A2(n_257_76_6777), .ZN(
      n_257_76_6778));
   NAND2_X1 i_257_76_6790 (.A1(n_257_76_6493), .A2(n_257_76_6494), .ZN(
      n_257_76_6779));
   INV_X1 i_257_76_6791 (.A(n_257_76_6779), .ZN(n_257_76_6780));
   NAND2_X1 i_257_76_6792 (.A1(n_257_76_6778), .A2(n_257_76_6780), .ZN(
      n_257_76_6781));
   NOR2_X1 i_257_76_6793 (.A1(n_257_76_6774), .A2(n_257_76_6781), .ZN(
      n_257_76_6782));
   NAND2_X1 i_257_76_6794 (.A1(n_257_76_6749), .A2(n_257_76_6782), .ZN(
      n_257_76_6783));
   NAND2_X1 i_257_76_6795 (.A1(n_257_76_6559), .A2(n_257_76_6469), .ZN(
      n_257_76_6784));
   NOR2_X1 i_257_76_6796 (.A1(n_257_76_6783), .A2(n_257_76_6784), .ZN(
      n_257_76_6785));
   NAND2_X1 i_257_76_6797 (.A1(n_257_76_18073), .A2(n_257_76_6785), .ZN(
      n_257_76_6786));
   NAND3_X1 i_257_76_6798 (.A1(n_257_76_6528), .A2(n_257_76_6460), .A3(
      n_257_76_6491), .ZN(n_257_76_6787));
   INV_X1 i_257_76_6799 (.A(n_257_76_6787), .ZN(n_257_76_6788));
   NAND4_X1 i_257_76_6800 (.A1(n_257_124), .A2(n_257_76_6479), .A3(n_257_76_6480), 
      .A4(n_257_76_6481), .ZN(n_257_76_6789));
   INV_X1 i_257_76_6801 (.A(n_257_76_6789), .ZN(n_257_76_6790));
   NAND3_X1 i_257_76_6802 (.A1(n_257_76_6538), .A2(n_257_76_6539), .A3(
      n_257_76_17925), .ZN(n_257_76_6791));
   INV_X1 i_257_76_6803 (.A(n_257_76_6791), .ZN(n_257_76_6792));
   NAND4_X1 i_257_76_6804 (.A1(n_257_76_6487), .A2(n_257_76_6488), .A3(
      n_257_76_6542), .A4(n_257_76_6792), .ZN(n_257_76_6793));
   NOR2_X1 i_257_76_6805 (.A1(n_257_76_6793), .A2(n_257_76_6597), .ZN(
      n_257_76_6794));
   NAND4_X1 i_257_76_6806 (.A1(n_257_76_6788), .A2(n_257_76_6790), .A3(
      n_257_76_6794), .A4(n_257_76_6495), .ZN(n_257_76_6795));
   NOR2_X1 i_257_76_6807 (.A1(n_257_76_6795), .A2(n_257_76_6600), .ZN(
      n_257_76_6796));
   NAND3_X1 i_257_76_6808 (.A1(n_257_76_6796), .A2(n_257_76_6459), .A3(
      n_257_76_6498), .ZN(n_257_76_6797));
   NOR2_X1 i_257_76_6809 (.A1(n_257_76_6797), .A2(n_257_76_6500), .ZN(
      n_257_76_6798));
   NAND2_X1 i_257_76_6810 (.A1(n_257_76_18068), .A2(n_257_76_6798), .ZN(
      n_257_76_6799));
   NAND3_X1 i_257_76_6811 (.A1(n_257_76_6745), .A2(n_257_76_6786), .A3(
      n_257_76_6799), .ZN(n_257_76_6800));
   INV_X1 i_257_76_6812 (.A(n_257_76_6800), .ZN(n_257_76_6801));
   NAND2_X1 i_257_76_6813 (.A1(n_257_776), .A2(n_257_442), .ZN(n_257_76_6802));
   NOR2_X1 i_257_76_6814 (.A1(n_257_1070), .A2(n_257_76_6802), .ZN(n_257_76_6803));
   NAND4_X1 i_257_76_6815 (.A1(n_257_447), .A2(n_257_76_6487), .A3(n_257_76_6488), 
      .A4(n_257_76_6803), .ZN(n_257_76_6804));
   INV_X1 i_257_76_6816 (.A(n_257_76_6804), .ZN(n_257_76_6805));
   NAND4_X1 i_257_76_6817 (.A1(n_257_76_6805), .A2(n_257_76_6460), .A3(
      n_257_76_6491), .A4(n_257_76_6479), .ZN(n_257_76_6806));
   NOR2_X1 i_257_76_6818 (.A1(n_257_76_6621), .A2(n_257_76_6806), .ZN(
      n_257_76_6807));
   NAND2_X1 i_257_76_6819 (.A1(n_257_76_6459), .A2(n_257_76_6807), .ZN(
      n_257_76_6808));
   INV_X1 i_257_76_6820 (.A(n_257_76_6808), .ZN(n_257_76_6809));
   NAND2_X1 i_257_76_6821 (.A1(n_257_76_6809), .A2(n_257_76_6469), .ZN(
      n_257_76_6810));
   INV_X1 i_257_76_6822 (.A(n_257_76_6810), .ZN(n_257_76_6811));
   NAND4_X1 i_257_76_6823 (.A1(n_257_76_6493), .A2(n_257_76_6494), .A3(
      n_257_76_6495), .A4(n_257_86), .ZN(n_257_76_6812));
   NAND3_X1 i_257_76_6824 (.A1(n_257_76_6538), .A2(n_257_76_6539), .A3(
      n_257_76_17932), .ZN(n_257_76_6813));
   INV_X1 i_257_76_6825 (.A(n_257_76_6813), .ZN(n_257_76_6814));
   NAND4_X1 i_257_76_6826 (.A1(n_257_76_6487), .A2(n_257_76_6488), .A3(
      n_257_76_6542), .A4(n_257_76_6814), .ZN(n_257_76_6815));
   NOR2_X1 i_257_76_6827 (.A1(n_257_76_6815), .A2(n_257_76_6597), .ZN(
      n_257_76_6816));
   NAND3_X1 i_257_76_6828 (.A1(n_257_76_6589), .A2(n_257_76_6651), .A3(
      n_257_76_6816), .ZN(n_257_76_6817));
   NOR2_X1 i_257_76_6829 (.A1(n_257_76_6812), .A2(n_257_76_6817), .ZN(
      n_257_76_6818));
   NAND3_X1 i_257_76_6830 (.A1(n_257_76_6818), .A2(n_257_76_6459), .A3(
      n_257_76_6498), .ZN(n_257_76_6819));
   NOR2_X1 i_257_76_6831 (.A1(n_257_76_6819), .A2(n_257_76_6500), .ZN(
      n_257_76_6820));
   AOI22_X1 i_257_76_6832 (.A1(n_257_76_18085), .A2(n_257_76_6811), .B1(
      n_257_76_18080), .B2(n_257_76_6820), .ZN(n_257_76_6821));
   NAND3_X1 i_257_76_6833 (.A1(n_257_76_6735), .A2(n_257_76_6801), .A3(
      n_257_76_6821), .ZN(n_257_76_6822));
   NAND3_X1 i_257_76_6834 (.A1(n_257_76_18043), .A2(n_257_76_6479), .A3(
      n_257_76_6481), .ZN(n_257_76_6823));
   INV_X1 i_257_76_6835 (.A(n_257_76_6823), .ZN(n_257_76_6824));
   INV_X1 i_257_76_6836 (.A(n_257_76_6484), .ZN(n_257_76_6825));
   NAND2_X1 i_257_76_6837 (.A1(n_257_76_6487), .A2(n_257_448), .ZN(n_257_76_6826));
   NOR2_X1 i_257_76_6838 (.A1(n_257_76_6825), .A2(n_257_76_6826), .ZN(
      n_257_76_6827));
   NAND4_X1 i_257_76_6839 (.A1(n_257_76_6824), .A2(n_257_76_6827), .A3(
      n_257_76_6460), .A4(n_257_76_6491), .ZN(n_257_76_6828));
   NOR2_X1 i_257_76_6840 (.A1(n_257_76_6828), .A2(n_257_76_6496), .ZN(
      n_257_76_6829));
   NAND3_X1 i_257_76_6841 (.A1(n_257_76_6829), .A2(n_257_76_6459), .A3(n_257_680), 
      .ZN(n_257_76_6830));
   NOR2_X1 i_257_76_6842 (.A1(n_257_76_6830), .A2(n_257_76_6500), .ZN(
      n_257_76_6831));
   NAND2_X1 i_257_76_6843 (.A1(n_257_76_18079), .A2(n_257_76_6831), .ZN(
      n_257_76_6832));
   NAND4_X1 i_257_76_6844 (.A1(n_257_76_6537), .A2(n_257_76_6538), .A3(
      n_257_76_6539), .A4(n_257_425), .ZN(n_257_76_6833));
   INV_X1 i_257_76_6845 (.A(n_257_76_6833), .ZN(n_257_76_6834));
   NAND3_X1 i_257_76_6846 (.A1(n_257_76_6834), .A2(n_257_76_6488), .A3(
      n_257_76_6542), .ZN(n_257_76_6835));
   NOR2_X1 i_257_76_6847 (.A1(n_257_76_6835), .A2(n_257_76_6757), .ZN(
      n_257_76_6836));
   NAND3_X1 i_257_76_6848 (.A1(n_257_76_6836), .A2(n_257_76_6483), .A3(
      n_257_76_6534), .ZN(n_257_76_6837));
   NAND4_X1 i_257_76_6849 (.A1(n_257_76_6527), .A2(n_257_76_6528), .A3(
      n_257_76_6460), .A4(n_257_76_6491), .ZN(n_257_76_6838));
   NOR2_X1 i_257_76_6850 (.A1(n_257_76_6837), .A2(n_257_76_6838), .ZN(
      n_257_76_6839));
   NAND2_X1 i_257_76_6851 (.A1(n_257_76_6552), .A2(n_257_243), .ZN(n_257_76_6840));
   INV_X1 i_257_76_6852 (.A(n_257_76_6840), .ZN(n_257_76_6841));
   INV_X1 i_257_76_6853 (.A(n_257_76_6496), .ZN(n_257_76_6842));
   NAND3_X1 i_257_76_6854 (.A1(n_257_76_6839), .A2(n_257_76_6841), .A3(
      n_257_76_6842), .ZN(n_257_76_6843));
   INV_X1 i_257_76_6855 (.A(n_257_76_6843), .ZN(n_257_76_6844));
   NAND2_X1 i_257_76_6856 (.A1(n_257_76_6469), .A2(n_257_76_6844), .ZN(
      n_257_76_6845));
   NAND3_X1 i_257_76_6857 (.A1(n_257_76_6557), .A2(n_257_76_6459), .A3(
      n_257_76_6498), .ZN(n_257_76_6846));
   NOR2_X1 i_257_76_6858 (.A1(n_257_76_6845), .A2(n_257_76_6846), .ZN(
      n_257_76_6847));
   NAND2_X1 i_257_76_6859 (.A1(n_257_76_18064), .A2(n_257_76_6847), .ZN(
      n_257_76_6848));
   NAND4_X1 i_257_76_6860 (.A1(n_257_76_6537), .A2(n_257_76_6538), .A3(
      n_257_76_6539), .A4(n_257_421), .ZN(n_257_76_6849));
   INV_X1 i_257_76_6861 (.A(n_257_76_6849), .ZN(n_257_76_6850));
   NAND4_X1 i_257_76_6862 (.A1(n_257_76_6850), .A2(n_257_76_6488), .A3(
      n_257_76_6542), .A4(n_257_76_6543), .ZN(n_257_76_6851));
   INV_X1 i_257_76_6863 (.A(n_257_76_6851), .ZN(n_257_76_6852));
   NAND3_X1 i_257_76_6864 (.A1(n_257_76_6755), .A2(n_257_76_6546), .A3(
      n_257_76_6487), .ZN(n_257_76_6853));
   INV_X1 i_257_76_6865 (.A(n_257_76_6853), .ZN(n_257_76_6854));
   NAND3_X1 i_257_76_6866 (.A1(n_257_76_6852), .A2(n_257_76_6623), .A3(
      n_257_76_6854), .ZN(n_257_76_6855));
   NAND4_X1 i_257_76_6867 (.A1(n_257_76_6479), .A2(n_257_76_6480), .A3(
      n_257_76_6481), .A4(n_257_76_6531), .ZN(n_257_76_6856));
   NOR2_X1 i_257_76_6868 (.A1(n_257_76_6855), .A2(n_257_76_6856), .ZN(
      n_257_76_6857));
   NAND3_X1 i_257_76_6869 (.A1(n_257_360), .A2(n_257_76_6491), .A3(n_257_76_6750), 
      .ZN(n_257_76_6858));
   NOR2_X1 i_257_76_6870 (.A1(n_257_76_6586), .A2(n_257_76_6858), .ZN(
      n_257_76_6859));
   NAND3_X1 i_257_76_6871 (.A1(n_257_76_6842), .A2(n_257_76_6857), .A3(
      n_257_76_6859), .ZN(n_257_76_6860));
   INV_X1 i_257_76_6872 (.A(n_257_76_6860), .ZN(n_257_76_6861));
   NAND2_X1 i_257_76_6873 (.A1(n_257_76_6469), .A2(n_257_76_6861), .ZN(
      n_257_76_6862));
   NAND4_X1 i_257_76_6874 (.A1(n_257_76_6557), .A2(n_257_76_6459), .A3(
      n_257_76_6498), .A4(n_257_76_6747), .ZN(n_257_76_6863));
   NOR2_X1 i_257_76_6875 (.A1(n_257_76_6862), .A2(n_257_76_6863), .ZN(
      n_257_76_6864));
   NAND2_X1 i_257_76_6876 (.A1(n_257_76_18082), .A2(n_257_76_6864), .ZN(
      n_257_76_6865));
   NAND3_X1 i_257_76_6877 (.A1(n_257_76_6832), .A2(n_257_76_6848), .A3(
      n_257_76_6865), .ZN(n_257_76_6866));
   INV_X1 i_257_76_6878 (.A(n_257_76_6866), .ZN(n_257_76_6867));
   NAND4_X1 i_257_76_6879 (.A1(n_257_76_6532), .A2(n_257_76_6487), .A3(
      n_257_76_6488), .A4(n_257_76_6542), .ZN(n_257_76_6868));
   NAND2_X1 i_257_76_6880 (.A1(n_257_76_6481), .A2(n_257_76_6484), .ZN(
      n_257_76_6869));
   NOR2_X1 i_257_76_6881 (.A1(n_257_76_6868), .A2(n_257_76_6869), .ZN(
      n_257_76_6870));
   NAND3_X1 i_257_76_6882 (.A1(n_257_76_6537), .A2(n_257_76_6538), .A3(
      n_257_76_6539), .ZN(n_257_76_6871));
   INV_X1 i_257_76_6883 (.A(n_257_76_6871), .ZN(n_257_76_6872));
   NAND3_X1 i_257_76_6884 (.A1(n_257_76_6872), .A2(n_257_203), .A3(n_257_427), 
      .ZN(n_257_76_6873));
   INV_X1 i_257_76_6885 (.A(n_257_76_6873), .ZN(n_257_76_6874));
   NAND4_X1 i_257_76_6886 (.A1(n_257_76_6491), .A2(n_257_76_6874), .A3(
      n_257_76_6479), .A4(n_257_76_6480), .ZN(n_257_76_6875));
   INV_X1 i_257_76_6887 (.A(n_257_76_6875), .ZN(n_257_76_6876));
   NAND4_X1 i_257_76_6888 (.A1(n_257_76_6587), .A2(n_257_76_6870), .A3(
      n_257_76_6495), .A4(n_257_76_6876), .ZN(n_257_76_6877));
   NOR2_X1 i_257_76_6889 (.A1(n_257_76_6877), .A2(n_257_76_6600), .ZN(
      n_257_76_6878));
   NAND4_X1 i_257_76_6890 (.A1(n_257_76_6878), .A2(n_257_76_6557), .A3(
      n_257_76_6459), .A4(n_257_76_6498), .ZN(n_257_76_6879));
   NOR2_X1 i_257_76_6891 (.A1(n_257_76_6879), .A2(n_257_76_6500), .ZN(
      n_257_76_6880));
   NAND2_X1 i_257_76_6892 (.A1(n_257_76_18065), .A2(n_257_76_6880), .ZN(
      n_257_76_6881));
   NAND2_X1 i_257_76_6893 (.A1(n_257_451), .A2(n_257_76_6484), .ZN(n_257_76_6882));
   INV_X1 i_257_76_6894 (.A(n_257_463), .ZN(n_257_76_6883));
   NOR2_X1 i_257_76_6895 (.A1(n_257_76_6504), .A2(n_257_76_6883), .ZN(
      n_257_76_6884));
   NAND4_X1 i_257_76_6896 (.A1(n_257_76_6884), .A2(n_257_76_6487), .A3(
      n_257_76_6488), .A4(n_257_76_6542), .ZN(n_257_76_6885));
   NOR2_X1 i_257_76_6897 (.A1(n_257_76_6882), .A2(n_257_76_6885), .ZN(
      n_257_76_6886));
   NAND2_X1 i_257_76_6898 (.A1(n_257_76_6460), .A2(n_257_76_6491), .ZN(
      n_257_76_6887));
   INV_X1 i_257_76_6899 (.A(n_257_76_6887), .ZN(n_257_76_6888));
   NAND3_X1 i_257_76_6900 (.A1(n_257_76_6886), .A2(n_257_76_6888), .A3(
      n_257_76_6483), .ZN(n_257_76_6889));
   NOR2_X1 i_257_76_6901 (.A1(n_257_76_6889), .A2(n_257_76_6496), .ZN(
      n_257_76_6890));
   NAND3_X1 i_257_76_6902 (.A1(n_257_76_6890), .A2(n_257_76_6459), .A3(
      n_257_76_6498), .ZN(n_257_76_6891));
   NOR2_X1 i_257_76_6903 (.A1(n_257_76_6891), .A2(n_257_76_6500), .ZN(
      n_257_76_6892));
   NAND2_X1 i_257_76_6904 (.A1(n_257_76_18063), .A2(n_257_76_6892), .ZN(
      n_257_76_6893));
   NAND4_X1 i_257_76_6905 (.A1(n_257_76_6546), .A2(n_257_76_6487), .A3(
      n_257_76_6488), .A4(n_257_76_6542), .ZN(n_257_76_6894));
   NOR2_X1 i_257_76_6906 (.A1(n_257_76_6533), .A2(n_257_76_6894), .ZN(
      n_257_76_6895));
   INV_X1 i_257_76_6907 (.A(n_257_76_6537), .ZN(n_257_76_6896));
   NOR2_X1 i_257_76_6908 (.A1(n_257_76_6896), .A2(n_257_1070), .ZN(n_257_76_6897));
   NAND2_X1 i_257_76_6909 (.A1(n_257_76_6539), .A2(n_257_424), .ZN(n_257_76_6898));
   INV_X1 i_257_76_6910 (.A(n_257_76_6898), .ZN(n_257_76_6899));
   NAND3_X1 i_257_76_6911 (.A1(n_257_76_6897), .A2(n_257_76_6899), .A3(n_257_512), 
      .ZN(n_257_76_6900));
   INV_X1 i_257_76_6912 (.A(n_257_76_6900), .ZN(n_257_76_6901));
   NAND4_X1 i_257_76_6913 (.A1(n_257_76_6479), .A2(n_257_76_6480), .A3(
      n_257_76_6481), .A4(n_257_76_6901), .ZN(n_257_76_6902));
   INV_X1 i_257_76_6914 (.A(n_257_76_6902), .ZN(n_257_76_6903));
   NAND3_X1 i_257_76_6915 (.A1(n_257_76_6895), .A2(n_257_76_6888), .A3(
      n_257_76_6903), .ZN(n_257_76_6904));
   NOR2_X1 i_257_76_6916 (.A1(n_257_76_6904), .A2(n_257_76_6725), .ZN(
      n_257_76_6905));
   NAND3_X1 i_257_76_6917 (.A1(n_257_76_6551), .A2(n_257_76_6552), .A3(
      n_257_76_6493), .ZN(n_257_76_6906));
   INV_X1 i_257_76_6918 (.A(n_257_76_6906), .ZN(n_257_76_6907));
   NAND3_X1 i_257_76_6919 (.A1(n_257_76_6905), .A2(n_257_76_6498), .A3(
      n_257_76_6907), .ZN(n_257_76_6908));
   INV_X1 i_257_76_6920 (.A(n_257_76_6908), .ZN(n_257_76_6909));
   NAND3_X1 i_257_76_6921 (.A1(n_257_76_6909), .A2(n_257_76_6559), .A3(
      n_257_76_6469), .ZN(n_257_76_6910));
   INV_X1 i_257_76_6922 (.A(n_257_76_6910), .ZN(n_257_76_6911));
   NAND2_X1 i_257_76_6923 (.A1(n_257_76_18062), .A2(n_257_76_6911), .ZN(
      n_257_76_6912));
   NAND3_X1 i_257_76_6924 (.A1(n_257_76_6881), .A2(n_257_76_6893), .A3(
      n_257_76_6912), .ZN(n_257_76_6913));
   INV_X1 i_257_76_6925 (.A(n_257_76_6913), .ZN(n_257_76_6914));
   NAND2_X1 i_257_76_6926 (.A1(n_257_76_6539), .A2(n_257_422), .ZN(n_257_76_6915));
   INV_X1 i_257_76_6927 (.A(n_257_76_6915), .ZN(n_257_76_6916));
   NAND4_X1 i_257_76_6928 (.A1(n_257_76_6543), .A2(n_257_76_6897), .A3(n_257_321), 
      .A4(n_257_76_6916), .ZN(n_257_76_6917));
   INV_X1 i_257_76_6929 (.A(n_257_76_6917), .ZN(n_257_76_6918));
   NAND3_X1 i_257_76_6930 (.A1(n_257_76_6460), .A2(n_257_76_6491), .A3(
      n_257_76_6918), .ZN(n_257_76_6919));
   INV_X1 i_257_76_6931 (.A(n_257_76_6919), .ZN(n_257_76_6920));
   NAND4_X1 i_257_76_6932 (.A1(n_257_76_6750), .A2(n_257_76_6479), .A3(
      n_257_76_6480), .A4(n_257_76_6481), .ZN(n_257_76_6921));
   INV_X1 i_257_76_6933 (.A(n_257_76_6921), .ZN(n_257_76_6922));
   NAND3_X1 i_257_76_6934 (.A1(n_257_76_6895), .A2(n_257_76_6920), .A3(
      n_257_76_6922), .ZN(n_257_76_6923));
   NOR2_X1 i_257_76_6935 (.A1(n_257_76_6923), .A2(n_257_76_6725), .ZN(
      n_257_76_6924));
   NAND3_X1 i_257_76_6936 (.A1(n_257_76_6924), .A2(n_257_76_6498), .A3(
      n_257_76_6907), .ZN(n_257_76_6925));
   INV_X1 i_257_76_6937 (.A(n_257_76_6925), .ZN(n_257_76_6926));
   NAND3_X1 i_257_76_6938 (.A1(n_257_76_6926), .A2(n_257_76_6559), .A3(
      n_257_76_6469), .ZN(n_257_76_6927));
   INV_X1 i_257_76_6939 (.A(n_257_76_6927), .ZN(n_257_76_6928));
   NAND2_X1 i_257_76_6940 (.A1(n_257_342), .A2(n_257_76_6928), .ZN(n_257_76_6929));
   NAND2_X1 i_257_76_6941 (.A1(n_257_420), .A2(n_257_664), .ZN(n_257_76_6930));
   NAND2_X1 i_257_76_6942 (.A1(n_257_76_6930), .A2(n_257_76_6538), .ZN(
      n_257_76_6931));
   INV_X1 i_257_76_6943 (.A(n_257_76_6931), .ZN(n_257_76_6932));
   INV_X1 i_257_76_6944 (.A(n_257_76_6539), .ZN(n_257_76_6933));
   NAND2_X1 i_257_76_6945 (.A1(n_257_428), .A2(n_257_576), .ZN(n_257_76_6934));
   NAND3_X1 i_257_76_6946 (.A1(n_257_484), .A2(n_257_399), .A3(n_257_442), 
      .ZN(n_257_76_6935));
   INV_X1 i_257_76_6947 (.A(n_257_76_6935), .ZN(n_257_76_6936));
   NAND2_X1 i_257_76_6948 (.A1(n_257_76_6934), .A2(n_257_76_6936), .ZN(
      n_257_76_6937));
   NOR2_X1 i_257_76_6949 (.A1(n_257_76_6933), .A2(n_257_76_6937), .ZN(
      n_257_76_6938));
   NAND4_X1 i_257_76_6950 (.A1(n_257_76_6932), .A2(n_257_76_6542), .A3(
      n_257_76_6938), .A4(n_257_76_6543), .ZN(n_257_76_6939));
   INV_X1 i_257_76_6951 (.A(n_257_76_6939), .ZN(n_257_76_6940));
   INV_X1 i_257_76_6952 (.A(n_257_76_6756), .ZN(n_257_76_6941));
   NAND3_X1 i_257_76_6953 (.A1(n_257_76_6546), .A2(n_257_76_6487), .A3(
      n_257_76_6488), .ZN(n_257_76_6942));
   INV_X1 i_257_76_6954 (.A(n_257_76_6942), .ZN(n_257_76_6943));
   NAND3_X1 i_257_76_6955 (.A1(n_257_76_6940), .A2(n_257_76_6941), .A3(
      n_257_76_6943), .ZN(n_257_76_6944));
   NAND4_X1 i_257_76_6956 (.A1(n_257_76_6480), .A2(n_257_76_6481), .A3(
      n_257_76_6531), .A4(n_257_76_6484), .ZN(n_257_76_6945));
   NOR2_X1 i_257_76_6957 (.A1(n_257_76_6944), .A2(n_257_76_6945), .ZN(
      n_257_76_6946));
   NAND3_X1 i_257_76_6958 (.A1(n_257_76_6946), .A2(n_257_76_6551), .A3(
      n_257_76_6552), .ZN(n_257_76_6947));
   NAND3_X1 i_257_76_6959 (.A1(n_257_76_6495), .A2(n_257_76_6775), .A3(
      n_257_76_6527), .ZN(n_257_76_6948));
   INV_X1 i_257_76_6960 (.A(n_257_76_6948), .ZN(n_257_76_6949));
   NAND3_X1 i_257_76_6961 (.A1(n_257_76_6491), .A2(n_257_76_6750), .A3(
      n_257_76_6479), .ZN(n_257_76_6950));
   NOR2_X1 i_257_76_6962 (.A1(n_257_76_6650), .A2(n_257_76_6950), .ZN(
      n_257_76_6951));
   NAND3_X1 i_257_76_6963 (.A1(n_257_76_6780), .A2(n_257_76_6949), .A3(
      n_257_76_6951), .ZN(n_257_76_6952));
   NOR2_X1 i_257_76_6964 (.A1(n_257_76_6947), .A2(n_257_76_6952), .ZN(
      n_257_76_6953));
   NAND4_X1 i_257_76_6965 (.A1(n_257_76_6953), .A2(n_257_76_6730), .A3(
      n_257_76_6469), .A4(n_257_76_6557), .ZN(n_257_76_6954));
   INV_X1 i_257_76_6966 (.A(n_257_76_6954), .ZN(n_257_76_6955));
   NAND2_X1 i_257_76_6967 (.A1(n_257_76_18060), .A2(n_257_76_6955), .ZN(
      n_257_76_6956));
   INV_X1 i_257_76_6968 (.A(Small_Packet_Data_Size[11]), .ZN(n_257_76_6957));
   NAND2_X1 i_257_76_6969 (.A1(n_257_76_6934), .A2(n_257_76_18044), .ZN(
      n_257_76_6958));
   INV_X1 i_257_76_6970 (.A(n_257_76_6958), .ZN(n_257_76_6959));
   NAND3_X1 i_257_76_6971 (.A1(n_257_76_6959), .A2(n_257_76_6930), .A3(
      n_257_76_6538), .ZN(n_257_76_6960));
   NAND2_X1 i_257_76_6972 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[11]), 
      .ZN(n_257_76_6961));
   NAND2_X1 i_257_76_6973 (.A1(n_257_76_6960), .A2(n_257_76_6961), .ZN(
      n_257_76_6962));
   INV_X1 i_257_76_6974 (.A(n_257_76_6802), .ZN(n_257_76_6963));
   NAND2_X1 i_257_76_6975 (.A1(n_257_447), .A2(n_257_76_6963), .ZN(n_257_76_6964));
   NAND2_X1 i_257_76_6976 (.A1(n_257_712), .A2(n_257_76_15655), .ZN(
      n_257_76_6965));
   NAND4_X1 i_257_76_6977 (.A1(n_257_76_6962), .A2(n_257_76_6964), .A3(
      n_257_76_6873), .A4(n_257_76_6965), .ZN(n_257_76_6966));
   INV_X1 i_257_76_6978 (.A(n_257_76_6966), .ZN(n_257_76_6967));
   NAND2_X1 i_257_76_6979 (.A1(n_257_840), .A2(n_257_442), .ZN(n_257_76_6968));
   INV_X1 i_257_76_6980 (.A(n_257_76_6968), .ZN(n_257_76_6969));
   NAND2_X1 i_257_76_6981 (.A1(n_257_446), .A2(n_257_76_6969), .ZN(n_257_76_6970));
   NAND2_X1 i_257_76_6982 (.A1(n_257_449), .A2(n_257_76_14266), .ZN(
      n_257_76_6971));
   NAND3_X1 i_257_76_6983 (.A1(n_257_76_6917), .A2(n_257_76_6970), .A3(
      n_257_76_6971), .ZN(n_257_76_6972));
   INV_X1 i_257_76_6984 (.A(n_257_76_6972), .ZN(n_257_76_6973));
   INV_X1 i_257_76_6985 (.A(n_257_76_6461), .ZN(n_257_76_6974));
   NAND2_X1 i_257_76_6986 (.A1(n_257_440), .A2(n_257_76_6974), .ZN(n_257_76_6975));
   NAND2_X1 i_257_76_6987 (.A1(n_257_438), .A2(n_257_76_9900), .ZN(n_257_76_6976));
   NAND2_X1 i_257_76_6988 (.A1(n_257_640), .A2(n_257_76_17928), .ZN(
      n_257_76_6977));
   NAND4_X1 i_257_76_6989 (.A1(n_257_76_6975), .A2(n_257_76_6976), .A3(
      n_257_76_6977), .A4(n_257_76_6654), .ZN(n_257_76_6978));
   NAND2_X1 i_257_76_6990 (.A1(n_257_46), .A2(n_257_76_17918), .ZN(n_257_76_6979));
   NAND2_X1 i_257_76_6991 (.A1(n_257_76_6979), .A2(n_257_76_6900), .ZN(
      n_257_76_6980));
   NOR2_X1 i_257_76_6992 (.A1(n_257_76_6978), .A2(n_257_76_6980), .ZN(
      n_257_76_6981));
   NAND2_X1 i_257_76_6993 (.A1(n_257_974), .A2(n_257_442), .ZN(n_257_76_6982));
   INV_X1 i_257_76_6994 (.A(n_257_76_6982), .ZN(n_257_76_6983));
   AOI22_X1 i_257_76_6995 (.A1(n_257_441), .A2(n_257_76_6983), .B1(n_257_910), 
      .B2(n_257_76_17940), .ZN(n_257_76_6984));
   NAND4_X1 i_257_76_6996 (.A1(n_257_76_6967), .A2(n_257_76_6973), .A3(
      n_257_76_6981), .A4(n_257_76_6984), .ZN(n_257_76_6985));
   NAND2_X1 i_257_76_6997 (.A1(n_257_463), .A2(n_257_442), .ZN(n_257_76_6986));
   INV_X1 i_257_76_6998 (.A(n_257_76_6986), .ZN(n_257_76_6987));
   AOI22_X1 i_257_76_6999 (.A1(n_257_124), .A2(n_257_76_17925), .B1(n_257_451), 
      .B2(n_257_76_6987), .ZN(n_257_76_6988));
   NAND2_X1 i_257_76_7000 (.A1(n_257_872), .A2(n_257_76_17903), .ZN(
      n_257_76_6989));
   NAND2_X1 i_257_76_7001 (.A1(n_257_808), .A2(n_257_76_17952), .ZN(
      n_257_76_6990));
   NAND3_X1 i_257_76_7002 (.A1(n_257_76_6988), .A2(n_257_76_6989), .A3(
      n_257_76_6990), .ZN(n_257_76_6991));
   NOR2_X1 i_257_76_7003 (.A1(n_257_76_6985), .A2(n_257_76_6991), .ZN(
      n_257_76_6992));
   NAND2_X1 i_257_76_7004 (.A1(n_257_680), .A2(n_257_76_17958), .ZN(
      n_257_76_6993));
   NAND2_X1 i_257_76_7005 (.A1(n_257_86), .A2(n_257_76_17932), .ZN(n_257_76_6994));
   NAND2_X1 i_257_76_7006 (.A1(n_257_744), .A2(n_257_76_17935), .ZN(
      n_257_76_6995));
   NAND4_X1 i_257_76_7007 (.A1(n_257_76_6549), .A2(n_257_76_6994), .A3(
      n_257_76_6630), .A4(n_257_76_6995), .ZN(n_257_76_6996));
   INV_X1 i_257_76_7008 (.A(n_257_76_6996), .ZN(n_257_76_6997));
   NAND3_X1 i_257_76_7009 (.A1(n_257_76_6992), .A2(n_257_76_6993), .A3(
      n_257_76_6997), .ZN(n_257_76_6998));
   INV_X1 i_257_76_7010 (.A(n_257_76_6998), .ZN(n_257_76_6999));
   NAND2_X1 i_257_76_7011 (.A1(n_257_163), .A2(n_257_76_17331), .ZN(
      n_257_76_7000));
   NAND2_X1 i_257_76_7012 (.A1(n_257_1006), .A2(n_257_76_17964), .ZN(
      n_257_76_7001));
   NAND3_X1 i_257_76_7013 (.A1(n_257_76_6860), .A2(n_257_76_7000), .A3(
      n_257_76_7001), .ZN(n_257_76_7002));
   INV_X1 i_257_76_7014 (.A(n_257_76_7002), .ZN(n_257_76_7003));
   NAND2_X1 i_257_76_7015 (.A1(n_257_1038), .A2(n_257_76_17969), .ZN(
      n_257_76_7004));
   NAND4_X1 i_257_76_7016 (.A1(n_257_76_6999), .A2(n_257_76_7003), .A3(
      n_257_76_7004), .A4(n_257_76_6843), .ZN(n_257_76_7005));
   NAND3_X1 i_257_76_7017 (.A1(n_257_76_6929), .A2(n_257_76_6956), .A3(
      n_257_76_7005), .ZN(n_257_76_7006));
   INV_X1 i_257_76_7018 (.A(n_257_76_7006), .ZN(n_257_76_7007));
   NAND3_X1 i_257_76_7019 (.A1(n_257_76_6867), .A2(n_257_76_6914), .A3(
      n_257_76_7007), .ZN(n_257_76_7008));
   NOR2_X1 i_257_76_7020 (.A1(n_257_76_6822), .A2(n_257_76_7008), .ZN(
      n_257_76_7009));
   NAND2_X1 i_257_76_7021 (.A1(n_257_76_6688), .A2(n_257_76_7009), .ZN(n_11));
   NAND2_X1 i_257_76_7022 (.A1(n_257_1007), .A2(n_257_444), .ZN(n_257_76_7010));
   NAND2_X1 i_257_76_7023 (.A1(n_257_441), .A2(n_257_975), .ZN(n_257_76_7011));
   INV_X1 i_257_76_7024 (.A(n_257_1071), .ZN(n_257_76_7012));
   NAND2_X1 i_257_76_7025 (.A1(n_257_943), .A2(n_257_442), .ZN(n_257_76_7013));
   INV_X1 i_257_76_7026 (.A(n_257_76_7013), .ZN(n_257_76_7014));
   NAND3_X1 i_257_76_7027 (.A1(n_257_440), .A2(n_257_76_7012), .A3(n_257_76_7014), 
      .ZN(n_257_76_7015));
   INV_X1 i_257_76_7028 (.A(n_257_76_7015), .ZN(n_257_76_7016));
   NAND2_X1 i_257_76_7029 (.A1(n_257_76_7011), .A2(n_257_76_7016), .ZN(
      n_257_76_7017));
   INV_X1 i_257_76_7030 (.A(n_257_76_7017), .ZN(n_257_76_7018));
   NAND2_X1 i_257_76_7031 (.A1(n_257_76_7010), .A2(n_257_76_7018), .ZN(
      n_257_76_7019));
   INV_X1 i_257_76_7032 (.A(n_257_76_7019), .ZN(n_257_76_7020));
   NAND2_X1 i_257_76_7033 (.A1(n_257_1039), .A2(n_257_443), .ZN(n_257_76_7021));
   NAND2_X1 i_257_76_7034 (.A1(n_257_76_7020), .A2(n_257_76_7021), .ZN(
      n_257_76_7022));
   INV_X1 i_257_76_7035 (.A(n_257_76_7022), .ZN(n_257_76_7023));
   NAND2_X1 i_257_76_7036 (.A1(n_257_17), .A2(n_257_76_7023), .ZN(n_257_76_7024));
   NOR2_X1 i_257_76_7037 (.A1(n_257_1071), .A2(n_257_76_17412), .ZN(
      n_257_76_7025));
   INV_X1 i_257_76_7038 (.A(n_257_76_7025), .ZN(n_257_76_7026));
   NOR2_X1 i_257_76_7039 (.A1(n_257_76_7026), .A2(n_257_76_15197), .ZN(
      n_257_76_7027));
   NAND2_X1 i_257_76_7040 (.A1(n_257_1039), .A2(n_257_76_7027), .ZN(
      n_257_76_7028));
   INV_X1 i_257_76_7041 (.A(n_257_76_7028), .ZN(n_257_76_7029));
   NAND2_X1 i_257_76_7042 (.A1(n_257_76_18072), .A2(n_257_76_7029), .ZN(
      n_257_76_7030));
   NAND2_X1 i_257_76_7043 (.A1(n_257_1077), .A2(n_257_438), .ZN(n_257_76_7031));
   NAND2_X1 i_257_76_7044 (.A1(n_257_440), .A2(n_257_943), .ZN(n_257_76_7032));
   NAND2_X1 i_257_76_7045 (.A1(n_257_76_7031), .A2(n_257_76_7032), .ZN(
      n_257_76_7033));
   INV_X1 i_257_76_7046 (.A(n_257_76_7033), .ZN(n_257_76_7034));
   NAND2_X1 i_257_76_7047 (.A1(n_257_447), .A2(n_257_777), .ZN(n_257_76_7035));
   NAND3_X1 i_257_76_7048 (.A1(n_257_641), .A2(n_257_76_17928), .A3(
      n_257_76_7012), .ZN(n_257_76_7036));
   INV_X1 i_257_76_7049 (.A(n_257_76_7036), .ZN(n_257_76_7037));
   NAND3_X1 i_257_76_7050 (.A1(n_257_76_7034), .A2(n_257_76_7035), .A3(
      n_257_76_7037), .ZN(n_257_76_7038));
   NAND2_X1 i_257_76_7051 (.A1(n_257_713), .A2(n_257_435), .ZN(n_257_76_7039));
   NAND2_X1 i_257_76_7052 (.A1(n_257_446), .A2(n_257_841), .ZN(n_257_76_7040));
   NAND2_X1 i_257_76_7053 (.A1(n_257_449), .A2(n_257_1085), .ZN(n_257_76_7041));
   NAND3_X1 i_257_76_7054 (.A1(n_257_76_7039), .A2(n_257_76_7040), .A3(
      n_257_76_7041), .ZN(n_257_76_7042));
   NOR2_X1 i_257_76_7055 (.A1(n_257_76_7038), .A2(n_257_76_7042), .ZN(
      n_257_76_7043));
   NAND2_X1 i_257_76_7056 (.A1(n_257_911), .A2(n_257_439), .ZN(n_257_76_7044));
   NAND2_X1 i_257_76_7057 (.A1(n_257_76_7044), .A2(n_257_76_7011), .ZN(
      n_257_76_7045));
   INV_X1 i_257_76_7058 (.A(n_257_76_7045), .ZN(n_257_76_7046));
   NAND2_X1 i_257_76_7059 (.A1(n_257_873), .A2(n_257_445), .ZN(n_257_76_7047));
   NAND3_X1 i_257_76_7060 (.A1(n_257_76_7043), .A2(n_257_76_7046), .A3(
      n_257_76_7047), .ZN(n_257_76_7048));
   NAND2_X1 i_257_76_7061 (.A1(n_257_745), .A2(n_257_436), .ZN(n_257_76_7049));
   NAND2_X1 i_257_76_7062 (.A1(n_257_809), .A2(n_257_437), .ZN(n_257_76_7050));
   NAND2_X1 i_257_76_7063 (.A1(n_257_76_7049), .A2(n_257_76_7050), .ZN(
      n_257_76_7051));
   NOR2_X1 i_257_76_7064 (.A1(n_257_76_7048), .A2(n_257_76_7051), .ZN(
      n_257_76_7052));
   NAND2_X1 i_257_76_7065 (.A1(n_257_76_7010), .A2(n_257_76_7052), .ZN(
      n_257_76_7053));
   INV_X1 i_257_76_7066 (.A(n_257_76_7053), .ZN(n_257_76_7054));
   NAND2_X1 i_257_76_7067 (.A1(n_257_681), .A2(n_257_448), .ZN(n_257_76_7055));
   NAND3_X1 i_257_76_7068 (.A1(n_257_76_7054), .A2(n_257_76_7021), .A3(
      n_257_76_7055), .ZN(n_257_76_7056));
   INV_X1 i_257_76_7069 (.A(n_257_76_7056), .ZN(n_257_76_7057));
   NAND2_X1 i_257_76_7070 (.A1(n_257_28), .A2(n_257_76_7057), .ZN(n_257_76_7058));
   NAND3_X1 i_257_76_7071 (.A1(n_257_76_7024), .A2(n_257_76_7030), .A3(
      n_257_76_7058), .ZN(n_257_76_7059));
   NAND3_X1 i_257_76_7072 (.A1(n_257_76_7025), .A2(n_257_76_7032), .A3(n_257_841), 
      .ZN(n_257_76_7060));
   NAND2_X1 i_257_76_7073 (.A1(n_257_76_7031), .A2(n_257_446), .ZN(n_257_76_7061));
   NOR2_X1 i_257_76_7074 (.A1(n_257_76_7060), .A2(n_257_76_7061), .ZN(
      n_257_76_7062));
   NAND3_X1 i_257_76_7075 (.A1(n_257_76_7062), .A2(n_257_76_7044), .A3(
      n_257_76_7011), .ZN(n_257_76_7063));
   INV_X1 i_257_76_7076 (.A(n_257_76_7047), .ZN(n_257_76_7064));
   NOR2_X1 i_257_76_7077 (.A1(n_257_76_7063), .A2(n_257_76_7064), .ZN(
      n_257_76_7065));
   NAND2_X1 i_257_76_7078 (.A1(n_257_76_7010), .A2(n_257_76_7065), .ZN(
      n_257_76_7066));
   INV_X1 i_257_76_7079 (.A(n_257_76_7066), .ZN(n_257_76_7067));
   NAND2_X1 i_257_76_7080 (.A1(n_257_76_7067), .A2(n_257_76_7021), .ZN(
      n_257_76_7068));
   INV_X1 i_257_76_7081 (.A(n_257_76_7068), .ZN(n_257_76_7069));
   NAND2_X1 i_257_76_7082 (.A1(n_257_76_18070), .A2(n_257_76_7069), .ZN(
      n_257_76_7070));
   NAND3_X1 i_257_76_7083 (.A1(n_257_76_7025), .A2(n_257_76_7032), .A3(n_257_439), 
      .ZN(n_257_76_7071));
   INV_X1 i_257_76_7084 (.A(n_257_76_7071), .ZN(n_257_76_7072));
   NAND3_X1 i_257_76_7085 (.A1(n_257_76_7011), .A2(n_257_911), .A3(n_257_76_7072), 
      .ZN(n_257_76_7073));
   INV_X1 i_257_76_7086 (.A(n_257_76_7073), .ZN(n_257_76_7074));
   NAND2_X1 i_257_76_7087 (.A1(n_257_76_7010), .A2(n_257_76_7074), .ZN(
      n_257_76_7075));
   INV_X1 i_257_76_7088 (.A(n_257_76_7075), .ZN(n_257_76_7076));
   NAND2_X1 i_257_76_7089 (.A1(n_257_76_7076), .A2(n_257_76_7021), .ZN(
      n_257_76_7077));
   INV_X1 i_257_76_7090 (.A(n_257_76_7077), .ZN(n_257_76_7078));
   NAND2_X1 i_257_76_7091 (.A1(n_257_76_18084), .A2(n_257_76_7078), .ZN(
      n_257_76_7079));
   NAND2_X1 i_257_76_7092 (.A1(n_257_87), .A2(n_257_431), .ZN(n_257_76_7080));
   NAND2_X1 i_257_76_7093 (.A1(n_257_451), .A2(n_257_464), .ZN(n_257_76_7081));
   NAND4_X1 i_257_76_7094 (.A1(n_257_76_7080), .A2(n_257_76_7049), .A3(
      n_257_76_7050), .A4(n_257_76_7081), .ZN(n_257_76_7082));
   NAND2_X1 i_257_76_7095 (.A1(n_257_164), .A2(n_257_429), .ZN(n_257_76_7083));
   INV_X1 i_257_76_7096 (.A(n_257_76_7083), .ZN(n_257_76_7084));
   NOR2_X1 i_257_76_7097 (.A1(n_257_76_7082), .A2(n_257_76_7084), .ZN(
      n_257_76_7085));
   NAND2_X1 i_257_76_7098 (.A1(n_257_47), .A2(n_257_433), .ZN(n_257_76_7086));
   NAND4_X1 i_257_76_7099 (.A1(n_257_76_7086), .A2(n_257_284), .A3(n_257_76_7039), 
      .A4(n_257_76_7040), .ZN(n_257_76_7087));
   NAND2_X1 i_257_76_7100 (.A1(n_257_545), .A2(n_257_426), .ZN(n_257_76_7088));
   NAND2_X1 i_257_76_7101 (.A1(n_257_76_7011), .A2(n_257_76_7088), .ZN(
      n_257_76_7089));
   NOR2_X1 i_257_76_7102 (.A1(n_257_76_7087), .A2(n_257_76_7089), .ZN(
      n_257_76_7090));
   NAND2_X1 i_257_76_7103 (.A1(n_257_125), .A2(n_257_430), .ZN(n_257_76_7091));
   NAND2_X1 i_257_76_7104 (.A1(n_257_76_7091), .A2(n_257_76_7044), .ZN(
      n_257_76_7092));
   INV_X1 i_257_76_7105 (.A(n_257_76_7092), .ZN(n_257_76_7093));
   NAND2_X1 i_257_76_7106 (.A1(n_257_513), .A2(n_257_424), .ZN(n_257_76_7094));
   NAND2_X1 i_257_76_7107 (.A1(n_257_76_7032), .A2(n_257_76_7094), .ZN(
      n_257_76_7095));
   INV_X1 i_257_76_7108 (.A(n_257_76_7095), .ZN(n_257_76_7096));
   INV_X1 i_257_76_7109 (.A(n_257_577), .ZN(n_257_76_7097));
   NAND2_X1 i_257_76_7110 (.A1(n_257_76_7097), .A2(n_257_442), .ZN(n_257_76_7098));
   OAI21_X1 i_257_76_7111 (.A(n_257_76_7098), .B1(n_257_428), .B2(n_257_76_17412), 
      .ZN(n_257_76_7099));
   NAND2_X1 i_257_76_7112 (.A1(n_257_432), .A2(n_257_609), .ZN(n_257_76_7100));
   NAND4_X1 i_257_76_7113 (.A1(n_257_76_7012), .A2(n_257_76_7099), .A3(
      n_257_76_7100), .A4(n_257_423), .ZN(n_257_76_7101));
   INV_X1 i_257_76_7114 (.A(n_257_76_7101), .ZN(n_257_76_7102));
   NAND2_X1 i_257_76_7115 (.A1(n_257_641), .A2(n_257_450), .ZN(n_257_76_7103));
   NAND4_X1 i_257_76_7116 (.A1(n_257_76_7096), .A2(n_257_76_7102), .A3(
      n_257_76_7103), .A4(n_257_76_7031), .ZN(n_257_76_7104));
   NAND2_X1 i_257_76_7117 (.A1(n_257_204), .A2(n_257_427), .ZN(n_257_76_7105));
   NAND3_X1 i_257_76_7118 (.A1(n_257_76_7041), .A2(n_257_76_7035), .A3(
      n_257_76_7105), .ZN(n_257_76_7106));
   NOR2_X1 i_257_76_7119 (.A1(n_257_76_7104), .A2(n_257_76_7106), .ZN(
      n_257_76_7107));
   NAND4_X1 i_257_76_7120 (.A1(n_257_76_7090), .A2(n_257_76_7093), .A3(
      n_257_76_7107), .A4(n_257_76_7047), .ZN(n_257_76_7108));
   INV_X1 i_257_76_7121 (.A(n_257_76_7108), .ZN(n_257_76_7109));
   NAND2_X1 i_257_76_7122 (.A1(n_257_244), .A2(n_257_425), .ZN(n_257_76_7110));
   NAND4_X1 i_257_76_7123 (.A1(n_257_76_7085), .A2(n_257_76_7010), .A3(
      n_257_76_7109), .A4(n_257_76_7110), .ZN(n_257_76_7111));
   NAND2_X1 i_257_76_7124 (.A1(n_257_76_7021), .A2(n_257_76_7055), .ZN(
      n_257_76_7112));
   NOR2_X1 i_257_76_7125 (.A1(n_257_76_7111), .A2(n_257_76_7112), .ZN(
      n_257_76_7113));
   NAND2_X1 i_257_76_7126 (.A1(n_257_76_18066), .A2(n_257_76_7113), .ZN(
      n_257_76_7114));
   NAND3_X1 i_257_76_7127 (.A1(n_257_76_7070), .A2(n_257_76_7079), .A3(
      n_257_76_7114), .ZN(n_257_76_7115));
   NOR2_X1 i_257_76_7128 (.A1(n_257_76_7059), .A2(n_257_76_7115), .ZN(
      n_257_76_7116));
   NAND2_X1 i_257_76_7129 (.A1(n_257_76_7025), .A2(n_257_975), .ZN(n_257_76_7117));
   NOR2_X1 i_257_76_7130 (.A1(n_257_76_13147), .A2(n_257_76_7117), .ZN(
      n_257_76_7118));
   NAND2_X1 i_257_76_7131 (.A1(n_257_76_7010), .A2(n_257_76_7118), .ZN(
      n_257_76_7119));
   INV_X1 i_257_76_7132 (.A(n_257_76_7119), .ZN(n_257_76_7120));
   NAND2_X1 i_257_76_7133 (.A1(n_257_76_7120), .A2(n_257_76_7021), .ZN(
      n_257_76_7121));
   INV_X1 i_257_76_7134 (.A(n_257_76_7121), .ZN(n_257_76_7122));
   NAND2_X1 i_257_76_7135 (.A1(n_257_76_18071), .A2(n_257_76_7122), .ZN(
      n_257_76_7123));
   INV_X1 i_257_76_7136 (.A(n_257_76_7021), .ZN(n_257_76_7124));
   NOR2_X1 i_257_76_7137 (.A1(n_257_1071), .A2(n_257_76_15289), .ZN(
      n_257_76_7125));
   NAND4_X1 i_257_76_7138 (.A1(n_257_713), .A2(n_257_76_7031), .A3(n_257_76_7032), 
      .A4(n_257_76_7125), .ZN(n_257_76_7126));
   NAND2_X1 i_257_76_7139 (.A1(n_257_76_7040), .A2(n_257_76_7035), .ZN(
      n_257_76_7127));
   NOR2_X1 i_257_76_7140 (.A1(n_257_76_7126), .A2(n_257_76_7127), .ZN(
      n_257_76_7128));
   NAND3_X1 i_257_76_7141 (.A1(n_257_76_7128), .A2(n_257_76_7046), .A3(
      n_257_76_7047), .ZN(n_257_76_7129));
   NOR2_X1 i_257_76_7142 (.A1(n_257_76_7129), .A2(n_257_76_7051), .ZN(
      n_257_76_7130));
   NAND2_X1 i_257_76_7143 (.A1(n_257_76_7010), .A2(n_257_76_7130), .ZN(
      n_257_76_7131));
   NOR2_X1 i_257_76_7144 (.A1(n_257_76_7124), .A2(n_257_76_7131), .ZN(
      n_257_76_7132));
   NAND2_X1 i_257_76_7145 (.A1(n_257_76_18078), .A2(n_257_76_7132), .ZN(
      n_257_76_7133));
   NAND3_X1 i_257_76_7146 (.A1(n_257_76_7040), .A2(n_257_76_7041), .A3(
      n_257_76_7035), .ZN(n_257_76_7134));
   INV_X1 i_257_76_7147 (.A(n_257_76_7134), .ZN(n_257_76_7135));
   NAND2_X1 i_257_76_7148 (.A1(n_257_76_7086), .A2(n_257_76_7039), .ZN(
      n_257_76_7136));
   INV_X1 i_257_76_7149 (.A(n_257_76_7136), .ZN(n_257_76_7137));
   NAND2_X1 i_257_76_7150 (.A1(n_257_442), .A2(n_257_577), .ZN(n_257_76_7138));
   INV_X1 i_257_76_7151 (.A(n_257_76_7138), .ZN(n_257_76_7139));
   NAND2_X1 i_257_76_7152 (.A1(n_257_428), .A2(n_257_76_7139), .ZN(n_257_76_7140));
   INV_X1 i_257_76_7153 (.A(n_257_76_7140), .ZN(n_257_76_7141));
   NAND2_X1 i_257_76_7154 (.A1(n_257_76_7141), .A2(n_257_76_7100), .ZN(
      n_257_76_7142));
   NOR2_X1 i_257_76_7155 (.A1(n_257_76_7142), .A2(n_257_1071), .ZN(n_257_76_7143));
   NAND4_X1 i_257_76_7156 (.A1(n_257_76_7143), .A2(n_257_76_7103), .A3(
      n_257_76_7031), .A4(n_257_76_7032), .ZN(n_257_76_7144));
   INV_X1 i_257_76_7157 (.A(n_257_76_7144), .ZN(n_257_76_7145));
   NAND3_X1 i_257_76_7158 (.A1(n_257_76_7135), .A2(n_257_76_7137), .A3(
      n_257_76_7145), .ZN(n_257_76_7146));
   NAND3_X1 i_257_76_7159 (.A1(n_257_76_7091), .A2(n_257_76_7044), .A3(
      n_257_76_7011), .ZN(n_257_76_7147));
   NOR2_X1 i_257_76_7160 (.A1(n_257_76_7146), .A2(n_257_76_7147), .ZN(
      n_257_76_7148));
   NAND2_X1 i_257_76_7161 (.A1(n_257_76_7080), .A2(n_257_76_7049), .ZN(
      n_257_76_7149));
   INV_X1 i_257_76_7162 (.A(n_257_76_7149), .ZN(n_257_76_7150));
   NAND3_X1 i_257_76_7163 (.A1(n_257_76_7050), .A2(n_257_76_7047), .A3(
      n_257_76_7081), .ZN(n_257_76_7151));
   INV_X1 i_257_76_7164 (.A(n_257_76_7151), .ZN(n_257_76_7152));
   NAND4_X1 i_257_76_7165 (.A1(n_257_76_7148), .A2(n_257_76_7150), .A3(
      n_257_76_7152), .A4(n_257_76_7083), .ZN(n_257_76_7153));
   INV_X1 i_257_76_7166 (.A(n_257_76_7153), .ZN(n_257_76_7154));
   NAND4_X1 i_257_76_7167 (.A1(n_257_76_7154), .A2(n_257_76_7021), .A3(
      n_257_76_7055), .A4(n_257_76_7010), .ZN(n_257_76_7155));
   INV_X1 i_257_76_7168 (.A(n_257_76_7155), .ZN(n_257_76_7156));
   NAND2_X1 i_257_76_7169 (.A1(n_257_76_18074), .A2(n_257_76_7156), .ZN(
      n_257_76_7157));
   NAND3_X1 i_257_76_7170 (.A1(n_257_76_7123), .A2(n_257_76_7133), .A3(
      n_257_76_7157), .ZN(n_257_76_7158));
   NAND2_X1 i_257_76_7171 (.A1(n_257_1071), .A2(n_257_442), .ZN(n_257_76_7159));
   INV_X1 i_257_76_7172 (.A(n_257_76_7159), .ZN(n_257_76_7160));
   NAND2_X1 i_257_76_7173 (.A1(n_257_13), .A2(n_257_76_7160), .ZN(n_257_76_7161));
   NOR2_X1 i_257_76_7174 (.A1(n_257_76_17902), .A2(n_257_1071), .ZN(
      n_257_76_7162));
   NAND3_X1 i_257_76_7175 (.A1(n_257_76_7031), .A2(n_257_76_7162), .A3(
      n_257_76_7032), .ZN(n_257_76_7163));
   INV_X1 i_257_76_7176 (.A(n_257_76_7163), .ZN(n_257_76_7164));
   NAND4_X1 i_257_76_7177 (.A1(n_257_873), .A2(n_257_76_7044), .A3(n_257_76_7011), 
      .A4(n_257_76_7164), .ZN(n_257_76_7165));
   INV_X1 i_257_76_7178 (.A(n_257_76_7165), .ZN(n_257_76_7166));
   NAND2_X1 i_257_76_7179 (.A1(n_257_76_7010), .A2(n_257_76_7166), .ZN(
      n_257_76_7167));
   INV_X1 i_257_76_7180 (.A(n_257_76_7167), .ZN(n_257_76_7168));
   NAND2_X1 i_257_76_7181 (.A1(n_257_76_7168), .A2(n_257_76_7021), .ZN(
      n_257_76_7169));
   INV_X1 i_257_76_7182 (.A(n_257_76_7169), .ZN(n_257_76_7170));
   NAND2_X1 i_257_76_7183 (.A1(n_257_76_18077), .A2(n_257_76_7170), .ZN(
      n_257_76_7171));
   NAND2_X1 i_257_76_7184 (.A1(n_257_76_7161), .A2(n_257_76_7171), .ZN(
      n_257_76_7172));
   NOR2_X1 i_257_76_7185 (.A1(n_257_76_7158), .A2(n_257_76_7172), .ZN(
      n_257_76_7173));
   INV_X1 i_257_76_7186 (.A(n_257_76_7080), .ZN(n_257_76_7174));
   INV_X1 i_257_76_7187 (.A(n_257_76_7099), .ZN(n_257_76_7175));
   NOR2_X1 i_257_76_7188 (.A1(n_257_76_7175), .A2(n_257_1071), .ZN(n_257_76_7176));
   NAND2_X1 i_257_76_7189 (.A1(n_257_76_7100), .A2(n_257_426), .ZN(n_257_76_7177));
   INV_X1 i_257_76_7190 (.A(n_257_76_7177), .ZN(n_257_76_7178));
   NAND4_X1 i_257_76_7191 (.A1(n_257_76_7031), .A2(n_257_76_7176), .A3(
      n_257_76_7032), .A4(n_257_76_7178), .ZN(n_257_76_7179));
   INV_X1 i_257_76_7192 (.A(n_257_76_7179), .ZN(n_257_76_7180));
   NAND3_X1 i_257_76_7193 (.A1(n_257_545), .A2(n_257_76_7105), .A3(n_257_76_7103), 
      .ZN(n_257_76_7181));
   INV_X1 i_257_76_7194 (.A(n_257_76_7181), .ZN(n_257_76_7182));
   NAND4_X1 i_257_76_7195 (.A1(n_257_76_7180), .A2(n_257_76_7182), .A3(
      n_257_76_7086), .A4(n_257_76_7039), .ZN(n_257_76_7183));
   NOR2_X1 i_257_76_7196 (.A1(n_257_76_7174), .A2(n_257_76_7183), .ZN(
      n_257_76_7184));
   NAND3_X1 i_257_76_7197 (.A1(n_257_76_7049), .A2(n_257_76_7050), .A3(
      n_257_76_7047), .ZN(n_257_76_7185));
   INV_X1 i_257_76_7198 (.A(n_257_76_7185), .ZN(n_257_76_7186));
   NAND3_X1 i_257_76_7199 (.A1(n_257_76_7135), .A2(n_257_76_7044), .A3(
      n_257_76_7011), .ZN(n_257_76_7187));
   NAND2_X1 i_257_76_7200 (.A1(n_257_76_7081), .A2(n_257_76_7091), .ZN(
      n_257_76_7188));
   NOR2_X1 i_257_76_7201 (.A1(n_257_76_7187), .A2(n_257_76_7188), .ZN(
      n_257_76_7189));
   NAND4_X1 i_257_76_7202 (.A1(n_257_76_7184), .A2(n_257_76_7186), .A3(
      n_257_76_7189), .A4(n_257_76_7083), .ZN(n_257_76_7190));
   INV_X1 i_257_76_7203 (.A(n_257_76_7190), .ZN(n_257_76_7191));
   NAND4_X1 i_257_76_7204 (.A1(n_257_76_7191), .A2(n_257_76_7021), .A3(
      n_257_76_7055), .A4(n_257_76_7010), .ZN(n_257_76_7192));
   INV_X1 i_257_76_7205 (.A(n_257_76_7192), .ZN(n_257_76_7193));
   NAND2_X1 i_257_76_7206 (.A1(n_257_76_18076), .A2(n_257_76_7193), .ZN(
      n_257_76_7194));
   NAND2_X1 i_257_76_7207 (.A1(n_257_76_7011), .A2(n_257_76_7040), .ZN(
      n_257_76_7195));
   INV_X1 i_257_76_7208 (.A(n_257_76_7195), .ZN(n_257_76_7196));
   NOR2_X1 i_257_76_7209 (.A1(n_257_1071), .A2(n_257_76_17934), .ZN(
      n_257_76_7197));
   NAND3_X1 i_257_76_7210 (.A1(n_257_76_7031), .A2(n_257_76_7032), .A3(
      n_257_76_7197), .ZN(n_257_76_7198));
   INV_X1 i_257_76_7211 (.A(n_257_76_7035), .ZN(n_257_76_7199));
   NOR2_X1 i_257_76_7212 (.A1(n_257_76_7198), .A2(n_257_76_7199), .ZN(
      n_257_76_7200));
   NAND4_X1 i_257_76_7213 (.A1(n_257_745), .A2(n_257_76_7196), .A3(n_257_76_7200), 
      .A4(n_257_76_7044), .ZN(n_257_76_7201));
   NAND2_X1 i_257_76_7214 (.A1(n_257_76_7050), .A2(n_257_76_7047), .ZN(
      n_257_76_7202));
   NOR2_X1 i_257_76_7215 (.A1(n_257_76_7201), .A2(n_257_76_7202), .ZN(
      n_257_76_7203));
   NAND2_X1 i_257_76_7216 (.A1(n_257_76_7010), .A2(n_257_76_7203), .ZN(
      n_257_76_7204));
   NOR2_X1 i_257_76_7217 (.A1(n_257_76_7124), .A2(n_257_76_7204), .ZN(
      n_257_76_7205));
   NAND2_X1 i_257_76_7218 (.A1(n_257_76_18069), .A2(n_257_76_7205), .ZN(
      n_257_76_7206));
   NAND2_X1 i_257_76_7219 (.A1(n_257_609), .A2(n_257_442), .ZN(n_257_76_7207));
   INV_X1 i_257_76_7220 (.A(n_257_76_7207), .ZN(n_257_76_7208));
   NAND2_X1 i_257_76_7221 (.A1(n_257_432), .A2(n_257_76_7208), .ZN(n_257_76_7209));
   NOR2_X1 i_257_76_7222 (.A1(n_257_1071), .A2(n_257_76_7209), .ZN(n_257_76_7210));
   NAND4_X1 i_257_76_7223 (.A1(n_257_76_7103), .A2(n_257_76_7031), .A3(
      n_257_76_7032), .A4(n_257_76_7210), .ZN(n_257_76_7211));
   NOR2_X1 i_257_76_7224 (.A1(n_257_76_7134), .A2(n_257_76_7211), .ZN(
      n_257_76_7212));
   NAND3_X1 i_257_76_7225 (.A1(n_257_76_7011), .A2(n_257_76_7086), .A3(
      n_257_76_7039), .ZN(n_257_76_7213));
   INV_X1 i_257_76_7226 (.A(n_257_76_7213), .ZN(n_257_76_7214));
   NAND4_X1 i_257_76_7227 (.A1(n_257_76_7212), .A2(n_257_76_7214), .A3(
      n_257_76_7081), .A4(n_257_76_7044), .ZN(n_257_76_7215));
   NOR2_X1 i_257_76_7228 (.A1(n_257_76_7215), .A2(n_257_76_7185), .ZN(
      n_257_76_7216));
   NAND2_X1 i_257_76_7229 (.A1(n_257_76_7010), .A2(n_257_76_7216), .ZN(
      n_257_76_7217));
   INV_X1 i_257_76_7230 (.A(n_257_76_7217), .ZN(n_257_76_7218));
   NAND3_X1 i_257_76_7231 (.A1(n_257_76_7218), .A2(n_257_76_7021), .A3(
      n_257_76_7055), .ZN(n_257_76_7219));
   INV_X1 i_257_76_7232 (.A(n_257_76_7219), .ZN(n_257_76_7220));
   NAND2_X1 i_257_76_7233 (.A1(n_257_68), .A2(n_257_76_7220), .ZN(n_257_76_7221));
   NAND3_X1 i_257_76_7234 (.A1(n_257_76_7194), .A2(n_257_76_7206), .A3(
      n_257_76_7221), .ZN(n_257_76_7222));
   NOR2_X1 i_257_76_7235 (.A1(n_257_1071), .A2(n_257_76_17951), .ZN(
      n_257_76_7223));
   NAND3_X1 i_257_76_7236 (.A1(n_257_76_7031), .A2(n_257_76_7032), .A3(
      n_257_76_7223), .ZN(n_257_76_7224));
   INV_X1 i_257_76_7237 (.A(n_257_76_7224), .ZN(n_257_76_7225));
   NAND3_X1 i_257_76_7238 (.A1(n_257_76_7011), .A2(n_257_76_7225), .A3(
      n_257_76_7040), .ZN(n_257_76_7226));
   INV_X1 i_257_76_7239 (.A(n_257_76_7226), .ZN(n_257_76_7227));
   NAND4_X1 i_257_76_7240 (.A1(n_257_76_7227), .A2(n_257_76_7047), .A3(n_257_809), 
      .A4(n_257_76_7044), .ZN(n_257_76_7228));
   INV_X1 i_257_76_7241 (.A(n_257_76_7228), .ZN(n_257_76_7229));
   NAND2_X1 i_257_76_7242 (.A1(n_257_76_7010), .A2(n_257_76_7229), .ZN(
      n_257_76_7230));
   INV_X1 i_257_76_7243 (.A(n_257_76_7230), .ZN(n_257_76_7231));
   NAND2_X1 i_257_76_7244 (.A1(n_257_76_7231), .A2(n_257_76_7021), .ZN(
      n_257_76_7232));
   INV_X1 i_257_76_7245 (.A(n_257_76_7232), .ZN(n_257_76_7233));
   NAND2_X1 i_257_76_7246 (.A1(n_257_22), .A2(n_257_76_7233), .ZN(n_257_76_7234));
   NAND2_X1 i_257_76_7247 (.A1(n_257_444), .A2(n_257_76_7025), .ZN(n_257_76_7235));
   INV_X1 i_257_76_7248 (.A(n_257_76_7235), .ZN(n_257_76_7236));
   NAND2_X1 i_257_76_7249 (.A1(n_257_1007), .A2(n_257_76_7236), .ZN(
      n_257_76_7237));
   INV_X1 i_257_76_7250 (.A(n_257_76_7237), .ZN(n_257_76_7238));
   NAND2_X1 i_257_76_7251 (.A1(n_257_76_7021), .A2(n_257_76_7238), .ZN(
      n_257_76_7239));
   INV_X1 i_257_76_7252 (.A(n_257_76_7239), .ZN(n_257_76_7240));
   NAND2_X1 i_257_76_7253 (.A1(n_257_76_18075), .A2(n_257_76_7240), .ZN(
      n_257_76_7241));
   NAND2_X1 i_257_76_7254 (.A1(n_257_76_7234), .A2(n_257_76_7241), .ZN(
      n_257_76_7242));
   NOR2_X1 i_257_76_7255 (.A1(n_257_76_7222), .A2(n_257_76_7242), .ZN(
      n_257_76_7243));
   NAND3_X1 i_257_76_7256 (.A1(n_257_76_7116), .A2(n_257_76_7173), .A3(
      n_257_76_7243), .ZN(n_257_76_7244));
   INV_X1 i_257_76_7257 (.A(n_257_76_7244), .ZN(n_257_76_7245));
   NAND3_X1 i_257_76_7258 (.A1(n_257_76_7041), .A2(n_257_76_7035), .A3(n_257_47), 
      .ZN(n_257_76_7246));
   NOR2_X1 i_257_76_7259 (.A1(n_257_1071), .A2(n_257_76_17633), .ZN(
      n_257_76_7247));
   NAND4_X1 i_257_76_7260 (.A1(n_257_76_7103), .A2(n_257_76_7031), .A3(
      n_257_76_7032), .A4(n_257_76_7247), .ZN(n_257_76_7248));
   NOR2_X1 i_257_76_7261 (.A1(n_257_76_7246), .A2(n_257_76_7248), .ZN(
      n_257_76_7249));
   NAND3_X1 i_257_76_7262 (.A1(n_257_76_7011), .A2(n_257_76_7039), .A3(
      n_257_76_7040), .ZN(n_257_76_7250));
   INV_X1 i_257_76_7263 (.A(n_257_76_7250), .ZN(n_257_76_7251));
   NAND4_X1 i_257_76_7264 (.A1(n_257_76_7249), .A2(n_257_76_7251), .A3(
      n_257_76_7081), .A4(n_257_76_7044), .ZN(n_257_76_7252));
   NOR2_X1 i_257_76_7265 (.A1(n_257_76_7252), .A2(n_257_76_7185), .ZN(
      n_257_76_7253));
   NAND2_X1 i_257_76_7266 (.A1(n_257_76_7010), .A2(n_257_76_7253), .ZN(
      n_257_76_7254));
   INV_X1 i_257_76_7267 (.A(n_257_76_7254), .ZN(n_257_76_7255));
   NAND3_X1 i_257_76_7268 (.A1(n_257_76_7255), .A2(n_257_76_7021), .A3(
      n_257_76_7055), .ZN(n_257_76_7256));
   INV_X1 i_257_76_7269 (.A(n_257_76_7256), .ZN(n_257_76_7257));
   NAND2_X1 i_257_76_7270 (.A1(n_257_76_18081), .A2(n_257_76_7257), .ZN(
      n_257_76_7258));
   NAND2_X1 i_257_76_7271 (.A1(n_257_76_7031), .A2(n_257_449), .ZN(n_257_76_7259));
   INV_X1 i_257_76_7272 (.A(n_257_76_7259), .ZN(n_257_76_7260));
   NAND3_X1 i_257_76_7273 (.A1(n_257_76_7025), .A2(n_257_76_7032), .A3(
      n_257_1085), .ZN(n_257_76_7261));
   INV_X1 i_257_76_7274 (.A(n_257_76_7261), .ZN(n_257_76_7262));
   NAND2_X1 i_257_76_7275 (.A1(n_257_76_7260), .A2(n_257_76_7262), .ZN(
      n_257_76_7263));
   NAND3_X1 i_257_76_7276 (.A1(n_257_76_7039), .A2(n_257_76_7040), .A3(
      n_257_76_7035), .ZN(n_257_76_7264));
   NOR2_X1 i_257_76_7277 (.A1(n_257_76_7263), .A2(n_257_76_7264), .ZN(
      n_257_76_7265));
   NAND3_X1 i_257_76_7278 (.A1(n_257_76_7265), .A2(n_257_76_7046), .A3(
      n_257_76_7047), .ZN(n_257_76_7266));
   NOR2_X1 i_257_76_7279 (.A1(n_257_76_7266), .A2(n_257_76_7051), .ZN(
      n_257_76_7267));
   NAND2_X1 i_257_76_7280 (.A1(n_257_76_7010), .A2(n_257_76_7267), .ZN(
      n_257_76_7268));
   INV_X1 i_257_76_7281 (.A(n_257_76_7268), .ZN(n_257_76_7269));
   NAND3_X1 i_257_76_7282 (.A1(n_257_76_7269), .A2(n_257_76_7021), .A3(
      n_257_76_7055), .ZN(n_257_76_7270));
   INV_X1 i_257_76_7283 (.A(n_257_76_7270), .ZN(n_257_76_7271));
   NAND2_X1 i_257_76_7284 (.A1(n_257_76_18083), .A2(n_257_76_7271), .ZN(
      n_257_76_7272));
   INV_X1 i_257_76_7285 (.A(n_257_609), .ZN(n_257_76_7273));
   NAND2_X1 i_257_76_7286 (.A1(n_257_76_7273), .A2(n_257_442), .ZN(n_257_76_7274));
   OAI21_X1 i_257_76_7287 (.A(n_257_76_7274), .B1(n_257_432), .B2(n_257_76_17412), 
      .ZN(n_257_76_7275));
   NAND3_X1 i_257_76_7288 (.A1(n_257_76_7012), .A2(n_257_76_7275), .A3(n_257_429), 
      .ZN(n_257_76_7276));
   INV_X1 i_257_76_7289 (.A(n_257_76_7032), .ZN(n_257_76_7277));
   NOR2_X1 i_257_76_7290 (.A1(n_257_76_7276), .A2(n_257_76_7277), .ZN(
      n_257_76_7278));
   NAND2_X1 i_257_76_7291 (.A1(n_257_76_7103), .A2(n_257_76_7031), .ZN(
      n_257_76_7279));
   INV_X1 i_257_76_7292 (.A(n_257_76_7279), .ZN(n_257_76_7280));
   NAND4_X1 i_257_76_7293 (.A1(n_257_76_7278), .A2(n_257_76_7280), .A3(
      n_257_76_7041), .A4(n_257_76_7035), .ZN(n_257_76_7281));
   NAND4_X1 i_257_76_7294 (.A1(n_257_76_7011), .A2(n_257_76_7086), .A3(
      n_257_76_7039), .A4(n_257_76_7040), .ZN(n_257_76_7282));
   NOR2_X1 i_257_76_7295 (.A1(n_257_76_7281), .A2(n_257_76_7282), .ZN(
      n_257_76_7283));
   NAND3_X1 i_257_76_7296 (.A1(n_257_76_7081), .A2(n_257_76_7091), .A3(
      n_257_76_7044), .ZN(n_257_76_7284));
   INV_X1 i_257_76_7297 (.A(n_257_76_7284), .ZN(n_257_76_7285));
   NAND3_X1 i_257_76_7298 (.A1(n_257_76_7283), .A2(n_257_76_7285), .A3(
      n_257_76_7047), .ZN(n_257_76_7286));
   NAND4_X1 i_257_76_7299 (.A1(n_257_76_7080), .A2(n_257_164), .A3(n_257_76_7049), 
      .A4(n_257_76_7050), .ZN(n_257_76_7287));
   NOR2_X1 i_257_76_7300 (.A1(n_257_76_7286), .A2(n_257_76_7287), .ZN(
      n_257_76_7288));
   NAND4_X1 i_257_76_7301 (.A1(n_257_76_7288), .A2(n_257_76_7021), .A3(
      n_257_76_7055), .A4(n_257_76_7010), .ZN(n_257_76_7289));
   INV_X1 i_257_76_7302 (.A(n_257_76_7289), .ZN(n_257_76_7290));
   NAND2_X1 i_257_76_7303 (.A1(n_257_76_18061), .A2(n_257_76_7290), .ZN(
      n_257_76_7291));
   NAND3_X1 i_257_76_7304 (.A1(n_257_76_7258), .A2(n_257_76_7272), .A3(
      n_257_76_7291), .ZN(n_257_76_7292));
   INV_X1 i_257_76_7305 (.A(n_257_76_7292), .ZN(n_257_76_7293));
   NAND4_X1 i_257_76_7306 (.A1(n_257_76_7025), .A2(n_257_76_7032), .A3(
      n_257_1077), .A4(n_257_438), .ZN(n_257_76_7294));
   INV_X1 i_257_76_7307 (.A(n_257_76_7294), .ZN(n_257_76_7295));
   NAND3_X1 i_257_76_7308 (.A1(n_257_76_7044), .A2(n_257_76_7011), .A3(
      n_257_76_7295), .ZN(n_257_76_7296));
   INV_X1 i_257_76_7309 (.A(n_257_76_7296), .ZN(n_257_76_7297));
   NAND2_X1 i_257_76_7310 (.A1(n_257_76_7010), .A2(n_257_76_7297), .ZN(
      n_257_76_7298));
   INV_X1 i_257_76_7311 (.A(n_257_76_7298), .ZN(n_257_76_7299));
   NAND2_X1 i_257_76_7312 (.A1(n_257_76_7299), .A2(n_257_76_7021), .ZN(
      n_257_76_7300));
   INV_X1 i_257_76_7313 (.A(n_257_76_7300), .ZN(n_257_76_7301));
   NAND2_X1 i_257_76_7314 (.A1(n_257_76_18067), .A2(n_257_76_7301), .ZN(
      n_257_76_7302));
   NAND3_X1 i_257_76_7315 (.A1(n_257_76_7080), .A2(n_257_76_7049), .A3(
      n_257_76_7050), .ZN(n_257_76_7303));
   NOR2_X1 i_257_76_7316 (.A1(n_257_76_7303), .A2(n_257_76_7084), .ZN(
      n_257_76_7304));
   NAND4_X1 i_257_76_7317 (.A1(n_257_76_7105), .A2(n_257_76_7103), .A3(
      n_257_76_7031), .A4(n_257_76_7032), .ZN(n_257_76_7305));
   NAND2_X1 i_257_76_7318 (.A1(n_257_322), .A2(n_257_422), .ZN(n_257_76_7306));
   NAND2_X1 i_257_76_7319 (.A1(n_257_76_7035), .A2(n_257_76_7306), .ZN(
      n_257_76_7307));
   NOR2_X1 i_257_76_7320 (.A1(n_257_76_7305), .A2(n_257_76_7307), .ZN(
      n_257_76_7308));
   NAND2_X1 i_257_76_7321 (.A1(n_257_284), .A2(n_257_423), .ZN(n_257_76_7309));
   NAND2_X1 i_257_76_7322 (.A1(n_257_76_7044), .A2(n_257_76_7309), .ZN(
      n_257_76_7310));
   INV_X1 i_257_76_7323 (.A(n_257_76_7310), .ZN(n_257_76_7311));
   NOR2_X1 i_257_76_7324 (.A1(n_257_76_15955), .A2(n_257_577), .ZN(n_257_76_7312));
   AOI21_X1 i_257_76_7325 (.A(n_257_76_7312), .B1(n_257_76_16810), .B2(
      n_257_76_16253), .ZN(n_257_76_7313));
   NOR2_X1 i_257_76_7326 (.A1(n_257_76_7313), .A2(n_257_1071), .ZN(n_257_76_7314));
   NAND2_X1 i_257_76_7327 (.A1(n_257_420), .A2(n_257_76_7100), .ZN(n_257_76_7315));
   INV_X1 i_257_76_7328 (.A(n_257_76_7315), .ZN(n_257_76_7316));
   NAND3_X1 i_257_76_7329 (.A1(n_257_76_7314), .A2(n_257_76_7094), .A3(
      n_257_76_7316), .ZN(n_257_76_7317));
   INV_X1 i_257_76_7330 (.A(n_257_76_7317), .ZN(n_257_76_7318));
   NAND3_X1 i_257_76_7331 (.A1(n_257_76_7318), .A2(n_257_76_7011), .A3(
      n_257_76_7088), .ZN(n_257_76_7319));
   INV_X1 i_257_76_7332 (.A(n_257_76_7319), .ZN(n_257_76_7320));
   NAND4_X1 i_257_76_7333 (.A1(n_257_76_7086), .A2(n_257_76_7039), .A3(
      n_257_76_7040), .A4(n_257_76_7041), .ZN(n_257_76_7321));
   INV_X1 i_257_76_7334 (.A(n_257_76_7321), .ZN(n_257_76_7322));
   NAND4_X1 i_257_76_7335 (.A1(n_257_76_7308), .A2(n_257_76_7311), .A3(
      n_257_76_7320), .A4(n_257_76_7322), .ZN(n_257_76_7323));
   NAND2_X1 i_257_76_7336 (.A1(n_257_361), .A2(n_257_421), .ZN(n_257_76_7324));
   NAND4_X1 i_257_76_7337 (.A1(n_257_76_7324), .A2(n_257_76_7047), .A3(
      n_257_76_7081), .A4(n_257_76_7091), .ZN(n_257_76_7325));
   NOR2_X1 i_257_76_7338 (.A1(n_257_76_7323), .A2(n_257_76_7325), .ZN(
      n_257_76_7326));
   NAND4_X1 i_257_76_7339 (.A1(n_257_76_7010), .A2(n_257_76_7304), .A3(
      n_257_76_7326), .A4(n_257_76_7110), .ZN(n_257_76_7327));
   NOR2_X1 i_257_76_7340 (.A1(n_257_76_7327), .A2(n_257_76_7112), .ZN(
      n_257_76_7328));
   NAND2_X1 i_257_76_7341 (.A1(n_257_76_18073), .A2(n_257_76_7328), .ZN(
      n_257_76_7329));
   NAND2_X1 i_257_76_7342 (.A1(n_257_76_7081), .A2(n_257_76_7044), .ZN(
      n_257_76_7330));
   INV_X1 i_257_76_7343 (.A(n_257_76_7330), .ZN(n_257_76_7331));
   NAND3_X1 i_257_76_7344 (.A1(n_257_76_7012), .A2(n_257_76_7275), .A3(n_257_430), 
      .ZN(n_257_76_7332));
   INV_X1 i_257_76_7345 (.A(n_257_76_7332), .ZN(n_257_76_7333));
   NAND4_X1 i_257_76_7346 (.A1(n_257_76_7333), .A2(n_257_76_7103), .A3(
      n_257_76_7031), .A4(n_257_76_7032), .ZN(n_257_76_7334));
   NOR2_X1 i_257_76_7347 (.A1(n_257_76_7134), .A2(n_257_76_7334), .ZN(
      n_257_76_7335));
   NAND4_X1 i_257_76_7348 (.A1(n_257_76_7011), .A2(n_257_125), .A3(n_257_76_7086), 
      .A4(n_257_76_7039), .ZN(n_257_76_7336));
   INV_X1 i_257_76_7349 (.A(n_257_76_7336), .ZN(n_257_76_7337));
   NAND4_X1 i_257_76_7350 (.A1(n_257_76_7331), .A2(n_257_76_7335), .A3(
      n_257_76_7337), .A4(n_257_76_7047), .ZN(n_257_76_7338));
   NOR2_X1 i_257_76_7351 (.A1(n_257_76_7338), .A2(n_257_76_7303), .ZN(
      n_257_76_7339));
   NAND3_X1 i_257_76_7352 (.A1(n_257_76_7339), .A2(n_257_76_7055), .A3(
      n_257_76_7010), .ZN(n_257_76_7340));
   NOR2_X1 i_257_76_7353 (.A1(n_257_76_7340), .A2(n_257_76_7124), .ZN(
      n_257_76_7341));
   NAND2_X1 i_257_76_7354 (.A1(n_257_76_18068), .A2(n_257_76_7341), .ZN(
      n_257_76_7342));
   NAND3_X1 i_257_76_7355 (.A1(n_257_76_7302), .A2(n_257_76_7329), .A3(
      n_257_76_7342), .ZN(n_257_76_7343));
   INV_X1 i_257_76_7356 (.A(n_257_76_7343), .ZN(n_257_76_7344));
   NAND2_X1 i_257_76_7357 (.A1(n_257_777), .A2(n_257_442), .ZN(n_257_76_7345));
   NOR2_X1 i_257_76_7358 (.A1(n_257_1071), .A2(n_257_76_7345), .ZN(n_257_76_7346));
   NAND4_X1 i_257_76_7359 (.A1(n_257_76_7031), .A2(n_257_447), .A3(n_257_76_7346), 
      .A4(n_257_76_7032), .ZN(n_257_76_7347));
   INV_X1 i_257_76_7360 (.A(n_257_76_7040), .ZN(n_257_76_7348));
   NOR2_X1 i_257_76_7361 (.A1(n_257_76_7347), .A2(n_257_76_7348), .ZN(
      n_257_76_7349));
   NAND4_X1 i_257_76_7362 (.A1(n_257_76_7050), .A2(n_257_76_7046), .A3(
      n_257_76_7349), .A4(n_257_76_7047), .ZN(n_257_76_7350));
   INV_X1 i_257_76_7363 (.A(n_257_76_7350), .ZN(n_257_76_7351));
   NAND2_X1 i_257_76_7364 (.A1(n_257_76_7010), .A2(n_257_76_7351), .ZN(
      n_257_76_7352));
   INV_X1 i_257_76_7365 (.A(n_257_76_7352), .ZN(n_257_76_7353));
   NAND2_X1 i_257_76_7366 (.A1(n_257_76_7353), .A2(n_257_76_7021), .ZN(
      n_257_76_7354));
   INV_X1 i_257_76_7367 (.A(n_257_76_7354), .ZN(n_257_76_7355));
   NAND3_X1 i_257_76_7368 (.A1(n_257_76_7012), .A2(n_257_76_7275), .A3(n_257_431), 
      .ZN(n_257_76_7356));
   INV_X1 i_257_76_7369 (.A(n_257_76_7356), .ZN(n_257_76_7357));
   NAND4_X1 i_257_76_7370 (.A1(n_257_76_7357), .A2(n_257_76_7103), .A3(
      n_257_76_7031), .A4(n_257_76_7032), .ZN(n_257_76_7358));
   NOR2_X1 i_257_76_7371 (.A1(n_257_76_7134), .A2(n_257_76_7358), .ZN(
      n_257_76_7359));
   NAND4_X1 i_257_76_7372 (.A1(n_257_76_7359), .A2(n_257_76_7214), .A3(
      n_257_76_7081), .A4(n_257_76_7044), .ZN(n_257_76_7360));
   NAND4_X1 i_257_76_7373 (.A1(n_257_76_7049), .A2(n_257_76_7050), .A3(
      n_257_76_7047), .A4(n_257_87), .ZN(n_257_76_7361));
   NOR2_X1 i_257_76_7374 (.A1(n_257_76_7360), .A2(n_257_76_7361), .ZN(
      n_257_76_7362));
   NAND3_X1 i_257_76_7375 (.A1(n_257_76_7362), .A2(n_257_76_7055), .A3(
      n_257_76_7010), .ZN(n_257_76_7363));
   NOR2_X1 i_257_76_7376 (.A1(n_257_76_7363), .A2(n_257_76_7124), .ZN(
      n_257_76_7364));
   AOI22_X1 i_257_76_7377 (.A1(n_257_76_18085), .A2(n_257_76_7355), .B1(
      n_257_76_18080), .B2(n_257_76_7364), .ZN(n_257_76_7365));
   NAND3_X1 i_257_76_7378 (.A1(n_257_76_7293), .A2(n_257_76_7344), .A3(
      n_257_76_7365), .ZN(n_257_76_7366));
   NAND3_X1 i_257_76_7379 (.A1(n_257_76_7105), .A2(n_257_76_7103), .A3(
      n_257_76_7031), .ZN(n_257_76_7367));
   NAND2_X1 i_257_76_7380 (.A1(n_257_76_7100), .A2(n_257_421), .ZN(n_257_76_7368));
   INV_X1 i_257_76_7381 (.A(n_257_76_7368), .ZN(n_257_76_7369));
   NAND4_X1 i_257_76_7382 (.A1(n_257_76_7176), .A2(n_257_76_7032), .A3(
      n_257_76_7094), .A4(n_257_76_7369), .ZN(n_257_76_7370));
   NOR2_X1 i_257_76_7383 (.A1(n_257_76_7367), .A2(n_257_76_7370), .ZN(
      n_257_76_7371));
   NAND3_X1 i_257_76_7384 (.A1(n_257_76_7088), .A2(n_257_76_7086), .A3(
      n_257_76_7039), .ZN(n_257_76_7372));
   INV_X1 i_257_76_7385 (.A(n_257_76_7372), .ZN(n_257_76_7373));
   NAND4_X1 i_257_76_7386 (.A1(n_257_76_7040), .A2(n_257_76_7041), .A3(
      n_257_76_7035), .A4(n_257_76_7306), .ZN(n_257_76_7374));
   INV_X1 i_257_76_7387 (.A(n_257_76_7374), .ZN(n_257_76_7375));
   NAND3_X1 i_257_76_7388 (.A1(n_257_76_7371), .A2(n_257_76_7373), .A3(
      n_257_76_7375), .ZN(n_257_76_7376));
   NAND4_X1 i_257_76_7389 (.A1(n_257_361), .A2(n_257_76_7044), .A3(n_257_76_7309), 
      .A4(n_257_76_7011), .ZN(n_257_76_7377));
   NOR2_X1 i_257_76_7390 (.A1(n_257_76_7376), .A2(n_257_76_7377), .ZN(
      n_257_76_7378));
   NAND4_X1 i_257_76_7391 (.A1(n_257_76_7050), .A2(n_257_76_7047), .A3(
      n_257_76_7081), .A4(n_257_76_7091), .ZN(n_257_76_7379));
   INV_X1 i_257_76_7392 (.A(n_257_76_7379), .ZN(n_257_76_7380));
   NAND3_X1 i_257_76_7393 (.A1(n_257_76_7378), .A2(n_257_76_7150), .A3(
      n_257_76_7380), .ZN(n_257_76_7381));
   INV_X1 i_257_76_7394 (.A(n_257_76_7381), .ZN(n_257_76_7382));
   NAND2_X1 i_257_76_7395 (.A1(n_257_76_7021), .A2(n_257_76_7382), .ZN(
      n_257_76_7383));
   NAND2_X1 i_257_76_7396 (.A1(n_257_76_7110), .A2(n_257_76_7083), .ZN(
      n_257_76_7384));
   INV_X1 i_257_76_7397 (.A(n_257_76_7384), .ZN(n_257_76_7385));
   NAND3_X1 i_257_76_7398 (.A1(n_257_76_7055), .A2(n_257_76_7385), .A3(
      n_257_76_7010), .ZN(n_257_76_7386));
   NOR2_X1 i_257_76_7399 (.A1(n_257_76_7383), .A2(n_257_76_7386), .ZN(
      n_257_76_7387));
   NAND2_X1 i_257_76_7400 (.A1(n_257_76_18082), .A2(n_257_76_7387), .ZN(
      n_257_76_7388));
   NAND4_X1 i_257_76_7401 (.A1(n_257_76_7031), .A2(n_257_76_7032), .A3(n_257_204), 
      .A4(n_257_427), .ZN(n_257_76_7389));
   INV_X1 i_257_76_7402 (.A(n_257_76_7389), .ZN(n_257_76_7390));
   NAND3_X1 i_257_76_7403 (.A1(n_257_76_7012), .A2(n_257_76_7099), .A3(
      n_257_76_7100), .ZN(n_257_76_7391));
   INV_X1 i_257_76_7404 (.A(n_257_76_7391), .ZN(n_257_76_7392));
   NAND2_X1 i_257_76_7405 (.A1(n_257_76_7103), .A2(n_257_76_7392), .ZN(
      n_257_76_7393));
   INV_X1 i_257_76_7406 (.A(n_257_76_7393), .ZN(n_257_76_7394));
   NAND4_X1 i_257_76_7407 (.A1(n_257_76_7390), .A2(n_257_76_7394), .A3(
      n_257_76_7086), .A4(n_257_76_7039), .ZN(n_257_76_7395));
   INV_X1 i_257_76_7408 (.A(n_257_76_7395), .ZN(n_257_76_7396));
   NAND2_X1 i_257_76_7409 (.A1(n_257_76_7080), .A2(n_257_76_7396), .ZN(
      n_257_76_7397));
   INV_X1 i_257_76_7410 (.A(n_257_76_7397), .ZN(n_257_76_7398));
   NAND4_X1 i_257_76_7411 (.A1(n_257_76_7398), .A2(n_257_76_7186), .A3(
      n_257_76_7189), .A4(n_257_76_7083), .ZN(n_257_76_7399));
   INV_X1 i_257_76_7412 (.A(n_257_76_7399), .ZN(n_257_76_7400));
   NAND4_X1 i_257_76_7413 (.A1(n_257_76_7400), .A2(n_257_76_7021), .A3(
      n_257_76_7055), .A4(n_257_76_7010), .ZN(n_257_76_7401));
   INV_X1 i_257_76_7414 (.A(n_257_76_7401), .ZN(n_257_76_7402));
   NAND2_X1 i_257_76_7415 (.A1(n_257_76_18065), .A2(n_257_76_7402), .ZN(
      n_257_76_7403));
   INV_X1 i_257_76_7416 (.A(n_257_76_7010), .ZN(n_257_76_7404));
   NAND2_X1 i_257_76_7417 (.A1(n_257_76_7035), .A2(n_257_76_7103), .ZN(
      n_257_76_7405));
   NAND4_X1 i_257_76_7418 (.A1(n_257_76_7031), .A2(n_257_76_7025), .A3(
      n_257_76_7032), .A4(n_257_464), .ZN(n_257_76_7406));
   NOR2_X1 i_257_76_7419 (.A1(n_257_76_7405), .A2(n_257_76_7406), .ZN(
      n_257_76_7407));
   NAND2_X1 i_257_76_7420 (.A1(n_257_451), .A2(n_257_76_7011), .ZN(n_257_76_7408));
   INV_X1 i_257_76_7421 (.A(n_257_76_7408), .ZN(n_257_76_7409));
   INV_X1 i_257_76_7422 (.A(n_257_76_7042), .ZN(n_257_76_7410));
   NAND4_X1 i_257_76_7423 (.A1(n_257_76_7407), .A2(n_257_76_7409), .A3(
      n_257_76_7044), .A4(n_257_76_7410), .ZN(n_257_76_7411));
   INV_X1 i_257_76_7424 (.A(n_257_76_7411), .ZN(n_257_76_7412));
   NAND2_X1 i_257_76_7425 (.A1(n_257_76_7186), .A2(n_257_76_7412), .ZN(
      n_257_76_7413));
   NOR2_X1 i_257_76_7426 (.A1(n_257_76_7404), .A2(n_257_76_7413), .ZN(
      n_257_76_7414));
   NAND3_X1 i_257_76_7427 (.A1(n_257_76_7414), .A2(n_257_76_7021), .A3(
      n_257_76_7055), .ZN(n_257_76_7415));
   INV_X1 i_257_76_7428 (.A(n_257_76_7415), .ZN(n_257_76_7416));
   NAND2_X1 i_257_76_7429 (.A1(n_257_76_18063), .A2(n_257_76_7416), .ZN(
      n_257_76_7417));
   NAND3_X1 i_257_76_7430 (.A1(n_257_76_7388), .A2(n_257_76_7403), .A3(
      n_257_76_7417), .ZN(n_257_76_7418));
   INV_X1 i_257_76_7431 (.A(n_257_76_7418), .ZN(n_257_76_7419));
   NAND4_X1 i_257_76_7432 (.A1(n_257_76_7047), .A2(n_257_76_7081), .A3(
      n_257_76_7091), .A4(n_257_76_7044), .ZN(n_257_76_7420));
   NAND3_X1 i_257_76_7433 (.A1(n_257_76_7011), .A2(n_257_76_7088), .A3(
      n_257_76_7086), .ZN(n_257_76_7421));
   INV_X1 i_257_76_7434 (.A(n_257_76_7421), .ZN(n_257_76_7422));
   NAND2_X1 i_257_76_7435 (.A1(n_257_76_7100), .A2(n_257_424), .ZN(n_257_76_7423));
   INV_X1 i_257_76_7436 (.A(n_257_76_7423), .ZN(n_257_76_7424));
   NAND4_X1 i_257_76_7437 (.A1(n_257_76_7424), .A2(n_257_76_7012), .A3(n_257_513), 
      .A4(n_257_76_7099), .ZN(n_257_76_7425));
   INV_X1 i_257_76_7438 (.A(n_257_76_7425), .ZN(n_257_76_7426));
   NAND4_X1 i_257_76_7439 (.A1(n_257_76_7426), .A2(n_257_76_7039), .A3(
      n_257_76_7040), .A4(n_257_76_7041), .ZN(n_257_76_7427));
   INV_X1 i_257_76_7440 (.A(n_257_76_7427), .ZN(n_257_76_7428));
   NAND2_X1 i_257_76_7441 (.A1(n_257_76_7035), .A2(n_257_76_7105), .ZN(
      n_257_76_7429));
   NAND3_X1 i_257_76_7442 (.A1(n_257_76_7103), .A2(n_257_76_7031), .A3(
      n_257_76_7032), .ZN(n_257_76_7430));
   NOR2_X1 i_257_76_7443 (.A1(n_257_76_7429), .A2(n_257_76_7430), .ZN(
      n_257_76_7431));
   NAND3_X1 i_257_76_7444 (.A1(n_257_76_7422), .A2(n_257_76_7428), .A3(
      n_257_76_7431), .ZN(n_257_76_7432));
   NOR2_X1 i_257_76_7445 (.A1(n_257_76_7420), .A2(n_257_76_7432), .ZN(
      n_257_76_7433));
   NAND4_X1 i_257_76_7446 (.A1(n_257_76_7304), .A2(n_257_76_7010), .A3(
      n_257_76_7433), .A4(n_257_76_7110), .ZN(n_257_76_7434));
   NOR2_X1 i_257_76_7447 (.A1(n_257_76_7434), .A2(n_257_76_7112), .ZN(
      n_257_76_7435));
   NAND2_X1 i_257_76_7448 (.A1(n_257_76_18062), .A2(n_257_76_7435), .ZN(
      n_257_76_7436));
   INV_X1 i_257_76_7449 (.A(n_257_76_7188), .ZN(n_257_76_7437));
   INV_X1 i_257_76_7450 (.A(n_257_76_7011), .ZN(n_257_76_7438));
   NOR2_X1 i_257_76_7451 (.A1(n_257_76_7134), .A2(n_257_76_7438), .ZN(
      n_257_76_7439));
   NAND4_X1 i_257_76_7452 (.A1(n_257_76_7437), .A2(n_257_76_7439), .A3(
      n_257_76_7047), .A4(n_257_76_7311), .ZN(n_257_76_7440));
   NOR2_X1 i_257_76_7453 (.A1(n_257_76_7440), .A2(n_257_76_7303), .ZN(
      n_257_76_7441));
   NAND4_X1 i_257_76_7454 (.A1(n_257_76_7032), .A2(n_257_76_7094), .A3(n_257_322), 
      .A4(n_257_422), .ZN(n_257_76_7442));
   NOR2_X1 i_257_76_7455 (.A1(n_257_76_7442), .A2(n_257_76_7279), .ZN(
      n_257_76_7443));
   NAND2_X1 i_257_76_7456 (.A1(n_257_76_7088), .A2(n_257_76_7086), .ZN(
      n_257_76_7444));
   INV_X1 i_257_76_7457 (.A(n_257_76_7444), .ZN(n_257_76_7445));
   NAND3_X1 i_257_76_7458 (.A1(n_257_76_7039), .A2(n_257_76_7105), .A3(
      n_257_76_7392), .ZN(n_257_76_7446));
   INV_X1 i_257_76_7459 (.A(n_257_76_7446), .ZN(n_257_76_7447));
   NAND3_X1 i_257_76_7460 (.A1(n_257_76_7443), .A2(n_257_76_7445), .A3(
      n_257_76_7447), .ZN(n_257_76_7448));
   INV_X1 i_257_76_7461 (.A(n_257_76_7448), .ZN(n_257_76_7449));
   NAND2_X1 i_257_76_7462 (.A1(n_257_76_7083), .A2(n_257_76_7449), .ZN(
      n_257_76_7450));
   INV_X1 i_257_76_7463 (.A(n_257_76_7450), .ZN(n_257_76_7451));
   NAND4_X1 i_257_76_7464 (.A1(n_257_76_7441), .A2(n_257_76_7010), .A3(
      n_257_76_7110), .A4(n_257_76_7451), .ZN(n_257_76_7452));
   NOR2_X1 i_257_76_7465 (.A1(n_257_76_7452), .A2(n_257_76_7112), .ZN(
      n_257_76_7453));
   NAND2_X1 i_257_76_7466 (.A1(n_257_342), .A2(n_257_76_7453), .ZN(n_257_76_7454));
   INV_X1 i_257_76_7467 (.A(n_257_1007), .ZN(n_257_76_7455));
   OAI21_X1 i_257_76_7468 (.A(n_257_76_7108), .B1(n_257_76_7455), .B2(
      n_257_76_17963), .ZN(n_257_76_7456));
   INV_X1 i_257_76_7469 (.A(n_257_76_7456), .ZN(n_257_76_7457));
   INV_X1 i_257_76_7470 (.A(n_257_76_7345), .ZN(n_257_76_7458));
   NAND2_X1 i_257_76_7471 (.A1(n_257_447), .A2(n_257_76_7458), .ZN(n_257_76_7459));
   NAND2_X1 i_257_76_7472 (.A1(n_257_76_7459), .A2(n_257_76_7425), .ZN(
      n_257_76_7460));
   NAND3_X1 i_257_76_7473 (.A1(n_257_1077), .A2(n_257_438), .A3(n_257_442), 
      .ZN(n_257_76_7461));
   NAND2_X1 i_257_76_7474 (.A1(n_257_641), .A2(n_257_76_17928), .ZN(
      n_257_76_7462));
   NAND2_X1 i_257_76_7475 (.A1(n_257_440), .A2(n_257_76_7014), .ZN(n_257_76_7463));
   NAND3_X1 i_257_76_7476 (.A1(n_257_76_7461), .A2(n_257_76_7462), .A3(
      n_257_76_7463), .ZN(n_257_76_7464));
   NOR2_X1 i_257_76_7477 (.A1(n_257_76_7460), .A2(n_257_76_7464), .ZN(
      n_257_76_7465));
   NAND2_X1 i_257_76_7478 (.A1(n_257_47), .A2(n_257_76_17918), .ZN(n_257_76_7466));
   INV_X1 i_257_76_7479 (.A(Small_Packet_Data_Size[12]), .ZN(n_257_76_7467));
   NAND2_X1 i_257_76_7480 (.A1(n_257_428), .A2(n_257_577), .ZN(n_257_76_7468));
   NAND4_X1 i_257_76_7481 (.A1(n_257_76_7012), .A2(n_257_76_18041), .A3(
      n_257_76_7100), .A4(n_257_76_7468), .ZN(n_257_76_7469));
   NAND2_X1 i_257_76_7482 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[12]), 
      .ZN(n_257_76_7470));
   NAND2_X1 i_257_76_7483 (.A1(n_257_76_7469), .A2(n_257_76_7470), .ZN(
      n_257_76_7471));
   NAND3_X1 i_257_76_7484 (.A1(n_257_76_7317), .A2(n_257_76_7466), .A3(
      n_257_76_7471), .ZN(n_257_76_7472));
   INV_X1 i_257_76_7485 (.A(n_257_76_7472), .ZN(n_257_76_7473));
   NAND2_X1 i_257_76_7486 (.A1(n_257_713), .A2(n_257_76_15655), .ZN(
      n_257_76_7474));
   NAND2_X1 i_257_76_7487 (.A1(n_257_841), .A2(n_257_442), .ZN(n_257_76_7475));
   INV_X1 i_257_76_7488 (.A(n_257_76_7475), .ZN(n_257_76_7476));
   NAND2_X1 i_257_76_7489 (.A1(n_257_446), .A2(n_257_76_7476), .ZN(n_257_76_7477));
   NAND2_X1 i_257_76_7490 (.A1(n_257_449), .A2(n_257_76_14798), .ZN(
      n_257_76_7478));
   NAND3_X1 i_257_76_7491 (.A1(n_257_76_7474), .A2(n_257_76_7477), .A3(
      n_257_76_7478), .ZN(n_257_76_7479));
   INV_X1 i_257_76_7492 (.A(n_257_76_7479), .ZN(n_257_76_7480));
   NAND3_X1 i_257_76_7493 (.A1(n_257_76_7465), .A2(n_257_76_7473), .A3(
      n_257_76_7480), .ZN(n_257_76_7481));
   NAND2_X1 i_257_76_7494 (.A1(n_257_464), .A2(n_257_442), .ZN(n_257_76_7482));
   INV_X1 i_257_76_7495 (.A(n_257_76_7482), .ZN(n_257_76_7483));
   NAND2_X1 i_257_76_7496 (.A1(n_257_451), .A2(n_257_76_7483), .ZN(n_257_76_7484));
   NAND2_X1 i_257_76_7497 (.A1(n_257_125), .A2(n_257_76_17925), .ZN(
      n_257_76_7485));
   NAND2_X1 i_257_76_7498 (.A1(n_257_911), .A2(n_257_76_17940), .ZN(
      n_257_76_7486));
   NAND2_X1 i_257_76_7499 (.A1(n_257_975), .A2(n_257_442), .ZN(n_257_76_7487));
   INV_X1 i_257_76_7500 (.A(n_257_76_7487), .ZN(n_257_76_7488));
   NAND2_X1 i_257_76_7501 (.A1(n_257_441), .A2(n_257_76_7488), .ZN(n_257_76_7489));
   NAND4_X1 i_257_76_7502 (.A1(n_257_76_7484), .A2(n_257_76_7485), .A3(
      n_257_76_7486), .A4(n_257_76_7489), .ZN(n_257_76_7490));
   NOR2_X1 i_257_76_7503 (.A1(n_257_76_7481), .A2(n_257_76_7490), .ZN(
      n_257_76_7491));
   NAND2_X1 i_257_76_7504 (.A1(n_257_87), .A2(n_257_76_17932), .ZN(n_257_76_7492));
   NAND3_X1 i_257_76_7505 (.A1(n_257_76_7448), .A2(n_257_76_7492), .A3(
      n_257_76_7183), .ZN(n_257_76_7493));
   INV_X1 i_257_76_7506 (.A(n_257_76_7493), .ZN(n_257_76_7494));
   NAND2_X1 i_257_76_7507 (.A1(n_257_745), .A2(n_257_76_17935), .ZN(
      n_257_76_7495));
   NAND2_X1 i_257_76_7508 (.A1(n_257_809), .A2(n_257_76_17952), .ZN(
      n_257_76_7496));
   NAND2_X1 i_257_76_7509 (.A1(n_257_873), .A2(n_257_76_17903), .ZN(
      n_257_76_7497));
   NAND4_X1 i_257_76_7510 (.A1(n_257_76_7495), .A2(n_257_76_7496), .A3(
      n_257_76_7395), .A4(n_257_76_7497), .ZN(n_257_76_7498));
   INV_X1 i_257_76_7511 (.A(n_257_76_7498), .ZN(n_257_76_7499));
   NAND2_X1 i_257_76_7512 (.A1(n_257_164), .A2(n_257_76_17331), .ZN(
      n_257_76_7500));
   NAND4_X1 i_257_76_7513 (.A1(n_257_76_7491), .A2(n_257_76_7494), .A3(
      n_257_76_7499), .A4(n_257_76_7500), .ZN(n_257_76_7501));
   INV_X1 i_257_76_7514 (.A(n_257_76_7501), .ZN(n_257_76_7502));
   NAND2_X1 i_257_76_7515 (.A1(n_257_76_7457), .A2(n_257_76_7502), .ZN(
      n_257_76_7503));
   NAND2_X1 i_257_76_7516 (.A1(n_257_1039), .A2(n_257_76_17969), .ZN(
      n_257_76_7504));
   NAND2_X1 i_257_76_7517 (.A1(n_257_681), .A2(n_257_76_17958), .ZN(
      n_257_76_7505));
   NAND2_X1 i_257_76_7518 (.A1(n_257_76_7504), .A2(n_257_76_7505), .ZN(
      n_257_76_7506));
   NAND2_X1 i_257_76_7519 (.A1(n_257_76_7100), .A2(n_257_425), .ZN(n_257_76_7507));
   INV_X1 i_257_76_7520 (.A(n_257_76_7507), .ZN(n_257_76_7508));
   NAND4_X1 i_257_76_7521 (.A1(n_257_76_7031), .A2(n_257_76_7176), .A3(
      n_257_76_7032), .A4(n_257_76_7508), .ZN(n_257_76_7509));
   NAND2_X1 i_257_76_7522 (.A1(n_257_76_7105), .A2(n_257_76_7103), .ZN(
      n_257_76_7510));
   NOR2_X1 i_257_76_7523 (.A1(n_257_76_7509), .A2(n_257_76_7510), .ZN(
      n_257_76_7511));
   NAND3_X1 i_257_76_7524 (.A1(n_257_76_7511), .A2(n_257_76_7135), .A3(
      n_257_76_7137), .ZN(n_257_76_7512));
   INV_X1 i_257_76_7525 (.A(n_257_76_7089), .ZN(n_257_76_7513));
   NAND4_X1 i_257_76_7526 (.A1(n_257_76_7513), .A2(n_257_76_7081), .A3(
      n_257_76_7091), .A4(n_257_76_7044), .ZN(n_257_76_7514));
   NOR2_X1 i_257_76_7527 (.A1(n_257_76_7512), .A2(n_257_76_7514), .ZN(
      n_257_76_7515));
   NAND2_X1 i_257_76_7528 (.A1(n_257_76_7083), .A2(n_257_244), .ZN(n_257_76_7516));
   INV_X1 i_257_76_7529 (.A(n_257_76_7516), .ZN(n_257_76_7517));
   NAND4_X1 i_257_76_7530 (.A1(n_257_76_7080), .A2(n_257_76_7049), .A3(
      n_257_76_7050), .A4(n_257_76_7047), .ZN(n_257_76_7518));
   INV_X1 i_257_76_7531 (.A(n_257_76_7518), .ZN(n_257_76_7519));
   NAND3_X1 i_257_76_7532 (.A1(n_257_76_7515), .A2(n_257_76_7517), .A3(
      n_257_76_7519), .ZN(n_257_76_7520));
   NAND2_X1 i_257_76_7533 (.A1(n_257_76_7520), .A2(n_257_76_7381), .ZN(
      n_257_76_7521));
   NOR3_X1 i_257_76_7534 (.A1(n_257_76_7503), .A2(n_257_76_7506), .A3(
      n_257_76_7521), .ZN(n_257_76_7522));
   INV_X1 i_257_76_7535 (.A(n_257_76_7100), .ZN(n_257_76_7523));
   NOR2_X1 i_257_76_7536 (.A1(n_257_1071), .A2(n_257_76_7523), .ZN(n_257_76_7524));
   NAND2_X1 i_257_76_7537 (.A1(n_257_420), .A2(n_257_665), .ZN(n_257_76_7525));
   NAND3_X1 i_257_76_7538 (.A1(n_257_400), .A2(n_257_484), .A3(n_257_442), 
      .ZN(n_257_76_7526));
   INV_X1 i_257_76_7539 (.A(n_257_76_7526), .ZN(n_257_76_7527));
   NAND2_X1 i_257_76_7540 (.A1(n_257_76_7527), .A2(n_257_76_7468), .ZN(
      n_257_76_7528));
   INV_X1 i_257_76_7541 (.A(n_257_76_7528), .ZN(n_257_76_7529));
   NAND3_X1 i_257_76_7542 (.A1(n_257_76_7524), .A2(n_257_76_7525), .A3(
      n_257_76_7529), .ZN(n_257_76_7530));
   NOR2_X1 i_257_76_7543 (.A1(n_257_76_7530), .A2(n_257_76_7095), .ZN(
      n_257_76_7531));
   INV_X1 i_257_76_7544 (.A(n_257_76_7307), .ZN(n_257_76_7532));
   INV_X1 i_257_76_7545 (.A(n_257_76_7367), .ZN(n_257_76_7533));
   NAND3_X1 i_257_76_7546 (.A1(n_257_76_7531), .A2(n_257_76_7532), .A3(
      n_257_76_7533), .ZN(n_257_76_7534));
   NOR2_X1 i_257_76_7547 (.A1(n_257_76_7534), .A2(n_257_76_7321), .ZN(
      n_257_76_7535));
   NAND3_X1 i_257_76_7548 (.A1(n_257_76_7535), .A2(n_257_76_7083), .A3(
      n_257_76_7080), .ZN(n_257_76_7536));
   INV_X1 i_257_76_7549 (.A(n_257_76_7536), .ZN(n_257_76_7537));
   NAND4_X1 i_257_76_7550 (.A1(n_257_76_7044), .A2(n_257_76_7309), .A3(
      n_257_76_7011), .A4(n_257_76_7088), .ZN(n_257_76_7538));
   INV_X1 i_257_76_7551 (.A(n_257_76_7538), .ZN(n_257_76_7539));
   NAND3_X1 i_257_76_7552 (.A1(n_257_76_7539), .A2(n_257_76_7437), .A3(
      n_257_76_7047), .ZN(n_257_76_7540));
   NAND3_X1 i_257_76_7553 (.A1(n_257_76_7049), .A2(n_257_76_7050), .A3(
      n_257_76_7324), .ZN(n_257_76_7541));
   NOR2_X1 i_257_76_7554 (.A1(n_257_76_7540), .A2(n_257_76_7541), .ZN(
      n_257_76_7542));
   NAND4_X1 i_257_76_7555 (.A1(n_257_76_7537), .A2(n_257_76_7542), .A3(
      n_257_76_7010), .A4(n_257_76_7110), .ZN(n_257_76_7543));
   NOR2_X1 i_257_76_7556 (.A1(n_257_76_7543), .A2(n_257_76_7112), .ZN(
      n_257_76_7544));
   AOI21_X1 i_257_76_7557 (.A(n_257_76_7522), .B1(n_257_76_18060), .B2(
      n_257_76_7544), .ZN(n_257_76_7545));
   NAND3_X1 i_257_76_7558 (.A1(n_257_76_7436), .A2(n_257_76_7454), .A3(
      n_257_76_7545), .ZN(n_257_76_7546));
   INV_X1 i_257_76_7559 (.A(n_257_76_7546), .ZN(n_257_76_7547));
   NAND3_X1 i_257_76_7560 (.A1(n_257_76_18042), .A2(n_257_76_7039), .A3(
      n_257_76_7040), .ZN(n_257_76_7548));
   NAND2_X1 i_257_76_7561 (.A1(n_257_448), .A2(n_257_76_7012), .ZN(n_257_76_7549));
   INV_X1 i_257_76_7562 (.A(n_257_76_7549), .ZN(n_257_76_7550));
   NAND3_X1 i_257_76_7563 (.A1(n_257_76_7550), .A2(n_257_76_7035), .A3(
      n_257_76_7032), .ZN(n_257_76_7551));
   NOR2_X1 i_257_76_7564 (.A1(n_257_76_7548), .A2(n_257_76_7551), .ZN(
      n_257_76_7552));
   NAND3_X1 i_257_76_7565 (.A1(n_257_76_7552), .A2(n_257_76_7046), .A3(
      n_257_76_7047), .ZN(n_257_76_7553));
   NOR2_X1 i_257_76_7566 (.A1(n_257_76_7553), .A2(n_257_76_7051), .ZN(
      n_257_76_7554));
   NAND3_X1 i_257_76_7567 (.A1(n_257_76_7554), .A2(n_257_76_7010), .A3(n_257_681), 
      .ZN(n_257_76_7555));
   NOR2_X1 i_257_76_7568 (.A1(n_257_76_7555), .A2(n_257_76_7124), .ZN(
      n_257_76_7556));
   NAND2_X1 i_257_76_7569 (.A1(n_257_76_7055), .A2(n_257_76_7010), .ZN(
      n_257_76_7557));
   INV_X1 i_257_76_7570 (.A(n_257_76_7557), .ZN(n_257_76_7558));
   INV_X1 i_257_76_7571 (.A(n_257_76_7520), .ZN(n_257_76_7559));
   NAND3_X1 i_257_76_7572 (.A1(n_257_76_7558), .A2(n_257_76_7559), .A3(
      n_257_76_7021), .ZN(n_257_76_7560));
   INV_X1 i_257_76_7573 (.A(n_257_76_7560), .ZN(n_257_76_7561));
   AOI22_X1 i_257_76_7574 (.A1(n_257_76_18079), .A2(n_257_76_7556), .B1(
      n_257_76_18064), .B2(n_257_76_7561), .ZN(n_257_76_7562));
   NAND3_X1 i_257_76_7575 (.A1(n_257_76_7419), .A2(n_257_76_7547), .A3(
      n_257_76_7562), .ZN(n_257_76_7563));
   NOR2_X1 i_257_76_7576 (.A1(n_257_76_7366), .A2(n_257_76_7563), .ZN(
      n_257_76_7564));
   NAND2_X1 i_257_76_7577 (.A1(n_257_76_7245), .A2(n_257_76_7564), .ZN(n_12));
   NAND2_X1 i_257_76_7578 (.A1(n_257_1008), .A2(n_257_444), .ZN(n_257_76_7565));
   NAND2_X1 i_257_76_7579 (.A1(n_257_441), .A2(n_257_976), .ZN(n_257_76_7566));
   NAND2_X1 i_257_76_7580 (.A1(n_257_944), .A2(n_257_442), .ZN(n_257_76_7567));
   NOR2_X1 i_257_76_7581 (.A1(n_257_1072), .A2(n_257_76_7567), .ZN(n_257_76_7568));
   NAND2_X1 i_257_76_7582 (.A1(n_257_440), .A2(n_257_76_7568), .ZN(n_257_76_7569));
   INV_X1 i_257_76_7583 (.A(n_257_76_7569), .ZN(n_257_76_7570));
   NAND2_X1 i_257_76_7584 (.A1(n_257_76_7566), .A2(n_257_76_7570), .ZN(
      n_257_76_7571));
   INV_X1 i_257_76_7585 (.A(n_257_76_7571), .ZN(n_257_76_7572));
   NAND2_X1 i_257_76_7586 (.A1(n_257_76_7565), .A2(n_257_76_7572), .ZN(
      n_257_76_7573));
   INV_X1 i_257_76_7587 (.A(n_257_76_7573), .ZN(n_257_76_7574));
   NAND2_X1 i_257_76_7588 (.A1(n_257_1040), .A2(n_257_443), .ZN(n_257_76_7575));
   NAND2_X1 i_257_76_7589 (.A1(n_257_76_7574), .A2(n_257_76_7575), .ZN(
      n_257_76_7576));
   INV_X1 i_257_76_7590 (.A(n_257_76_7576), .ZN(n_257_76_7577));
   NAND2_X1 i_257_76_7591 (.A1(n_257_17), .A2(n_257_76_7577), .ZN(n_257_76_7578));
   NOR2_X1 i_257_76_7592 (.A1(n_257_1072), .A2(n_257_76_17412), .ZN(
      n_257_76_7579));
   NAND2_X1 i_257_76_7593 (.A1(n_257_443), .A2(n_257_76_7579), .ZN(n_257_76_7580));
   INV_X1 i_257_76_7594 (.A(n_257_76_7580), .ZN(n_257_76_7581));
   NAND2_X1 i_257_76_7595 (.A1(n_257_1040), .A2(n_257_76_7581), .ZN(
      n_257_76_7582));
   INV_X1 i_257_76_7596 (.A(n_257_76_7582), .ZN(n_257_76_7583));
   NAND2_X1 i_257_76_7597 (.A1(n_257_76_18072), .A2(n_257_76_7583), .ZN(
      n_257_76_7584));
   NAND2_X1 i_257_76_7598 (.A1(n_257_912), .A2(n_257_439), .ZN(n_257_76_7585));
   NAND2_X1 i_257_76_7599 (.A1(n_257_446), .A2(n_257_842), .ZN(n_257_76_7586));
   NAND2_X1 i_257_76_7600 (.A1(n_257_76_7585), .A2(n_257_76_7586), .ZN(
      n_257_76_7587));
   INV_X1 i_257_76_7601 (.A(n_257_76_7587), .ZN(n_257_76_7588));
   NAND2_X1 i_257_76_7602 (.A1(n_257_76_7579), .A2(n_257_450), .ZN(n_257_76_7589));
   INV_X1 i_257_76_7603 (.A(n_257_642), .ZN(n_257_76_7590));
   NOR2_X1 i_257_76_7604 (.A1(n_257_76_7589), .A2(n_257_76_7590), .ZN(
      n_257_76_7591));
   NAND2_X1 i_257_76_7605 (.A1(n_257_714), .A2(n_257_435), .ZN(n_257_76_7592));
   NAND2_X1 i_257_76_7606 (.A1(n_257_440), .A2(n_257_944), .ZN(n_257_76_7593));
   NAND2_X1 i_257_76_7607 (.A1(n_257_438), .A2(n_257_1078), .ZN(n_257_76_7594));
   NAND4_X1 i_257_76_7608 (.A1(n_257_76_7591), .A2(n_257_76_7592), .A3(
      n_257_76_7593), .A4(n_257_76_7594), .ZN(n_257_76_7595));
   INV_X1 i_257_76_7609 (.A(n_257_76_7595), .ZN(n_257_76_7596));
   NAND2_X1 i_257_76_7610 (.A1(n_257_449), .A2(n_257_1086), .ZN(n_257_76_7597));
   NAND2_X1 i_257_76_7611 (.A1(n_257_447), .A2(n_257_778), .ZN(n_257_76_7598));
   NAND2_X1 i_257_76_7612 (.A1(n_257_76_7597), .A2(n_257_76_7598), .ZN(
      n_257_76_7599));
   INV_X1 i_257_76_7613 (.A(n_257_76_7599), .ZN(n_257_76_7600));
   NAND4_X1 i_257_76_7614 (.A1(n_257_76_7588), .A2(n_257_76_7596), .A3(
      n_257_76_7600), .A4(n_257_76_7566), .ZN(n_257_76_7601));
   NAND2_X1 i_257_76_7615 (.A1(n_257_746), .A2(n_257_436), .ZN(n_257_76_7602));
   NAND2_X1 i_257_76_7616 (.A1(n_257_810), .A2(n_257_437), .ZN(n_257_76_7603));
   NAND2_X1 i_257_76_7617 (.A1(n_257_874), .A2(n_257_445), .ZN(n_257_76_7604));
   NAND3_X1 i_257_76_7618 (.A1(n_257_76_7602), .A2(n_257_76_7603), .A3(
      n_257_76_7604), .ZN(n_257_76_7605));
   NOR2_X1 i_257_76_7619 (.A1(n_257_76_7601), .A2(n_257_76_7605), .ZN(
      n_257_76_7606));
   NAND2_X1 i_257_76_7620 (.A1(n_257_682), .A2(n_257_448), .ZN(n_257_76_7607));
   NAND3_X1 i_257_76_7621 (.A1(n_257_76_7606), .A2(n_257_76_7607), .A3(
      n_257_76_7565), .ZN(n_257_76_7608));
   INV_X1 i_257_76_7622 (.A(n_257_76_7575), .ZN(n_257_76_7609));
   NOR2_X1 i_257_76_7623 (.A1(n_257_76_7608), .A2(n_257_76_7609), .ZN(
      n_257_76_7610));
   NAND2_X1 i_257_76_7624 (.A1(n_257_28), .A2(n_257_76_7610), .ZN(n_257_76_7611));
   NAND3_X1 i_257_76_7625 (.A1(n_257_76_7578), .A2(n_257_76_7584), .A3(
      n_257_76_7611), .ZN(n_257_76_7612));
   NAND2_X1 i_257_76_7626 (.A1(n_257_842), .A2(n_257_76_7579), .ZN(n_257_76_7613));
   INV_X1 i_257_76_7627 (.A(n_257_76_7613), .ZN(n_257_76_7614));
   NAND4_X1 i_257_76_7628 (.A1(n_257_446), .A2(n_257_76_7593), .A3(n_257_76_7594), 
      .A4(n_257_76_7614), .ZN(n_257_76_7615));
   INV_X1 i_257_76_7629 (.A(n_257_76_7615), .ZN(n_257_76_7616));
   NAND4_X1 i_257_76_7630 (.A1(n_257_76_7604), .A2(n_257_76_7616), .A3(
      n_257_76_7566), .A4(n_257_76_7585), .ZN(n_257_76_7617));
   INV_X1 i_257_76_7631 (.A(n_257_76_7617), .ZN(n_257_76_7618));
   NAND2_X1 i_257_76_7632 (.A1(n_257_76_7565), .A2(n_257_76_7618), .ZN(
      n_257_76_7619));
   INV_X1 i_257_76_7633 (.A(n_257_76_7619), .ZN(n_257_76_7620));
   NAND2_X1 i_257_76_7634 (.A1(n_257_76_7620), .A2(n_257_76_7575), .ZN(
      n_257_76_7621));
   INV_X1 i_257_76_7635 (.A(n_257_76_7621), .ZN(n_257_76_7622));
   NAND2_X1 i_257_76_7636 (.A1(n_257_76_18070), .A2(n_257_76_7622), .ZN(
      n_257_76_7623));
   NAND2_X1 i_257_76_7637 (.A1(n_257_439), .A2(n_257_76_7579), .ZN(n_257_76_7624));
   INV_X1 i_257_76_7638 (.A(n_257_76_7624), .ZN(n_257_76_7625));
   NAND3_X1 i_257_76_7639 (.A1(n_257_912), .A2(n_257_76_7593), .A3(n_257_76_7625), 
      .ZN(n_257_76_7626));
   INV_X1 i_257_76_7640 (.A(n_257_76_7626), .ZN(n_257_76_7627));
   NAND2_X1 i_257_76_7641 (.A1(n_257_76_7627), .A2(n_257_76_7566), .ZN(
      n_257_76_7628));
   INV_X1 i_257_76_7642 (.A(n_257_76_7628), .ZN(n_257_76_7629));
   NAND2_X1 i_257_76_7643 (.A1(n_257_76_7565), .A2(n_257_76_7629), .ZN(
      n_257_76_7630));
   INV_X1 i_257_76_7644 (.A(n_257_76_7630), .ZN(n_257_76_7631));
   NAND2_X1 i_257_76_7645 (.A1(n_257_76_7631), .A2(n_257_76_7575), .ZN(
      n_257_76_7632));
   INV_X1 i_257_76_7646 (.A(n_257_76_7632), .ZN(n_257_76_7633));
   NAND2_X1 i_257_76_7647 (.A1(n_257_76_18084), .A2(n_257_76_7633), .ZN(
      n_257_76_7634));
   NAND2_X1 i_257_76_7648 (.A1(n_257_165), .A2(n_257_429), .ZN(n_257_76_7635));
   NOR2_X1 i_257_76_7649 (.A1(n_257_1072), .A2(n_257_76_17476), .ZN(
      n_257_76_7636));
   NAND2_X1 i_257_76_7650 (.A1(n_257_432), .A2(n_257_610), .ZN(n_257_76_7637));
   INV_X1 i_257_76_7651 (.A(n_257_578), .ZN(n_257_76_7638));
   NAND2_X1 i_257_76_7652 (.A1(n_257_76_7638), .A2(n_257_442), .ZN(n_257_76_7639));
   OAI21_X1 i_257_76_7653 (.A(n_257_76_7639), .B1(n_257_428), .B2(n_257_76_17412), 
      .ZN(n_257_76_7640));
   NAND3_X1 i_257_76_7654 (.A1(n_257_76_7636), .A2(n_257_76_7637), .A3(
      n_257_76_7640), .ZN(n_257_76_7641));
   INV_X1 i_257_76_7655 (.A(n_257_76_7641), .ZN(n_257_76_7642));
   NAND2_X1 i_257_76_7656 (.A1(n_257_642), .A2(n_257_450), .ZN(n_257_76_7643));
   NAND2_X1 i_257_76_7657 (.A1(n_257_514), .A2(n_257_424), .ZN(n_257_76_7644));
   NAND3_X1 i_257_76_7658 (.A1(n_257_76_7642), .A2(n_257_76_7643), .A3(
      n_257_76_7644), .ZN(n_257_76_7645));
   NAND2_X1 i_257_76_7659 (.A1(n_257_76_7593), .A2(n_257_76_7594), .ZN(
      n_257_76_7646));
   NOR2_X1 i_257_76_7660 (.A1(n_257_76_7645), .A2(n_257_76_7646), .ZN(
      n_257_76_7647));
   NAND2_X1 i_257_76_7661 (.A1(n_257_546), .A2(n_257_426), .ZN(n_257_76_7648));
   NAND2_X1 i_257_76_7662 (.A1(n_257_48), .A2(n_257_433), .ZN(n_257_76_7649));
   NAND2_X1 i_257_76_7663 (.A1(n_257_76_7648), .A2(n_257_76_7649), .ZN(
      n_257_76_7650));
   INV_X1 i_257_76_7664 (.A(n_257_76_7650), .ZN(n_257_76_7651));
   NAND2_X1 i_257_76_7665 (.A1(n_257_205), .A2(n_257_427), .ZN(n_257_76_7652));
   NAND3_X1 i_257_76_7666 (.A1(n_257_285), .A2(n_257_76_7592), .A3(n_257_76_7652), 
      .ZN(n_257_76_7653));
   INV_X1 i_257_76_7667 (.A(n_257_76_7653), .ZN(n_257_76_7654));
   NAND4_X1 i_257_76_7668 (.A1(n_257_76_7647), .A2(n_257_76_7651), .A3(
      n_257_76_7654), .A4(n_257_76_7585), .ZN(n_257_76_7655));
   INV_X1 i_257_76_7669 (.A(n_257_76_7655), .ZN(n_257_76_7656));
   NAND2_X1 i_257_76_7670 (.A1(n_257_245), .A2(n_257_425), .ZN(n_257_76_7657));
   NAND3_X1 i_257_76_7671 (.A1(n_257_76_7635), .A2(n_257_76_7656), .A3(
      n_257_76_7657), .ZN(n_257_76_7658));
   NAND2_X1 i_257_76_7672 (.A1(n_257_76_7602), .A2(n_257_76_7603), .ZN(
      n_257_76_7659));
   INV_X1 i_257_76_7673 (.A(n_257_76_7659), .ZN(n_257_76_7660));
   NAND2_X1 i_257_76_7674 (.A1(n_257_126), .A2(n_257_430), .ZN(n_257_76_7661));
   NAND3_X1 i_257_76_7675 (.A1(n_257_76_7604), .A2(n_257_76_7661), .A3(
      n_257_76_7566), .ZN(n_257_76_7662));
   INV_X1 i_257_76_7676 (.A(n_257_76_7662), .ZN(n_257_76_7663));
   NAND3_X1 i_257_76_7677 (.A1(n_257_76_7586), .A2(n_257_76_7597), .A3(
      n_257_76_7598), .ZN(n_257_76_7664));
   NAND2_X1 i_257_76_7678 (.A1(n_257_451), .A2(n_257_465), .ZN(n_257_76_7665));
   INV_X1 i_257_76_7679 (.A(n_257_76_7665), .ZN(n_257_76_7666));
   NOR2_X1 i_257_76_7680 (.A1(n_257_76_7664), .A2(n_257_76_7666), .ZN(
      n_257_76_7667));
   NAND2_X1 i_257_76_7681 (.A1(n_257_88), .A2(n_257_431), .ZN(n_257_76_7668));
   NAND4_X1 i_257_76_7682 (.A1(n_257_76_7660), .A2(n_257_76_7663), .A3(
      n_257_76_7667), .A4(n_257_76_7668), .ZN(n_257_76_7669));
   NOR2_X1 i_257_76_7683 (.A1(n_257_76_7658), .A2(n_257_76_7669), .ZN(
      n_257_76_7670));
   NAND2_X1 i_257_76_7684 (.A1(n_257_76_7607), .A2(n_257_76_7565), .ZN(
      n_257_76_7671));
   INV_X1 i_257_76_7685 (.A(n_257_76_7671), .ZN(n_257_76_7672));
   NAND3_X1 i_257_76_7686 (.A1(n_257_76_7670), .A2(n_257_76_7672), .A3(
      n_257_76_7575), .ZN(n_257_76_7673));
   INV_X1 i_257_76_7687 (.A(n_257_76_7673), .ZN(n_257_76_7674));
   NAND2_X1 i_257_76_7688 (.A1(n_257_76_18066), .A2(n_257_76_7674), .ZN(
      n_257_76_7675));
   NAND3_X1 i_257_76_7689 (.A1(n_257_76_7623), .A2(n_257_76_7634), .A3(
      n_257_76_7675), .ZN(n_257_76_7676));
   NOR2_X1 i_257_76_7690 (.A1(n_257_76_7612), .A2(n_257_76_7676), .ZN(
      n_257_76_7677));
   NAND2_X1 i_257_76_7691 (.A1(n_257_976), .A2(n_257_76_7579), .ZN(n_257_76_7678));
   INV_X1 i_257_76_7692 (.A(n_257_76_7678), .ZN(n_257_76_7679));
   NAND2_X1 i_257_76_7693 (.A1(n_257_441), .A2(n_257_76_7679), .ZN(n_257_76_7680));
   INV_X1 i_257_76_7694 (.A(n_257_76_7680), .ZN(n_257_76_7681));
   NAND2_X1 i_257_76_7695 (.A1(n_257_76_7565), .A2(n_257_76_7681), .ZN(
      n_257_76_7682));
   INV_X1 i_257_76_7696 (.A(n_257_76_7682), .ZN(n_257_76_7683));
   NAND2_X1 i_257_76_7697 (.A1(n_257_76_7683), .A2(n_257_76_7575), .ZN(
      n_257_76_7684));
   INV_X1 i_257_76_7698 (.A(n_257_76_7684), .ZN(n_257_76_7685));
   NAND2_X1 i_257_76_7699 (.A1(n_257_76_18071), .A2(n_257_76_7685), .ZN(
      n_257_76_7686));
   NAND2_X1 i_257_76_7700 (.A1(n_257_76_7586), .A2(n_257_76_7598), .ZN(
      n_257_76_7687));
   INV_X1 i_257_76_7701 (.A(n_257_76_7687), .ZN(n_257_76_7688));
   INV_X1 i_257_76_7702 (.A(n_257_76_7579), .ZN(n_257_76_7689));
   NOR2_X1 i_257_76_7703 (.A1(n_257_76_7689), .A2(n_257_76_17760), .ZN(
      n_257_76_7690));
   NAND4_X1 i_257_76_7704 (.A1(n_257_76_7593), .A2(n_257_76_7594), .A3(n_257_714), 
      .A4(n_257_76_7690), .ZN(n_257_76_7691));
   INV_X1 i_257_76_7705 (.A(n_257_76_7691), .ZN(n_257_76_7692));
   NAND4_X1 i_257_76_7706 (.A1(n_257_76_7688), .A2(n_257_76_7692), .A3(
      n_257_76_7566), .A4(n_257_76_7585), .ZN(n_257_76_7693));
   NOR2_X1 i_257_76_7707 (.A1(n_257_76_7605), .A2(n_257_76_7693), .ZN(
      n_257_76_7694));
   NAND2_X1 i_257_76_7708 (.A1(n_257_76_7565), .A2(n_257_76_7694), .ZN(
      n_257_76_7695));
   NOR2_X1 i_257_76_7709 (.A1(n_257_76_7609), .A2(n_257_76_7695), .ZN(
      n_257_76_7696));
   NAND2_X1 i_257_76_7710 (.A1(n_257_76_18078), .A2(n_257_76_7696), .ZN(
      n_257_76_7697));
   NAND4_X1 i_257_76_7711 (.A1(n_257_76_7665), .A2(n_257_76_7585), .A3(
      n_257_76_7586), .A4(n_257_76_7597), .ZN(n_257_76_7698));
   NAND2_X1 i_257_76_7712 (.A1(n_257_76_7592), .A2(n_257_76_7593), .ZN(
      n_257_76_7699));
   INV_X1 i_257_76_7713 (.A(n_257_76_7699), .ZN(n_257_76_7700));
   NAND2_X1 i_257_76_7714 (.A1(n_257_442), .A2(n_257_578), .ZN(n_257_76_7701));
   INV_X1 i_257_76_7715 (.A(n_257_76_7701), .ZN(n_257_76_7702));
   NAND2_X1 i_257_76_7716 (.A1(n_257_428), .A2(n_257_76_7702), .ZN(n_257_76_7703));
   INV_X1 i_257_76_7717 (.A(n_257_76_7703), .ZN(n_257_76_7704));
   INV_X1 i_257_76_7718 (.A(n_257_1072), .ZN(n_257_76_7705));
   NAND2_X1 i_257_76_7719 (.A1(n_257_76_7704), .A2(n_257_76_7705), .ZN(
      n_257_76_7706));
   INV_X1 i_257_76_7720 (.A(n_257_76_7637), .ZN(n_257_76_7707));
   NOR2_X1 i_257_76_7721 (.A1(n_257_76_7706), .A2(n_257_76_7707), .ZN(
      n_257_76_7708));
   NAND3_X1 i_257_76_7722 (.A1(n_257_76_7594), .A2(n_257_76_7708), .A3(
      n_257_76_7643), .ZN(n_257_76_7709));
   INV_X1 i_257_76_7723 (.A(n_257_76_7709), .ZN(n_257_76_7710));
   NAND4_X1 i_257_76_7724 (.A1(n_257_76_7700), .A2(n_257_76_7710), .A3(
      n_257_76_7598), .A4(n_257_76_7649), .ZN(n_257_76_7711));
   NOR2_X1 i_257_76_7725 (.A1(n_257_76_7698), .A2(n_257_76_7711), .ZN(
      n_257_76_7712));
   NAND2_X1 i_257_76_7726 (.A1(n_257_76_7668), .A2(n_257_76_7602), .ZN(
      n_257_76_7713));
   INV_X1 i_257_76_7727 (.A(n_257_76_7713), .ZN(n_257_76_7714));
   NAND4_X1 i_257_76_7728 (.A1(n_257_76_7603), .A2(n_257_76_7604), .A3(
      n_257_76_7661), .A4(n_257_76_7566), .ZN(n_257_76_7715));
   INV_X1 i_257_76_7729 (.A(n_257_76_7715), .ZN(n_257_76_7716));
   NAND4_X1 i_257_76_7730 (.A1(n_257_76_7712), .A2(n_257_76_7714), .A3(
      n_257_76_7635), .A4(n_257_76_7716), .ZN(n_257_76_7717));
   INV_X1 i_257_76_7731 (.A(n_257_76_7717), .ZN(n_257_76_7718));
   NAND3_X1 i_257_76_7732 (.A1(n_257_76_7718), .A2(n_257_76_7672), .A3(
      n_257_76_7575), .ZN(n_257_76_7719));
   INV_X1 i_257_76_7733 (.A(n_257_76_7719), .ZN(n_257_76_7720));
   NAND2_X1 i_257_76_7734 (.A1(n_257_76_18074), .A2(n_257_76_7720), .ZN(
      n_257_76_7721));
   NAND3_X1 i_257_76_7735 (.A1(n_257_76_7686), .A2(n_257_76_7697), .A3(
      n_257_76_7721), .ZN(n_257_76_7722));
   NAND2_X1 i_257_76_7736 (.A1(n_257_1072), .A2(n_257_442), .ZN(n_257_76_7723));
   INV_X1 i_257_76_7737 (.A(n_257_76_7723), .ZN(n_257_76_7724));
   NAND2_X1 i_257_76_7738 (.A1(n_257_13), .A2(n_257_76_7724), .ZN(n_257_76_7725));
   NAND2_X1 i_257_76_7739 (.A1(n_257_445), .A2(n_257_76_7579), .ZN(n_257_76_7726));
   INV_X1 i_257_76_7740 (.A(n_257_76_7726), .ZN(n_257_76_7727));
   NAND3_X1 i_257_76_7741 (.A1(n_257_76_7593), .A2(n_257_76_7594), .A3(
      n_257_76_7727), .ZN(n_257_76_7728));
   INV_X1 i_257_76_7742 (.A(n_257_76_7728), .ZN(n_257_76_7729));
   NAND4_X1 i_257_76_7743 (.A1(n_257_76_7566), .A2(n_257_76_7729), .A3(n_257_874), 
      .A4(n_257_76_7585), .ZN(n_257_76_7730));
   INV_X1 i_257_76_7744 (.A(n_257_76_7730), .ZN(n_257_76_7731));
   NAND2_X1 i_257_76_7745 (.A1(n_257_76_7565), .A2(n_257_76_7731), .ZN(
      n_257_76_7732));
   INV_X1 i_257_76_7746 (.A(n_257_76_7732), .ZN(n_257_76_7733));
   NAND2_X1 i_257_76_7747 (.A1(n_257_76_7733), .A2(n_257_76_7575), .ZN(
      n_257_76_7734));
   INV_X1 i_257_76_7748 (.A(n_257_76_7734), .ZN(n_257_76_7735));
   NAND2_X1 i_257_76_7749 (.A1(n_257_76_18077), .A2(n_257_76_7735), .ZN(
      n_257_76_7736));
   NAND2_X1 i_257_76_7750 (.A1(n_257_76_7725), .A2(n_257_76_7736), .ZN(
      n_257_76_7737));
   NOR2_X1 i_257_76_7751 (.A1(n_257_76_7722), .A2(n_257_76_7737), .ZN(
      n_257_76_7738));
   INV_X1 i_257_76_7752 (.A(n_257_76_7668), .ZN(n_257_76_7739));
   NAND2_X1 i_257_76_7753 (.A1(n_257_76_7649), .A2(n_257_76_7592), .ZN(
      n_257_76_7740));
   INV_X1 i_257_76_7754 (.A(n_257_76_7740), .ZN(n_257_76_7741));
   NAND3_X1 i_257_76_7755 (.A1(n_257_76_7652), .A2(n_257_76_7593), .A3(
      n_257_76_7594), .ZN(n_257_76_7742));
   INV_X1 i_257_76_7756 (.A(n_257_76_7742), .ZN(n_257_76_7743));
   NOR2_X1 i_257_76_7757 (.A1(n_257_1072), .A2(n_257_76_17564), .ZN(
      n_257_76_7744));
   NAND3_X1 i_257_76_7758 (.A1(n_257_76_7744), .A2(n_257_76_7637), .A3(
      n_257_76_7640), .ZN(n_257_76_7745));
   INV_X1 i_257_76_7759 (.A(n_257_76_7745), .ZN(n_257_76_7746));
   NAND3_X1 i_257_76_7760 (.A1(n_257_546), .A2(n_257_76_7746), .A3(n_257_76_7643), 
      .ZN(n_257_76_7747));
   INV_X1 i_257_76_7761 (.A(n_257_76_7747), .ZN(n_257_76_7748));
   NAND4_X1 i_257_76_7762 (.A1(n_257_76_7741), .A2(n_257_76_7743), .A3(
      n_257_76_7748), .A4(n_257_76_7585), .ZN(n_257_76_7749));
   NOR2_X1 i_257_76_7763 (.A1(n_257_76_7739), .A2(n_257_76_7749), .ZN(
      n_257_76_7750));
   INV_X1 i_257_76_7764 (.A(n_257_76_7605), .ZN(n_257_76_7751));
   NAND3_X1 i_257_76_7765 (.A1(n_257_76_7661), .A2(n_257_76_7566), .A3(
      n_257_76_7665), .ZN(n_257_76_7752));
   NOR2_X1 i_257_76_7766 (.A1(n_257_76_7752), .A2(n_257_76_7664), .ZN(
      n_257_76_7753));
   NAND4_X1 i_257_76_7767 (.A1(n_257_76_7750), .A2(n_257_76_7635), .A3(
      n_257_76_7751), .A4(n_257_76_7753), .ZN(n_257_76_7754));
   INV_X1 i_257_76_7768 (.A(n_257_76_7754), .ZN(n_257_76_7755));
   NAND3_X1 i_257_76_7769 (.A1(n_257_76_7755), .A2(n_257_76_7672), .A3(
      n_257_76_7575), .ZN(n_257_76_7756));
   INV_X1 i_257_76_7770 (.A(n_257_76_7756), .ZN(n_257_76_7757));
   NAND2_X1 i_257_76_7771 (.A1(n_257_76_18076), .A2(n_257_76_7757), .ZN(
      n_257_76_7758));
   NAND3_X1 i_257_76_7772 (.A1(n_257_76_7603), .A2(n_257_76_7604), .A3(n_257_746), 
      .ZN(n_257_76_7759));
   NOR2_X1 i_257_76_7773 (.A1(n_257_76_7689), .A2(n_257_76_8311), .ZN(
      n_257_76_7760));
   NAND3_X1 i_257_76_7774 (.A1(n_257_76_7593), .A2(n_257_76_7594), .A3(
      n_257_76_7760), .ZN(n_257_76_7761));
   INV_X1 i_257_76_7775 (.A(n_257_76_7761), .ZN(n_257_76_7762));
   NAND4_X1 i_257_76_7776 (.A1(n_257_76_7688), .A2(n_257_76_7566), .A3(
      n_257_76_7585), .A4(n_257_76_7762), .ZN(n_257_76_7763));
   NOR2_X1 i_257_76_7777 (.A1(n_257_76_7759), .A2(n_257_76_7763), .ZN(
      n_257_76_7764));
   NAND2_X1 i_257_76_7778 (.A1(n_257_76_7565), .A2(n_257_76_7764), .ZN(
      n_257_76_7765));
   NOR2_X1 i_257_76_7779 (.A1(n_257_76_7609), .A2(n_257_76_7765), .ZN(
      n_257_76_7766));
   NAND2_X1 i_257_76_7780 (.A1(n_257_76_18069), .A2(n_257_76_7766), .ZN(
      n_257_76_7767));
   NAND4_X1 i_257_76_7781 (.A1(n_257_76_7585), .A2(n_257_76_7586), .A3(
      n_257_76_7597), .A4(n_257_76_7598), .ZN(n_257_76_7768));
   INV_X1 i_257_76_7782 (.A(n_257_76_7768), .ZN(n_257_76_7769));
   NAND2_X1 i_257_76_7783 (.A1(n_257_76_7566), .A2(n_257_76_7665), .ZN(
      n_257_76_7770));
   INV_X1 i_257_76_7784 (.A(n_257_76_7770), .ZN(n_257_76_7771));
   NAND2_X1 i_257_76_7785 (.A1(n_257_610), .A2(n_257_442), .ZN(n_257_76_7772));
   INV_X1 i_257_76_7786 (.A(n_257_76_7772), .ZN(n_257_76_7773));
   NAND3_X1 i_257_76_7787 (.A1(n_257_76_7705), .A2(n_257_432), .A3(n_257_76_7773), 
      .ZN(n_257_76_7774));
   INV_X1 i_257_76_7788 (.A(n_257_76_7774), .ZN(n_257_76_7775));
   NAND4_X1 i_257_76_7789 (.A1(n_257_76_7593), .A2(n_257_76_7594), .A3(
      n_257_76_7643), .A4(n_257_76_7775), .ZN(n_257_76_7776));
   NOR2_X1 i_257_76_7790 (.A1(n_257_76_7776), .A2(n_257_76_7740), .ZN(
      n_257_76_7777));
   NAND3_X1 i_257_76_7791 (.A1(n_257_76_7769), .A2(n_257_76_7771), .A3(
      n_257_76_7777), .ZN(n_257_76_7778));
   NOR2_X1 i_257_76_7792 (.A1(n_257_76_7778), .A2(n_257_76_7605), .ZN(
      n_257_76_7779));
   NAND3_X1 i_257_76_7793 (.A1(n_257_76_7779), .A2(n_257_76_7607), .A3(
      n_257_76_7565), .ZN(n_257_76_7780));
   NOR2_X1 i_257_76_7794 (.A1(n_257_76_7780), .A2(n_257_76_7609), .ZN(
      n_257_76_7781));
   NAND2_X1 i_257_76_7795 (.A1(n_257_68), .A2(n_257_76_7781), .ZN(n_257_76_7782));
   NAND3_X1 i_257_76_7796 (.A1(n_257_76_7758), .A2(n_257_76_7767), .A3(
      n_257_76_7782), .ZN(n_257_76_7783));
   NOR2_X1 i_257_76_7797 (.A1(n_257_76_7689), .A2(n_257_76_15924), .ZN(
      n_257_76_7784));
   NAND3_X1 i_257_76_7798 (.A1(n_257_76_7593), .A2(n_257_76_7594), .A3(
      n_257_76_7784), .ZN(n_257_76_7785));
   INV_X1 i_257_76_7799 (.A(n_257_76_7785), .ZN(n_257_76_7786));
   NAND4_X1 i_257_76_7800 (.A1(n_257_810), .A2(n_257_76_7786), .A3(n_257_76_7585), 
      .A4(n_257_76_7586), .ZN(n_257_76_7787));
   NAND2_X1 i_257_76_7801 (.A1(n_257_76_7604), .A2(n_257_76_7566), .ZN(
      n_257_76_7788));
   NOR2_X1 i_257_76_7802 (.A1(n_257_76_7787), .A2(n_257_76_7788), .ZN(
      n_257_76_7789));
   NAND2_X1 i_257_76_7803 (.A1(n_257_76_7565), .A2(n_257_76_7789), .ZN(
      n_257_76_7790));
   INV_X1 i_257_76_7804 (.A(n_257_76_7790), .ZN(n_257_76_7791));
   NAND2_X1 i_257_76_7805 (.A1(n_257_76_7791), .A2(n_257_76_7575), .ZN(
      n_257_76_7792));
   INV_X1 i_257_76_7806 (.A(n_257_76_7792), .ZN(n_257_76_7793));
   NAND2_X1 i_257_76_7807 (.A1(n_257_22), .A2(n_257_76_7793), .ZN(n_257_76_7794));
   NAND2_X1 i_257_76_7808 (.A1(n_257_444), .A2(n_257_76_7579), .ZN(n_257_76_7795));
   INV_X1 i_257_76_7809 (.A(n_257_76_7795), .ZN(n_257_76_7796));
   NAND2_X1 i_257_76_7810 (.A1(n_257_1008), .A2(n_257_76_7796), .ZN(
      n_257_76_7797));
   INV_X1 i_257_76_7811 (.A(n_257_76_7797), .ZN(n_257_76_7798));
   NAND2_X1 i_257_76_7812 (.A1(n_257_76_7575), .A2(n_257_76_7798), .ZN(
      n_257_76_7799));
   INV_X1 i_257_76_7813 (.A(n_257_76_7799), .ZN(n_257_76_7800));
   NAND2_X1 i_257_76_7814 (.A1(n_257_76_18075), .A2(n_257_76_7800), .ZN(
      n_257_76_7801));
   NAND2_X1 i_257_76_7815 (.A1(n_257_76_7794), .A2(n_257_76_7801), .ZN(
      n_257_76_7802));
   NOR2_X1 i_257_76_7816 (.A1(n_257_76_7783), .A2(n_257_76_7802), .ZN(
      n_257_76_7803));
   NAND3_X1 i_257_76_7817 (.A1(n_257_76_7677), .A2(n_257_76_7738), .A3(
      n_257_76_7803), .ZN(n_257_76_7804));
   INV_X1 i_257_76_7818 (.A(n_257_76_7804), .ZN(n_257_76_7805));
   NOR2_X1 i_257_76_7819 (.A1(n_257_76_17633), .A2(n_257_1072), .ZN(
      n_257_76_7806));
   NAND4_X1 i_257_76_7820 (.A1(n_257_76_7594), .A2(n_257_76_7643), .A3(n_257_48), 
      .A4(n_257_76_7806), .ZN(n_257_76_7807));
   NOR2_X1 i_257_76_7821 (.A1(n_257_76_7807), .A2(n_257_76_7699), .ZN(
      n_257_76_7808));
   NAND3_X1 i_257_76_7822 (.A1(n_257_76_7769), .A2(n_257_76_7771), .A3(
      n_257_76_7808), .ZN(n_257_76_7809));
   NOR2_X1 i_257_76_7823 (.A1(n_257_76_7809), .A2(n_257_76_7605), .ZN(
      n_257_76_7810));
   NAND3_X1 i_257_76_7824 (.A1(n_257_76_7810), .A2(n_257_76_7607), .A3(
      n_257_76_7565), .ZN(n_257_76_7811));
   NOR2_X1 i_257_76_7825 (.A1(n_257_76_7811), .A2(n_257_76_7609), .ZN(
      n_257_76_7812));
   NAND2_X1 i_257_76_7826 (.A1(n_257_76_18081), .A2(n_257_76_7812), .ZN(
      n_257_76_7813));
   NAND2_X1 i_257_76_7827 (.A1(n_257_1086), .A2(n_257_76_7579), .ZN(
      n_257_76_7814));
   INV_X1 i_257_76_7828 (.A(n_257_76_7814), .ZN(n_257_76_7815));
   NAND3_X1 i_257_76_7829 (.A1(n_257_76_7593), .A2(n_257_76_7594), .A3(
      n_257_76_7815), .ZN(n_257_76_7816));
   NAND2_X1 i_257_76_7830 (.A1(n_257_76_7592), .A2(n_257_449), .ZN(n_257_76_7817));
   NOR2_X1 i_257_76_7831 (.A1(n_257_76_7816), .A2(n_257_76_7817), .ZN(
      n_257_76_7818));
   NAND4_X1 i_257_76_7832 (.A1(n_257_76_7818), .A2(n_257_76_7688), .A3(
      n_257_76_7566), .A4(n_257_76_7585), .ZN(n_257_76_7819));
   NOR2_X1 i_257_76_7833 (.A1(n_257_76_7819), .A2(n_257_76_7605), .ZN(
      n_257_76_7820));
   NAND3_X1 i_257_76_7834 (.A1(n_257_76_7820), .A2(n_257_76_7607), .A3(
      n_257_76_7565), .ZN(n_257_76_7821));
   NOR2_X1 i_257_76_7835 (.A1(n_257_76_7821), .A2(n_257_76_7609), .ZN(
      n_257_76_7822));
   NAND2_X1 i_257_76_7836 (.A1(n_257_76_18083), .A2(n_257_76_7822), .ZN(
      n_257_76_7823));
   NAND2_X1 i_257_76_7837 (.A1(n_257_76_7603), .A2(n_257_76_7604), .ZN(
      n_257_76_7824));
   INV_X1 i_257_76_7838 (.A(n_257_76_7824), .ZN(n_257_76_7825));
   INV_X1 i_257_76_7839 (.A(n_257_76_7646), .ZN(n_257_76_7826));
   NAND3_X1 i_257_76_7840 (.A1(n_257_76_7637), .A2(n_257_76_17331), .A3(
      n_257_76_7705), .ZN(n_257_76_7827));
   INV_X1 i_257_76_7841 (.A(n_257_76_7827), .ZN(n_257_76_7828));
   NAND2_X1 i_257_76_7842 (.A1(n_257_76_7643), .A2(n_257_76_7828), .ZN(
      n_257_76_7829));
   INV_X1 i_257_76_7843 (.A(n_257_76_7829), .ZN(n_257_76_7830));
   NAND4_X1 i_257_76_7844 (.A1(n_257_76_7826), .A2(n_257_76_7830), .A3(
      n_257_76_7649), .A4(n_257_76_7592), .ZN(n_257_76_7831));
   NOR2_X1 i_257_76_7845 (.A1(n_257_76_7831), .A2(n_257_76_7664), .ZN(
      n_257_76_7832));
   NAND4_X1 i_257_76_7846 (.A1(n_257_76_7661), .A2(n_257_76_7566), .A3(
      n_257_76_7665), .A4(n_257_76_7585), .ZN(n_257_76_7833));
   INV_X1 i_257_76_7847 (.A(n_257_76_7833), .ZN(n_257_76_7834));
   NAND3_X1 i_257_76_7848 (.A1(n_257_76_7825), .A2(n_257_76_7832), .A3(
      n_257_76_7834), .ZN(n_257_76_7835));
   NAND3_X1 i_257_76_7849 (.A1(n_257_165), .A2(n_257_76_7668), .A3(n_257_76_7602), 
      .ZN(n_257_76_7836));
   NOR2_X1 i_257_76_7850 (.A1(n_257_76_7835), .A2(n_257_76_7836), .ZN(
      n_257_76_7837));
   NAND4_X1 i_257_76_7851 (.A1(n_257_76_7837), .A2(n_257_76_7575), .A3(
      n_257_76_7607), .A4(n_257_76_7565), .ZN(n_257_76_7838));
   INV_X1 i_257_76_7852 (.A(n_257_76_7838), .ZN(n_257_76_7839));
   NAND2_X1 i_257_76_7853 (.A1(n_257_76_18061), .A2(n_257_76_7839), .ZN(
      n_257_76_7840));
   NAND3_X1 i_257_76_7854 (.A1(n_257_76_7813), .A2(n_257_76_7823), .A3(
      n_257_76_7840), .ZN(n_257_76_7841));
   INV_X1 i_257_76_7855 (.A(n_257_76_7841), .ZN(n_257_76_7842));
   NAND2_X1 i_257_76_7856 (.A1(n_257_1078), .A2(n_257_76_7579), .ZN(
      n_257_76_7843));
   INV_X1 i_257_76_7857 (.A(n_257_76_7843), .ZN(n_257_76_7844));
   NAND3_X1 i_257_76_7858 (.A1(n_257_76_7593), .A2(n_257_76_7844), .A3(n_257_438), 
      .ZN(n_257_76_7845));
   INV_X1 i_257_76_7859 (.A(n_257_76_7845), .ZN(n_257_76_7846));
   NAND3_X1 i_257_76_7860 (.A1(n_257_76_7566), .A2(n_257_76_7585), .A3(
      n_257_76_7846), .ZN(n_257_76_7847));
   INV_X1 i_257_76_7861 (.A(n_257_76_7847), .ZN(n_257_76_7848));
   NAND2_X1 i_257_76_7862 (.A1(n_257_76_7565), .A2(n_257_76_7848), .ZN(
      n_257_76_7849));
   INV_X1 i_257_76_7863 (.A(n_257_76_7849), .ZN(n_257_76_7850));
   NAND2_X1 i_257_76_7864 (.A1(n_257_76_7850), .A2(n_257_76_7575), .ZN(
      n_257_76_7851));
   INV_X1 i_257_76_7865 (.A(n_257_76_7851), .ZN(n_257_76_7852));
   NAND2_X1 i_257_76_7866 (.A1(n_257_76_18067), .A2(n_257_76_7852), .ZN(
      n_257_76_7853));
   NAND2_X1 i_257_76_7867 (.A1(n_257_76_7657), .A2(n_257_76_7668), .ZN(
      n_257_76_7854));
   INV_X1 i_257_76_7868 (.A(n_257_76_7635), .ZN(n_257_76_7855));
   NOR2_X1 i_257_76_7869 (.A1(n_257_76_7854), .A2(n_257_76_7855), .ZN(
      n_257_76_7856));
   INV_X1 i_257_76_7870 (.A(n_257_76_7652), .ZN(n_257_76_7857));
   NOR2_X1 i_257_76_7871 (.A1(n_257_76_7646), .A2(n_257_76_7857), .ZN(
      n_257_76_7858));
   NAND2_X1 i_257_76_7872 (.A1(n_257_76_16781), .A2(n_257_76_7638), .ZN(
      n_257_76_7859));
   OAI21_X1 i_257_76_7873 (.A(n_257_76_7859), .B1(n_257_428), .B2(n_257_76_16526), 
      .ZN(n_257_76_7860));
   NAND2_X1 i_257_76_7874 (.A1(n_257_76_7637), .A2(n_257_76_7860), .ZN(
      n_257_76_7861));
   NAND2_X1 i_257_76_7875 (.A1(n_257_420), .A2(n_257_76_7705), .ZN(n_257_76_7862));
   NOR2_X1 i_257_76_7876 (.A1(n_257_76_7861), .A2(n_257_76_7862), .ZN(
      n_257_76_7863));
   NAND2_X1 i_257_76_7877 (.A1(n_257_76_7863), .A2(n_257_76_7644), .ZN(
      n_257_76_7864));
   NAND2_X1 i_257_76_7878 (.A1(n_257_323), .A2(n_257_422), .ZN(n_257_76_7865));
   NAND2_X1 i_257_76_7879 (.A1(n_257_76_7865), .A2(n_257_76_7643), .ZN(
      n_257_76_7866));
   NOR2_X1 i_257_76_7880 (.A1(n_257_76_7864), .A2(n_257_76_7866), .ZN(
      n_257_76_7867));
   NAND2_X1 i_257_76_7881 (.A1(n_257_76_7858), .A2(n_257_76_7867), .ZN(
      n_257_76_7868));
   NAND2_X1 i_257_76_7882 (.A1(n_257_76_7598), .A2(n_257_76_7648), .ZN(
      n_257_76_7869));
   INV_X1 i_257_76_7883 (.A(n_257_76_7869), .ZN(n_257_76_7870));
   NAND2_X1 i_257_76_7884 (.A1(n_257_76_7870), .A2(n_257_76_7741), .ZN(
      n_257_76_7871));
   NOR2_X1 i_257_76_7885 (.A1(n_257_76_7868), .A2(n_257_76_7871), .ZN(
      n_257_76_7872));
   NAND2_X1 i_257_76_7886 (.A1(n_257_76_7586), .A2(n_257_76_7597), .ZN(
      n_257_76_7873));
   INV_X1 i_257_76_7887 (.A(n_257_76_7873), .ZN(n_257_76_7874));
   NAND2_X1 i_257_76_7888 (.A1(n_257_285), .A2(n_257_423), .ZN(n_257_76_7875));
   NAND2_X1 i_257_76_7889 (.A1(n_257_76_7874), .A2(n_257_76_7875), .ZN(
      n_257_76_7876));
   NAND2_X1 i_257_76_7890 (.A1(n_257_76_7665), .A2(n_257_76_7585), .ZN(
      n_257_76_7877));
   NOR2_X1 i_257_76_7891 (.A1(n_257_76_7876), .A2(n_257_76_7877), .ZN(
      n_257_76_7878));
   NAND2_X1 i_257_76_7892 (.A1(n_257_76_7872), .A2(n_257_76_7878), .ZN(
      n_257_76_7879));
   NAND2_X1 i_257_76_7893 (.A1(n_257_362), .A2(n_257_421), .ZN(n_257_76_7880));
   NAND2_X1 i_257_76_7894 (.A1(n_257_76_7604), .A2(n_257_76_7880), .ZN(
      n_257_76_7881));
   NAND2_X1 i_257_76_7895 (.A1(n_257_76_7661), .A2(n_257_76_7566), .ZN(
      n_257_76_7882));
   NOR2_X1 i_257_76_7896 (.A1(n_257_76_7881), .A2(n_257_76_7882), .ZN(
      n_257_76_7883));
   NAND2_X1 i_257_76_7897 (.A1(n_257_76_7660), .A2(n_257_76_7883), .ZN(
      n_257_76_7884));
   NOR2_X1 i_257_76_7898 (.A1(n_257_76_7879), .A2(n_257_76_7884), .ZN(
      n_257_76_7885));
   NAND2_X1 i_257_76_7899 (.A1(n_257_76_7856), .A2(n_257_76_7885), .ZN(
      n_257_76_7886));
   NAND2_X1 i_257_76_7900 (.A1(n_257_76_7672), .A2(n_257_76_7575), .ZN(
      n_257_76_7887));
   NOR2_X1 i_257_76_7901 (.A1(n_257_76_7886), .A2(n_257_76_7887), .ZN(
      n_257_76_7888));
   NAND2_X1 i_257_76_7902 (.A1(n_257_76_18073), .A2(n_257_76_7888), .ZN(
      n_257_76_7889));
   NOR2_X1 i_257_76_7903 (.A1(n_257_76_7605), .A2(n_257_76_7739), .ZN(
      n_257_76_7890));
   NAND2_X1 i_257_76_7904 (.A1(n_257_76_17925), .A2(n_257_76_7705), .ZN(
      n_257_76_7891));
   NOR2_X1 i_257_76_7905 (.A1(n_257_76_7707), .A2(n_257_76_7891), .ZN(
      n_257_76_7892));
   NAND3_X1 i_257_76_7906 (.A1(n_257_76_7594), .A2(n_257_76_7892), .A3(
      n_257_76_7643), .ZN(n_257_76_7893));
   NOR2_X1 i_257_76_7907 (.A1(n_257_76_7893), .A2(n_257_76_7699), .ZN(
      n_257_76_7894));
   NAND2_X1 i_257_76_7908 (.A1(n_257_76_7598), .A2(n_257_76_7649), .ZN(
      n_257_76_7895));
   INV_X1 i_257_76_7909 (.A(n_257_76_7895), .ZN(n_257_76_7896));
   NAND3_X1 i_257_76_7910 (.A1(n_257_76_7894), .A2(n_257_76_7874), .A3(
      n_257_76_7896), .ZN(n_257_76_7897));
   NAND4_X1 i_257_76_7911 (.A1(n_257_76_7566), .A2(n_257_76_7665), .A3(
      n_257_76_7585), .A4(n_257_126), .ZN(n_257_76_7898));
   NOR2_X1 i_257_76_7912 (.A1(n_257_76_7897), .A2(n_257_76_7898), .ZN(
      n_257_76_7899));
   NAND4_X1 i_257_76_7913 (.A1(n_257_76_7607), .A2(n_257_76_7565), .A3(
      n_257_76_7890), .A4(n_257_76_7899), .ZN(n_257_76_7900));
   NOR2_X1 i_257_76_7914 (.A1(n_257_76_7900), .A2(n_257_76_7609), .ZN(
      n_257_76_7901));
   NAND2_X1 i_257_76_7915 (.A1(n_257_76_18068), .A2(n_257_76_7901), .ZN(
      n_257_76_7902));
   NAND3_X1 i_257_76_7916 (.A1(n_257_76_7853), .A2(n_257_76_7889), .A3(
      n_257_76_7902), .ZN(n_257_76_7903));
   INV_X1 i_257_76_7917 (.A(n_257_76_7903), .ZN(n_257_76_7904));
   NAND2_X1 i_257_76_7918 (.A1(n_257_778), .A2(n_257_442), .ZN(n_257_76_7905));
   NOR2_X1 i_257_76_7919 (.A1(n_257_76_7905), .A2(n_257_1072), .ZN(n_257_76_7906));
   NAND4_X1 i_257_76_7920 (.A1(n_257_447), .A2(n_257_76_7593), .A3(n_257_76_7594), 
      .A4(n_257_76_7906), .ZN(n_257_76_7907));
   INV_X1 i_257_76_7921 (.A(n_257_76_7907), .ZN(n_257_76_7908));
   NAND4_X1 i_257_76_7922 (.A1(n_257_76_7908), .A2(n_257_76_7566), .A3(
      n_257_76_7585), .A4(n_257_76_7586), .ZN(n_257_76_7909));
   NOR2_X1 i_257_76_7923 (.A1(n_257_76_7909), .A2(n_257_76_7824), .ZN(
      n_257_76_7910));
   NAND2_X1 i_257_76_7924 (.A1(n_257_76_7565), .A2(n_257_76_7910), .ZN(
      n_257_76_7911));
   INV_X1 i_257_76_7925 (.A(n_257_76_7911), .ZN(n_257_76_7912));
   NAND2_X1 i_257_76_7926 (.A1(n_257_76_7912), .A2(n_257_76_7575), .ZN(
      n_257_76_7913));
   INV_X1 i_257_76_7927 (.A(n_257_76_7913), .ZN(n_257_76_7914));
   NAND2_X1 i_257_76_7928 (.A1(n_257_76_7705), .A2(n_257_76_17932), .ZN(
      n_257_76_7915));
   NOR2_X1 i_257_76_7929 (.A1(n_257_76_7707), .A2(n_257_76_7915), .ZN(
      n_257_76_7916));
   NAND4_X1 i_257_76_7930 (.A1(n_257_76_7593), .A2(n_257_76_7594), .A3(
      n_257_76_7916), .A4(n_257_76_7643), .ZN(n_257_76_7917));
   NOR2_X1 i_257_76_7931 (.A1(n_257_76_7917), .A2(n_257_76_7740), .ZN(
      n_257_76_7918));
   NAND3_X1 i_257_76_7932 (.A1(n_257_76_7769), .A2(n_257_76_7771), .A3(
      n_257_76_7918), .ZN(n_257_76_7919));
   NAND4_X1 i_257_76_7933 (.A1(n_257_76_7602), .A2(n_257_76_7603), .A3(n_257_88), 
      .A4(n_257_76_7604), .ZN(n_257_76_7920));
   NOR2_X1 i_257_76_7934 (.A1(n_257_76_7919), .A2(n_257_76_7920), .ZN(
      n_257_76_7921));
   NAND3_X1 i_257_76_7935 (.A1(n_257_76_7921), .A2(n_257_76_7607), .A3(
      n_257_76_7565), .ZN(n_257_76_7922));
   NOR2_X1 i_257_76_7936 (.A1(n_257_76_7922), .A2(n_257_76_7609), .ZN(
      n_257_76_7923));
   AOI22_X1 i_257_76_7937 (.A1(n_257_76_18085), .A2(n_257_76_7914), .B1(
      n_257_76_18080), .B2(n_257_76_7923), .ZN(n_257_76_7924));
   NAND3_X1 i_257_76_7938 (.A1(n_257_76_7842), .A2(n_257_76_7904), .A3(
      n_257_76_7924), .ZN(n_257_76_7925));
   INV_X1 i_257_76_7939 (.A(n_257_76_7598), .ZN(n_257_76_7926));
   NAND3_X1 i_257_76_7940 (.A1(n_257_76_7593), .A2(n_257_76_7594), .A3(n_257_448), 
      .ZN(n_257_76_7927));
   NOR2_X1 i_257_76_7941 (.A1(n_257_76_7926), .A2(n_257_76_7927), .ZN(
      n_257_76_7928));
   NAND2_X1 i_257_76_7942 (.A1(n_257_76_7579), .A2(n_257_76_17760), .ZN(
      n_257_76_7929));
   OAI21_X1 i_257_76_7943 (.A(n_257_76_7929), .B1(n_257_714), .B2(n_257_76_7689), 
      .ZN(n_257_76_7930));
   NAND2_X1 i_257_76_7944 (.A1(n_257_76_7586), .A2(n_257_76_7930), .ZN(
      n_257_76_7931));
   INV_X1 i_257_76_7945 (.A(n_257_76_7931), .ZN(n_257_76_7932));
   NAND4_X1 i_257_76_7946 (.A1(n_257_76_7928), .A2(n_257_76_7932), .A3(
      n_257_76_7566), .A4(n_257_76_7585), .ZN(n_257_76_7933));
   NOR2_X1 i_257_76_7947 (.A1(n_257_76_7933), .A2(n_257_76_7605), .ZN(
      n_257_76_7934));
   NAND3_X1 i_257_76_7948 (.A1(n_257_76_7934), .A2(n_257_76_7565), .A3(n_257_682), 
      .ZN(n_257_76_7935));
   NOR2_X1 i_257_76_7949 (.A1(n_257_76_7935), .A2(n_257_76_7609), .ZN(
      n_257_76_7936));
   NAND2_X1 i_257_76_7950 (.A1(n_257_76_18079), .A2(n_257_76_7936), .ZN(
      n_257_76_7937));
   NOR2_X1 i_257_76_7951 (.A1(n_257_76_7659), .A2(n_257_76_7662), .ZN(
      n_257_76_7938));
   NAND2_X1 i_257_76_7952 (.A1(n_257_76_7668), .A2(n_257_245), .ZN(n_257_76_7939));
   INV_X1 i_257_76_7953 (.A(n_257_76_7939), .ZN(n_257_76_7940));
   NOR2_X1 i_257_76_7954 (.A1(n_257_1072), .A2(n_257_76_17778), .ZN(
      n_257_76_7941));
   NAND3_X1 i_257_76_7955 (.A1(n_257_76_7941), .A2(n_257_76_7637), .A3(
      n_257_76_7640), .ZN(n_257_76_7942));
   INV_X1 i_257_76_7956 (.A(n_257_76_7942), .ZN(n_257_76_7943));
   NAND4_X1 i_257_76_7957 (.A1(n_257_76_7593), .A2(n_257_76_7594), .A3(
      n_257_76_7943), .A4(n_257_76_7643), .ZN(n_257_76_7944));
   INV_X1 i_257_76_7958 (.A(n_257_76_7944), .ZN(n_257_76_7945));
   NAND3_X1 i_257_76_7959 (.A1(n_257_76_7649), .A2(n_257_76_7592), .A3(
      n_257_76_7652), .ZN(n_257_76_7946));
   INV_X1 i_257_76_7960 (.A(n_257_76_7946), .ZN(n_257_76_7947));
   NAND3_X1 i_257_76_7961 (.A1(n_257_76_7870), .A2(n_257_76_7945), .A3(
      n_257_76_7947), .ZN(n_257_76_7948));
   NOR2_X1 i_257_76_7962 (.A1(n_257_76_7948), .A2(n_257_76_7698), .ZN(
      n_257_76_7949));
   NAND4_X1 i_257_76_7963 (.A1(n_257_76_7938), .A2(n_257_76_7940), .A3(
      n_257_76_7949), .A4(n_257_76_7635), .ZN(n_257_76_7950));
   INV_X1 i_257_76_7964 (.A(n_257_76_7950), .ZN(n_257_76_7951));
   NAND3_X1 i_257_76_7965 (.A1(n_257_76_7951), .A2(n_257_76_7672), .A3(
      n_257_76_7575), .ZN(n_257_76_7952));
   INV_X1 i_257_76_7966 (.A(n_257_76_7952), .ZN(n_257_76_7953));
   NAND2_X1 i_257_76_7967 (.A1(n_257_76_18064), .A2(n_257_76_7953), .ZN(
      n_257_76_7954));
   NAND3_X1 i_257_76_7968 (.A1(n_257_362), .A2(n_257_76_7585), .A3(n_257_76_7875), 
      .ZN(n_257_76_7955));
   NOR2_X1 i_257_76_7969 (.A1(n_257_76_7955), .A2(n_257_76_7664), .ZN(
      n_257_76_7956));
   INV_X1 i_257_76_7970 (.A(n_257_76_7866), .ZN(n_257_76_7957));
   NOR2_X1 i_257_76_7971 (.A1(n_257_1072), .A2(n_257_76_17792), .ZN(
      n_257_76_7958));
   NAND3_X1 i_257_76_7972 (.A1(n_257_76_7958), .A2(n_257_76_7637), .A3(
      n_257_76_7640), .ZN(n_257_76_7959));
   INV_X1 i_257_76_7973 (.A(n_257_76_7644), .ZN(n_257_76_7960));
   NOR2_X1 i_257_76_7974 (.A1(n_257_76_7959), .A2(n_257_76_7960), .ZN(
      n_257_76_7961));
   NAND3_X1 i_257_76_7975 (.A1(n_257_76_7826), .A2(n_257_76_7957), .A3(
      n_257_76_7961), .ZN(n_257_76_7962));
   NAND4_X1 i_257_76_7976 (.A1(n_257_76_7648), .A2(n_257_76_7649), .A3(
      n_257_76_7592), .A4(n_257_76_7652), .ZN(n_257_76_7963));
   NOR2_X1 i_257_76_7977 (.A1(n_257_76_7962), .A2(n_257_76_7963), .ZN(
      n_257_76_7964));
   NAND3_X1 i_257_76_7978 (.A1(n_257_76_7604), .A2(n_257_76_7661), .A3(
      n_257_76_7665), .ZN(n_257_76_7965));
   INV_X1 i_257_76_7979 (.A(n_257_76_7965), .ZN(n_257_76_7966));
   NAND4_X1 i_257_76_7980 (.A1(n_257_76_7660), .A2(n_257_76_7956), .A3(
      n_257_76_7964), .A4(n_257_76_7966), .ZN(n_257_76_7967));
   INV_X1 i_257_76_7981 (.A(n_257_76_7967), .ZN(n_257_76_7968));
   NAND2_X1 i_257_76_7982 (.A1(n_257_76_7575), .A2(n_257_76_7968), .ZN(
      n_257_76_7969));
   NAND2_X1 i_257_76_7983 (.A1(n_257_76_7635), .A2(n_257_76_7657), .ZN(
      n_257_76_7970));
   INV_X1 i_257_76_7984 (.A(n_257_76_7970), .ZN(n_257_76_7971));
   NAND2_X1 i_257_76_7985 (.A1(n_257_76_7668), .A2(n_257_76_7566), .ZN(
      n_257_76_7972));
   INV_X1 i_257_76_7986 (.A(n_257_76_7972), .ZN(n_257_76_7973));
   NAND4_X1 i_257_76_7987 (.A1(n_257_76_7971), .A2(n_257_76_7607), .A3(
      n_257_76_7565), .A4(n_257_76_7973), .ZN(n_257_76_7974));
   NOR2_X1 i_257_76_7988 (.A1(n_257_76_7969), .A2(n_257_76_7974), .ZN(
      n_257_76_7975));
   NAND2_X1 i_257_76_7989 (.A1(n_257_76_18082), .A2(n_257_76_7975), .ZN(
      n_257_76_7976));
   NAND3_X1 i_257_76_7990 (.A1(n_257_76_7937), .A2(n_257_76_7954), .A3(
      n_257_76_7976), .ZN(n_257_76_7977));
   INV_X1 i_257_76_7991 (.A(n_257_76_7977), .ZN(n_257_76_7978));
   NAND3_X1 i_257_76_7992 (.A1(n_257_76_7593), .A2(n_257_76_7594), .A3(
      n_257_76_7643), .ZN(n_257_76_7979));
   NOR2_X1 i_257_76_7993 (.A1(n_257_76_7740), .A2(n_257_76_7979), .ZN(
      n_257_76_7980));
   NAND3_X1 i_257_76_7994 (.A1(n_257_76_7637), .A2(n_257_76_7640), .A3(
      n_257_76_7705), .ZN(n_257_76_7981));
   INV_X1 i_257_76_7995 (.A(n_257_76_7981), .ZN(n_257_76_7982));
   NAND3_X1 i_257_76_7996 (.A1(n_257_76_7982), .A2(n_257_205), .A3(n_257_427), 
      .ZN(n_257_76_7983));
   INV_X1 i_257_76_7997 (.A(n_257_76_7983), .ZN(n_257_76_7984));
   NAND2_X1 i_257_76_7998 (.A1(n_257_76_7586), .A2(n_257_76_7984), .ZN(
      n_257_76_7985));
   INV_X1 i_257_76_7999 (.A(n_257_76_7985), .ZN(n_257_76_7986));
   NAND3_X1 i_257_76_8000 (.A1(n_257_76_7980), .A2(n_257_76_7600), .A3(
      n_257_76_7986), .ZN(n_257_76_7987));
   NOR2_X1 i_257_76_8001 (.A1(n_257_76_7987), .A2(n_257_76_7833), .ZN(
      n_257_76_7988));
   NAND4_X1 i_257_76_8002 (.A1(n_257_76_7988), .A2(n_257_76_7635), .A3(
      n_257_76_7668), .A4(n_257_76_7751), .ZN(n_257_76_7989));
   INV_X1 i_257_76_8003 (.A(n_257_76_7989), .ZN(n_257_76_7990));
   NAND3_X1 i_257_76_8004 (.A1(n_257_76_7990), .A2(n_257_76_7672), .A3(
      n_257_76_7575), .ZN(n_257_76_7991));
   INV_X1 i_257_76_8005 (.A(n_257_76_7991), .ZN(n_257_76_7992));
   NAND2_X1 i_257_76_8006 (.A1(n_257_76_18065), .A2(n_257_76_7992), .ZN(
      n_257_76_7993));
   NAND2_X1 i_257_76_8007 (.A1(n_257_465), .A2(n_257_76_7579), .ZN(n_257_76_7994));
   INV_X1 i_257_76_8008 (.A(n_257_76_7994), .ZN(n_257_76_7995));
   NAND3_X1 i_257_76_8009 (.A1(n_257_76_7594), .A2(n_257_76_7643), .A3(
      n_257_76_7995), .ZN(n_257_76_7996));
   NOR2_X1 i_257_76_8010 (.A1(n_257_76_7699), .A2(n_257_76_7996), .ZN(
      n_257_76_7997));
   NAND3_X1 i_257_76_8011 (.A1(n_257_76_7597), .A2(n_257_76_7598), .A3(n_257_451), 
      .ZN(n_257_76_7998));
   INV_X1 i_257_76_8012 (.A(n_257_76_7998), .ZN(n_257_76_7999));
   NAND4_X1 i_257_76_8013 (.A1(n_257_76_7997), .A2(n_257_76_7999), .A3(
      n_257_76_7588), .A4(n_257_76_7566), .ZN(n_257_76_8000));
   NOR2_X1 i_257_76_8014 (.A1(n_257_76_8000), .A2(n_257_76_7605), .ZN(
      n_257_76_8001));
   NAND3_X1 i_257_76_8015 (.A1(n_257_76_8001), .A2(n_257_76_7607), .A3(
      n_257_76_7565), .ZN(n_257_76_8002));
   NOR2_X1 i_257_76_8016 (.A1(n_257_76_8002), .A2(n_257_76_7609), .ZN(
      n_257_76_8003));
   NAND2_X1 i_257_76_8017 (.A1(n_257_76_18063), .A2(n_257_76_8003), .ZN(
      n_257_76_8004));
   NOR2_X1 i_257_76_8018 (.A1(n_257_76_16145), .A2(n_257_1072), .ZN(
      n_257_76_8005));
   NAND4_X1 i_257_76_8019 (.A1(n_257_76_8005), .A2(n_257_514), .A3(n_257_76_7640), 
      .A4(n_257_76_7637), .ZN(n_257_76_8006));
   INV_X1 i_257_76_8020 (.A(n_257_76_8006), .ZN(n_257_76_8007));
   NAND3_X1 i_257_76_8021 (.A1(n_257_76_8007), .A2(n_257_76_7594), .A3(
      n_257_76_7643), .ZN(n_257_76_8008));
   INV_X1 i_257_76_8022 (.A(n_257_76_8008), .ZN(n_257_76_8009));
   NAND3_X1 i_257_76_8023 (.A1(n_257_76_7592), .A2(n_257_76_7652), .A3(
      n_257_76_7593), .ZN(n_257_76_8010));
   INV_X1 i_257_76_8024 (.A(n_257_76_8010), .ZN(n_257_76_8011));
   NAND3_X1 i_257_76_8025 (.A1(n_257_76_7651), .A2(n_257_76_8009), .A3(
      n_257_76_8011), .ZN(n_257_76_8012));
   NOR2_X1 i_257_76_8026 (.A1(n_257_76_8012), .A2(n_257_76_7768), .ZN(
      n_257_76_8013));
   NAND4_X1 i_257_76_8027 (.A1(n_257_76_7604), .A2(n_257_76_7661), .A3(
      n_257_76_7566), .A4(n_257_76_7665), .ZN(n_257_76_8014));
   INV_X1 i_257_76_8028 (.A(n_257_76_8014), .ZN(n_257_76_8015));
   NAND3_X1 i_257_76_8029 (.A1(n_257_76_8013), .A2(n_257_76_7660), .A3(
      n_257_76_8015), .ZN(n_257_76_8016));
   NAND3_X1 i_257_76_8030 (.A1(n_257_76_7635), .A2(n_257_76_7657), .A3(
      n_257_76_7668), .ZN(n_257_76_8017));
   NOR2_X1 i_257_76_8031 (.A1(n_257_76_8016), .A2(n_257_76_8017), .ZN(
      n_257_76_8018));
   NAND3_X1 i_257_76_8032 (.A1(n_257_76_8018), .A2(n_257_76_7672), .A3(
      n_257_76_7575), .ZN(n_257_76_8019));
   INV_X1 i_257_76_8033 (.A(n_257_76_8019), .ZN(n_257_76_8020));
   NAND2_X1 i_257_76_8034 (.A1(n_257_76_18062), .A2(n_257_76_8020), .ZN(
      n_257_76_8021));
   NAND3_X1 i_257_76_8035 (.A1(n_257_76_7993), .A2(n_257_76_8004), .A3(
      n_257_76_8021), .ZN(n_257_76_8022));
   INV_X1 i_257_76_8036 (.A(n_257_76_8022), .ZN(n_257_76_8023));
   NAND4_X1 i_257_76_8037 (.A1(n_257_76_7652), .A2(n_257_76_7593), .A3(
      n_257_76_7594), .A4(n_257_76_7643), .ZN(n_257_76_8024));
   NOR2_X1 i_257_76_8038 (.A1(n_257_76_8024), .A2(n_257_76_7740), .ZN(
      n_257_76_8025));
   NAND2_X1 i_257_76_8039 (.A1(n_257_76_7637), .A2(n_257_76_7640), .ZN(
      n_257_76_8026));
   INV_X1 i_257_76_8040 (.A(n_257_76_8026), .ZN(n_257_76_8027));
   NAND2_X1 i_257_76_8041 (.A1(n_257_422), .A2(n_257_76_7705), .ZN(n_257_76_8028));
   INV_X1 i_257_76_8042 (.A(n_257_76_8028), .ZN(n_257_76_8029));
   NAND4_X1 i_257_76_8043 (.A1(n_257_76_8027), .A2(n_257_76_7644), .A3(n_257_323), 
      .A4(n_257_76_8029), .ZN(n_257_76_8030));
   INV_X1 i_257_76_8044 (.A(n_257_76_8030), .ZN(n_257_76_8031));
   NAND3_X1 i_257_76_8045 (.A1(n_257_76_7875), .A2(n_257_76_7586), .A3(
      n_257_76_8031), .ZN(n_257_76_8032));
   INV_X1 i_257_76_8046 (.A(n_257_76_8032), .ZN(n_257_76_8033));
   NAND3_X1 i_257_76_8047 (.A1(n_257_76_7597), .A2(n_257_76_7598), .A3(
      n_257_76_7648), .ZN(n_257_76_8034));
   INV_X1 i_257_76_8048 (.A(n_257_76_8034), .ZN(n_257_76_8035));
   NAND3_X1 i_257_76_8049 (.A1(n_257_76_8025), .A2(n_257_76_8033), .A3(
      n_257_76_8035), .ZN(n_257_76_8036));
   INV_X1 i_257_76_8050 (.A(n_257_76_8036), .ZN(n_257_76_8037));
   NAND2_X1 i_257_76_8051 (.A1(n_257_76_7604), .A2(n_257_76_7661), .ZN(
      n_257_76_8038));
   NAND3_X1 i_257_76_8052 (.A1(n_257_76_7566), .A2(n_257_76_7665), .A3(
      n_257_76_7585), .ZN(n_257_76_8039));
   NOR2_X1 i_257_76_8053 (.A1(n_257_76_8038), .A2(n_257_76_8039), .ZN(
      n_257_76_8040));
   NAND3_X1 i_257_76_8054 (.A1(n_257_76_7660), .A2(n_257_76_8037), .A3(
      n_257_76_8040), .ZN(n_257_76_8041));
   NOR2_X1 i_257_76_8055 (.A1(n_257_76_8041), .A2(n_257_76_8017), .ZN(
      n_257_76_8042));
   NAND3_X1 i_257_76_8056 (.A1(n_257_76_8042), .A2(n_257_76_7672), .A3(
      n_257_76_7575), .ZN(n_257_76_8043));
   INV_X1 i_257_76_8057 (.A(n_257_76_8043), .ZN(n_257_76_8044));
   NAND2_X1 i_257_76_8058 (.A1(n_257_342), .A2(n_257_76_8044), .ZN(n_257_76_8045));
   NAND3_X1 i_257_76_8059 (.A1(n_257_76_7585), .A2(n_257_76_7875), .A3(
      n_257_76_7586), .ZN(n_257_76_8046));
   NOR2_X1 i_257_76_8060 (.A1(n_257_76_7770), .A2(n_257_76_8046), .ZN(
      n_257_76_8047));
   NAND3_X1 i_257_76_8061 (.A1(n_257_76_7604), .A2(n_257_76_7880), .A3(
      n_257_76_7661), .ZN(n_257_76_8048));
   INV_X1 i_257_76_8062 (.A(n_257_76_8048), .ZN(n_257_76_8049));
   NAND4_X1 i_257_76_8063 (.A1(n_257_76_8047), .A2(n_257_76_7660), .A3(
      n_257_76_8049), .A4(n_257_76_7668), .ZN(n_257_76_8050));
   NAND2_X1 i_257_76_8064 (.A1(n_257_428), .A2(n_257_578), .ZN(n_257_76_8051));
   NAND3_X1 i_257_76_8065 (.A1(n_257_484), .A2(n_257_401), .A3(n_257_442), 
      .ZN(n_257_76_8052));
   INV_X1 i_257_76_8066 (.A(n_257_76_8052), .ZN(n_257_76_8053));
   NAND3_X1 i_257_76_8067 (.A1(n_257_76_7705), .A2(n_257_76_8051), .A3(
      n_257_76_8053), .ZN(n_257_76_8054));
   NOR2_X1 i_257_76_8068 (.A1(n_257_76_8054), .A2(n_257_76_7707), .ZN(
      n_257_76_8055));
   NAND2_X1 i_257_76_8069 (.A1(n_257_420), .A2(n_257_666), .ZN(n_257_76_8056));
   NAND4_X1 i_257_76_8070 (.A1(n_257_76_8055), .A2(n_257_76_7643), .A3(
      n_257_76_7644), .A4(n_257_76_8056), .ZN(n_257_76_8057));
   INV_X1 i_257_76_8071 (.A(n_257_76_8057), .ZN(n_257_76_8058));
   NAND2_X1 i_257_76_8072 (.A1(n_257_76_7592), .A2(n_257_76_7652), .ZN(
      n_257_76_8059));
   INV_X1 i_257_76_8073 (.A(n_257_76_8059), .ZN(n_257_76_8060));
   NAND3_X1 i_257_76_8074 (.A1(n_257_76_7593), .A2(n_257_76_7594), .A3(
      n_257_76_7865), .ZN(n_257_76_8061));
   INV_X1 i_257_76_8075 (.A(n_257_76_8061), .ZN(n_257_76_8062));
   NAND3_X1 i_257_76_8076 (.A1(n_257_76_8058), .A2(n_257_76_8060), .A3(
      n_257_76_8062), .ZN(n_257_76_8063));
   NAND4_X1 i_257_76_8077 (.A1(n_257_76_7597), .A2(n_257_76_7598), .A3(
      n_257_76_7648), .A4(n_257_76_7649), .ZN(n_257_76_8064));
   NOR2_X1 i_257_76_8078 (.A1(n_257_76_8063), .A2(n_257_76_8064), .ZN(
      n_257_76_8065));
   NAND3_X1 i_257_76_8079 (.A1(n_257_76_7635), .A2(n_257_76_8065), .A3(
      n_257_76_7657), .ZN(n_257_76_8066));
   NOR2_X1 i_257_76_8080 (.A1(n_257_76_8050), .A2(n_257_76_8066), .ZN(
      n_257_76_8067));
   NAND3_X1 i_257_76_8081 (.A1(n_257_76_8067), .A2(n_257_76_7672), .A3(
      n_257_76_7575), .ZN(n_257_76_8068));
   INV_X1 i_257_76_8082 (.A(n_257_76_8068), .ZN(n_257_76_8069));
   NAND2_X1 i_257_76_8083 (.A1(n_257_76_18060), .A2(n_257_76_8069), .ZN(
      n_257_76_8070));
   NAND2_X1 i_257_76_8084 (.A1(n_257_88), .A2(n_257_76_17932), .ZN(n_257_76_8071));
   NAND2_X1 i_257_76_8085 (.A1(n_257_76_7749), .A2(n_257_76_8071), .ZN(
      n_257_76_8072));
   INV_X1 i_257_76_8086 (.A(n_257_76_8072), .ZN(n_257_76_8073));
   NAND2_X1 i_257_76_8087 (.A1(n_257_165), .A2(n_257_76_17331), .ZN(
      n_257_76_8074));
   NAND3_X1 i_257_76_8088 (.A1(n_257_76_8073), .A2(n_257_76_8074), .A3(
      n_257_76_7655), .ZN(n_257_76_8075));
   NAND2_X1 i_257_76_8089 (.A1(n_257_874), .A2(n_257_76_17903), .ZN(
      n_257_76_8076));
   NAND2_X1 i_257_76_8090 (.A1(n_257_126), .A2(n_257_76_17925), .ZN(
      n_257_76_8077));
   NAND2_X1 i_257_76_8091 (.A1(n_257_76_8076), .A2(n_257_76_8077), .ZN(
      n_257_76_8078));
   NAND2_X1 i_257_76_8092 (.A1(n_257_976), .A2(n_257_442), .ZN(n_257_76_8079));
   INV_X1 i_257_76_8093 (.A(n_257_76_8079), .ZN(n_257_76_8080));
   NAND2_X1 i_257_76_8094 (.A1(n_257_441), .A2(n_257_76_8080), .ZN(n_257_76_8081));
   NAND2_X1 i_257_76_8095 (.A1(n_257_465), .A2(n_257_442), .ZN(n_257_76_8082));
   INV_X1 i_257_76_8096 (.A(n_257_76_8082), .ZN(n_257_76_8083));
   NAND2_X1 i_257_76_8097 (.A1(n_257_451), .A2(n_257_76_8083), .ZN(n_257_76_8084));
   NAND2_X1 i_257_76_8098 (.A1(n_257_912), .A2(n_257_76_17940), .ZN(
      n_257_76_8085));
   NAND3_X1 i_257_76_8099 (.A1(n_257_76_8081), .A2(n_257_76_8084), .A3(
      n_257_76_8085), .ZN(n_257_76_8086));
   NOR2_X1 i_257_76_8100 (.A1(n_257_76_8078), .A2(n_257_76_8086), .ZN(
      n_257_76_8087));
   NAND2_X1 i_257_76_8101 (.A1(n_257_48), .A2(n_257_76_17918), .ZN(n_257_76_8088));
   NAND2_X1 i_257_76_8102 (.A1(n_257_714), .A2(n_257_76_15655), .ZN(
      n_257_76_8089));
   NAND3_X1 i_257_76_8103 (.A1(n_257_438), .A2(n_257_1078), .A3(n_257_442), 
      .ZN(n_257_76_8090));
   NAND3_X1 i_257_76_8104 (.A1(n_257_76_8088), .A2(n_257_76_8089), .A3(
      n_257_76_8090), .ZN(n_257_76_8091));
   INV_X1 i_257_76_8105 (.A(n_257_76_8091), .ZN(n_257_76_8092));
   NAND2_X1 i_257_76_8106 (.A1(n_257_76_7983), .A2(n_257_76_8030), .ZN(
      n_257_76_8093));
   INV_X1 i_257_76_8107 (.A(n_257_76_8093), .ZN(n_257_76_8094));
   INV_X1 i_257_76_8108 (.A(n_257_76_7567), .ZN(n_257_76_8095));
   NAND2_X1 i_257_76_8109 (.A1(n_257_440), .A2(n_257_76_8095), .ZN(n_257_76_8096));
   NAND2_X1 i_257_76_8110 (.A1(n_257_642), .A2(n_257_76_17928), .ZN(
      n_257_76_8097));
   NAND2_X1 i_257_76_8111 (.A1(n_257_432), .A2(n_257_76_7773), .ZN(n_257_76_8098));
   NAND3_X1 i_257_76_8112 (.A1(n_257_76_8096), .A2(n_257_76_8097), .A3(
      n_257_76_8098), .ZN(n_257_76_8099));
   INV_X1 i_257_76_8113 (.A(n_257_76_8099), .ZN(n_257_76_8100));
   NAND3_X1 i_257_76_8114 (.A1(n_257_76_8092), .A2(n_257_76_8094), .A3(
      n_257_76_8100), .ZN(n_257_76_8101));
   INV_X1 i_257_76_8115 (.A(Small_Packet_Data_Size[13]), .ZN(n_257_76_8102));
   NAND3_X1 i_257_76_8116 (.A1(n_257_76_18040), .A2(n_257_76_7705), .A3(
      n_257_76_8051), .ZN(n_257_76_8103));
   INV_X1 i_257_76_8117 (.A(n_257_76_8103), .ZN(n_257_76_8104));
   NAND3_X1 i_257_76_8118 (.A1(n_257_76_8104), .A2(n_257_76_7644), .A3(
      n_257_76_8056), .ZN(n_257_76_8105));
   NAND2_X1 i_257_76_8119 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[13]), 
      .ZN(n_257_76_8106));
   NAND2_X1 i_257_76_8120 (.A1(n_257_76_8105), .A2(n_257_76_8106), .ZN(
      n_257_76_8107));
   NAND2_X1 i_257_76_8121 (.A1(n_257_842), .A2(n_257_442), .ZN(n_257_76_8108));
   INV_X1 i_257_76_8122 (.A(n_257_76_8108), .ZN(n_257_76_8109));
   NAND2_X1 i_257_76_8123 (.A1(n_257_446), .A2(n_257_76_8109), .ZN(n_257_76_8110));
   NAND2_X1 i_257_76_8124 (.A1(n_257_449), .A2(n_257_76_15320), .ZN(
      n_257_76_8111));
   INV_X1 i_257_76_8125 (.A(n_257_76_7905), .ZN(n_257_76_8112));
   NAND2_X1 i_257_76_8126 (.A1(n_257_447), .A2(n_257_76_8112), .ZN(n_257_76_8113));
   NAND4_X1 i_257_76_8127 (.A1(n_257_76_8107), .A2(n_257_76_8110), .A3(
      n_257_76_8111), .A4(n_257_76_8113), .ZN(n_257_76_8114));
   NOR2_X1 i_257_76_8128 (.A1(n_257_76_8101), .A2(n_257_76_8114), .ZN(
      n_257_76_8115));
   AOI22_X1 i_257_76_8129 (.A1(n_257_746), .A2(n_257_76_17935), .B1(n_257_810), 
      .B2(n_257_76_17952), .ZN(n_257_76_8116));
   NAND3_X1 i_257_76_8130 (.A1(n_257_76_8087), .A2(n_257_76_8115), .A3(
      n_257_76_8116), .ZN(n_257_76_8117));
   NOR2_X1 i_257_76_8131 (.A1(n_257_76_8075), .A2(n_257_76_8117), .ZN(
      n_257_76_8118));
   NAND2_X1 i_257_76_8132 (.A1(n_257_682), .A2(n_257_76_17958), .ZN(
      n_257_76_8119));
   NAND2_X1 i_257_76_8133 (.A1(n_257_1008), .A2(n_257_76_17964), .ZN(
      n_257_76_8120));
   NAND3_X1 i_257_76_8134 (.A1(n_257_76_8119), .A2(n_257_76_7967), .A3(
      n_257_76_8120), .ZN(n_257_76_8121));
   INV_X1 i_257_76_8135 (.A(n_257_76_8121), .ZN(n_257_76_8122));
   NAND2_X1 i_257_76_8136 (.A1(n_257_1040), .A2(n_257_76_17969), .ZN(
      n_257_76_8123));
   NAND4_X1 i_257_76_8137 (.A1(n_257_76_8118), .A2(n_257_76_8122), .A3(
      n_257_76_7950), .A4(n_257_76_8123), .ZN(n_257_76_8124));
   NAND3_X1 i_257_76_8138 (.A1(n_257_76_8045), .A2(n_257_76_8070), .A3(
      n_257_76_8124), .ZN(n_257_76_8125));
   INV_X1 i_257_76_8139 (.A(n_257_76_8125), .ZN(n_257_76_8126));
   NAND3_X1 i_257_76_8140 (.A1(n_257_76_7978), .A2(n_257_76_8023), .A3(
      n_257_76_8126), .ZN(n_257_76_8127));
   NOR2_X1 i_257_76_8141 (.A1(n_257_76_7925), .A2(n_257_76_8127), .ZN(
      n_257_76_8128));
   NAND2_X1 i_257_76_8142 (.A1(n_257_76_7805), .A2(n_257_76_8128), .ZN(n_13));
   NAND2_X1 i_257_76_8143 (.A1(n_257_1041), .A2(n_257_443), .ZN(n_257_76_8129));
   NAND2_X1 i_257_76_8144 (.A1(n_257_1009), .A2(n_257_444), .ZN(n_257_76_8130));
   NAND2_X1 i_257_76_8145 (.A1(n_257_441), .A2(n_257_977), .ZN(n_257_76_8131));
   NAND2_X1 i_257_76_8146 (.A1(n_257_945), .A2(n_257_442), .ZN(n_257_76_8132));
   NOR2_X1 i_257_76_8147 (.A1(n_257_1073), .A2(n_257_76_8132), .ZN(n_257_76_8133));
   NAND2_X1 i_257_76_8148 (.A1(n_257_440), .A2(n_257_76_8133), .ZN(n_257_76_8134));
   INV_X1 i_257_76_8149 (.A(n_257_76_8134), .ZN(n_257_76_8135));
   NAND2_X1 i_257_76_8150 (.A1(n_257_76_8131), .A2(n_257_76_8135), .ZN(
      n_257_76_8136));
   INV_X1 i_257_76_8151 (.A(n_257_76_8136), .ZN(n_257_76_8137));
   NAND2_X1 i_257_76_8152 (.A1(n_257_76_8130), .A2(n_257_76_8137), .ZN(
      n_257_76_8138));
   INV_X1 i_257_76_8153 (.A(n_257_76_8138), .ZN(n_257_76_8139));
   NAND2_X1 i_257_76_8154 (.A1(n_257_76_8129), .A2(n_257_76_8139), .ZN(
      n_257_76_8140));
   INV_X1 i_257_76_8155 (.A(n_257_76_8140), .ZN(n_257_76_8141));
   NAND2_X1 i_257_76_8156 (.A1(n_257_17), .A2(n_257_76_8141), .ZN(n_257_76_8142));
   NOR2_X1 i_257_76_8157 (.A1(n_257_1073), .A2(n_257_76_17412), .ZN(
      n_257_76_8143));
   NAND2_X1 i_257_76_8158 (.A1(n_257_443), .A2(n_257_76_8143), .ZN(n_257_76_8144));
   INV_X1 i_257_76_8159 (.A(n_257_76_8144), .ZN(n_257_76_8145));
   NAND2_X1 i_257_76_8160 (.A1(n_257_1041), .A2(n_257_76_8145), .ZN(
      n_257_76_8146));
   INV_X1 i_257_76_8161 (.A(n_257_76_8146), .ZN(n_257_76_8147));
   NAND2_X1 i_257_76_8162 (.A1(n_257_76_18072), .A2(n_257_76_8147), .ZN(
      n_257_76_8148));
   NAND2_X1 i_257_76_8163 (.A1(n_257_446), .A2(n_257_843), .ZN(n_257_76_8149));
   NAND2_X1 i_257_76_8164 (.A1(n_257_449), .A2(n_257_1087), .ZN(n_257_76_8150));
   NAND2_X1 i_257_76_8165 (.A1(n_257_76_8149), .A2(n_257_76_8150), .ZN(
      n_257_76_8151));
   INV_X1 i_257_76_8166 (.A(n_257_76_8151), .ZN(n_257_76_8152));
   NAND2_X1 i_257_76_8167 (.A1(n_257_913), .A2(n_257_439), .ZN(n_257_76_8153));
   NAND2_X1 i_257_76_8168 (.A1(n_257_447), .A2(n_257_779), .ZN(n_257_76_8154));
   NAND2_X1 i_257_76_8169 (.A1(n_257_76_8153), .A2(n_257_76_8154), .ZN(
      n_257_76_8155));
   INV_X1 i_257_76_8170 (.A(n_257_76_8155), .ZN(n_257_76_8156));
   NAND3_X1 i_257_76_8171 (.A1(n_257_76_8143), .A2(n_257_643), .A3(n_257_450), 
      .ZN(n_257_76_8157));
   INV_X1 i_257_76_8172 (.A(n_257_76_8157), .ZN(n_257_76_8158));
   NAND2_X1 i_257_76_8173 (.A1(n_257_440), .A2(n_257_945), .ZN(n_257_76_8159));
   NAND2_X1 i_257_76_8174 (.A1(n_257_438), .A2(n_257_1079), .ZN(n_257_76_8160));
   NAND2_X1 i_257_76_8175 (.A1(n_257_715), .A2(n_257_435), .ZN(n_257_76_8161));
   NAND4_X1 i_257_76_8176 (.A1(n_257_76_8158), .A2(n_257_76_8159), .A3(
      n_257_76_8160), .A4(n_257_76_8161), .ZN(n_257_76_8162));
   INV_X1 i_257_76_8177 (.A(n_257_76_8162), .ZN(n_257_76_8163));
   NAND4_X1 i_257_76_8178 (.A1(n_257_76_8152), .A2(n_257_76_8156), .A3(
      n_257_76_8163), .A4(n_257_76_8131), .ZN(n_257_76_8164));
   NAND2_X1 i_257_76_8179 (.A1(n_257_747), .A2(n_257_436), .ZN(n_257_76_8165));
   NAND2_X1 i_257_76_8180 (.A1(n_257_811), .A2(n_257_437), .ZN(n_257_76_8166));
   NAND2_X1 i_257_76_8181 (.A1(n_257_875), .A2(n_257_445), .ZN(n_257_76_8167));
   NAND3_X1 i_257_76_8182 (.A1(n_257_76_8165), .A2(n_257_76_8166), .A3(
      n_257_76_8167), .ZN(n_257_76_8168));
   NOR2_X1 i_257_76_8183 (.A1(n_257_76_8164), .A2(n_257_76_8168), .ZN(
      n_257_76_8169));
   NAND2_X1 i_257_76_8184 (.A1(n_257_683), .A2(n_257_448), .ZN(n_257_76_8170));
   NAND3_X1 i_257_76_8185 (.A1(n_257_76_8169), .A2(n_257_76_8170), .A3(
      n_257_76_8130), .ZN(n_257_76_8171));
   INV_X1 i_257_76_8186 (.A(n_257_76_8129), .ZN(n_257_76_8172));
   NOR2_X1 i_257_76_8187 (.A1(n_257_76_8171), .A2(n_257_76_8172), .ZN(
      n_257_76_8173));
   NAND2_X1 i_257_76_8188 (.A1(n_257_28), .A2(n_257_76_8173), .ZN(n_257_76_8174));
   NAND3_X1 i_257_76_8189 (.A1(n_257_76_8142), .A2(n_257_76_8148), .A3(
      n_257_76_8174), .ZN(n_257_76_8175));
   INV_X1 i_257_76_8190 (.A(n_257_76_8143), .ZN(n_257_76_8176));
   INV_X1 i_257_76_8191 (.A(n_257_843), .ZN(n_257_76_8177));
   NOR2_X1 i_257_76_8192 (.A1(n_257_76_8176), .A2(n_257_76_8177), .ZN(
      n_257_76_8178));
   NAND4_X1 i_257_76_8193 (.A1(n_257_446), .A2(n_257_76_8178), .A3(n_257_76_8159), 
      .A4(n_257_76_8160), .ZN(n_257_76_8179));
   INV_X1 i_257_76_8194 (.A(n_257_76_8179), .ZN(n_257_76_8180));
   NAND4_X1 i_257_76_8195 (.A1(n_257_76_8180), .A2(n_257_76_8167), .A3(
      n_257_76_8131), .A4(n_257_76_8153), .ZN(n_257_76_8181));
   INV_X1 i_257_76_8196 (.A(n_257_76_8181), .ZN(n_257_76_8182));
   NAND2_X1 i_257_76_8197 (.A1(n_257_76_8130), .A2(n_257_76_8182), .ZN(
      n_257_76_8183));
   INV_X1 i_257_76_8198 (.A(n_257_76_8183), .ZN(n_257_76_8184));
   NAND2_X1 i_257_76_8199 (.A1(n_257_76_8129), .A2(n_257_76_8184), .ZN(
      n_257_76_8185));
   INV_X1 i_257_76_8200 (.A(n_257_76_8185), .ZN(n_257_76_8186));
   NAND2_X1 i_257_76_8201 (.A1(n_257_76_18070), .A2(n_257_76_8186), .ZN(
      n_257_76_8187));
   NAND2_X1 i_257_76_8202 (.A1(n_257_439), .A2(n_257_76_8143), .ZN(n_257_76_8188));
   INV_X1 i_257_76_8203 (.A(n_257_76_8188), .ZN(n_257_76_8189));
   NAND3_X1 i_257_76_8204 (.A1(n_257_913), .A2(n_257_76_8189), .A3(n_257_76_8159), 
      .ZN(n_257_76_8190));
   INV_X1 i_257_76_8205 (.A(n_257_76_8190), .ZN(n_257_76_8191));
   NAND2_X1 i_257_76_8206 (.A1(n_257_76_8131), .A2(n_257_76_8191), .ZN(
      n_257_76_8192));
   INV_X1 i_257_76_8207 (.A(n_257_76_8192), .ZN(n_257_76_8193));
   NAND2_X1 i_257_76_8208 (.A1(n_257_76_8130), .A2(n_257_76_8193), .ZN(
      n_257_76_8194));
   INV_X1 i_257_76_8209 (.A(n_257_76_8194), .ZN(n_257_76_8195));
   NAND2_X1 i_257_76_8210 (.A1(n_257_76_8129), .A2(n_257_76_8195), .ZN(
      n_257_76_8196));
   INV_X1 i_257_76_8211 (.A(n_257_76_8196), .ZN(n_257_76_8197));
   NAND2_X1 i_257_76_8212 (.A1(n_257_76_18084), .A2(n_257_76_8197), .ZN(
      n_257_76_8198));
   NAND2_X1 i_257_76_8213 (.A1(n_257_127), .A2(n_257_430), .ZN(n_257_76_8199));
   NAND2_X1 i_257_76_8214 (.A1(n_257_451), .A2(n_257_466), .ZN(n_257_76_8200));
   NAND4_X1 i_257_76_8215 (.A1(n_257_76_8131), .A2(n_257_76_8199), .A3(n_257_286), 
      .A4(n_257_76_8200), .ZN(n_257_76_8201));
   NAND2_X1 i_257_76_8216 (.A1(n_257_76_8166), .A2(n_257_76_8167), .ZN(
      n_257_76_8202));
   NOR2_X1 i_257_76_8217 (.A1(n_257_76_8201), .A2(n_257_76_8202), .ZN(
      n_257_76_8203));
   NAND2_X1 i_257_76_8218 (.A1(n_257_89), .A2(n_257_431), .ZN(n_257_76_8204));
   NAND2_X1 i_257_76_8219 (.A1(n_257_76_8204), .A2(n_257_76_8165), .ZN(
      n_257_76_8205));
   INV_X1 i_257_76_8220 (.A(n_257_76_8205), .ZN(n_257_76_8206));
   NAND2_X1 i_257_76_8221 (.A1(n_257_643), .A2(n_257_450), .ZN(n_257_76_8207));
   NAND3_X1 i_257_76_8222 (.A1(n_257_76_8160), .A2(n_257_76_8161), .A3(
      n_257_76_8207), .ZN(n_257_76_8208));
   INV_X1 i_257_76_8223 (.A(n_257_76_8208), .ZN(n_257_76_8209));
   NAND2_X1 i_257_76_8224 (.A1(n_257_49), .A2(n_257_433), .ZN(n_257_76_8210));
   NAND2_X1 i_257_76_8225 (.A1(n_257_76_8210), .A2(n_257_76_8159), .ZN(
      n_257_76_8211));
   INV_X1 i_257_76_8226 (.A(n_257_76_8211), .ZN(n_257_76_8212));
   NAND2_X1 i_257_76_8227 (.A1(n_257_427), .A2(n_257_206), .ZN(n_257_76_8213));
   NAND2_X1 i_257_76_8228 (.A1(n_257_432), .A2(n_257_611), .ZN(n_257_76_8214));
   INV_X1 i_257_76_8229 (.A(n_257_1073), .ZN(n_257_76_8215));
   NAND2_X1 i_257_76_8230 (.A1(n_257_76_8214), .A2(n_257_76_8215), .ZN(
      n_257_76_8216));
   INV_X1 i_257_76_8231 (.A(n_257_76_8216), .ZN(n_257_76_8217));
   NAND2_X1 i_257_76_8232 (.A1(n_257_515), .A2(n_257_424), .ZN(n_257_76_8218));
   INV_X1 i_257_76_8233 (.A(n_257_579), .ZN(n_257_76_8219));
   NAND2_X1 i_257_76_8234 (.A1(n_257_76_8219), .A2(n_257_442), .ZN(n_257_76_8220));
   OAI21_X1 i_257_76_8235 (.A(n_257_76_8220), .B1(n_257_428), .B2(n_257_76_17412), 
      .ZN(n_257_76_8221));
   NAND2_X1 i_257_76_8236 (.A1(n_257_76_8221), .A2(n_257_423), .ZN(n_257_76_8222));
   INV_X1 i_257_76_8237 (.A(n_257_76_8222), .ZN(n_257_76_8223));
   NAND4_X1 i_257_76_8238 (.A1(n_257_76_8213), .A2(n_257_76_8217), .A3(
      n_257_76_8218), .A4(n_257_76_8223), .ZN(n_257_76_8224));
   INV_X1 i_257_76_8239 (.A(n_257_76_8224), .ZN(n_257_76_8225));
   NAND2_X1 i_257_76_8240 (.A1(n_257_547), .A2(n_257_426), .ZN(n_257_76_8226));
   NAND4_X1 i_257_76_8241 (.A1(n_257_76_8209), .A2(n_257_76_8212), .A3(
      n_257_76_8225), .A4(n_257_76_8226), .ZN(n_257_76_8227));
   NAND4_X1 i_257_76_8242 (.A1(n_257_76_8149), .A2(n_257_76_8150), .A3(
      n_257_76_8153), .A4(n_257_76_8154), .ZN(n_257_76_8228));
   NOR2_X1 i_257_76_8243 (.A1(n_257_76_8227), .A2(n_257_76_8228), .ZN(
      n_257_76_8229));
   NAND3_X1 i_257_76_8244 (.A1(n_257_76_8203), .A2(n_257_76_8206), .A3(
      n_257_76_8229), .ZN(n_257_76_8230));
   INV_X1 i_257_76_8245 (.A(n_257_76_8230), .ZN(n_257_76_8231));
   NAND2_X1 i_257_76_8246 (.A1(n_257_76_8129), .A2(n_257_76_8231), .ZN(
      n_257_76_8232));
   NAND2_X1 i_257_76_8247 (.A1(n_257_166), .A2(n_257_429), .ZN(n_257_76_8233));
   NAND2_X1 i_257_76_8248 (.A1(n_257_246), .A2(n_257_425), .ZN(n_257_76_8234));
   NAND4_X1 i_257_76_8249 (.A1(n_257_76_8170), .A2(n_257_76_8233), .A3(
      n_257_76_8130), .A4(n_257_76_8234), .ZN(n_257_76_8235));
   NOR2_X1 i_257_76_8250 (.A1(n_257_76_8232), .A2(n_257_76_8235), .ZN(
      n_257_76_8236));
   NAND2_X1 i_257_76_8251 (.A1(n_257_76_18066), .A2(n_257_76_8236), .ZN(
      n_257_76_8237));
   NAND3_X1 i_257_76_8252 (.A1(n_257_76_8187), .A2(n_257_76_8198), .A3(
      n_257_76_8237), .ZN(n_257_76_8238));
   NOR2_X1 i_257_76_8253 (.A1(n_257_76_8175), .A2(n_257_76_8238), .ZN(
      n_257_76_8239));
   INV_X1 i_257_76_8254 (.A(n_257_977), .ZN(n_257_76_8240));
   NOR2_X1 i_257_76_8255 (.A1(n_257_76_8176), .A2(n_257_76_8240), .ZN(
      n_257_76_8241));
   NAND2_X1 i_257_76_8256 (.A1(n_257_441), .A2(n_257_76_8241), .ZN(n_257_76_8242));
   INV_X1 i_257_76_8257 (.A(n_257_76_8242), .ZN(n_257_76_8243));
   NAND2_X1 i_257_76_8258 (.A1(n_257_76_8130), .A2(n_257_76_8243), .ZN(
      n_257_76_8244));
   INV_X1 i_257_76_8259 (.A(n_257_76_8244), .ZN(n_257_76_8245));
   NAND2_X1 i_257_76_8260 (.A1(n_257_76_8129), .A2(n_257_76_8245), .ZN(
      n_257_76_8246));
   INV_X1 i_257_76_8261 (.A(n_257_76_8246), .ZN(n_257_76_8247));
   NAND2_X1 i_257_76_8262 (.A1(n_257_76_18071), .A2(n_257_76_8247), .ZN(
      n_257_76_8248));
   NOR2_X1 i_257_76_8263 (.A1(n_257_76_8176), .A2(n_257_76_17760), .ZN(
      n_257_76_8249));
   NAND4_X1 i_257_76_8264 (.A1(n_257_76_8249), .A2(n_257_76_8159), .A3(
      n_257_76_8160), .A4(n_257_715), .ZN(n_257_76_8250));
   INV_X1 i_257_76_8265 (.A(n_257_76_8250), .ZN(n_257_76_8251));
   NAND4_X1 i_257_76_8266 (.A1(n_257_76_8156), .A2(n_257_76_8251), .A3(
      n_257_76_8131), .A4(n_257_76_8149), .ZN(n_257_76_8252));
   NOR2_X1 i_257_76_8267 (.A1(n_257_76_8168), .A2(n_257_76_8252), .ZN(
      n_257_76_8253));
   NAND2_X1 i_257_76_8268 (.A1(n_257_76_8130), .A2(n_257_76_8253), .ZN(
      n_257_76_8254));
   NOR2_X1 i_257_76_8269 (.A1(n_257_76_8172), .A2(n_257_76_8254), .ZN(
      n_257_76_8255));
   NAND2_X1 i_257_76_8270 (.A1(n_257_76_18078), .A2(n_257_76_8255), .ZN(
      n_257_76_8256));
   NAND3_X1 i_257_76_8271 (.A1(n_257_76_8210), .A2(n_257_76_8159), .A3(
      n_257_76_8160), .ZN(n_257_76_8257));
   NAND2_X1 i_257_76_8272 (.A1(n_257_442), .A2(n_257_579), .ZN(n_257_76_8258));
   INV_X1 i_257_76_8273 (.A(n_257_76_8258), .ZN(n_257_76_8259));
   NAND2_X1 i_257_76_8274 (.A1(n_257_428), .A2(n_257_76_8259), .ZN(n_257_76_8260));
   INV_X1 i_257_76_8275 (.A(n_257_76_8260), .ZN(n_257_76_8261));
   NAND3_X1 i_257_76_8276 (.A1(n_257_76_8214), .A2(n_257_76_8215), .A3(
      n_257_76_8261), .ZN(n_257_76_8262));
   INV_X1 i_257_76_8277 (.A(n_257_76_8262), .ZN(n_257_76_8263));
   NAND3_X1 i_257_76_8278 (.A1(n_257_76_8161), .A2(n_257_76_8207), .A3(
      n_257_76_8263), .ZN(n_257_76_8264));
   NOR2_X1 i_257_76_8279 (.A1(n_257_76_8257), .A2(n_257_76_8264), .ZN(
      n_257_76_8265));
   NAND3_X1 i_257_76_8280 (.A1(n_257_76_8265), .A2(n_257_76_8152), .A3(
      n_257_76_8156), .ZN(n_257_76_8266));
   NAND4_X1 i_257_76_8281 (.A1(n_257_76_8167), .A2(n_257_76_8131), .A3(
      n_257_76_8199), .A4(n_257_76_8200), .ZN(n_257_76_8267));
   NOR2_X1 i_257_76_8282 (.A1(n_257_76_8266), .A2(n_257_76_8267), .ZN(
      n_257_76_8268));
   NAND3_X1 i_257_76_8283 (.A1(n_257_76_8204), .A2(n_257_76_8165), .A3(
      n_257_76_8166), .ZN(n_257_76_8269));
   INV_X1 i_257_76_8284 (.A(n_257_76_8269), .ZN(n_257_76_8270));
   NAND3_X1 i_257_76_8285 (.A1(n_257_76_8268), .A2(n_257_76_8130), .A3(
      n_257_76_8270), .ZN(n_257_76_8271));
   INV_X1 i_257_76_8286 (.A(n_257_76_8271), .ZN(n_257_76_8272));
   NAND2_X1 i_257_76_8287 (.A1(n_257_76_8170), .A2(n_257_76_8233), .ZN(
      n_257_76_8273));
   INV_X1 i_257_76_8288 (.A(n_257_76_8273), .ZN(n_257_76_8274));
   NAND3_X1 i_257_76_8289 (.A1(n_257_76_8272), .A2(n_257_76_8274), .A3(
      n_257_76_8129), .ZN(n_257_76_8275));
   INV_X1 i_257_76_8290 (.A(n_257_76_8275), .ZN(n_257_76_8276));
   NAND2_X1 i_257_76_8291 (.A1(n_257_76_18074), .A2(n_257_76_8276), .ZN(
      n_257_76_8277));
   NAND3_X1 i_257_76_8292 (.A1(n_257_76_8248), .A2(n_257_76_8256), .A3(
      n_257_76_8277), .ZN(n_257_76_8278));
   NAND2_X1 i_257_76_8293 (.A1(n_257_1073), .A2(n_257_442), .ZN(n_257_76_8279));
   INV_X1 i_257_76_8294 (.A(n_257_76_8279), .ZN(n_257_76_8280));
   NAND2_X1 i_257_76_8295 (.A1(n_257_13), .A2(n_257_76_8280), .ZN(n_257_76_8281));
   NOR2_X1 i_257_76_8296 (.A1(n_257_76_8176), .A2(n_257_76_11918), .ZN(
      n_257_76_8282));
   NAND3_X1 i_257_76_8297 (.A1(n_257_76_8282), .A2(n_257_76_8159), .A3(
      n_257_76_8160), .ZN(n_257_76_8283));
   INV_X1 i_257_76_8298 (.A(n_257_76_8283), .ZN(n_257_76_8284));
   NAND4_X1 i_257_76_8299 (.A1(n_257_76_8131), .A2(n_257_76_8284), .A3(n_257_875), 
      .A4(n_257_76_8153), .ZN(n_257_76_8285));
   INV_X1 i_257_76_8300 (.A(n_257_76_8285), .ZN(n_257_76_8286));
   NAND2_X1 i_257_76_8301 (.A1(n_257_76_8130), .A2(n_257_76_8286), .ZN(
      n_257_76_8287));
   INV_X1 i_257_76_8302 (.A(n_257_76_8287), .ZN(n_257_76_8288));
   NAND2_X1 i_257_76_8303 (.A1(n_257_76_8129), .A2(n_257_76_8288), .ZN(
      n_257_76_8289));
   INV_X1 i_257_76_8304 (.A(n_257_76_8289), .ZN(n_257_76_8290));
   NAND2_X1 i_257_76_8305 (.A1(n_257_76_18077), .A2(n_257_76_8290), .ZN(
      n_257_76_8291));
   NAND2_X1 i_257_76_8306 (.A1(n_257_76_8281), .A2(n_257_76_8291), .ZN(
      n_257_76_8292));
   NOR2_X1 i_257_76_8307 (.A1(n_257_76_8278), .A2(n_257_76_8292), .ZN(
      n_257_76_8293));
   NAND4_X1 i_257_76_8308 (.A1(n_257_76_8210), .A2(n_257_76_8159), .A3(
      n_257_76_8160), .A4(n_257_76_8161), .ZN(n_257_76_8294));
   INV_X1 i_257_76_8309 (.A(n_257_76_8294), .ZN(n_257_76_8295));
   NAND4_X1 i_257_76_8310 (.A1(n_257_76_8214), .A2(n_257_76_8215), .A3(
      n_257_76_8221), .A4(n_257_426), .ZN(n_257_76_8296));
   INV_X1 i_257_76_8311 (.A(n_257_76_8296), .ZN(n_257_76_8297));
   NAND4_X1 i_257_76_8312 (.A1(n_257_76_8297), .A2(n_257_547), .A3(n_257_76_8207), 
      .A4(n_257_76_8213), .ZN(n_257_76_8298));
   INV_X1 i_257_76_8313 (.A(n_257_76_8298), .ZN(n_257_76_8299));
   NAND4_X1 i_257_76_8314 (.A1(n_257_76_8295), .A2(n_257_76_8299), .A3(
      n_257_76_8199), .A4(n_257_76_8153), .ZN(n_257_76_8300));
   NOR2_X1 i_257_76_8315 (.A1(n_257_76_8205), .A2(n_257_76_8300), .ZN(
      n_257_76_8301));
   NAND3_X1 i_257_76_8316 (.A1(n_257_76_8166), .A2(n_257_76_8167), .A3(
      n_257_76_8131), .ZN(n_257_76_8302));
   NAND4_X1 i_257_76_8317 (.A1(n_257_76_8200), .A2(n_257_76_8149), .A3(
      n_257_76_8150), .A4(n_257_76_8154), .ZN(n_257_76_8303));
   NOR2_X1 i_257_76_8318 (.A1(n_257_76_8302), .A2(n_257_76_8303), .ZN(
      n_257_76_8304));
   NAND3_X1 i_257_76_8319 (.A1(n_257_76_8301), .A2(n_257_76_8130), .A3(
      n_257_76_8304), .ZN(n_257_76_8305));
   INV_X1 i_257_76_8320 (.A(n_257_76_8305), .ZN(n_257_76_8306));
   NAND3_X1 i_257_76_8321 (.A1(n_257_76_8306), .A2(n_257_76_8274), .A3(
      n_257_76_8129), .ZN(n_257_76_8307));
   INV_X1 i_257_76_8322 (.A(n_257_76_8307), .ZN(n_257_76_8308));
   NAND2_X1 i_257_76_8323 (.A1(n_257_76_18076), .A2(n_257_76_8308), .ZN(
      n_257_76_8309));
   INV_X1 i_257_76_8324 (.A(n_257_76_8154), .ZN(n_257_76_8310));
   INV_X1 i_257_76_8325 (.A(n_257_436), .ZN(n_257_76_8311));
   NOR2_X1 i_257_76_8326 (.A1(n_257_76_8176), .A2(n_257_76_8311), .ZN(
      n_257_76_8312));
   NAND3_X1 i_257_76_8327 (.A1(n_257_76_8312), .A2(n_257_76_8159), .A3(
      n_257_76_8160), .ZN(n_257_76_8313));
   NOR2_X1 i_257_76_8328 (.A1(n_257_76_8310), .A2(n_257_76_8313), .ZN(
      n_257_76_8314));
   NAND2_X1 i_257_76_8329 (.A1(n_257_76_8149), .A2(n_257_76_8153), .ZN(
      n_257_76_8315));
   INV_X1 i_257_76_8330 (.A(n_257_76_8315), .ZN(n_257_76_8316));
   NAND3_X1 i_257_76_8331 (.A1(n_257_76_8314), .A2(n_257_76_8316), .A3(
      n_257_76_8131), .ZN(n_257_76_8317));
   NAND3_X1 i_257_76_8332 (.A1(n_257_76_8166), .A2(n_257_76_8167), .A3(n_257_747), 
      .ZN(n_257_76_8318));
   NOR2_X1 i_257_76_8333 (.A1(n_257_76_8317), .A2(n_257_76_8318), .ZN(
      n_257_76_8319));
   NAND2_X1 i_257_76_8334 (.A1(n_257_76_8130), .A2(n_257_76_8319), .ZN(
      n_257_76_8320));
   NOR2_X1 i_257_76_8335 (.A1(n_257_76_8172), .A2(n_257_76_8320), .ZN(
      n_257_76_8321));
   NAND2_X1 i_257_76_8336 (.A1(n_257_76_18069), .A2(n_257_76_8321), .ZN(
      n_257_76_8322));
   NAND2_X1 i_257_76_8337 (.A1(n_257_611), .A2(n_257_442), .ZN(n_257_76_8323));
   INV_X1 i_257_76_8338 (.A(n_257_76_8323), .ZN(n_257_76_8324));
   NAND2_X1 i_257_76_8339 (.A1(n_257_432), .A2(n_257_76_8324), .ZN(n_257_76_8325));
   NOR2_X1 i_257_76_8340 (.A1(n_257_76_8325), .A2(n_257_1073), .ZN(n_257_76_8326));
   NAND3_X1 i_257_76_8341 (.A1(n_257_76_8161), .A2(n_257_76_8207), .A3(
      n_257_76_8326), .ZN(n_257_76_8327));
   NOR2_X1 i_257_76_8342 (.A1(n_257_76_8257), .A2(n_257_76_8327), .ZN(
      n_257_76_8328));
   NAND3_X1 i_257_76_8343 (.A1(n_257_76_8150), .A2(n_257_76_8153), .A3(
      n_257_76_8154), .ZN(n_257_76_8329));
   INV_X1 i_257_76_8344 (.A(n_257_76_8329), .ZN(n_257_76_8330));
   NAND2_X1 i_257_76_8345 (.A1(n_257_76_8200), .A2(n_257_76_8149), .ZN(
      n_257_76_8331));
   INV_X1 i_257_76_8346 (.A(n_257_76_8331), .ZN(n_257_76_8332));
   NAND4_X1 i_257_76_8347 (.A1(n_257_76_8328), .A2(n_257_76_8330), .A3(
      n_257_76_8332), .A4(n_257_76_8131), .ZN(n_257_76_8333));
   NOR2_X1 i_257_76_8348 (.A1(n_257_76_8333), .A2(n_257_76_8168), .ZN(
      n_257_76_8334));
   NAND3_X1 i_257_76_8349 (.A1(n_257_76_8334), .A2(n_257_76_8170), .A3(
      n_257_76_8130), .ZN(n_257_76_8335));
   NOR2_X1 i_257_76_8350 (.A1(n_257_76_8335), .A2(n_257_76_8172), .ZN(
      n_257_76_8336));
   NAND2_X1 i_257_76_8351 (.A1(n_257_68), .A2(n_257_76_8336), .ZN(n_257_76_8337));
   NAND3_X1 i_257_76_8352 (.A1(n_257_76_8309), .A2(n_257_76_8322), .A3(
      n_257_76_8337), .ZN(n_257_76_8338));
   NOR2_X1 i_257_76_8353 (.A1(n_257_76_8176), .A2(n_257_76_15924), .ZN(
      n_257_76_8339));
   NAND3_X1 i_257_76_8354 (.A1(n_257_76_8339), .A2(n_257_76_8159), .A3(
      n_257_76_8160), .ZN(n_257_76_8340));
   INV_X1 i_257_76_8355 (.A(n_257_76_8340), .ZN(n_257_76_8341));
   NAND4_X1 i_257_76_8356 (.A1(n_257_76_8341), .A2(n_257_811), .A3(n_257_76_8149), 
      .A4(n_257_76_8153), .ZN(n_257_76_8342));
   NAND2_X1 i_257_76_8357 (.A1(n_257_76_8167), .A2(n_257_76_8131), .ZN(
      n_257_76_8343));
   NOR2_X1 i_257_76_8358 (.A1(n_257_76_8342), .A2(n_257_76_8343), .ZN(
      n_257_76_8344));
   NAND2_X1 i_257_76_8359 (.A1(n_257_76_8130), .A2(n_257_76_8344), .ZN(
      n_257_76_8345));
   INV_X1 i_257_76_8360 (.A(n_257_76_8345), .ZN(n_257_76_8346));
   NAND2_X1 i_257_76_8361 (.A1(n_257_76_8129), .A2(n_257_76_8346), .ZN(
      n_257_76_8347));
   INV_X1 i_257_76_8362 (.A(n_257_76_8347), .ZN(n_257_76_8348));
   NAND2_X1 i_257_76_8363 (.A1(n_257_22), .A2(n_257_76_8348), .ZN(n_257_76_8349));
   NAND2_X1 i_257_76_8364 (.A1(n_257_444), .A2(n_257_76_8143), .ZN(n_257_76_8350));
   INV_X1 i_257_76_8365 (.A(n_257_76_8350), .ZN(n_257_76_8351));
   NAND2_X1 i_257_76_8366 (.A1(n_257_1009), .A2(n_257_76_8351), .ZN(
      n_257_76_8352));
   INV_X1 i_257_76_8367 (.A(n_257_76_8352), .ZN(n_257_76_8353));
   NAND2_X1 i_257_76_8368 (.A1(n_257_76_8129), .A2(n_257_76_8353), .ZN(
      n_257_76_8354));
   INV_X1 i_257_76_8369 (.A(n_257_76_8354), .ZN(n_257_76_8355));
   NAND2_X1 i_257_76_8370 (.A1(n_257_76_18075), .A2(n_257_76_8355), .ZN(
      n_257_76_8356));
   NAND2_X1 i_257_76_8371 (.A1(n_257_76_8349), .A2(n_257_76_8356), .ZN(
      n_257_76_8357));
   NOR2_X1 i_257_76_8372 (.A1(n_257_76_8338), .A2(n_257_76_8357), .ZN(
      n_257_76_8358));
   NAND3_X1 i_257_76_8373 (.A1(n_257_76_8239), .A2(n_257_76_8293), .A3(
      n_257_76_8358), .ZN(n_257_76_8359));
   INV_X1 i_257_76_8374 (.A(n_257_76_8359), .ZN(n_257_76_8360));
   NAND3_X1 i_257_76_8375 (.A1(n_257_76_8159), .A2(n_257_76_8160), .A3(
      n_257_76_8161), .ZN(n_257_76_8361));
   NOR2_X1 i_257_76_8376 (.A1(n_257_1073), .A2(n_257_76_17633), .ZN(
      n_257_76_8362));
   NAND3_X1 i_257_76_8377 (.A1(n_257_76_8207), .A2(n_257_49), .A3(n_257_76_8362), 
      .ZN(n_257_76_8363));
   NOR2_X1 i_257_76_8378 (.A1(n_257_76_8361), .A2(n_257_76_8363), .ZN(
      n_257_76_8364));
   NAND4_X1 i_257_76_8379 (.A1(n_257_76_8330), .A2(n_257_76_8332), .A3(
      n_257_76_8364), .A4(n_257_76_8131), .ZN(n_257_76_8365));
   NOR2_X1 i_257_76_8380 (.A1(n_257_76_8365), .A2(n_257_76_8168), .ZN(
      n_257_76_8366));
   NAND3_X1 i_257_76_8381 (.A1(n_257_76_8366), .A2(n_257_76_8170), .A3(
      n_257_76_8130), .ZN(n_257_76_8367));
   NOR2_X1 i_257_76_8382 (.A1(n_257_76_8367), .A2(n_257_76_8172), .ZN(
      n_257_76_8368));
   NAND2_X1 i_257_76_8383 (.A1(n_257_76_18081), .A2(n_257_76_8368), .ZN(
      n_257_76_8369));
   INV_X1 i_257_76_8384 (.A(n_257_76_8168), .ZN(n_257_76_8370));
   NAND3_X1 i_257_76_8385 (.A1(n_257_76_8149), .A2(n_257_76_8153), .A3(
      n_257_76_8154), .ZN(n_257_76_8371));
   INV_X1 i_257_76_8386 (.A(n_257_76_8371), .ZN(n_257_76_8372));
   NOR2_X1 i_257_76_8387 (.A1(n_257_76_8176), .A2(n_257_76_15906), .ZN(
      n_257_76_8373));
   NAND3_X1 i_257_76_8388 (.A1(n_257_76_8373), .A2(n_257_76_8160), .A3(
      n_257_76_8161), .ZN(n_257_76_8374));
   NAND2_X1 i_257_76_8389 (.A1(n_257_449), .A2(n_257_76_8159), .ZN(n_257_76_8375));
   NOR2_X1 i_257_76_8390 (.A1(n_257_76_8374), .A2(n_257_76_8375), .ZN(
      n_257_76_8376));
   NAND3_X1 i_257_76_8391 (.A1(n_257_76_8372), .A2(n_257_76_8376), .A3(
      n_257_76_8131), .ZN(n_257_76_8377));
   INV_X1 i_257_76_8392 (.A(n_257_76_8377), .ZN(n_257_76_8378));
   NAND2_X1 i_257_76_8393 (.A1(n_257_76_8370), .A2(n_257_76_8378), .ZN(
      n_257_76_8379));
   INV_X1 i_257_76_8394 (.A(n_257_76_8130), .ZN(n_257_76_8380));
   NOR2_X1 i_257_76_8395 (.A1(n_257_76_8379), .A2(n_257_76_8380), .ZN(
      n_257_76_8381));
   NAND3_X1 i_257_76_8396 (.A1(n_257_76_8381), .A2(n_257_76_8129), .A3(
      n_257_76_8170), .ZN(n_257_76_8382));
   INV_X1 i_257_76_8397 (.A(n_257_76_8382), .ZN(n_257_76_8383));
   NAND2_X1 i_257_76_8398 (.A1(n_257_76_18083), .A2(n_257_76_8383), .ZN(
      n_257_76_8384));
   NAND4_X1 i_257_76_8399 (.A1(n_257_76_8204), .A2(n_257_76_8165), .A3(
      n_257_76_8166), .A4(n_257_76_8167), .ZN(n_257_76_8385));
   NAND4_X1 i_257_76_8400 (.A1(n_257_76_8200), .A2(n_257_76_8149), .A3(
      n_257_76_8150), .A4(n_257_76_8153), .ZN(n_257_76_8386));
   INV_X1 i_257_76_8401 (.A(n_257_76_8386), .ZN(n_257_76_8387));
   NAND2_X1 i_257_76_8402 (.A1(n_257_76_8131), .A2(n_257_76_8199), .ZN(
      n_257_76_8388));
   INV_X1 i_257_76_8403 (.A(n_257_76_8388), .ZN(n_257_76_8389));
   INV_X1 i_257_76_8404 (.A(n_257_76_8257), .ZN(n_257_76_8390));
   NAND3_X1 i_257_76_8405 (.A1(n_257_76_8214), .A2(n_257_76_8215), .A3(
      n_257_76_17331), .ZN(n_257_76_8391));
   INV_X1 i_257_76_8406 (.A(n_257_76_8391), .ZN(n_257_76_8392));
   NAND3_X1 i_257_76_8407 (.A1(n_257_76_8161), .A2(n_257_76_8207), .A3(
      n_257_76_8392), .ZN(n_257_76_8393));
   INV_X1 i_257_76_8408 (.A(n_257_76_8393), .ZN(n_257_76_8394));
   NAND3_X1 i_257_76_8409 (.A1(n_257_76_8390), .A2(n_257_76_8154), .A3(
      n_257_76_8394), .ZN(n_257_76_8395));
   INV_X1 i_257_76_8410 (.A(n_257_76_8395), .ZN(n_257_76_8396));
   NAND3_X1 i_257_76_8411 (.A1(n_257_76_8387), .A2(n_257_76_8389), .A3(
      n_257_76_8396), .ZN(n_257_76_8397));
   NOR2_X1 i_257_76_8412 (.A1(n_257_76_8385), .A2(n_257_76_8397), .ZN(
      n_257_76_8398));
   NAND2_X1 i_257_76_8413 (.A1(n_257_76_8130), .A2(n_257_166), .ZN(n_257_76_8399));
   INV_X1 i_257_76_8414 (.A(n_257_76_8399), .ZN(n_257_76_8400));
   NAND4_X1 i_257_76_8415 (.A1(n_257_76_8129), .A2(n_257_76_8398), .A3(
      n_257_76_8400), .A4(n_257_76_8170), .ZN(n_257_76_8401));
   INV_X1 i_257_76_8416 (.A(n_257_76_8401), .ZN(n_257_76_8402));
   NAND2_X1 i_257_76_8417 (.A1(n_257_76_18061), .A2(n_257_76_8402), .ZN(
      n_257_76_8403));
   NAND3_X1 i_257_76_8418 (.A1(n_257_76_8369), .A2(n_257_76_8384), .A3(
      n_257_76_8403), .ZN(n_257_76_8404));
   INV_X1 i_257_76_8419 (.A(n_257_76_8404), .ZN(n_257_76_8405));
   NAND2_X1 i_257_76_8420 (.A1(n_257_1079), .A2(n_257_76_8143), .ZN(
      n_257_76_8406));
   INV_X1 i_257_76_8421 (.A(n_257_76_8406), .ZN(n_257_76_8407));
   NAND3_X1 i_257_76_8422 (.A1(n_257_76_8407), .A2(n_257_76_8159), .A3(n_257_438), 
      .ZN(n_257_76_8408));
   INV_X1 i_257_76_8423 (.A(n_257_76_8408), .ZN(n_257_76_8409));
   NAND3_X1 i_257_76_8424 (.A1(n_257_76_8131), .A2(n_257_76_8409), .A3(
      n_257_76_8153), .ZN(n_257_76_8410));
   INV_X1 i_257_76_8425 (.A(n_257_76_8410), .ZN(n_257_76_8411));
   NAND2_X1 i_257_76_8426 (.A1(n_257_76_8130), .A2(n_257_76_8411), .ZN(
      n_257_76_8412));
   INV_X1 i_257_76_8427 (.A(n_257_76_8412), .ZN(n_257_76_8413));
   NAND2_X1 i_257_76_8428 (.A1(n_257_76_8129), .A2(n_257_76_8413), .ZN(
      n_257_76_8414));
   INV_X1 i_257_76_8429 (.A(n_257_76_8414), .ZN(n_257_76_8415));
   NAND2_X1 i_257_76_8430 (.A1(n_257_76_18067), .A2(n_257_76_8415), .ZN(
      n_257_76_8416));
   NAND2_X1 i_257_76_8431 (.A1(n_257_76_8234), .A2(n_257_76_8204), .ZN(
      n_257_76_8417));
   INV_X1 i_257_76_8432 (.A(n_257_76_8417), .ZN(n_257_76_8418));
   NAND2_X1 i_257_76_8433 (.A1(n_257_76_8418), .A2(n_257_76_8130), .ZN(
      n_257_76_8419));
   INV_X1 i_257_76_8434 (.A(n_257_76_8419), .ZN(n_257_76_8420));
   NAND2_X1 i_257_76_8435 (.A1(n_257_76_8159), .A2(n_257_76_8160), .ZN(
      n_257_76_8421));
   NAND2_X1 i_257_76_8436 (.A1(n_257_76_8161), .A2(n_257_76_8207), .ZN(
      n_257_76_8422));
   NOR2_X1 i_257_76_8437 (.A1(n_257_76_8421), .A2(n_257_76_8422), .ZN(
      n_257_76_8423));
   NAND2_X1 i_257_76_8438 (.A1(n_257_76_17354), .A2(n_257_76_8219), .ZN(
      n_257_76_8424));
   OAI21_X1 i_257_76_8439 (.A(n_257_76_8424), .B1(n_257_428), .B2(n_257_76_17090), 
      .ZN(n_257_76_8425));
   NAND2_X1 i_257_76_8440 (.A1(n_257_76_8425), .A2(n_257_420), .ZN(n_257_76_8426));
   NOR2_X1 i_257_76_8441 (.A1(n_257_76_8216), .A2(n_257_76_8426), .ZN(
      n_257_76_8427));
   NAND2_X1 i_257_76_8442 (.A1(n_257_76_8427), .A2(n_257_76_8218), .ZN(
      n_257_76_8428));
   NAND2_X1 i_257_76_8443 (.A1(n_257_324), .A2(n_257_422), .ZN(n_257_76_8429));
   NAND2_X1 i_257_76_8444 (.A1(n_257_76_8213), .A2(n_257_76_8429), .ZN(
      n_257_76_8430));
   NOR2_X1 i_257_76_8445 (.A1(n_257_76_8428), .A2(n_257_76_8430), .ZN(
      n_257_76_8431));
   NAND2_X1 i_257_76_8446 (.A1(n_257_76_8423), .A2(n_257_76_8431), .ZN(
      n_257_76_8432));
   NAND2_X1 i_257_76_8447 (.A1(n_257_76_8226), .A2(n_257_76_8210), .ZN(
      n_257_76_8433));
   INV_X1 i_257_76_8448 (.A(n_257_76_8433), .ZN(n_257_76_8434));
   NAND2_X1 i_257_76_8449 (.A1(n_257_76_8156), .A2(n_257_76_8434), .ZN(
      n_257_76_8435));
   NOR2_X1 i_257_76_8450 (.A1(n_257_76_8432), .A2(n_257_76_8435), .ZN(
      n_257_76_8436));
   NAND2_X1 i_257_76_8451 (.A1(n_257_76_8152), .A2(n_257_76_8200), .ZN(
      n_257_76_8437));
   NOR2_X1 i_257_76_8452 (.A1(n_257_76_8437), .A2(n_257_76_8388), .ZN(
      n_257_76_8438));
   NAND2_X1 i_257_76_8453 (.A1(n_257_76_8436), .A2(n_257_76_8438), .ZN(
      n_257_76_8439));
   NAND2_X1 i_257_76_8454 (.A1(n_257_286), .A2(n_257_423), .ZN(n_257_76_8440));
   NAND2_X1 i_257_76_8455 (.A1(n_257_76_8165), .A2(n_257_76_8440), .ZN(
      n_257_76_8441));
   INV_X1 i_257_76_8456 (.A(n_257_76_8441), .ZN(n_257_76_8442));
   NAND2_X1 i_257_76_8457 (.A1(n_257_363), .A2(n_257_421), .ZN(n_257_76_8443));
   NAND2_X1 i_257_76_8458 (.A1(n_257_76_8167), .A2(n_257_76_8443), .ZN(
      n_257_76_8444));
   INV_X1 i_257_76_8459 (.A(n_257_76_8166), .ZN(n_257_76_8445));
   NOR2_X1 i_257_76_8460 (.A1(n_257_76_8444), .A2(n_257_76_8445), .ZN(
      n_257_76_8446));
   NAND2_X1 i_257_76_8461 (.A1(n_257_76_8442), .A2(n_257_76_8446), .ZN(
      n_257_76_8447));
   NOR2_X1 i_257_76_8462 (.A1(n_257_76_8439), .A2(n_257_76_8447), .ZN(
      n_257_76_8448));
   NAND2_X1 i_257_76_8463 (.A1(n_257_76_8420), .A2(n_257_76_8448), .ZN(
      n_257_76_8449));
   NAND2_X1 i_257_76_8464 (.A1(n_257_76_8274), .A2(n_257_76_8129), .ZN(
      n_257_76_8450));
   NOR2_X1 i_257_76_8465 (.A1(n_257_76_8449), .A2(n_257_76_8450), .ZN(
      n_257_76_8451));
   NAND2_X1 i_257_76_8466 (.A1(n_257_76_18073), .A2(n_257_76_8451), .ZN(
      n_257_76_8452));
   NAND3_X1 i_257_76_8467 (.A1(n_257_76_8214), .A2(n_257_76_8215), .A3(
      n_257_76_17925), .ZN(n_257_76_8453));
   INV_X1 i_257_76_8468 (.A(n_257_76_8453), .ZN(n_257_76_8454));
   NAND3_X1 i_257_76_8469 (.A1(n_257_76_8161), .A2(n_257_76_8207), .A3(
      n_257_76_8454), .ZN(n_257_76_8455));
   INV_X1 i_257_76_8470 (.A(n_257_76_8455), .ZN(n_257_76_8456));
   NAND4_X1 i_257_76_8471 (.A1(n_257_76_8390), .A2(n_257_76_8456), .A3(
      n_257_76_8154), .A4(n_257_127), .ZN(n_257_76_8457));
   INV_X1 i_257_76_8472 (.A(n_257_76_8457), .ZN(n_257_76_8458));
   INV_X1 i_257_76_8473 (.A(n_257_76_8343), .ZN(n_257_76_8459));
   NAND3_X1 i_257_76_8474 (.A1(n_257_76_8458), .A2(n_257_76_8459), .A3(
      n_257_76_8387), .ZN(n_257_76_8460));
   NOR2_X1 i_257_76_8475 (.A1(n_257_76_8460), .A2(n_257_76_8269), .ZN(
      n_257_76_8461));
   NAND3_X1 i_257_76_8476 (.A1(n_257_76_8461), .A2(n_257_76_8170), .A3(
      n_257_76_8130), .ZN(n_257_76_8462));
   NOR2_X1 i_257_76_8477 (.A1(n_257_76_8462), .A2(n_257_76_8172), .ZN(
      n_257_76_8463));
   NAND2_X1 i_257_76_8478 (.A1(n_257_76_18068), .A2(n_257_76_8463), .ZN(
      n_257_76_8464));
   NAND3_X1 i_257_76_8479 (.A1(n_257_76_8416), .A2(n_257_76_8452), .A3(
      n_257_76_8464), .ZN(n_257_76_8465));
   INV_X1 i_257_76_8480 (.A(n_257_76_8465), .ZN(n_257_76_8466));
   NAND2_X1 i_257_76_8481 (.A1(n_257_779), .A2(n_257_442), .ZN(n_257_76_8467));
   NOR2_X1 i_257_76_8482 (.A1(n_257_1073), .A2(n_257_76_8467), .ZN(n_257_76_8468));
   NAND4_X1 i_257_76_8483 (.A1(n_257_447), .A2(n_257_76_8159), .A3(n_257_76_8160), 
      .A4(n_257_76_8468), .ZN(n_257_76_8469));
   INV_X1 i_257_76_8484 (.A(n_257_76_8469), .ZN(n_257_76_8470));
   NAND3_X1 i_257_76_8485 (.A1(n_257_76_8316), .A2(n_257_76_8470), .A3(
      n_257_76_8131), .ZN(n_257_76_8471));
   NOR2_X1 i_257_76_8486 (.A1(n_257_76_8471), .A2(n_257_76_8202), .ZN(
      n_257_76_8472));
   NAND2_X1 i_257_76_8487 (.A1(n_257_76_8130), .A2(n_257_76_8472), .ZN(
      n_257_76_8473));
   INV_X1 i_257_76_8488 (.A(n_257_76_8473), .ZN(n_257_76_8474));
   NAND2_X1 i_257_76_8489 (.A1(n_257_76_8129), .A2(n_257_76_8474), .ZN(
      n_257_76_8475));
   INV_X1 i_257_76_8490 (.A(n_257_76_8475), .ZN(n_257_76_8476));
   NAND3_X1 i_257_76_8491 (.A1(n_257_76_8214), .A2(n_257_76_8215), .A3(
      n_257_76_17932), .ZN(n_257_76_8477));
   INV_X1 i_257_76_8492 (.A(n_257_76_8477), .ZN(n_257_76_8478));
   NAND3_X1 i_257_76_8493 (.A1(n_257_76_8161), .A2(n_257_76_8207), .A3(
      n_257_76_8478), .ZN(n_257_76_8479));
   NOR2_X1 i_257_76_8494 (.A1(n_257_76_8257), .A2(n_257_76_8479), .ZN(
      n_257_76_8480));
   NAND4_X1 i_257_76_8495 (.A1(n_257_76_8480), .A2(n_257_76_8330), .A3(
      n_257_76_8332), .A4(n_257_76_8131), .ZN(n_257_76_8481));
   NAND4_X1 i_257_76_8496 (.A1(n_257_76_8165), .A2(n_257_76_8166), .A3(n_257_89), 
      .A4(n_257_76_8167), .ZN(n_257_76_8482));
   NOR2_X1 i_257_76_8497 (.A1(n_257_76_8481), .A2(n_257_76_8482), .ZN(
      n_257_76_8483));
   NAND3_X1 i_257_76_8498 (.A1(n_257_76_8483), .A2(n_257_76_8170), .A3(
      n_257_76_8130), .ZN(n_257_76_8484));
   NOR2_X1 i_257_76_8499 (.A1(n_257_76_8484), .A2(n_257_76_8172), .ZN(
      n_257_76_8485));
   AOI22_X1 i_257_76_8500 (.A1(n_257_76_18085), .A2(n_257_76_8476), .B1(
      n_257_76_18080), .B2(n_257_76_8485), .ZN(n_257_76_8486));
   NAND3_X1 i_257_76_8501 (.A1(n_257_76_8405), .A2(n_257_76_8466), .A3(
      n_257_76_8486), .ZN(n_257_76_8487));
   NAND3_X1 i_257_76_8502 (.A1(n_257_76_8159), .A2(n_257_76_8160), .A3(n_257_448), 
      .ZN(n_257_76_8488));
   NOR2_X1 i_257_76_8503 (.A1(n_257_76_8310), .A2(n_257_76_8488), .ZN(
      n_257_76_8489));
   NAND2_X1 i_257_76_8504 (.A1(n_257_76_8143), .A2(n_257_76_17760), .ZN(
      n_257_76_8490));
   OAI21_X1 i_257_76_8505 (.A(n_257_76_8490), .B1(n_257_715), .B2(n_257_76_8176), 
      .ZN(n_257_76_8491));
   NAND3_X1 i_257_76_8506 (.A1(n_257_76_8149), .A2(n_257_76_8153), .A3(
      n_257_76_8491), .ZN(n_257_76_8492));
   INV_X1 i_257_76_8507 (.A(n_257_76_8492), .ZN(n_257_76_8493));
   NAND3_X1 i_257_76_8508 (.A1(n_257_76_8489), .A2(n_257_76_8493), .A3(
      n_257_76_8131), .ZN(n_257_76_8494));
   NOR2_X1 i_257_76_8509 (.A1(n_257_76_8494), .A2(n_257_76_8168), .ZN(
      n_257_76_8495));
   NAND3_X1 i_257_76_8510 (.A1(n_257_76_8495), .A2(n_257_76_8130), .A3(n_257_683), 
      .ZN(n_257_76_8496));
   NOR2_X1 i_257_76_8511 (.A1(n_257_76_8496), .A2(n_257_76_8172), .ZN(
      n_257_76_8497));
   NAND2_X1 i_257_76_8512 (.A1(n_257_76_18079), .A2(n_257_76_8497), .ZN(
      n_257_76_8498));
   NAND4_X1 i_257_76_8513 (.A1(n_257_76_8214), .A2(n_257_76_8215), .A3(
      n_257_76_8221), .A4(n_257_425), .ZN(n_257_76_8499));
   INV_X1 i_257_76_8514 (.A(n_257_76_8499), .ZN(n_257_76_8500));
   NAND3_X1 i_257_76_8515 (.A1(n_257_76_8500), .A2(n_257_76_8207), .A3(
      n_257_76_8213), .ZN(n_257_76_8501));
   NOR2_X1 i_257_76_8516 (.A1(n_257_76_8361), .A2(n_257_76_8501), .ZN(
      n_257_76_8502));
   NAND3_X1 i_257_76_8517 (.A1(n_257_76_8149), .A2(n_257_76_8150), .A3(
      n_257_76_8153), .ZN(n_257_76_8503));
   INV_X1 i_257_76_8518 (.A(n_257_76_8503), .ZN(n_257_76_8504));
   NAND3_X1 i_257_76_8519 (.A1(n_257_76_8154), .A2(n_257_76_8226), .A3(
      n_257_76_8210), .ZN(n_257_76_8505));
   INV_X1 i_257_76_8520 (.A(n_257_76_8505), .ZN(n_257_76_8506));
   NAND3_X1 i_257_76_8521 (.A1(n_257_76_8502), .A2(n_257_76_8504), .A3(
      n_257_76_8506), .ZN(n_257_76_8507));
   NOR2_X1 i_257_76_8522 (.A1(n_257_76_8507), .A2(n_257_76_8267), .ZN(
      n_257_76_8508));
   NAND4_X1 i_257_76_8523 (.A1(n_257_76_8204), .A2(n_257_246), .A3(n_257_76_8165), 
      .A4(n_257_76_8166), .ZN(n_257_76_8509));
   INV_X1 i_257_76_8524 (.A(n_257_76_8509), .ZN(n_257_76_8510));
   NAND3_X1 i_257_76_8525 (.A1(n_257_76_8508), .A2(n_257_76_8233), .A3(
      n_257_76_8510), .ZN(n_257_76_8511));
   INV_X1 i_257_76_8526 (.A(n_257_76_8511), .ZN(n_257_76_8512));
   NAND2_X1 i_257_76_8527 (.A1(n_257_76_8170), .A2(n_257_76_8130), .ZN(
      n_257_76_8513));
   INV_X1 i_257_76_8528 (.A(n_257_76_8513), .ZN(n_257_76_8514));
   NAND3_X1 i_257_76_8529 (.A1(n_257_76_8512), .A2(n_257_76_8514), .A3(
      n_257_76_8129), .ZN(n_257_76_8515));
   INV_X1 i_257_76_8530 (.A(n_257_76_8515), .ZN(n_257_76_8516));
   NAND2_X1 i_257_76_8531 (.A1(n_257_76_18064), .A2(n_257_76_8516), .ZN(
      n_257_76_8517));
   INV_X1 i_257_76_8532 (.A(n_257_76_8303), .ZN(n_257_76_8518));
   NAND3_X1 i_257_76_8533 (.A1(n_257_76_8459), .A2(n_257_76_8518), .A3(
      n_257_76_8166), .ZN(n_257_76_8519));
   NAND3_X1 i_257_76_8534 (.A1(n_257_76_8204), .A2(n_257_76_8165), .A3(
      n_257_76_8440), .ZN(n_257_76_8520));
   NOR2_X1 i_257_76_8535 (.A1(n_257_76_8519), .A2(n_257_76_8520), .ZN(
      n_257_76_8521));
   NAND2_X1 i_257_76_8536 (.A1(n_257_363), .A2(n_257_76_8153), .ZN(n_257_76_8522));
   INV_X1 i_257_76_8537 (.A(n_257_76_8522), .ZN(n_257_76_8523));
   INV_X1 i_257_76_8538 (.A(n_257_76_8226), .ZN(n_257_76_8524));
   NOR2_X1 i_257_76_8539 (.A1(n_257_76_8257), .A2(n_257_76_8524), .ZN(
      n_257_76_8525));
   NAND3_X1 i_257_76_8540 (.A1(n_257_76_8161), .A2(n_257_76_8207), .A3(
      n_257_76_8213), .ZN(n_257_76_8526));
   NAND2_X1 i_257_76_8541 (.A1(n_257_76_8221), .A2(n_257_421), .ZN(n_257_76_8527));
   INV_X1 i_257_76_8542 (.A(n_257_76_8527), .ZN(n_257_76_8528));
   NAND4_X1 i_257_76_8543 (.A1(n_257_76_8429), .A2(n_257_76_8217), .A3(
      n_257_76_8218), .A4(n_257_76_8528), .ZN(n_257_76_8529));
   NOR2_X1 i_257_76_8544 (.A1(n_257_76_8526), .A2(n_257_76_8529), .ZN(
      n_257_76_8530));
   NAND4_X1 i_257_76_8545 (.A1(n_257_76_8523), .A2(n_257_76_8525), .A3(
      n_257_76_8530), .A4(n_257_76_8199), .ZN(n_257_76_8531));
   INV_X1 i_257_76_8546 (.A(n_257_76_8234), .ZN(n_257_76_8532));
   NOR2_X1 i_257_76_8547 (.A1(n_257_76_8531), .A2(n_257_76_8532), .ZN(
      n_257_76_8533));
   NAND4_X1 i_257_76_8548 (.A1(n_257_76_8521), .A2(n_257_76_8533), .A3(
      n_257_76_8233), .A4(n_257_76_8130), .ZN(n_257_76_8534));
   NAND2_X1 i_257_76_8549 (.A1(n_257_76_8129), .A2(n_257_76_8170), .ZN(
      n_257_76_8535));
   NOR2_X1 i_257_76_8550 (.A1(n_257_76_8534), .A2(n_257_76_8535), .ZN(
      n_257_76_8536));
   NAND2_X1 i_257_76_8551 (.A1(n_257_76_18082), .A2(n_257_76_8536), .ZN(
      n_257_76_8537));
   NAND3_X1 i_257_76_8552 (.A1(n_257_76_8498), .A2(n_257_76_8517), .A3(
      n_257_76_8537), .ZN(n_257_76_8538));
   INV_X1 i_257_76_8553 (.A(n_257_76_8538), .ZN(n_257_76_8539));
   NOR2_X1 i_257_76_8554 (.A1(n_257_76_8208), .A2(n_257_76_8211), .ZN(
      n_257_76_8540));
   NAND3_X1 i_257_76_8555 (.A1(n_257_76_8540), .A2(n_257_76_8152), .A3(
      n_257_76_8156), .ZN(n_257_76_8541));
   INV_X1 i_257_76_8556 (.A(n_257_76_8221), .ZN(n_257_76_8542));
   NOR2_X1 i_257_76_8557 (.A1(n_257_76_8542), .A2(n_257_1073), .ZN(n_257_76_8543));
   NAND4_X1 i_257_76_8558 (.A1(n_257_76_8543), .A2(n_257_427), .A3(n_257_206), 
      .A4(n_257_76_8214), .ZN(n_257_76_8544));
   INV_X1 i_257_76_8559 (.A(n_257_76_8544), .ZN(n_257_76_8545));
   NAND4_X1 i_257_76_8560 (.A1(n_257_76_8131), .A2(n_257_76_8199), .A3(
      n_257_76_8200), .A4(n_257_76_8545), .ZN(n_257_76_8546));
   NOR2_X1 i_257_76_8561 (.A1(n_257_76_8541), .A2(n_257_76_8546), .ZN(
      n_257_76_8547));
   INV_X1 i_257_76_8562 (.A(n_257_76_8385), .ZN(n_257_76_8548));
   NAND3_X1 i_257_76_8563 (.A1(n_257_76_8547), .A2(n_257_76_8130), .A3(
      n_257_76_8548), .ZN(n_257_76_8549));
   INV_X1 i_257_76_8564 (.A(n_257_76_8549), .ZN(n_257_76_8550));
   NAND3_X1 i_257_76_8565 (.A1(n_257_76_8550), .A2(n_257_76_8274), .A3(
      n_257_76_8129), .ZN(n_257_76_8551));
   INV_X1 i_257_76_8566 (.A(n_257_76_8551), .ZN(n_257_76_8552));
   NAND2_X1 i_257_76_8567 (.A1(n_257_76_18065), .A2(n_257_76_8552), .ZN(
      n_257_76_8553));
   INV_X1 i_257_76_8568 (.A(n_257_466), .ZN(n_257_76_8554));
   NOR2_X1 i_257_76_8569 (.A1(n_257_76_8176), .A2(n_257_76_8554), .ZN(
      n_257_76_8555));
   NAND3_X1 i_257_76_8570 (.A1(n_257_76_8555), .A2(n_257_76_8161), .A3(
      n_257_76_8207), .ZN(n_257_76_8556));
   NOR2_X1 i_257_76_8571 (.A1(n_257_76_8556), .A2(n_257_76_8421), .ZN(
      n_257_76_8557));
   NAND3_X1 i_257_76_8572 (.A1(n_257_76_8153), .A2(n_257_76_8154), .A3(n_257_451), 
      .ZN(n_257_76_8558));
   INV_X1 i_257_76_8573 (.A(n_257_76_8558), .ZN(n_257_76_8559));
   NAND4_X1 i_257_76_8574 (.A1(n_257_76_8557), .A2(n_257_76_8559), .A3(
      n_257_76_8152), .A4(n_257_76_8131), .ZN(n_257_76_8560));
   NOR2_X1 i_257_76_8575 (.A1(n_257_76_8560), .A2(n_257_76_8168), .ZN(
      n_257_76_8561));
   NAND3_X1 i_257_76_8576 (.A1(n_257_76_8561), .A2(n_257_76_8170), .A3(
      n_257_76_8130), .ZN(n_257_76_8562));
   NOR2_X1 i_257_76_8577 (.A1(n_257_76_8562), .A2(n_257_76_8172), .ZN(
      n_257_76_8563));
   NAND2_X1 i_257_76_8578 (.A1(n_257_76_18063), .A2(n_257_76_8563), .ZN(
      n_257_76_8564));
   NAND3_X1 i_257_76_8579 (.A1(n_257_76_8215), .A2(n_257_76_8221), .A3(n_257_424), 
      .ZN(n_257_76_8565));
   NAND2_X1 i_257_76_8580 (.A1(n_257_515), .A2(n_257_76_8214), .ZN(n_257_76_8566));
   NOR2_X1 i_257_76_8581 (.A1(n_257_76_8565), .A2(n_257_76_8566), .ZN(
      n_257_76_8567));
   NAND4_X1 i_257_76_8582 (.A1(n_257_76_8567), .A2(n_257_76_8161), .A3(
      n_257_76_8207), .A4(n_257_76_8213), .ZN(n_257_76_8568));
   NOR2_X1 i_257_76_8583 (.A1(n_257_76_8568), .A2(n_257_76_8257), .ZN(
      n_257_76_8569));
   NAND3_X1 i_257_76_8584 (.A1(n_257_76_8200), .A2(n_257_76_8149), .A3(
      n_257_76_8150), .ZN(n_257_76_8570));
   INV_X1 i_257_76_8585 (.A(n_257_76_8570), .ZN(n_257_76_8571));
   NAND3_X1 i_257_76_8586 (.A1(n_257_76_8153), .A2(n_257_76_8154), .A3(
      n_257_76_8226), .ZN(n_257_76_8572));
   INV_X1 i_257_76_8587 (.A(n_257_76_8572), .ZN(n_257_76_8573));
   NAND3_X1 i_257_76_8588 (.A1(n_257_76_8569), .A2(n_257_76_8571), .A3(
      n_257_76_8573), .ZN(n_257_76_8574));
   NAND4_X1 i_257_76_8589 (.A1(n_257_76_8166), .A2(n_257_76_8167), .A3(
      n_257_76_8131), .A4(n_257_76_8199), .ZN(n_257_76_8575));
   NOR2_X1 i_257_76_8590 (.A1(n_257_76_8574), .A2(n_257_76_8575), .ZN(
      n_257_76_8576));
   NOR2_X1 i_257_76_8591 (.A1(n_257_76_8532), .A2(n_257_76_8205), .ZN(
      n_257_76_8577));
   NAND3_X1 i_257_76_8592 (.A1(n_257_76_8576), .A2(n_257_76_8577), .A3(
      n_257_76_8130), .ZN(n_257_76_8578));
   NOR3_X1 i_257_76_8593 (.A1(n_257_76_8578), .A2(n_257_76_8172), .A3(
      n_257_76_8273), .ZN(n_257_76_8579));
   NAND2_X1 i_257_76_8594 (.A1(n_257_76_18062), .A2(n_257_76_8579), .ZN(
      n_257_76_8580));
   NAND3_X1 i_257_76_8595 (.A1(n_257_76_8553), .A2(n_257_76_8564), .A3(
      n_257_76_8580), .ZN(n_257_76_8581));
   INV_X1 i_257_76_8596 (.A(n_257_76_8581), .ZN(n_257_76_8582));
   NAND3_X1 i_257_76_8597 (.A1(n_257_76_8226), .A2(n_257_76_8210), .A3(
      n_257_76_8159), .ZN(n_257_76_8583));
   NAND4_X1 i_257_76_8598 (.A1(n_257_76_8160), .A2(n_257_76_8161), .A3(
      n_257_76_8207), .A4(n_257_76_8213), .ZN(n_257_76_8584));
   NOR2_X1 i_257_76_8599 (.A1(n_257_76_8583), .A2(n_257_76_8584), .ZN(
      n_257_76_8585));
   NAND2_X1 i_257_76_8600 (.A1(n_257_76_8221), .A2(n_257_422), .ZN(n_257_76_8586));
   INV_X1 i_257_76_8601 (.A(n_257_76_8586), .ZN(n_257_76_8587));
   NAND4_X1 i_257_76_8602 (.A1(n_257_76_8217), .A2(n_257_76_8218), .A3(
      n_257_76_8587), .A4(n_257_324), .ZN(n_257_76_8588));
   INV_X1 i_257_76_8603 (.A(n_257_76_8588), .ZN(n_257_76_8589));
   NAND3_X1 i_257_76_8604 (.A1(n_257_76_8200), .A2(n_257_76_8589), .A3(
      n_257_76_8149), .ZN(n_257_76_8590));
   INV_X1 i_257_76_8605 (.A(n_257_76_8590), .ZN(n_257_76_8591));
   NAND3_X1 i_257_76_8606 (.A1(n_257_76_8585), .A2(n_257_76_8591), .A3(
      n_257_76_8330), .ZN(n_257_76_8592));
   NOR2_X1 i_257_76_8607 (.A1(n_257_76_8592), .A2(n_257_76_8575), .ZN(
      n_257_76_8593));
   NOR2_X1 i_257_76_8608 (.A1(n_257_76_8520), .A2(n_257_76_8532), .ZN(
      n_257_76_8594));
   NAND4_X1 i_257_76_8609 (.A1(n_257_76_8593), .A2(n_257_76_8594), .A3(
      n_257_76_8233), .A4(n_257_76_8130), .ZN(n_257_76_8595));
   NOR2_X1 i_257_76_8610 (.A1(n_257_76_8595), .A2(n_257_76_8535), .ZN(
      n_257_76_8596));
   NAND2_X1 i_257_76_8611 (.A1(n_257_342), .A2(n_257_76_8596), .ZN(n_257_76_8597));
   NAND4_X1 i_257_76_8612 (.A1(n_257_76_8204), .A2(n_257_76_8165), .A3(
      n_257_76_8440), .A4(n_257_76_8166), .ZN(n_257_76_8598));
   INV_X1 i_257_76_8613 (.A(n_257_76_8444), .ZN(n_257_76_8599));
   NAND3_X1 i_257_76_8614 (.A1(n_257_76_8599), .A2(n_257_76_8389), .A3(
      n_257_76_8571), .ZN(n_257_76_8600));
   NOR2_X1 i_257_76_8615 (.A1(n_257_76_8598), .A2(n_257_76_8600), .ZN(
      n_257_76_8601));
   INV_X1 i_257_76_8616 (.A(n_257_76_8526), .ZN(n_257_76_8602));
   INV_X1 i_257_76_8617 (.A(n_257_76_8421), .ZN(n_257_76_8603));
   NAND2_X1 i_257_76_8618 (.A1(n_257_420), .A2(n_257_667), .ZN(n_257_76_8604));
   NAND2_X1 i_257_76_8619 (.A1(n_257_76_8604), .A2(n_257_76_8214), .ZN(
      n_257_76_8605));
   INV_X1 i_257_76_8620 (.A(n_257_76_8605), .ZN(n_257_76_8606));
   NAND2_X1 i_257_76_8621 (.A1(n_257_428), .A2(n_257_579), .ZN(n_257_76_8607));
   NAND3_X1 i_257_76_8622 (.A1(n_257_484), .A2(n_257_402), .A3(n_257_442), 
      .ZN(n_257_76_8608));
   INV_X1 i_257_76_8623 (.A(n_257_76_8608), .ZN(n_257_76_8609));
   NAND2_X1 i_257_76_8624 (.A1(n_257_76_8607), .A2(n_257_76_8609), .ZN(
      n_257_76_8610));
   NOR2_X1 i_257_76_8625 (.A1(n_257_76_8610), .A2(n_257_1073), .ZN(n_257_76_8611));
   NAND4_X1 i_257_76_8626 (.A1(n_257_76_8606), .A2(n_257_76_8429), .A3(
      n_257_76_8611), .A4(n_257_76_8218), .ZN(n_257_76_8612));
   INV_X1 i_257_76_8627 (.A(n_257_76_8612), .ZN(n_257_76_8613));
   NAND3_X1 i_257_76_8628 (.A1(n_257_76_8602), .A2(n_257_76_8603), .A3(
      n_257_76_8613), .ZN(n_257_76_8614));
   INV_X1 i_257_76_8629 (.A(n_257_76_8614), .ZN(n_257_76_8615));
   NAND4_X1 i_257_76_8630 (.A1(n_257_76_8153), .A2(n_257_76_8154), .A3(
      n_257_76_8226), .A4(n_257_76_8210), .ZN(n_257_76_8616));
   INV_X1 i_257_76_8631 (.A(n_257_76_8616), .ZN(n_257_76_8617));
   NAND2_X1 i_257_76_8632 (.A1(n_257_76_8615), .A2(n_257_76_8617), .ZN(
      n_257_76_8618));
   NOR2_X1 i_257_76_8633 (.A1(n_257_76_8532), .A2(n_257_76_8618), .ZN(
      n_257_76_8619));
   NAND4_X1 i_257_76_8634 (.A1(n_257_76_8601), .A2(n_257_76_8233), .A3(
      n_257_76_8619), .A4(n_257_76_8130), .ZN(n_257_76_8620));
   NOR2_X1 i_257_76_8635 (.A1(n_257_76_8620), .A2(n_257_76_8535), .ZN(
      n_257_76_8621));
   NAND2_X1 i_257_76_8636 (.A1(n_257_76_18060), .A2(n_257_76_8621), .ZN(
      n_257_76_8622));
   INV_X1 i_257_76_8637 (.A(Small_Packet_Data_Size[14]), .ZN(n_257_76_8623));
   NAND2_X1 i_257_76_8638 (.A1(n_257_76_8607), .A2(n_257_76_18039), .ZN(
      n_257_76_8624));
   NOR2_X1 i_257_76_8639 (.A1(n_257_76_8624), .A2(n_257_1073), .ZN(n_257_76_8625));
   NAND3_X1 i_257_76_8640 (.A1(n_257_76_8625), .A2(n_257_76_8218), .A3(
      n_257_76_8604), .ZN(n_257_76_8626));
   NAND2_X1 i_257_76_8641 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[14]), 
      .ZN(n_257_76_8627));
   NAND2_X1 i_257_76_8642 (.A1(n_257_76_8626), .A2(n_257_76_8627), .ZN(
      n_257_76_8628));
   NAND2_X1 i_257_76_8643 (.A1(n_257_466), .A2(n_257_442), .ZN(n_257_76_8629));
   INV_X1 i_257_76_8644 (.A(n_257_76_8629), .ZN(n_257_76_8630));
   NAND2_X1 i_257_76_8645 (.A1(n_257_451), .A2(n_257_76_8630), .ZN(n_257_76_8631));
   NAND2_X1 i_257_76_8646 (.A1(n_257_843), .A2(n_257_442), .ZN(n_257_76_8632));
   INV_X1 i_257_76_8647 (.A(n_257_76_8632), .ZN(n_257_76_8633));
   NAND2_X1 i_257_76_8648 (.A1(n_257_446), .A2(n_257_76_8633), .ZN(n_257_76_8634));
   NAND3_X1 i_257_76_8649 (.A1(n_257_76_8628), .A2(n_257_76_8631), .A3(
      n_257_76_8634), .ZN(n_257_76_8635));
   INV_X1 i_257_76_8650 (.A(n_257_76_8635), .ZN(n_257_76_8636));
   NAND2_X1 i_257_76_8651 (.A1(n_257_913), .A2(n_257_76_17940), .ZN(
      n_257_76_8637));
   NAND2_X1 i_257_76_8652 (.A1(n_257_449), .A2(n_257_76_15863), .ZN(
      n_257_76_8638));
   INV_X1 i_257_76_8653 (.A(n_257_76_8467), .ZN(n_257_76_8639));
   NAND2_X1 i_257_76_8654 (.A1(n_257_447), .A2(n_257_76_8639), .ZN(n_257_76_8640));
   NAND4_X1 i_257_76_8655 (.A1(n_257_76_8637), .A2(n_257_76_8638), .A3(
      n_257_76_8640), .A4(n_257_76_8588), .ZN(n_257_76_8641));
   INV_X1 i_257_76_8656 (.A(n_257_76_8641), .ZN(n_257_76_8642));
   INV_X1 i_257_76_8657 (.A(n_257_76_8132), .ZN(n_257_76_8643));
   NAND2_X1 i_257_76_8658 (.A1(n_257_440), .A2(n_257_76_8643), .ZN(n_257_76_8644));
   NAND2_X1 i_257_76_8659 (.A1(n_257_715), .A2(n_257_76_15655), .ZN(
      n_257_76_8645));
   NAND2_X1 i_257_76_8660 (.A1(n_257_643), .A2(n_257_76_17928), .ZN(
      n_257_76_8646));
   NAND4_X1 i_257_76_8661 (.A1(n_257_76_8644), .A2(n_257_76_8645), .A3(
      n_257_76_8646), .A4(n_257_76_8325), .ZN(n_257_76_8647));
   NAND2_X1 i_257_76_8662 (.A1(n_257_49), .A2(n_257_76_17918), .ZN(n_257_76_8648));
   NAND3_X1 i_257_76_8663 (.A1(n_257_438), .A2(n_257_1079), .A3(n_257_442), 
      .ZN(n_257_76_8649));
   NAND3_X1 i_257_76_8664 (.A1(n_257_76_8544), .A2(n_257_76_8648), .A3(
      n_257_76_8649), .ZN(n_257_76_8650));
   NOR2_X1 i_257_76_8665 (.A1(n_257_76_8647), .A2(n_257_76_8650), .ZN(
      n_257_76_8651));
   NAND3_X1 i_257_76_8666 (.A1(n_257_76_8636), .A2(n_257_76_8642), .A3(
      n_257_76_8651), .ZN(n_257_76_8652));
   NAND2_X1 i_257_76_8667 (.A1(n_257_811), .A2(n_257_76_17952), .ZN(
      n_257_76_8653));
   NAND2_X1 i_257_76_8668 (.A1(n_257_875), .A2(n_257_76_17903), .ZN(
      n_257_76_8654));
   NAND2_X1 i_257_76_8669 (.A1(n_257_977), .A2(n_257_442), .ZN(n_257_76_8655));
   INV_X1 i_257_76_8670 (.A(n_257_76_8655), .ZN(n_257_76_8656));
   NAND2_X1 i_257_76_8671 (.A1(n_257_441), .A2(n_257_76_8656), .ZN(n_257_76_8657));
   NAND2_X1 i_257_76_8672 (.A1(n_257_127), .A2(n_257_76_17925), .ZN(
      n_257_76_8658));
   NAND4_X1 i_257_76_8673 (.A1(n_257_76_8653), .A2(n_257_76_8654), .A3(
      n_257_76_8657), .A4(n_257_76_8658), .ZN(n_257_76_8659));
   NOR2_X1 i_257_76_8674 (.A1(n_257_76_8652), .A2(n_257_76_8659), .ZN(
      n_257_76_8660));
   NAND2_X1 i_257_76_8675 (.A1(n_257_89), .A2(n_257_76_17932), .ZN(n_257_76_8661));
   NAND2_X1 i_257_76_8676 (.A1(n_257_747), .A2(n_257_76_17935), .ZN(
      n_257_76_8662));
   NAND3_X1 i_257_76_8677 (.A1(n_257_76_8300), .A2(n_257_76_8661), .A3(
      n_257_76_8662), .ZN(n_257_76_8663));
   INV_X1 i_257_76_8678 (.A(n_257_76_8663), .ZN(n_257_76_8664));
   NAND2_X1 i_257_76_8679 (.A1(n_257_1009), .A2(n_257_76_17964), .ZN(
      n_257_76_8665));
   NAND4_X1 i_257_76_8680 (.A1(n_257_76_8660), .A2(n_257_76_8664), .A3(
      n_257_76_8665), .A4(n_257_76_8531), .ZN(n_257_76_8666));
   INV_X1 i_257_76_8681 (.A(n_257_76_8666), .ZN(n_257_76_8667));
   NAND2_X1 i_257_76_8682 (.A1(n_257_683), .A2(n_257_76_17958), .ZN(
      n_257_76_8668));
   NAND2_X1 i_257_76_8683 (.A1(n_257_166), .A2(n_257_76_17331), .ZN(
      n_257_76_8669));
   NAND3_X1 i_257_76_8684 (.A1(n_257_76_8230), .A2(n_257_76_8668), .A3(
      n_257_76_8669), .ZN(n_257_76_8670));
   INV_X1 i_257_76_8685 (.A(n_257_76_8670), .ZN(n_257_76_8671));
   NAND2_X1 i_257_76_8686 (.A1(n_257_1041), .A2(n_257_76_17969), .ZN(
      n_257_76_8672));
   NAND4_X1 i_257_76_8687 (.A1(n_257_76_8667), .A2(n_257_76_8671), .A3(
      n_257_76_8511), .A4(n_257_76_8672), .ZN(n_257_76_8673));
   NAND3_X1 i_257_76_8688 (.A1(n_257_76_8597), .A2(n_257_76_8622), .A3(
      n_257_76_8673), .ZN(n_257_76_8674));
   INV_X1 i_257_76_8689 (.A(n_257_76_8674), .ZN(n_257_76_8675));
   NAND3_X1 i_257_76_8690 (.A1(n_257_76_8539), .A2(n_257_76_8582), .A3(
      n_257_76_8675), .ZN(n_257_76_8676));
   NOR2_X1 i_257_76_8691 (.A1(n_257_76_8487), .A2(n_257_76_8676), .ZN(
      n_257_76_8677));
   NAND2_X1 i_257_76_8692 (.A1(n_257_76_8360), .A2(n_257_76_8677), .ZN(n_14));
   NAND2_X1 i_257_76_8693 (.A1(n_257_1010), .A2(n_257_444), .ZN(n_257_76_8678));
   NAND2_X1 i_257_76_8694 (.A1(n_257_441), .A2(n_257_978), .ZN(n_257_76_8679));
   INV_X1 i_257_76_8695 (.A(n_257_1074), .ZN(n_257_76_8680));
   NAND2_X1 i_257_76_8696 (.A1(n_257_946), .A2(n_257_442), .ZN(n_257_76_8681));
   INV_X1 i_257_76_8697 (.A(n_257_76_8681), .ZN(n_257_76_8682));
   NAND3_X1 i_257_76_8698 (.A1(n_257_440), .A2(n_257_76_8680), .A3(n_257_76_8682), 
      .ZN(n_257_76_8683));
   INV_X1 i_257_76_8699 (.A(n_257_76_8683), .ZN(n_257_76_8684));
   NAND2_X1 i_257_76_8700 (.A1(n_257_76_8679), .A2(n_257_76_8684), .ZN(
      n_257_76_8685));
   INV_X1 i_257_76_8701 (.A(n_257_76_8685), .ZN(n_257_76_8686));
   NAND2_X1 i_257_76_8702 (.A1(n_257_76_8678), .A2(n_257_76_8686), .ZN(
      n_257_76_8687));
   INV_X1 i_257_76_8703 (.A(n_257_76_8687), .ZN(n_257_76_8688));
   NAND2_X1 i_257_76_8704 (.A1(n_257_1042), .A2(n_257_443), .ZN(n_257_76_8689));
   NAND2_X1 i_257_76_8705 (.A1(n_257_76_8688), .A2(n_257_76_8689), .ZN(
      n_257_76_8690));
   INV_X1 i_257_76_8706 (.A(n_257_76_8690), .ZN(n_257_76_8691));
   NAND2_X1 i_257_76_8707 (.A1(n_257_17), .A2(n_257_76_8691), .ZN(n_257_76_8692));
   NOR2_X1 i_257_76_8708 (.A1(n_257_1074), .A2(n_257_76_17412), .ZN(
      n_257_76_8693));
   INV_X1 i_257_76_8709 (.A(n_257_76_8693), .ZN(n_257_76_8694));
   NOR2_X1 i_257_76_8710 (.A1(n_257_76_8694), .A2(n_257_76_15197), .ZN(
      n_257_76_8695));
   NAND2_X1 i_257_76_8711 (.A1(n_257_1042), .A2(n_257_76_8695), .ZN(
      n_257_76_8696));
   INV_X1 i_257_76_8712 (.A(n_257_76_8696), .ZN(n_257_76_8697));
   NAND2_X1 i_257_76_8713 (.A1(n_257_76_18072), .A2(n_257_76_8697), .ZN(
      n_257_76_8698));
   NAND2_X1 i_257_76_8714 (.A1(n_257_440), .A2(n_257_946), .ZN(n_257_76_8699));
   NAND2_X1 i_257_76_8715 (.A1(n_257_76_8699), .A2(n_257_644), .ZN(n_257_76_8700));
   INV_X1 i_257_76_8716 (.A(n_257_76_8700), .ZN(n_257_76_8701));
   NAND2_X1 i_257_76_8717 (.A1(n_257_447), .A2(n_257_780), .ZN(n_257_76_8702));
   NAND2_X1 i_257_76_8718 (.A1(n_257_1080), .A2(n_257_438), .ZN(n_257_76_8703));
   NOR2_X1 i_257_76_8719 (.A1(n_257_1074), .A2(n_257_76_17927), .ZN(
      n_257_76_8704));
   NAND4_X1 i_257_76_8720 (.A1(n_257_76_8701), .A2(n_257_76_8702), .A3(
      n_257_76_8703), .A4(n_257_76_8704), .ZN(n_257_76_8705));
   NAND2_X1 i_257_76_8721 (.A1(n_257_716), .A2(n_257_435), .ZN(n_257_76_8706));
   NAND2_X1 i_257_76_8722 (.A1(n_257_446), .A2(n_257_844), .ZN(n_257_76_8707));
   NAND2_X1 i_257_76_8723 (.A1(n_257_449), .A2(n_257_1088), .ZN(n_257_76_8708));
   NAND3_X1 i_257_76_8724 (.A1(n_257_76_8706), .A2(n_257_76_8707), .A3(
      n_257_76_8708), .ZN(n_257_76_8709));
   NOR2_X1 i_257_76_8725 (.A1(n_257_76_8705), .A2(n_257_76_8709), .ZN(
      n_257_76_8710));
   NAND2_X1 i_257_76_8726 (.A1(n_257_914), .A2(n_257_439), .ZN(n_257_76_8711));
   NAND2_X1 i_257_76_8727 (.A1(n_257_76_8711), .A2(n_257_76_8679), .ZN(
      n_257_76_8712));
   INV_X1 i_257_76_8728 (.A(n_257_76_8712), .ZN(n_257_76_8713));
   NAND2_X1 i_257_76_8729 (.A1(n_257_876), .A2(n_257_445), .ZN(n_257_76_8714));
   NAND3_X1 i_257_76_8730 (.A1(n_257_76_8710), .A2(n_257_76_8713), .A3(
      n_257_76_8714), .ZN(n_257_76_8715));
   NAND2_X1 i_257_76_8731 (.A1(n_257_748), .A2(n_257_436), .ZN(n_257_76_8716));
   NAND2_X1 i_257_76_8732 (.A1(n_257_812), .A2(n_257_437), .ZN(n_257_76_8717));
   NAND2_X1 i_257_76_8733 (.A1(n_257_76_8716), .A2(n_257_76_8717), .ZN(
      n_257_76_8718));
   NOR2_X1 i_257_76_8734 (.A1(n_257_76_8715), .A2(n_257_76_8718), .ZN(
      n_257_76_8719));
   NAND2_X1 i_257_76_8735 (.A1(n_257_684), .A2(n_257_448), .ZN(n_257_76_8720));
   NAND3_X1 i_257_76_8736 (.A1(n_257_76_8719), .A2(n_257_76_8720), .A3(
      n_257_76_8678), .ZN(n_257_76_8721));
   INV_X1 i_257_76_8737 (.A(n_257_76_8689), .ZN(n_257_76_8722));
   NOR2_X1 i_257_76_8738 (.A1(n_257_76_8721), .A2(n_257_76_8722), .ZN(
      n_257_76_8723));
   NAND2_X1 i_257_76_8739 (.A1(n_257_28), .A2(n_257_76_8723), .ZN(n_257_76_8724));
   NAND3_X1 i_257_76_8740 (.A1(n_257_76_8692), .A2(n_257_76_8698), .A3(
      n_257_76_8724), .ZN(n_257_76_8725));
   NAND3_X1 i_257_76_8741 (.A1(n_257_76_8693), .A2(n_257_76_8699), .A3(n_257_844), 
      .ZN(n_257_76_8726));
   NAND2_X1 i_257_76_8742 (.A1(n_257_76_8703), .A2(n_257_446), .ZN(n_257_76_8727));
   NOR2_X1 i_257_76_8743 (.A1(n_257_76_8726), .A2(n_257_76_8727), .ZN(
      n_257_76_8728));
   NAND3_X1 i_257_76_8744 (.A1(n_257_76_8728), .A2(n_257_76_8711), .A3(
      n_257_76_8679), .ZN(n_257_76_8729));
   INV_X1 i_257_76_8745 (.A(n_257_76_8714), .ZN(n_257_76_8730));
   NOR2_X1 i_257_76_8746 (.A1(n_257_76_8729), .A2(n_257_76_8730), .ZN(
      n_257_76_8731));
   NAND2_X1 i_257_76_8747 (.A1(n_257_76_8678), .A2(n_257_76_8731), .ZN(
      n_257_76_8732));
   INV_X1 i_257_76_8748 (.A(n_257_76_8732), .ZN(n_257_76_8733));
   NAND2_X1 i_257_76_8749 (.A1(n_257_76_8733), .A2(n_257_76_8689), .ZN(
      n_257_76_8734));
   INV_X1 i_257_76_8750 (.A(n_257_76_8734), .ZN(n_257_76_8735));
   NAND2_X1 i_257_76_8751 (.A1(n_257_76_18070), .A2(n_257_76_8735), .ZN(
      n_257_76_8736));
   NAND3_X1 i_257_76_8752 (.A1(n_257_76_8693), .A2(n_257_76_8699), .A3(n_257_439), 
      .ZN(n_257_76_8737));
   INV_X1 i_257_76_8753 (.A(n_257_76_8737), .ZN(n_257_76_8738));
   NAND3_X1 i_257_76_8754 (.A1(n_257_76_8679), .A2(n_257_914), .A3(n_257_76_8738), 
      .ZN(n_257_76_8739));
   INV_X1 i_257_76_8755 (.A(n_257_76_8739), .ZN(n_257_76_8740));
   NAND2_X1 i_257_76_8756 (.A1(n_257_76_8678), .A2(n_257_76_8740), .ZN(
      n_257_76_8741));
   INV_X1 i_257_76_8757 (.A(n_257_76_8741), .ZN(n_257_76_8742));
   NAND2_X1 i_257_76_8758 (.A1(n_257_76_8742), .A2(n_257_76_8689), .ZN(
      n_257_76_8743));
   INV_X1 i_257_76_8759 (.A(n_257_76_8743), .ZN(n_257_76_8744));
   NAND2_X1 i_257_76_8760 (.A1(n_257_76_18084), .A2(n_257_76_8744), .ZN(
      n_257_76_8745));
   NAND2_X1 i_257_76_8761 (.A1(n_257_128), .A2(n_257_430), .ZN(n_257_76_8746));
   NAND2_X1 i_257_76_8762 (.A1(n_257_76_8746), .A2(n_257_76_8711), .ZN(
      n_257_76_8747));
   INV_X1 i_257_76_8763 (.A(n_257_76_8747), .ZN(n_257_76_8748));
   NAND3_X1 i_257_76_8764 (.A1(n_257_76_8707), .A2(n_257_76_8708), .A3(
      n_257_76_8702), .ZN(n_257_76_8749));
   INV_X1 i_257_76_8765 (.A(n_257_76_8679), .ZN(n_257_76_8750));
   NOR2_X1 i_257_76_8766 (.A1(n_257_76_8749), .A2(n_257_76_8750), .ZN(
      n_257_76_8751));
   NAND2_X1 i_257_76_8767 (.A1(n_257_451), .A2(n_257_467), .ZN(n_257_76_8752));
   NAND4_X1 i_257_76_8768 (.A1(n_257_76_8748), .A2(n_257_76_8751), .A3(
      n_257_76_8714), .A4(n_257_76_8752), .ZN(n_257_76_8753));
   NAND2_X1 i_257_76_8769 (.A1(n_257_90), .A2(n_257_431), .ZN(n_257_76_8754));
   NAND3_X1 i_257_76_8770 (.A1(n_257_76_8754), .A2(n_257_76_8716), .A3(
      n_257_76_8717), .ZN(n_257_76_8755));
   NOR2_X1 i_257_76_8771 (.A1(n_257_76_8753), .A2(n_257_76_8755), .ZN(
      n_257_76_8756));
   NAND2_X1 i_257_76_8772 (.A1(n_257_247), .A2(n_257_425), .ZN(n_257_76_8757));
   NAND2_X1 i_257_76_8773 (.A1(n_257_167), .A2(n_257_429), .ZN(n_257_76_8758));
   NAND2_X1 i_257_76_8774 (.A1(n_257_644), .A2(n_257_450), .ZN(n_257_76_8759));
   NAND3_X1 i_257_76_8775 (.A1(n_257_76_8759), .A2(n_257_76_8703), .A3(
      n_257_76_8699), .ZN(n_257_76_8760));
   INV_X1 i_257_76_8776 (.A(n_257_580), .ZN(n_257_76_8761));
   NAND2_X1 i_257_76_8777 (.A1(n_257_76_8761), .A2(n_257_442), .ZN(n_257_76_8762));
   OAI21_X1 i_257_76_8778 (.A(n_257_76_8762), .B1(n_257_428), .B2(n_257_76_17412), 
      .ZN(n_257_76_8763));
   INV_X1 i_257_76_8779 (.A(n_257_76_8763), .ZN(n_257_76_8764));
   NOR2_X1 i_257_76_8780 (.A1(n_257_1074), .A2(n_257_76_8764), .ZN(n_257_76_8765));
   NAND2_X1 i_257_76_8781 (.A1(n_257_516), .A2(n_257_424), .ZN(n_257_76_8766));
   NAND2_X1 i_257_76_8782 (.A1(n_257_432), .A2(n_257_612), .ZN(n_257_76_8767));
   NAND2_X1 i_257_76_8783 (.A1(n_257_76_8767), .A2(n_257_423), .ZN(n_257_76_8768));
   INV_X1 i_257_76_8784 (.A(n_257_76_8768), .ZN(n_257_76_8769));
   NAND3_X1 i_257_76_8785 (.A1(n_257_76_8765), .A2(n_257_76_8766), .A3(
      n_257_76_8769), .ZN(n_257_76_8770));
   NOR2_X1 i_257_76_8786 (.A1(n_257_76_8760), .A2(n_257_76_8770), .ZN(
      n_257_76_8771));
   NAND2_X1 i_257_76_8787 (.A1(n_257_50), .A2(n_257_433), .ZN(n_257_76_8772));
   NAND2_X1 i_257_76_8788 (.A1(n_257_548), .A2(n_257_426), .ZN(n_257_76_8773));
   NAND2_X1 i_257_76_8789 (.A1(n_257_76_8772), .A2(n_257_76_8773), .ZN(
      n_257_76_8774));
   INV_X1 i_257_76_8790 (.A(n_257_76_8774), .ZN(n_257_76_8775));
   NAND2_X1 i_257_76_8791 (.A1(n_257_207), .A2(n_257_427), .ZN(n_257_76_8776));
   NAND3_X1 i_257_76_8792 (.A1(n_257_287), .A2(n_257_76_8706), .A3(n_257_76_8776), 
      .ZN(n_257_76_8777));
   INV_X1 i_257_76_8793 (.A(n_257_76_8777), .ZN(n_257_76_8778));
   NAND3_X1 i_257_76_8794 (.A1(n_257_76_8771), .A2(n_257_76_8775), .A3(
      n_257_76_8778), .ZN(n_257_76_8779));
   INV_X1 i_257_76_8795 (.A(n_257_76_8779), .ZN(n_257_76_8780));
   NAND3_X1 i_257_76_8796 (.A1(n_257_76_8757), .A2(n_257_76_8758), .A3(
      n_257_76_8780), .ZN(n_257_76_8781));
   INV_X1 i_257_76_8797 (.A(n_257_76_8781), .ZN(n_257_76_8782));
   NAND4_X1 i_257_76_8798 (.A1(n_257_76_8756), .A2(n_257_76_8720), .A3(
      n_257_76_8678), .A4(n_257_76_8782), .ZN(n_257_76_8783));
   NOR2_X1 i_257_76_8799 (.A1(n_257_76_8783), .A2(n_257_76_8722), .ZN(
      n_257_76_8784));
   NAND2_X1 i_257_76_8800 (.A1(n_257_76_18066), .A2(n_257_76_8784), .ZN(
      n_257_76_8785));
   NAND3_X1 i_257_76_8801 (.A1(n_257_76_8736), .A2(n_257_76_8745), .A3(
      n_257_76_8785), .ZN(n_257_76_8786));
   NOR2_X1 i_257_76_8802 (.A1(n_257_76_8725), .A2(n_257_76_8786), .ZN(
      n_257_76_8787));
   NAND2_X1 i_257_76_8803 (.A1(n_257_76_8693), .A2(n_257_978), .ZN(n_257_76_8788));
   NOR2_X1 i_257_76_8804 (.A1(n_257_76_13147), .A2(n_257_76_8788), .ZN(
      n_257_76_8789));
   NAND2_X1 i_257_76_8805 (.A1(n_257_76_8678), .A2(n_257_76_8789), .ZN(
      n_257_76_8790));
   INV_X1 i_257_76_8806 (.A(n_257_76_8790), .ZN(n_257_76_8791));
   NAND2_X1 i_257_76_8807 (.A1(n_257_76_8791), .A2(n_257_76_8689), .ZN(
      n_257_76_8792));
   INV_X1 i_257_76_8808 (.A(n_257_76_8792), .ZN(n_257_76_8793));
   NAND2_X1 i_257_76_8809 (.A1(n_257_76_18071), .A2(n_257_76_8793), .ZN(
      n_257_76_8794));
   NOR2_X1 i_257_76_8810 (.A1(n_257_1074), .A2(n_257_76_15289), .ZN(
      n_257_76_8795));
   NAND4_X1 i_257_76_8811 (.A1(n_257_76_8703), .A2(n_257_716), .A3(n_257_76_8795), 
      .A4(n_257_76_8699), .ZN(n_257_76_8796));
   NAND2_X1 i_257_76_8812 (.A1(n_257_76_8707), .A2(n_257_76_8702), .ZN(
      n_257_76_8797));
   NOR2_X1 i_257_76_8813 (.A1(n_257_76_8796), .A2(n_257_76_8797), .ZN(
      n_257_76_8798));
   NAND3_X1 i_257_76_8814 (.A1(n_257_76_8798), .A2(n_257_76_8713), .A3(
      n_257_76_8714), .ZN(n_257_76_8799));
   NOR2_X1 i_257_76_8815 (.A1(n_257_76_8799), .A2(n_257_76_8718), .ZN(
      n_257_76_8800));
   NAND2_X1 i_257_76_8816 (.A1(n_257_76_8678), .A2(n_257_76_8800), .ZN(
      n_257_76_8801));
   INV_X1 i_257_76_8817 (.A(n_257_76_8801), .ZN(n_257_76_8802));
   NAND2_X1 i_257_76_8818 (.A1(n_257_76_8802), .A2(n_257_76_8689), .ZN(
      n_257_76_8803));
   INV_X1 i_257_76_8819 (.A(n_257_76_8803), .ZN(n_257_76_8804));
   NAND2_X1 i_257_76_8820 (.A1(n_257_76_18078), .A2(n_257_76_8804), .ZN(
      n_257_76_8805));
   NAND2_X1 i_257_76_8821 (.A1(n_257_442), .A2(n_257_580), .ZN(n_257_76_8806));
   INV_X1 i_257_76_8822 (.A(n_257_76_8806), .ZN(n_257_76_8807));
   NAND2_X1 i_257_76_8823 (.A1(n_257_428), .A2(n_257_76_8807), .ZN(n_257_76_8808));
   INV_X1 i_257_76_8824 (.A(n_257_76_8808), .ZN(n_257_76_8809));
   NAND2_X1 i_257_76_8825 (.A1(n_257_76_8809), .A2(n_257_76_8767), .ZN(
      n_257_76_8810));
   NOR2_X1 i_257_76_8826 (.A1(n_257_76_8810), .A2(n_257_1074), .ZN(n_257_76_8811));
   NAND4_X1 i_257_76_8827 (.A1(n_257_76_8811), .A2(n_257_76_8759), .A3(
      n_257_76_8703), .A4(n_257_76_8699), .ZN(n_257_76_8812));
   NAND2_X1 i_257_76_8828 (.A1(n_257_76_8708), .A2(n_257_76_8702), .ZN(
      n_257_76_8813));
   NOR2_X1 i_257_76_8829 (.A1(n_257_76_8812), .A2(n_257_76_8813), .ZN(
      n_257_76_8814));
   NAND3_X1 i_257_76_8830 (.A1(n_257_76_8772), .A2(n_257_76_8706), .A3(
      n_257_76_8707), .ZN(n_257_76_8815));
   INV_X1 i_257_76_8831 (.A(n_257_76_8815), .ZN(n_257_76_8816));
   NAND4_X1 i_257_76_8832 (.A1(n_257_76_8814), .A2(n_257_76_8713), .A3(
      n_257_76_8746), .A4(n_257_76_8816), .ZN(n_257_76_8817));
   NAND3_X1 i_257_76_8833 (.A1(n_257_76_8717), .A2(n_257_76_8714), .A3(
      n_257_76_8752), .ZN(n_257_76_8818));
   NOR2_X1 i_257_76_8834 (.A1(n_257_76_8817), .A2(n_257_76_8818), .ZN(
      n_257_76_8819));
   INV_X1 i_257_76_8835 (.A(n_257_76_8758), .ZN(n_257_76_8820));
   NAND2_X1 i_257_76_8836 (.A1(n_257_76_8754), .A2(n_257_76_8716), .ZN(
      n_257_76_8821));
   NOR2_X1 i_257_76_8837 (.A1(n_257_76_8820), .A2(n_257_76_8821), .ZN(
      n_257_76_8822));
   NAND4_X1 i_257_76_8838 (.A1(n_257_76_8720), .A2(n_257_76_8678), .A3(
      n_257_76_8819), .A4(n_257_76_8822), .ZN(n_257_76_8823));
   NOR2_X1 i_257_76_8839 (.A1(n_257_76_8823), .A2(n_257_76_8722), .ZN(
      n_257_76_8824));
   NAND2_X1 i_257_76_8840 (.A1(n_257_76_18074), .A2(n_257_76_8824), .ZN(
      n_257_76_8825));
   NAND3_X1 i_257_76_8841 (.A1(n_257_76_8794), .A2(n_257_76_8805), .A3(
      n_257_76_8825), .ZN(n_257_76_8826));
   NAND2_X1 i_257_76_8842 (.A1(n_257_1074), .A2(n_257_442), .ZN(n_257_76_8827));
   INV_X1 i_257_76_8843 (.A(n_257_76_8827), .ZN(n_257_76_8828));
   NAND2_X1 i_257_76_8844 (.A1(n_257_13), .A2(n_257_76_8828), .ZN(n_257_76_8829));
   NOR2_X1 i_257_76_8845 (.A1(n_257_76_17902), .A2(n_257_1074), .ZN(
      n_257_76_8830));
   NAND3_X1 i_257_76_8846 (.A1(n_257_76_8703), .A2(n_257_76_8830), .A3(
      n_257_76_8699), .ZN(n_257_76_8831));
   INV_X1 i_257_76_8847 (.A(n_257_76_8831), .ZN(n_257_76_8832));
   NAND4_X1 i_257_76_8848 (.A1(n_257_876), .A2(n_257_76_8711), .A3(n_257_76_8832), 
      .A4(n_257_76_8679), .ZN(n_257_76_8833));
   INV_X1 i_257_76_8849 (.A(n_257_76_8833), .ZN(n_257_76_8834));
   NAND2_X1 i_257_76_8850 (.A1(n_257_76_8678), .A2(n_257_76_8834), .ZN(
      n_257_76_8835));
   INV_X1 i_257_76_8851 (.A(n_257_76_8835), .ZN(n_257_76_8836));
   NAND2_X1 i_257_76_8852 (.A1(n_257_76_8836), .A2(n_257_76_8689), .ZN(
      n_257_76_8837));
   INV_X1 i_257_76_8853 (.A(n_257_76_8837), .ZN(n_257_76_8838));
   NAND2_X1 i_257_76_8854 (.A1(n_257_76_18077), .A2(n_257_76_8838), .ZN(
      n_257_76_8839));
   NAND2_X1 i_257_76_8855 (.A1(n_257_76_8829), .A2(n_257_76_8839), .ZN(
      n_257_76_8840));
   NOR2_X1 i_257_76_8856 (.A1(n_257_76_8826), .A2(n_257_76_8840), .ZN(
      n_257_76_8841));
   NAND4_X1 i_257_76_8857 (.A1(n_257_76_8751), .A2(n_257_76_8752), .A3(
      n_257_76_8746), .A4(n_257_76_8711), .ZN(n_257_76_8842));
   NAND3_X1 i_257_76_8858 (.A1(n_257_76_8716), .A2(n_257_76_8717), .A3(
      n_257_76_8714), .ZN(n_257_76_8843));
   NOR2_X1 i_257_76_8859 (.A1(n_257_76_8842), .A2(n_257_76_8843), .ZN(
      n_257_76_8844));
   NAND2_X1 i_257_76_8860 (.A1(n_257_76_8767), .A2(n_257_426), .ZN(n_257_76_8845));
   INV_X1 i_257_76_8861 (.A(n_257_76_8845), .ZN(n_257_76_8846));
   NAND4_X1 i_257_76_8862 (.A1(n_257_76_8703), .A2(n_257_76_8765), .A3(
      n_257_76_8699), .A4(n_257_76_8846), .ZN(n_257_76_8847));
   INV_X1 i_257_76_8863 (.A(n_257_76_8847), .ZN(n_257_76_8848));
   NAND3_X1 i_257_76_8864 (.A1(n_257_548), .A2(n_257_76_8776), .A3(n_257_76_8759), 
      .ZN(n_257_76_8849));
   INV_X1 i_257_76_8865 (.A(n_257_76_8849), .ZN(n_257_76_8850));
   NAND4_X1 i_257_76_8866 (.A1(n_257_76_8848), .A2(n_257_76_8850), .A3(
      n_257_76_8772), .A4(n_257_76_8706), .ZN(n_257_76_8851));
   INV_X1 i_257_76_8867 (.A(n_257_76_8851), .ZN(n_257_76_8852));
   NAND3_X1 i_257_76_8868 (.A1(n_257_76_8758), .A2(n_257_76_8852), .A3(
      n_257_76_8754), .ZN(n_257_76_8853));
   INV_X1 i_257_76_8869 (.A(n_257_76_8853), .ZN(n_257_76_8854));
   NAND4_X1 i_257_76_8870 (.A1(n_257_76_8844), .A2(n_257_76_8720), .A3(
      n_257_76_8678), .A4(n_257_76_8854), .ZN(n_257_76_8855));
   NOR2_X1 i_257_76_8871 (.A1(n_257_76_8855), .A2(n_257_76_8722), .ZN(
      n_257_76_8856));
   NAND2_X1 i_257_76_8872 (.A1(n_257_76_18076), .A2(n_257_76_8856), .ZN(
      n_257_76_8857));
   NAND2_X1 i_257_76_8873 (.A1(n_257_76_8679), .A2(n_257_76_8707), .ZN(
      n_257_76_8858));
   INV_X1 i_257_76_8874 (.A(n_257_76_8858), .ZN(n_257_76_8859));
   NOR2_X1 i_257_76_8875 (.A1(n_257_1074), .A2(n_257_76_17934), .ZN(
      n_257_76_8860));
   NAND3_X1 i_257_76_8876 (.A1(n_257_76_8703), .A2(n_257_76_8699), .A3(
      n_257_76_8860), .ZN(n_257_76_8861));
   INV_X1 i_257_76_8877 (.A(n_257_76_8702), .ZN(n_257_76_8862));
   NOR2_X1 i_257_76_8878 (.A1(n_257_76_8861), .A2(n_257_76_8862), .ZN(
      n_257_76_8863));
   NAND4_X1 i_257_76_8879 (.A1(n_257_76_8859), .A2(n_257_748), .A3(n_257_76_8863), 
      .A4(n_257_76_8711), .ZN(n_257_76_8864));
   NAND2_X1 i_257_76_8880 (.A1(n_257_76_8717), .A2(n_257_76_8714), .ZN(
      n_257_76_8865));
   NOR2_X1 i_257_76_8881 (.A1(n_257_76_8864), .A2(n_257_76_8865), .ZN(
      n_257_76_8866));
   NAND2_X1 i_257_76_8882 (.A1(n_257_76_8678), .A2(n_257_76_8866), .ZN(
      n_257_76_8867));
   INV_X1 i_257_76_8883 (.A(n_257_76_8867), .ZN(n_257_76_8868));
   NAND2_X1 i_257_76_8884 (.A1(n_257_76_8868), .A2(n_257_76_8689), .ZN(
      n_257_76_8869));
   INV_X1 i_257_76_8885 (.A(n_257_76_8869), .ZN(n_257_76_8870));
   NAND2_X1 i_257_76_8886 (.A1(n_257_76_18069), .A2(n_257_76_8870), .ZN(
      n_257_76_8871));
   NAND2_X1 i_257_76_8887 (.A1(n_257_612), .A2(n_257_442), .ZN(n_257_76_8872));
   INV_X1 i_257_76_8888 (.A(n_257_76_8872), .ZN(n_257_76_8873));
   NAND2_X1 i_257_76_8889 (.A1(n_257_432), .A2(n_257_76_8873), .ZN(n_257_76_8874));
   NOR2_X1 i_257_76_8890 (.A1(n_257_1074), .A2(n_257_76_8874), .ZN(n_257_76_8875));
   NAND4_X1 i_257_76_8891 (.A1(n_257_76_8759), .A2(n_257_76_8703), .A3(
      n_257_76_8699), .A4(n_257_76_8875), .ZN(n_257_76_8876));
   NOR2_X1 i_257_76_8892 (.A1(n_257_76_8876), .A2(n_257_76_8813), .ZN(
      n_257_76_8877));
   NAND4_X1 i_257_76_8893 (.A1(n_257_76_8877), .A2(n_257_76_8713), .A3(
      n_257_76_8752), .A4(n_257_76_8816), .ZN(n_257_76_8878));
   NOR2_X1 i_257_76_8894 (.A1(n_257_76_8878), .A2(n_257_76_8843), .ZN(
      n_257_76_8879));
   NAND3_X1 i_257_76_8895 (.A1(n_257_76_8720), .A2(n_257_76_8879), .A3(
      n_257_76_8678), .ZN(n_257_76_8880));
   NOR2_X1 i_257_76_8896 (.A1(n_257_76_8880), .A2(n_257_76_8722), .ZN(
      n_257_76_8881));
   NAND2_X1 i_257_76_8897 (.A1(n_257_68), .A2(n_257_76_8881), .ZN(n_257_76_8882));
   NAND3_X1 i_257_76_8898 (.A1(n_257_76_8857), .A2(n_257_76_8871), .A3(
      n_257_76_8882), .ZN(n_257_76_8883));
   NOR2_X1 i_257_76_8899 (.A1(n_257_1074), .A2(n_257_76_17951), .ZN(
      n_257_76_8884));
   NAND3_X1 i_257_76_8900 (.A1(n_257_76_8703), .A2(n_257_76_8699), .A3(
      n_257_76_8884), .ZN(n_257_76_8885));
   INV_X1 i_257_76_8901 (.A(n_257_76_8707), .ZN(n_257_76_8886));
   NOR2_X1 i_257_76_8902 (.A1(n_257_76_8885), .A2(n_257_76_8886), .ZN(
      n_257_76_8887));
   NAND4_X1 i_257_76_8903 (.A1(n_257_76_8713), .A2(n_257_76_8714), .A3(n_257_812), 
      .A4(n_257_76_8887), .ZN(n_257_76_8888));
   INV_X1 i_257_76_8904 (.A(n_257_76_8888), .ZN(n_257_76_8889));
   NAND2_X1 i_257_76_8905 (.A1(n_257_76_8678), .A2(n_257_76_8889), .ZN(
      n_257_76_8890));
   INV_X1 i_257_76_8906 (.A(n_257_76_8890), .ZN(n_257_76_8891));
   NAND2_X1 i_257_76_8907 (.A1(n_257_76_8891), .A2(n_257_76_8689), .ZN(
      n_257_76_8892));
   INV_X1 i_257_76_8908 (.A(n_257_76_8892), .ZN(n_257_76_8893));
   NAND2_X1 i_257_76_8909 (.A1(n_257_22), .A2(n_257_76_8893), .ZN(n_257_76_8894));
   NAND2_X1 i_257_76_8910 (.A1(n_257_444), .A2(n_257_76_8693), .ZN(n_257_76_8895));
   INV_X1 i_257_76_8911 (.A(n_257_76_8895), .ZN(n_257_76_8896));
   NAND2_X1 i_257_76_8912 (.A1(n_257_1010), .A2(n_257_76_8896), .ZN(
      n_257_76_8897));
   INV_X1 i_257_76_8913 (.A(n_257_76_8897), .ZN(n_257_76_8898));
   NAND2_X1 i_257_76_8914 (.A1(n_257_76_8689), .A2(n_257_76_8898), .ZN(
      n_257_76_8899));
   INV_X1 i_257_76_8915 (.A(n_257_76_8899), .ZN(n_257_76_8900));
   NAND2_X1 i_257_76_8916 (.A1(n_257_76_18075), .A2(n_257_76_8900), .ZN(
      n_257_76_8901));
   NAND2_X1 i_257_76_8917 (.A1(n_257_76_8894), .A2(n_257_76_8901), .ZN(
      n_257_76_8902));
   NOR2_X1 i_257_76_8918 (.A1(n_257_76_8883), .A2(n_257_76_8902), .ZN(
      n_257_76_8903));
   NAND3_X1 i_257_76_8919 (.A1(n_257_76_8787), .A2(n_257_76_8841), .A3(
      n_257_76_8903), .ZN(n_257_76_8904));
   INV_X1 i_257_76_8920 (.A(n_257_76_8904), .ZN(n_257_76_8905));
   NOR2_X1 i_257_76_8921 (.A1(n_257_76_8709), .A2(n_257_76_8750), .ZN(
      n_257_76_8906));
   NOR2_X1 i_257_76_8922 (.A1(n_257_1074), .A2(n_257_76_17633), .ZN(
      n_257_76_8907));
   NAND4_X1 i_257_76_8923 (.A1(n_257_76_8759), .A2(n_257_76_8703), .A3(
      n_257_76_8699), .A4(n_257_76_8907), .ZN(n_257_76_8908));
   NAND2_X1 i_257_76_8924 (.A1(n_257_76_8702), .A2(n_257_50), .ZN(n_257_76_8909));
   NOR2_X1 i_257_76_8925 (.A1(n_257_76_8908), .A2(n_257_76_8909), .ZN(
      n_257_76_8910));
   NAND4_X1 i_257_76_8926 (.A1(n_257_76_8906), .A2(n_257_76_8910), .A3(
      n_257_76_8752), .A4(n_257_76_8711), .ZN(n_257_76_8911));
   NOR2_X1 i_257_76_8927 (.A1(n_257_76_8911), .A2(n_257_76_8843), .ZN(
      n_257_76_8912));
   NAND3_X1 i_257_76_8928 (.A1(n_257_76_8912), .A2(n_257_76_8720), .A3(
      n_257_76_8678), .ZN(n_257_76_8913));
   NOR2_X1 i_257_76_8929 (.A1(n_257_76_8913), .A2(n_257_76_8722), .ZN(
      n_257_76_8914));
   NAND2_X1 i_257_76_8930 (.A1(n_257_76_18081), .A2(n_257_76_8914), .ZN(
      n_257_76_8915));
   NAND2_X1 i_257_76_8931 (.A1(n_257_449), .A2(n_257_76_8693), .ZN(n_257_76_8916));
   INV_X1 i_257_76_8932 (.A(n_257_76_8916), .ZN(n_257_76_8917));
   NAND2_X1 i_257_76_8933 (.A1(n_257_76_8699), .A2(n_257_1088), .ZN(
      n_257_76_8918));
   INV_X1 i_257_76_8934 (.A(n_257_76_8918), .ZN(n_257_76_8919));
   NAND3_X1 i_257_76_8935 (.A1(n_257_76_8917), .A2(n_257_76_8703), .A3(
      n_257_76_8919), .ZN(n_257_76_8920));
   NAND3_X1 i_257_76_8936 (.A1(n_257_76_8706), .A2(n_257_76_8707), .A3(
      n_257_76_8702), .ZN(n_257_76_8921));
   NOR2_X1 i_257_76_8937 (.A1(n_257_76_8920), .A2(n_257_76_8921), .ZN(
      n_257_76_8922));
   NAND3_X1 i_257_76_8938 (.A1(n_257_76_8922), .A2(n_257_76_8713), .A3(
      n_257_76_8714), .ZN(n_257_76_8923));
   NOR2_X1 i_257_76_8939 (.A1(n_257_76_8923), .A2(n_257_76_8718), .ZN(
      n_257_76_8924));
   NAND3_X1 i_257_76_8940 (.A1(n_257_76_8720), .A2(n_257_76_8924), .A3(
      n_257_76_8678), .ZN(n_257_76_8925));
   NOR2_X1 i_257_76_8941 (.A1(n_257_76_8925), .A2(n_257_76_8722), .ZN(
      n_257_76_8926));
   NAND2_X1 i_257_76_8942 (.A1(n_257_76_18083), .A2(n_257_76_8926), .ZN(
      n_257_76_8927));
   NAND2_X1 i_257_76_8943 (.A1(n_257_76_8759), .A2(n_257_76_8703), .ZN(
      n_257_76_8928));
   INV_X1 i_257_76_8944 (.A(n_257_76_8928), .ZN(n_257_76_8929));
   INV_X1 i_257_76_8945 (.A(n_257_612), .ZN(n_257_76_8930));
   NAND2_X1 i_257_76_8946 (.A1(n_257_76_8930), .A2(n_257_442), .ZN(n_257_76_8931));
   OAI21_X1 i_257_76_8947 (.A(n_257_76_8931), .B1(n_257_432), .B2(n_257_76_17412), 
      .ZN(n_257_76_8932));
   NAND2_X1 i_257_76_8948 (.A1(n_257_76_8932), .A2(n_257_429), .ZN(n_257_76_8933));
   INV_X1 i_257_76_8949 (.A(n_257_76_8933), .ZN(n_257_76_8934));
   NAND3_X1 i_257_76_8950 (.A1(n_257_76_8934), .A2(n_257_76_8699), .A3(
      n_257_76_8680), .ZN(n_257_76_8935));
   INV_X1 i_257_76_8951 (.A(n_257_76_8935), .ZN(n_257_76_8936));
   NAND3_X1 i_257_76_8952 (.A1(n_257_76_8929), .A2(n_257_76_8936), .A3(
      n_257_76_8702), .ZN(n_257_76_8937));
   NOR2_X1 i_257_76_8953 (.A1(n_257_76_8937), .A2(n_257_76_8709), .ZN(
      n_257_76_8938));
   NAND2_X1 i_257_76_8954 (.A1(n_257_76_8752), .A2(n_257_76_8746), .ZN(
      n_257_76_8939));
   INV_X1 i_257_76_8955 (.A(n_257_76_8939), .ZN(n_257_76_8940));
   NAND3_X1 i_257_76_8956 (.A1(n_257_76_8711), .A2(n_257_76_8679), .A3(
      n_257_76_8772), .ZN(n_257_76_8941));
   INV_X1 i_257_76_8957 (.A(n_257_76_8941), .ZN(n_257_76_8942));
   NAND4_X1 i_257_76_8958 (.A1(n_257_76_8938), .A2(n_257_76_8940), .A3(
      n_257_76_8714), .A4(n_257_76_8942), .ZN(n_257_76_8943));
   NAND4_X1 i_257_76_8959 (.A1(n_257_76_8754), .A2(n_257_167), .A3(n_257_76_8716), 
      .A4(n_257_76_8717), .ZN(n_257_76_8944));
   NOR2_X1 i_257_76_8960 (.A1(n_257_76_8943), .A2(n_257_76_8944), .ZN(
      n_257_76_8945));
   NAND3_X1 i_257_76_8961 (.A1(n_257_76_8945), .A2(n_257_76_8720), .A3(
      n_257_76_8678), .ZN(n_257_76_8946));
   NOR2_X1 i_257_76_8962 (.A1(n_257_76_8946), .A2(n_257_76_8722), .ZN(
      n_257_76_8947));
   NAND2_X1 i_257_76_8963 (.A1(n_257_76_18061), .A2(n_257_76_8947), .ZN(
      n_257_76_8948));
   NAND3_X1 i_257_76_8964 (.A1(n_257_76_8915), .A2(n_257_76_8927), .A3(
      n_257_76_8948), .ZN(n_257_76_8949));
   NAND2_X1 i_257_76_8965 (.A1(n_257_780), .A2(n_257_442), .ZN(n_257_76_8950));
   NOR2_X1 i_257_76_8966 (.A1(n_257_1074), .A2(n_257_76_8950), .ZN(n_257_76_8951));
   NAND4_X1 i_257_76_8967 (.A1(n_257_76_8703), .A2(n_257_447), .A3(n_257_76_8951), 
      .A4(n_257_76_8699), .ZN(n_257_76_8952));
   NOR2_X1 i_257_76_8968 (.A1(n_257_76_8952), .A2(n_257_76_8886), .ZN(
      n_257_76_8953));
   NAND4_X1 i_257_76_8969 (.A1(n_257_76_8717), .A2(n_257_76_8713), .A3(
      n_257_76_8953), .A4(n_257_76_8714), .ZN(n_257_76_8954));
   INV_X1 i_257_76_8970 (.A(n_257_76_8954), .ZN(n_257_76_8955));
   NAND2_X1 i_257_76_8971 (.A1(n_257_76_8678), .A2(n_257_76_8955), .ZN(
      n_257_76_8956));
   INV_X1 i_257_76_8972 (.A(n_257_76_8956), .ZN(n_257_76_8957));
   NAND2_X1 i_257_76_8973 (.A1(n_257_76_8957), .A2(n_257_76_8689), .ZN(
      n_257_76_8958));
   INV_X1 i_257_76_8974 (.A(n_257_76_8958), .ZN(n_257_76_8959));
   NAND2_X1 i_257_76_8975 (.A1(n_257_76_18085), .A2(n_257_76_8959), .ZN(
      n_257_76_8960));
   NAND4_X1 i_257_76_8976 (.A1(n_257_76_8716), .A2(n_257_76_8717), .A3(
      n_257_76_8714), .A4(n_257_90), .ZN(n_257_76_8961));
   NAND3_X1 i_257_76_8977 (.A1(n_257_76_8680), .A2(n_257_76_8932), .A3(n_257_431), 
      .ZN(n_257_76_8962));
   INV_X1 i_257_76_8978 (.A(n_257_76_8962), .ZN(n_257_76_8963));
   NAND4_X1 i_257_76_8979 (.A1(n_257_76_8963), .A2(n_257_76_8759), .A3(
      n_257_76_8703), .A4(n_257_76_8699), .ZN(n_257_76_8964));
   NOR2_X1 i_257_76_8980 (.A1(n_257_76_8964), .A2(n_257_76_8813), .ZN(
      n_257_76_8965));
   NAND4_X1 i_257_76_8981 (.A1(n_257_76_8965), .A2(n_257_76_8713), .A3(
      n_257_76_8752), .A4(n_257_76_8816), .ZN(n_257_76_8966));
   NOR2_X1 i_257_76_8982 (.A1(n_257_76_8961), .A2(n_257_76_8966), .ZN(
      n_257_76_8967));
   NAND3_X1 i_257_76_8983 (.A1(n_257_76_8967), .A2(n_257_76_8720), .A3(
      n_257_76_8678), .ZN(n_257_76_8968));
   NOR2_X1 i_257_76_8984 (.A1(n_257_76_8968), .A2(n_257_76_8722), .ZN(
      n_257_76_8969));
   NAND2_X1 i_257_76_8985 (.A1(n_257_76_18080), .A2(n_257_76_8969), .ZN(
      n_257_76_8970));
   NAND2_X1 i_257_76_8986 (.A1(n_257_76_8960), .A2(n_257_76_8970), .ZN(
      n_257_76_8971));
   NOR2_X1 i_257_76_8987 (.A1(n_257_76_8949), .A2(n_257_76_8971), .ZN(
      n_257_76_8972));
   NAND2_X1 i_257_76_8988 (.A1(n_257_76_8752), .A2(n_257_76_8711), .ZN(
      n_257_76_8973));
   INV_X1 i_257_76_8989 (.A(n_257_76_8973), .ZN(n_257_76_8974));
   NAND3_X1 i_257_76_8990 (.A1(n_257_76_8680), .A2(n_257_76_8932), .A3(n_257_430), 
      .ZN(n_257_76_8975));
   INV_X1 i_257_76_8991 (.A(n_257_76_8975), .ZN(n_257_76_8976));
   NAND4_X1 i_257_76_8992 (.A1(n_257_76_8976), .A2(n_257_76_8759), .A3(
      n_257_76_8703), .A4(n_257_76_8699), .ZN(n_257_76_8977));
   NOR2_X1 i_257_76_8993 (.A1(n_257_76_8749), .A2(n_257_76_8977), .ZN(
      n_257_76_8978));
   NAND4_X1 i_257_76_8994 (.A1(n_257_76_8679), .A2(n_257_128), .A3(n_257_76_8772), 
      .A4(n_257_76_8706), .ZN(n_257_76_8979));
   INV_X1 i_257_76_8995 (.A(n_257_76_8979), .ZN(n_257_76_8980));
   NAND4_X1 i_257_76_8996 (.A1(n_257_76_8974), .A2(n_257_76_8978), .A3(
      n_257_76_8980), .A4(n_257_76_8714), .ZN(n_257_76_8981));
   NOR2_X1 i_257_76_8997 (.A1(n_257_76_8981), .A2(n_257_76_8755), .ZN(
      n_257_76_8982));
   NAND3_X1 i_257_76_8998 (.A1(n_257_76_8982), .A2(n_257_76_8720), .A3(
      n_257_76_8678), .ZN(n_257_76_8983));
   NOR2_X1 i_257_76_8999 (.A1(n_257_76_8983), .A2(n_257_76_8722), .ZN(
      n_257_76_8984));
   NAND2_X1 i_257_76_9000 (.A1(n_257_76_18068), .A2(n_257_76_8984), .ZN(
      n_257_76_8985));
   NAND3_X1 i_257_76_9001 (.A1(n_257_76_18037), .A2(n_257_76_8706), .A3(
      n_257_76_8707), .ZN(n_257_76_8986));
   NAND2_X1 i_257_76_9002 (.A1(n_257_448), .A2(n_257_76_8680), .ZN(n_257_76_8987));
   INV_X1 i_257_76_9003 (.A(n_257_76_8987), .ZN(n_257_76_8988));
   NAND3_X1 i_257_76_9004 (.A1(n_257_76_8988), .A2(n_257_76_8702), .A3(
      n_257_76_8699), .ZN(n_257_76_8989));
   NOR2_X1 i_257_76_9005 (.A1(n_257_76_8986), .A2(n_257_76_8989), .ZN(
      n_257_76_8990));
   NAND3_X1 i_257_76_9006 (.A1(n_257_76_8990), .A2(n_257_76_8713), .A3(
      n_257_76_8714), .ZN(n_257_76_8991));
   NOR2_X1 i_257_76_9007 (.A1(n_257_76_8991), .A2(n_257_76_8718), .ZN(
      n_257_76_8992));
   NAND3_X1 i_257_76_9008 (.A1(n_257_76_8992), .A2(n_257_76_8678), .A3(n_257_684), 
      .ZN(n_257_76_8993));
   NOR2_X1 i_257_76_9009 (.A1(n_257_76_8722), .A2(n_257_76_8993), .ZN(
      n_257_76_8994));
   NAND2_X1 i_257_76_9010 (.A1(n_257_76_18079), .A2(n_257_76_8994), .ZN(
      n_257_76_8995));
   NAND2_X1 i_257_76_9011 (.A1(n_257_76_8720), .A2(n_257_76_8678), .ZN(
      n_257_76_8996));
   INV_X1 i_257_76_9012 (.A(n_257_76_8996), .ZN(n_257_76_8997));
   NAND3_X1 i_257_76_9013 (.A1(n_257_76_8754), .A2(n_257_247), .A3(n_257_76_8716), 
      .ZN(n_257_76_8998));
   INV_X1 i_257_76_9014 (.A(n_257_76_8998), .ZN(n_257_76_8999));
   NAND3_X1 i_257_76_9015 (.A1(n_257_76_8708), .A2(n_257_76_8702), .A3(
      n_257_76_8776), .ZN(n_257_76_9000));
   INV_X1 i_257_76_9016 (.A(n_257_76_9000), .ZN(n_257_76_9001));
   NAND2_X1 i_257_76_9017 (.A1(n_257_76_8706), .A2(n_257_76_8707), .ZN(
      n_257_76_9002));
   INV_X1 i_257_76_9018 (.A(n_257_76_9002), .ZN(n_257_76_9003));
   NAND2_X1 i_257_76_9019 (.A1(n_257_76_8767), .A2(n_257_425), .ZN(n_257_76_9004));
   INV_X1 i_257_76_9020 (.A(n_257_76_9004), .ZN(n_257_76_9005));
   NAND3_X1 i_257_76_9021 (.A1(n_257_76_9005), .A2(n_257_76_8680), .A3(
      n_257_76_8763), .ZN(n_257_76_9006));
   INV_X1 i_257_76_9022 (.A(n_257_76_9006), .ZN(n_257_76_9007));
   NAND4_X1 i_257_76_9023 (.A1(n_257_76_9007), .A2(n_257_76_8759), .A3(
      n_257_76_8703), .A4(n_257_76_8699), .ZN(n_257_76_9008));
   INV_X1 i_257_76_9024 (.A(n_257_76_9008), .ZN(n_257_76_9009));
   NAND3_X1 i_257_76_9025 (.A1(n_257_76_9001), .A2(n_257_76_9003), .A3(
      n_257_76_9009), .ZN(n_257_76_9010));
   NAND4_X1 i_257_76_9026 (.A1(n_257_76_8711), .A2(n_257_76_8679), .A3(
      n_257_76_8772), .A4(n_257_76_8773), .ZN(n_257_76_9011));
   NOR2_X1 i_257_76_9027 (.A1(n_257_76_9010), .A2(n_257_76_9011), .ZN(
      n_257_76_9012));
   NAND4_X1 i_257_76_9028 (.A1(n_257_76_8717), .A2(n_257_76_8714), .A3(
      n_257_76_8752), .A4(n_257_76_8746), .ZN(n_257_76_9013));
   INV_X1 i_257_76_9029 (.A(n_257_76_9013), .ZN(n_257_76_9014));
   NAND4_X1 i_257_76_9030 (.A1(n_257_76_8999), .A2(n_257_76_9012), .A3(
      n_257_76_9014), .A4(n_257_76_8758), .ZN(n_257_76_9015));
   INV_X1 i_257_76_9031 (.A(n_257_76_9015), .ZN(n_257_76_9016));
   NAND3_X1 i_257_76_9032 (.A1(n_257_76_8997), .A2(n_257_76_9016), .A3(
      n_257_76_8689), .ZN(n_257_76_9017));
   INV_X1 i_257_76_9033 (.A(n_257_76_9017), .ZN(n_257_76_9018));
   NAND2_X1 i_257_76_9034 (.A1(n_257_76_18064), .A2(n_257_76_9018), .ZN(
      n_257_76_9019));
   NAND3_X1 i_257_76_9035 (.A1(n_257_76_8985), .A2(n_257_76_8995), .A3(
      n_257_76_9019), .ZN(n_257_76_9020));
   NAND4_X1 i_257_76_9036 (.A1(n_257_76_8693), .A2(n_257_76_8699), .A3(
      n_257_1080), .A4(n_257_438), .ZN(n_257_76_9021));
   INV_X1 i_257_76_9037 (.A(n_257_76_9021), .ZN(n_257_76_9022));
   NAND3_X1 i_257_76_9038 (.A1(n_257_76_8711), .A2(n_257_76_9022), .A3(
      n_257_76_8679), .ZN(n_257_76_9023));
   INV_X1 i_257_76_9039 (.A(n_257_76_9023), .ZN(n_257_76_9024));
   NAND2_X1 i_257_76_9040 (.A1(n_257_76_8678), .A2(n_257_76_9024), .ZN(
      n_257_76_9025));
   INV_X1 i_257_76_9041 (.A(n_257_76_9025), .ZN(n_257_76_9026));
   NAND2_X1 i_257_76_9042 (.A1(n_257_76_9026), .A2(n_257_76_8689), .ZN(
      n_257_76_9027));
   INV_X1 i_257_76_9043 (.A(n_257_76_9027), .ZN(n_257_76_9028));
   NAND2_X1 i_257_76_9044 (.A1(n_257_76_18067), .A2(n_257_76_9028), .ZN(
      n_257_76_9029));
   NAND2_X1 i_257_76_9045 (.A1(n_257_325), .A2(n_257_422), .ZN(n_257_76_9030));
   NAND3_X1 i_257_76_9046 (.A1(n_257_76_8708), .A2(n_257_76_8702), .A3(
      n_257_76_9030), .ZN(n_257_76_9031));
   NAND4_X1 i_257_76_9047 (.A1(n_257_76_8776), .A2(n_257_76_8759), .A3(
      n_257_76_8703), .A4(n_257_76_8699), .ZN(n_257_76_9032));
   NOR2_X1 i_257_76_9048 (.A1(n_257_76_9031), .A2(n_257_76_9032), .ZN(
      n_257_76_9033));
   NAND2_X1 i_257_76_9049 (.A1(n_257_287), .A2(n_257_423), .ZN(n_257_76_9034));
   NOR2_X1 i_257_76_9050 (.A1(n_257_76_17646), .A2(n_257_580), .ZN(n_257_76_9035));
   AOI21_X1 i_257_76_9051 (.A(n_257_76_9035), .B1(n_257_76_16810), .B2(
      n_257_76_17944), .ZN(n_257_76_9036));
   NOR2_X1 i_257_76_9052 (.A1(n_257_1074), .A2(n_257_76_9036), .ZN(n_257_76_9037));
   NAND2_X1 i_257_76_9053 (.A1(n_257_420), .A2(n_257_76_8767), .ZN(n_257_76_9038));
   INV_X1 i_257_76_9054 (.A(n_257_76_9038), .ZN(n_257_76_9039));
   NAND3_X1 i_257_76_9055 (.A1(n_257_76_9037), .A2(n_257_76_8766), .A3(
      n_257_76_9039), .ZN(n_257_76_9040));
   INV_X1 i_257_76_9056 (.A(n_257_76_9040), .ZN(n_257_76_9041));
   NAND3_X1 i_257_76_9057 (.A1(n_257_76_9034), .A2(n_257_76_8679), .A3(
      n_257_76_9041), .ZN(n_257_76_9042));
   INV_X1 i_257_76_9058 (.A(n_257_76_9042), .ZN(n_257_76_9043));
   NAND4_X1 i_257_76_9059 (.A1(n_257_76_8772), .A2(n_257_76_8773), .A3(
      n_257_76_8706), .A4(n_257_76_8707), .ZN(n_257_76_9044));
   INV_X1 i_257_76_9060 (.A(n_257_76_9044), .ZN(n_257_76_9045));
   NAND3_X1 i_257_76_9061 (.A1(n_257_76_9033), .A2(n_257_76_9043), .A3(
      n_257_76_9045), .ZN(n_257_76_9046));
   INV_X1 i_257_76_9062 (.A(n_257_76_9046), .ZN(n_257_76_9047));
   INV_X1 i_257_76_9063 (.A(n_257_76_8718), .ZN(n_257_76_9048));
   NAND3_X1 i_257_76_9064 (.A1(n_257_76_8752), .A2(n_257_76_8746), .A3(
      n_257_76_8711), .ZN(n_257_76_9049));
   NOR2_X1 i_257_76_9065 (.A1(n_257_76_9049), .A2(n_257_76_8730), .ZN(
      n_257_76_9050));
   NAND3_X1 i_257_76_9066 (.A1(n_257_76_9047), .A2(n_257_76_9048), .A3(
      n_257_76_9050), .ZN(n_257_76_9051));
   NAND2_X1 i_257_76_9067 (.A1(n_257_364), .A2(n_257_421), .ZN(n_257_76_9052));
   NAND4_X1 i_257_76_9068 (.A1(n_257_76_8757), .A2(n_257_76_8758), .A3(
      n_257_76_9052), .A4(n_257_76_8754), .ZN(n_257_76_9053));
   NOR2_X1 i_257_76_9069 (.A1(n_257_76_9051), .A2(n_257_76_9053), .ZN(
      n_257_76_9054));
   NAND3_X1 i_257_76_9070 (.A1(n_257_76_9054), .A2(n_257_76_8997), .A3(
      n_257_76_8689), .ZN(n_257_76_9055));
   INV_X1 i_257_76_9071 (.A(n_257_76_9055), .ZN(n_257_76_9056));
   NAND2_X1 i_257_76_9072 (.A1(n_257_76_18073), .A2(n_257_76_9056), .ZN(
      n_257_76_9057));
   NAND2_X1 i_257_76_9073 (.A1(n_257_76_9029), .A2(n_257_76_9057), .ZN(
      n_257_76_9058));
   NOR2_X1 i_257_76_9074 (.A1(n_257_76_9020), .A2(n_257_76_9058), .ZN(
      n_257_76_9059));
   NAND2_X1 i_257_76_9075 (.A1(n_257_76_8773), .A2(n_257_76_8706), .ZN(
      n_257_76_9060));
   NOR2_X1 i_257_76_9076 (.A1(n_257_76_9060), .A2(n_257_76_8749), .ZN(
      n_257_76_9061));
   NAND3_X1 i_257_76_9077 (.A1(n_257_76_9034), .A2(n_257_76_8679), .A3(
      n_257_76_8772), .ZN(n_257_76_9062));
   INV_X1 i_257_76_9078 (.A(n_257_76_9062), .ZN(n_257_76_9063));
   NAND2_X1 i_257_76_9079 (.A1(n_257_76_8767), .A2(n_257_421), .ZN(n_257_76_9064));
   INV_X1 i_257_76_9080 (.A(n_257_76_9064), .ZN(n_257_76_9065));
   NAND3_X1 i_257_76_9081 (.A1(n_257_76_9065), .A2(n_257_76_8680), .A3(
      n_257_76_8763), .ZN(n_257_76_9066));
   INV_X1 i_257_76_9082 (.A(n_257_76_9066), .ZN(n_257_76_9067));
   NAND4_X1 i_257_76_9083 (.A1(n_257_76_9067), .A2(n_257_76_8703), .A3(
      n_257_76_8699), .A4(n_257_76_8766), .ZN(n_257_76_9068));
   NAND3_X1 i_257_76_9084 (.A1(n_257_76_9030), .A2(n_257_76_8776), .A3(
      n_257_76_8759), .ZN(n_257_76_9069));
   NOR2_X1 i_257_76_9085 (.A1(n_257_76_9068), .A2(n_257_76_9069), .ZN(
      n_257_76_9070));
   NAND3_X1 i_257_76_9086 (.A1(n_257_76_9061), .A2(n_257_76_9063), .A3(
      n_257_76_9070), .ZN(n_257_76_9071));
   NAND4_X1 i_257_76_9087 (.A1(n_257_76_8714), .A2(n_257_76_8752), .A3(
      n_257_76_8746), .A4(n_257_76_8711), .ZN(n_257_76_9072));
   NOR2_X1 i_257_76_9088 (.A1(n_257_76_9071), .A2(n_257_76_9072), .ZN(
      n_257_76_9073));
   NAND2_X1 i_257_76_9089 (.A1(n_257_76_8757), .A2(n_257_76_8758), .ZN(
      n_257_76_9074));
   INV_X1 i_257_76_9090 (.A(n_257_76_9074), .ZN(n_257_76_9075));
   NAND4_X1 i_257_76_9091 (.A1(n_257_76_8754), .A2(n_257_76_8716), .A3(n_257_364), 
      .A4(n_257_76_8717), .ZN(n_257_76_9076));
   INV_X1 i_257_76_9092 (.A(n_257_76_9076), .ZN(n_257_76_9077));
   NAND3_X1 i_257_76_9093 (.A1(n_257_76_9073), .A2(n_257_76_9075), .A3(
      n_257_76_9077), .ZN(n_257_76_9078));
   NOR3_X1 i_257_76_9094 (.A1(n_257_76_8722), .A2(n_257_76_9078), .A3(
      n_257_76_8996), .ZN(n_257_76_9079));
   NAND2_X1 i_257_76_9095 (.A1(n_257_76_18082), .A2(n_257_76_9079), .ZN(
      n_257_76_9080));
   NAND2_X1 i_257_76_9096 (.A1(n_257_427), .A2(n_257_76_8767), .ZN(n_257_76_9081));
   INV_X1 i_257_76_9097 (.A(n_257_76_9081), .ZN(n_257_76_9082));
   NAND3_X1 i_257_76_9098 (.A1(n_257_76_8765), .A2(n_257_207), .A3(n_257_76_9082), 
      .ZN(n_257_76_9083));
   INV_X1 i_257_76_9099 (.A(n_257_76_9083), .ZN(n_257_76_9084));
   NAND4_X1 i_257_76_9100 (.A1(n_257_76_8679), .A2(n_257_76_9084), .A3(
      n_257_76_8772), .A4(n_257_76_8706), .ZN(n_257_76_9085));
   INV_X1 i_257_76_9101 (.A(n_257_76_9085), .ZN(n_257_76_9086));
   NOR2_X1 i_257_76_9102 (.A1(n_257_76_8749), .A2(n_257_76_8760), .ZN(
      n_257_76_9087));
   NAND3_X1 i_257_76_9103 (.A1(n_257_76_9086), .A2(n_257_76_8748), .A3(
      n_257_76_9087), .ZN(n_257_76_9088));
   NOR2_X1 i_257_76_9104 (.A1(n_257_76_9088), .A2(n_257_76_8818), .ZN(
      n_257_76_9089));
   NAND4_X1 i_257_76_9105 (.A1(n_257_76_8720), .A2(n_257_76_8678), .A3(
      n_257_76_8822), .A4(n_257_76_9089), .ZN(n_257_76_9090));
   NOR2_X1 i_257_76_9106 (.A1(n_257_76_9090), .A2(n_257_76_8722), .ZN(
      n_257_76_9091));
   NAND2_X1 i_257_76_9107 (.A1(n_257_76_18065), .A2(n_257_76_9091), .ZN(
      n_257_76_9092));
   NAND4_X1 i_257_76_9108 (.A1(n_257_76_8703), .A2(n_257_76_8693), .A3(
      n_257_76_8699), .A4(n_257_467), .ZN(n_257_76_9093));
   NAND2_X1 i_257_76_9109 (.A1(n_257_76_8702), .A2(n_257_76_8759), .ZN(
      n_257_76_9094));
   NOR2_X1 i_257_76_9110 (.A1(n_257_76_9093), .A2(n_257_76_9094), .ZN(
      n_257_76_9095));
   NAND2_X1 i_257_76_9111 (.A1(n_257_76_8679), .A2(n_257_451), .ZN(n_257_76_9096));
   INV_X1 i_257_76_9112 (.A(n_257_76_9096), .ZN(n_257_76_9097));
   INV_X1 i_257_76_9113 (.A(n_257_76_8709), .ZN(n_257_76_9098));
   NAND4_X1 i_257_76_9114 (.A1(n_257_76_9095), .A2(n_257_76_9097), .A3(
      n_257_76_8711), .A4(n_257_76_9098), .ZN(n_257_76_9099));
   NOR2_X1 i_257_76_9115 (.A1(n_257_76_9099), .A2(n_257_76_8843), .ZN(
      n_257_76_9100));
   NAND3_X1 i_257_76_9116 (.A1(n_257_76_8720), .A2(n_257_76_9100), .A3(
      n_257_76_8678), .ZN(n_257_76_9101));
   NOR2_X1 i_257_76_9117 (.A1(n_257_76_9101), .A2(n_257_76_8722), .ZN(
      n_257_76_9102));
   NAND2_X1 i_257_76_9118 (.A1(n_257_76_18063), .A2(n_257_76_9102), .ZN(
      n_257_76_9103));
   NAND3_X1 i_257_76_9119 (.A1(n_257_76_9080), .A2(n_257_76_9092), .A3(
      n_257_76_9103), .ZN(n_257_76_9104));
   NAND4_X1 i_257_76_9120 (.A1(n_257_76_8706), .A2(n_257_76_8707), .A3(
      n_257_76_8708), .A4(n_257_76_8702), .ZN(n_257_76_9105));
   NOR2_X1 i_257_76_9121 (.A1(n_257_76_9105), .A2(n_257_76_9032), .ZN(
      n_257_76_9106));
   NAND2_X1 i_257_76_9122 (.A1(n_257_76_8767), .A2(n_257_424), .ZN(n_257_76_9107));
   INV_X1 i_257_76_9123 (.A(n_257_76_9107), .ZN(n_257_76_9108));
   NAND4_X1 i_257_76_9124 (.A1(n_257_76_9108), .A2(n_257_76_8680), .A3(n_257_516), 
      .A4(n_257_76_8763), .ZN(n_257_76_9109));
   INV_X1 i_257_76_9125 (.A(n_257_76_9109), .ZN(n_257_76_9110));
   NAND4_X1 i_257_76_9126 (.A1(n_257_76_8679), .A2(n_257_76_8772), .A3(
      n_257_76_8773), .A4(n_257_76_9110), .ZN(n_257_76_9111));
   INV_X1 i_257_76_9127 (.A(n_257_76_9111), .ZN(n_257_76_9112));
   NAND3_X1 i_257_76_9128 (.A1(n_257_76_9106), .A2(n_257_76_8748), .A3(
      n_257_76_9112), .ZN(n_257_76_9113));
   NAND4_X1 i_257_76_9129 (.A1(n_257_76_8716), .A2(n_257_76_8717), .A3(
      n_257_76_8714), .A4(n_257_76_8752), .ZN(n_257_76_9114));
   NOR2_X1 i_257_76_9130 (.A1(n_257_76_9113), .A2(n_257_76_9114), .ZN(
      n_257_76_9115));
   NAND3_X1 i_257_76_9131 (.A1(n_257_76_8757), .A2(n_257_76_8758), .A3(
      n_257_76_8754), .ZN(n_257_76_9116));
   INV_X1 i_257_76_9132 (.A(n_257_76_9116), .ZN(n_257_76_9117));
   NAND4_X1 i_257_76_9133 (.A1(n_257_76_9115), .A2(n_257_76_8720), .A3(
      n_257_76_8678), .A4(n_257_76_9117), .ZN(n_257_76_9118));
   NOR2_X1 i_257_76_9134 (.A1(n_257_76_9118), .A2(n_257_76_8722), .ZN(
      n_257_76_9119));
   NAND2_X1 i_257_76_9135 (.A1(n_257_76_18062), .A2(n_257_76_9119), .ZN(
      n_257_76_9120));
   INV_X1 i_257_76_9136 (.A(n_257_76_8749), .ZN(n_257_76_9121));
   NAND3_X1 i_257_76_9137 (.A1(n_257_76_9121), .A2(n_257_76_8711), .A3(
      n_257_76_8679), .ZN(n_257_76_9122));
   NOR2_X1 i_257_76_9138 (.A1(n_257_76_9122), .A2(n_257_76_8939), .ZN(
      n_257_76_9123));
   INV_X1 i_257_76_9139 (.A(n_257_76_8865), .ZN(n_257_76_9124));
   NAND4_X1 i_257_76_9140 (.A1(n_257_76_9123), .A2(n_257_76_9124), .A3(
      n_257_76_8754), .A4(n_257_76_8716), .ZN(n_257_76_9125));
   NAND3_X1 i_257_76_9141 (.A1(n_257_76_8703), .A2(n_257_76_8699), .A3(n_257_325), 
      .ZN(n_257_76_9126));
   NAND2_X1 i_257_76_9142 (.A1(n_257_422), .A2(n_257_76_8767), .ZN(n_257_76_9127));
   INV_X1 i_257_76_9143 (.A(n_257_76_9127), .ZN(n_257_76_9128));
   NAND3_X1 i_257_76_9144 (.A1(n_257_76_8765), .A2(n_257_76_8766), .A3(
      n_257_76_9128), .ZN(n_257_76_9129));
   NOR2_X1 i_257_76_9145 (.A1(n_257_76_9126), .A2(n_257_76_9129), .ZN(
      n_257_76_9130));
   NAND3_X1 i_257_76_9146 (.A1(n_257_76_8706), .A2(n_257_76_8776), .A3(
      n_257_76_8759), .ZN(n_257_76_9131));
   INV_X1 i_257_76_9147 (.A(n_257_76_9131), .ZN(n_257_76_9132));
   NAND4_X1 i_257_76_9148 (.A1(n_257_76_9130), .A2(n_257_76_8775), .A3(
      n_257_76_9034), .A4(n_257_76_9132), .ZN(n_257_76_9133));
   INV_X1 i_257_76_9149 (.A(n_257_76_9133), .ZN(n_257_76_9134));
   NAND3_X1 i_257_76_9150 (.A1(n_257_76_9134), .A2(n_257_76_8757), .A3(
      n_257_76_8758), .ZN(n_257_76_9135));
   NOR2_X1 i_257_76_9151 (.A1(n_257_76_9125), .A2(n_257_76_9135), .ZN(
      n_257_76_9136));
   NAND3_X1 i_257_76_9152 (.A1(n_257_76_9136), .A2(n_257_76_8997), .A3(
      n_257_76_8689), .ZN(n_257_76_9137));
   INV_X1 i_257_76_9153 (.A(n_257_76_9137), .ZN(n_257_76_9138));
   NAND2_X1 i_257_76_9154 (.A1(n_257_342), .A2(n_257_76_9138), .ZN(n_257_76_9139));
   NAND2_X1 i_257_76_9155 (.A1(n_257_748), .A2(n_257_76_17935), .ZN(
      n_257_76_9140));
   NAND2_X1 i_257_76_9156 (.A1(n_257_812), .A2(n_257_76_17952), .ZN(
      n_257_76_9141));
   NAND2_X1 i_257_76_9157 (.A1(n_257_876), .A2(n_257_76_17903), .ZN(
      n_257_76_9142));
   NAND4_X1 i_257_76_9158 (.A1(n_257_76_8851), .A2(n_257_76_9140), .A3(
      n_257_76_9141), .A4(n_257_76_9142), .ZN(n_257_76_9143));
   NAND2_X1 i_257_76_9159 (.A1(n_257_716), .A2(n_257_76_15655), .ZN(
      n_257_76_9144));
   NAND2_X1 i_257_76_9160 (.A1(n_257_844), .A2(n_257_442), .ZN(n_257_76_9145));
   INV_X1 i_257_76_9161 (.A(n_257_76_9145), .ZN(n_257_76_9146));
   NAND2_X1 i_257_76_9162 (.A1(n_257_446), .A2(n_257_76_9146), .ZN(n_257_76_9147));
   NAND2_X1 i_257_76_9163 (.A1(n_257_449), .A2(n_257_76_16422), .ZN(
      n_257_76_9148));
   INV_X1 i_257_76_9164 (.A(n_257_76_8950), .ZN(n_257_76_9149));
   NAND2_X1 i_257_76_9165 (.A1(n_257_447), .A2(n_257_76_9149), .ZN(n_257_76_9150));
   NAND4_X1 i_257_76_9166 (.A1(n_257_76_9144), .A2(n_257_76_9147), .A3(
      n_257_76_9148), .A4(n_257_76_9150), .ZN(n_257_76_9151));
   NAND3_X1 i_257_76_9167 (.A1(n_257_1080), .A2(n_257_438), .A3(n_257_442), 
      .ZN(n_257_76_9152));
   NAND2_X1 i_257_76_9168 (.A1(n_257_644), .A2(n_257_76_17928), .ZN(
      n_257_76_9153));
   NAND2_X1 i_257_76_9169 (.A1(n_257_440), .A2(n_257_76_8682), .ZN(n_257_76_9154));
   NAND4_X1 i_257_76_9170 (.A1(n_257_76_9109), .A2(n_257_76_9152), .A3(
      n_257_76_9153), .A4(n_257_76_9154), .ZN(n_257_76_9155));
   NOR2_X1 i_257_76_9171 (.A1(n_257_76_9151), .A2(n_257_76_9155), .ZN(
      n_257_76_9156));
   NAND2_X1 i_257_76_9172 (.A1(n_257_467), .A2(n_257_442), .ZN(n_257_76_9157));
   INV_X1 i_257_76_9173 (.A(n_257_76_9157), .ZN(n_257_76_9158));
   NAND2_X1 i_257_76_9174 (.A1(n_257_451), .A2(n_257_76_9158), .ZN(n_257_76_9159));
   NAND2_X1 i_257_76_9175 (.A1(n_257_128), .A2(n_257_76_17925), .ZN(
      n_257_76_9160));
   NAND2_X1 i_257_76_9176 (.A1(n_257_914), .A2(n_257_76_17940), .ZN(
      n_257_76_9161));
   NAND3_X1 i_257_76_9177 (.A1(n_257_76_9159), .A2(n_257_76_9160), .A3(
      n_257_76_9161), .ZN(n_257_76_9162));
   INV_X1 i_257_76_9178 (.A(n_257_76_9162), .ZN(n_257_76_9163));
   NAND2_X1 i_257_76_9179 (.A1(n_257_978), .A2(n_257_442), .ZN(n_257_76_9164));
   INV_X1 i_257_76_9180 (.A(n_257_76_9164), .ZN(n_257_76_9165));
   NAND2_X1 i_257_76_9181 (.A1(n_257_441), .A2(n_257_76_9165), .ZN(n_257_76_9166));
   NAND2_X1 i_257_76_9182 (.A1(n_257_50), .A2(n_257_76_17918), .ZN(n_257_76_9167));
   NAND2_X1 i_257_76_9183 (.A1(n_257_76_9166), .A2(n_257_76_9167), .ZN(
      n_257_76_9168));
   NAND2_X1 i_257_76_9184 (.A1(n_257_428), .A2(n_257_580), .ZN(n_257_76_9169));
   NAND2_X1 i_257_76_9185 (.A1(n_257_76_8767), .A2(n_257_76_9169), .ZN(
      n_257_76_9170));
   INV_X1 i_257_76_9186 (.A(n_257_76_9170), .ZN(n_257_76_9171));
   INV_X1 i_257_76_9187 (.A(Small_Packet_Data_Size[15]), .ZN(n_257_76_9172));
   NAND3_X1 i_257_76_9188 (.A1(n_257_76_9171), .A2(n_257_76_8680), .A3(
      n_257_76_18038), .ZN(n_257_76_9173));
   NAND2_X1 i_257_76_9189 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[15]), 
      .ZN(n_257_76_9174));
   NAND2_X1 i_257_76_9190 (.A1(n_257_76_9173), .A2(n_257_76_9174), .ZN(
      n_257_76_9175));
   NAND3_X1 i_257_76_9191 (.A1(n_257_76_9175), .A2(n_257_76_9040), .A3(
      n_257_76_9083), .ZN(n_257_76_9176));
   NOR2_X1 i_257_76_9192 (.A1(n_257_76_9168), .A2(n_257_76_9176), .ZN(
      n_257_76_9177));
   NAND3_X1 i_257_76_9193 (.A1(n_257_76_9156), .A2(n_257_76_9163), .A3(
      n_257_76_9177), .ZN(n_257_76_9178));
   NOR2_X1 i_257_76_9194 (.A1(n_257_76_9143), .A2(n_257_76_9178), .ZN(
      n_257_76_9179));
   NAND2_X1 i_257_76_9195 (.A1(n_257_167), .A2(n_257_76_17331), .ZN(
      n_257_76_9180));
   NAND2_X1 i_257_76_9196 (.A1(n_257_90), .A2(n_257_76_17932), .ZN(n_257_76_9181));
   NAND4_X1 i_257_76_9197 (.A1(n_257_76_9180), .A2(n_257_76_9133), .A3(
      n_257_76_8779), .A4(n_257_76_9181), .ZN(n_257_76_9182));
   INV_X1 i_257_76_9198 (.A(n_257_76_9182), .ZN(n_257_76_9183));
   NAND2_X1 i_257_76_9199 (.A1(n_257_1010), .A2(n_257_76_17964), .ZN(
      n_257_76_9184));
   NAND3_X1 i_257_76_9200 (.A1(n_257_76_9179), .A2(n_257_76_9183), .A3(
      n_257_76_9184), .ZN(n_257_76_9185));
   INV_X1 i_257_76_9201 (.A(n_257_76_9185), .ZN(n_257_76_9186));
   NAND2_X1 i_257_76_9202 (.A1(n_257_684), .A2(n_257_76_17958), .ZN(
      n_257_76_9187));
   NAND2_X1 i_257_76_9203 (.A1(n_257_76_9015), .A2(n_257_76_9187), .ZN(
      n_257_76_9188));
   INV_X1 i_257_76_9204 (.A(n_257_76_9188), .ZN(n_257_76_9189));
   NAND2_X1 i_257_76_9205 (.A1(n_257_1042), .A2(n_257_76_17969), .ZN(
      n_257_76_9190));
   NAND4_X1 i_257_76_9206 (.A1(n_257_76_9186), .A2(n_257_76_9189), .A3(
      n_257_76_9078), .A4(n_257_76_9190), .ZN(n_257_76_9191));
   INV_X1 i_257_76_9207 (.A(n_257_76_9191), .ZN(n_257_76_9192));
   NAND4_X1 i_257_76_9208 (.A1(n_257_76_8711), .A2(n_257_76_9034), .A3(
      n_257_76_8679), .A4(n_257_76_8772), .ZN(n_257_76_9193));
   NOR2_X1 i_257_76_9209 (.A1(n_257_76_9193), .A2(n_257_76_8939), .ZN(
      n_257_76_9194));
   NAND4_X1 i_257_76_9210 (.A1(n_257_76_9194), .A2(n_257_76_9124), .A3(
      n_257_76_8754), .A4(n_257_76_8716), .ZN(n_257_76_9195));
   NAND2_X1 i_257_76_9211 (.A1(n_257_76_8699), .A2(n_257_76_8766), .ZN(
      n_257_76_9196));
   NAND3_X1 i_257_76_9212 (.A1(n_257_403), .A2(n_257_484), .A3(n_257_442), 
      .ZN(n_257_76_9197));
   INV_X1 i_257_76_9213 (.A(n_257_76_9197), .ZN(n_257_76_9198));
   NAND3_X1 i_257_76_9214 (.A1(n_257_76_8767), .A2(n_257_76_9169), .A3(
      n_257_76_9198), .ZN(n_257_76_9199));
   INV_X1 i_257_76_9215 (.A(n_257_76_9199), .ZN(n_257_76_9200));
   NAND2_X1 i_257_76_9216 (.A1(n_257_420), .A2(n_257_668), .ZN(n_257_76_9201));
   NAND3_X1 i_257_76_9217 (.A1(n_257_76_9200), .A2(n_257_76_9201), .A3(
      n_257_76_8680), .ZN(n_257_76_9202));
   NOR2_X1 i_257_76_9218 (.A1(n_257_76_9196), .A2(n_257_76_9202), .ZN(
      n_257_76_9203));
   NAND2_X1 i_257_76_9219 (.A1(n_257_76_8702), .A2(n_257_76_9030), .ZN(
      n_257_76_9204));
   INV_X1 i_257_76_9220 (.A(n_257_76_9204), .ZN(n_257_76_9205));
   NAND3_X1 i_257_76_9221 (.A1(n_257_76_8776), .A2(n_257_76_8759), .A3(
      n_257_76_8703), .ZN(n_257_76_9206));
   INV_X1 i_257_76_9222 (.A(n_257_76_9206), .ZN(n_257_76_9207));
   NAND3_X1 i_257_76_9223 (.A1(n_257_76_9203), .A2(n_257_76_9205), .A3(
      n_257_76_9207), .ZN(n_257_76_9208));
   NAND4_X1 i_257_76_9224 (.A1(n_257_76_8773), .A2(n_257_76_8706), .A3(
      n_257_76_8707), .A4(n_257_76_8708), .ZN(n_257_76_9209));
   NOR2_X1 i_257_76_9225 (.A1(n_257_76_9208), .A2(n_257_76_9209), .ZN(
      n_257_76_9210));
   NAND4_X1 i_257_76_9226 (.A1(n_257_76_9210), .A2(n_257_76_8757), .A3(
      n_257_76_8758), .A4(n_257_76_9052), .ZN(n_257_76_9211));
   NOR2_X1 i_257_76_9227 (.A1(n_257_76_9195), .A2(n_257_76_9211), .ZN(
      n_257_76_9212));
   NAND3_X1 i_257_76_9228 (.A1(n_257_76_9212), .A2(n_257_76_8997), .A3(
      n_257_76_8689), .ZN(n_257_76_9213));
   INV_X1 i_257_76_9229 (.A(n_257_76_9213), .ZN(n_257_76_9214));
   AOI21_X1 i_257_76_9230 (.A(n_257_76_9192), .B1(n_257_76_18060), .B2(
      n_257_76_9214), .ZN(n_257_76_9215));
   NAND3_X1 i_257_76_9231 (.A1(n_257_76_9120), .A2(n_257_76_9139), .A3(
      n_257_76_9215), .ZN(n_257_76_9216));
   NOR2_X1 i_257_76_9232 (.A1(n_257_76_9104), .A2(n_257_76_9216), .ZN(
      n_257_76_9217));
   NAND3_X1 i_257_76_9233 (.A1(n_257_76_8972), .A2(n_257_76_9059), .A3(
      n_257_76_9217), .ZN(n_257_76_9218));
   INV_X1 i_257_76_9234 (.A(n_257_76_9218), .ZN(n_257_76_9219));
   NAND2_X1 i_257_76_9235 (.A1(n_257_76_8905), .A2(n_257_76_9219), .ZN(n_15));
   NAND2_X1 i_257_76_9236 (.A1(n_257_1011), .A2(n_257_444), .ZN(n_257_76_9220));
   NAND2_X1 i_257_76_9237 (.A1(n_257_1043), .A2(n_257_443), .ZN(n_257_76_9221));
   NAND2_X1 i_257_76_9238 (.A1(n_257_441), .A2(n_257_979), .ZN(n_257_76_9222));
   INV_X1 i_257_76_9239 (.A(n_257_1075), .ZN(n_257_76_9223));
   NAND2_X1 i_257_76_9240 (.A1(n_257_947), .A2(n_257_442), .ZN(n_257_76_9224));
   INV_X1 i_257_76_9241 (.A(n_257_76_9224), .ZN(n_257_76_9225));
   NAND3_X1 i_257_76_9242 (.A1(n_257_76_9223), .A2(n_257_440), .A3(n_257_76_9225), 
      .ZN(n_257_76_9226));
   INV_X1 i_257_76_9243 (.A(n_257_76_9226), .ZN(n_257_76_9227));
   NAND2_X1 i_257_76_9244 (.A1(n_257_76_9222), .A2(n_257_76_9227), .ZN(
      n_257_76_9228));
   INV_X1 i_257_76_9245 (.A(n_257_76_9228), .ZN(n_257_76_9229));
   NAND3_X1 i_257_76_9246 (.A1(n_257_76_9220), .A2(n_257_76_9221), .A3(
      n_257_76_9229), .ZN(n_257_76_9230));
   INV_X1 i_257_76_9247 (.A(n_257_76_9230), .ZN(n_257_76_9231));
   NAND2_X1 i_257_76_9248 (.A1(n_257_17), .A2(n_257_76_9231), .ZN(n_257_76_9232));
   NAND2_X1 i_257_76_9249 (.A1(n_257_446), .A2(n_257_845), .ZN(n_257_76_9233));
   NAND2_X1 i_257_76_9250 (.A1(n_257_449), .A2(n_257_1089), .ZN(n_257_76_9234));
   NAND2_X1 i_257_76_9251 (.A1(n_257_447), .A2(n_257_781), .ZN(n_257_76_9235));
   NAND3_X1 i_257_76_9252 (.A1(n_257_76_9233), .A2(n_257_76_9234), .A3(
      n_257_76_9235), .ZN(n_257_76_9236));
   INV_X1 i_257_76_9253 (.A(n_257_76_9236), .ZN(n_257_76_9237));
   NAND2_X1 i_257_76_9254 (.A1(n_257_51), .A2(n_257_433), .ZN(n_257_76_9238));
   NAND3_X1 i_257_76_9255 (.A1(n_257_432), .A2(n_257_613), .A3(n_257_442), 
      .ZN(n_257_76_9239));
   NOR2_X1 i_257_76_9256 (.A1(n_257_1075), .A2(n_257_76_9239), .ZN(n_257_76_9240));
   NAND2_X1 i_257_76_9257 (.A1(n_257_717), .A2(n_257_435), .ZN(n_257_76_9241));
   NAND2_X1 i_257_76_9258 (.A1(n_257_1081), .A2(n_257_438), .ZN(n_257_76_9242));
   NAND2_X1 i_257_76_9259 (.A1(n_257_440), .A2(n_257_947), .ZN(n_257_76_9243));
   NAND4_X1 i_257_76_9260 (.A1(n_257_76_9240), .A2(n_257_76_9241), .A3(
      n_257_76_9242), .A4(n_257_76_9243), .ZN(n_257_76_9244));
   INV_X1 i_257_76_9261 (.A(n_257_76_9244), .ZN(n_257_76_9245));
   NAND3_X1 i_257_76_9262 (.A1(n_257_76_9237), .A2(n_257_76_9238), .A3(
      n_257_76_9245), .ZN(n_257_76_9246));
   NAND2_X1 i_257_76_9263 (.A1(n_257_451), .A2(n_257_468), .ZN(n_257_76_9247));
   NAND2_X1 i_257_76_9264 (.A1(n_257_645), .A2(n_257_450), .ZN(n_257_76_9248));
   NAND3_X1 i_257_76_9265 (.A1(n_257_76_9247), .A2(n_257_76_9248), .A3(
      n_257_76_9222), .ZN(n_257_76_9249));
   NOR2_X1 i_257_76_9266 (.A1(n_257_76_9246), .A2(n_257_76_9249), .ZN(
      n_257_76_9250));
   NAND2_X1 i_257_76_9267 (.A1(n_257_685), .A2(n_257_448), .ZN(n_257_76_9251));
   NAND2_X1 i_257_76_9268 (.A1(n_257_749), .A2(n_257_436), .ZN(n_257_76_9252));
   NAND2_X1 i_257_76_9269 (.A1(n_257_813), .A2(n_257_437), .ZN(n_257_76_9253));
   NAND2_X1 i_257_76_9270 (.A1(n_257_877), .A2(n_257_445), .ZN(n_257_76_9254));
   NAND2_X1 i_257_76_9271 (.A1(n_257_915), .A2(n_257_439), .ZN(n_257_76_9255));
   NAND3_X1 i_257_76_9272 (.A1(n_257_76_9253), .A2(n_257_76_9254), .A3(
      n_257_76_9255), .ZN(n_257_76_9256));
   INV_X1 i_257_76_9273 (.A(n_257_76_9256), .ZN(n_257_76_9257));
   NAND4_X1 i_257_76_9274 (.A1(n_257_76_9250), .A2(n_257_76_9251), .A3(
      n_257_76_9252), .A4(n_257_76_9257), .ZN(n_257_76_9258));
   INV_X1 i_257_76_9275 (.A(n_257_76_9258), .ZN(n_257_76_9259));
   NAND3_X1 i_257_76_9276 (.A1(n_257_76_9220), .A2(n_257_76_9259), .A3(
      n_257_76_9221), .ZN(n_257_76_9260));
   INV_X1 i_257_76_9277 (.A(n_257_76_9260), .ZN(n_257_76_9261));
   NAND2_X1 i_257_76_9278 (.A1(n_257_68), .A2(n_257_76_9261), .ZN(n_257_76_9262));
   NOR2_X1 i_257_76_9279 (.A1(n_257_1075), .A2(n_257_76_17927), .ZN(
      n_257_76_9263));
   NAND4_X1 i_257_76_9280 (.A1(n_257_76_9263), .A2(n_257_76_9241), .A3(
      n_257_76_9242), .A4(n_257_76_9243), .ZN(n_257_76_9264));
   NOR2_X1 i_257_76_9281 (.A1(n_257_76_9236), .A2(n_257_76_9264), .ZN(
      n_257_76_9265));
   NAND2_X1 i_257_76_9282 (.A1(n_257_76_9222), .A2(n_257_645), .ZN(n_257_76_9266));
   INV_X1 i_257_76_9283 (.A(n_257_76_9266), .ZN(n_257_76_9267));
   NAND4_X1 i_257_76_9284 (.A1(n_257_76_9265), .A2(n_257_76_9254), .A3(
      n_257_76_9267), .A4(n_257_76_9255), .ZN(n_257_76_9268));
   INV_X1 i_257_76_9285 (.A(n_257_76_9268), .ZN(n_257_76_9269));
   NAND2_X1 i_257_76_9286 (.A1(n_257_76_9252), .A2(n_257_76_9253), .ZN(
      n_257_76_9270));
   INV_X1 i_257_76_9287 (.A(n_257_76_9270), .ZN(n_257_76_9271));
   NAND3_X1 i_257_76_9288 (.A1(n_257_76_9269), .A2(n_257_76_9271), .A3(
      n_257_76_9251), .ZN(n_257_76_9272));
   INV_X1 i_257_76_9289 (.A(n_257_76_9272), .ZN(n_257_76_9273));
   NAND3_X1 i_257_76_9290 (.A1(n_257_76_9220), .A2(n_257_76_9273), .A3(
      n_257_76_9221), .ZN(n_257_76_9274));
   INV_X1 i_257_76_9291 (.A(n_257_76_9274), .ZN(n_257_76_9275));
   NAND2_X1 i_257_76_9292 (.A1(n_257_28), .A2(n_257_76_9275), .ZN(n_257_76_9276));
   NAND3_X1 i_257_76_9293 (.A1(n_257_76_9232), .A2(n_257_76_9262), .A3(
      n_257_76_9276), .ZN(n_257_76_9277));
   NOR2_X1 i_257_76_9294 (.A1(n_257_1075), .A2(n_257_76_17412), .ZN(
      n_257_76_9278));
   NAND3_X1 i_257_76_9295 (.A1(n_257_76_9278), .A2(n_257_76_9243), .A3(n_257_439), 
      .ZN(n_257_76_9279));
   INV_X1 i_257_76_9296 (.A(n_257_76_9279), .ZN(n_257_76_9280));
   NAND3_X1 i_257_76_9297 (.A1(n_257_76_9280), .A2(n_257_76_9222), .A3(n_257_915), 
      .ZN(n_257_76_9281));
   INV_X1 i_257_76_9298 (.A(n_257_76_9281), .ZN(n_257_76_9282));
   NAND3_X1 i_257_76_9299 (.A1(n_257_76_9220), .A2(n_257_76_9221), .A3(
      n_257_76_9282), .ZN(n_257_76_9283));
   INV_X1 i_257_76_9300 (.A(n_257_76_9283), .ZN(n_257_76_9284));
   NAND2_X1 i_257_76_9301 (.A1(n_257_76_18084), .A2(n_257_76_9284), .ZN(
      n_257_76_9285));
   NAND2_X1 i_257_76_9302 (.A1(n_257_845), .A2(n_257_442), .ZN(n_257_76_9286));
   NOR2_X1 i_257_76_9303 (.A1(n_257_1075), .A2(n_257_76_9286), .ZN(n_257_76_9287));
   NAND4_X1 i_257_76_9304 (.A1(n_257_76_9287), .A2(n_257_446), .A3(n_257_76_9242), 
      .A4(n_257_76_9243), .ZN(n_257_76_9288));
   INV_X1 i_257_76_9305 (.A(n_257_76_9288), .ZN(n_257_76_9289));
   NAND3_X1 i_257_76_9306 (.A1(n_257_76_9255), .A2(n_257_76_9289), .A3(
      n_257_76_9222), .ZN(n_257_76_9290));
   INV_X1 i_257_76_9307 (.A(n_257_76_9254), .ZN(n_257_76_9291));
   NOR2_X1 i_257_76_9308 (.A1(n_257_76_9290), .A2(n_257_76_9291), .ZN(
      n_257_76_9292));
   NAND3_X1 i_257_76_9309 (.A1(n_257_76_9220), .A2(n_257_76_9221), .A3(
      n_257_76_9292), .ZN(n_257_76_9293));
   INV_X1 i_257_76_9310 (.A(n_257_76_9293), .ZN(n_257_76_9294));
   NAND2_X1 i_257_76_9311 (.A1(n_257_76_18070), .A2(n_257_76_9294), .ZN(
      n_257_76_9295));
   INV_X1 i_257_76_9312 (.A(n_257_76_18031), .ZN(n_257_76_9296));
   NAND2_X1 i_257_76_9313 (.A1(n_257_432), .A2(n_257_613), .ZN(n_257_76_9297));
   NAND2_X1 i_257_76_9314 (.A1(n_257_76_9297), .A2(n_257_423), .ZN(n_257_76_9298));
   NOR2_X1 i_257_76_9315 (.A1(n_257_76_9296), .A2(n_257_76_9298), .ZN(
      n_257_76_9299));
   NAND3_X1 i_257_76_9316 (.A1(n_257_76_9299), .A2(n_257_76_9243), .A3(
      n_257_76_9223), .ZN(n_257_76_9300));
   NAND2_X1 i_257_76_9317 (.A1(n_257_208), .A2(n_257_427), .ZN(n_257_76_9301));
   NAND3_X1 i_257_76_9318 (.A1(n_257_76_9241), .A2(n_257_76_9301), .A3(
      n_257_76_9242), .ZN(n_257_76_9302));
   NOR2_X1 i_257_76_9319 (.A1(n_257_76_9300), .A2(n_257_76_9302), .ZN(
      n_257_76_9303));
   NAND2_X1 i_257_76_9320 (.A1(n_257_76_9237), .A2(n_257_76_9303), .ZN(
      n_257_76_9304));
   NAND2_X1 i_257_76_9321 (.A1(n_257_517), .A2(n_257_424), .ZN(n_257_76_9305));
   NAND4_X1 i_257_76_9322 (.A1(n_257_76_9222), .A2(n_257_76_9238), .A3(
      n_257_76_9305), .A4(n_257_288), .ZN(n_257_76_9306));
   NOR2_X1 i_257_76_9323 (.A1(n_257_76_9304), .A2(n_257_76_9306), .ZN(
      n_257_76_9307));
   NAND2_X1 i_257_76_9324 (.A1(n_257_549), .A2(n_257_426), .ZN(n_257_76_9308));
   NAND2_X1 i_257_76_9325 (.A1(n_257_129), .A2(n_257_430), .ZN(n_257_76_9309));
   NAND4_X1 i_257_76_9326 (.A1(n_257_76_9308), .A2(n_257_76_9309), .A3(
      n_257_76_9255), .A4(n_257_76_9248), .ZN(n_257_76_9310));
   INV_X1 i_257_76_9327 (.A(n_257_76_9310), .ZN(n_257_76_9311));
   NAND2_X1 i_257_76_9328 (.A1(n_257_76_9253), .A2(n_257_76_9254), .ZN(
      n_257_76_9312));
   INV_X1 i_257_76_9329 (.A(n_257_76_9312), .ZN(n_257_76_9313));
   NAND3_X1 i_257_76_9330 (.A1(n_257_76_9307), .A2(n_257_76_9311), .A3(
      n_257_76_9313), .ZN(n_257_76_9314));
   INV_X1 i_257_76_9331 (.A(n_257_76_9314), .ZN(n_257_76_9315));
   NAND2_X1 i_257_76_9332 (.A1(n_257_168), .A2(n_257_429), .ZN(n_257_76_9316));
   NAND2_X1 i_257_76_9333 (.A1(n_257_91), .A2(n_257_431), .ZN(n_257_76_9317));
   NAND4_X1 i_257_76_9334 (.A1(n_257_76_9316), .A2(n_257_76_9252), .A3(
      n_257_76_9317), .A4(n_257_76_9247), .ZN(n_257_76_9318));
   NAND2_X1 i_257_76_9335 (.A1(n_257_248), .A2(n_257_425), .ZN(n_257_76_9319));
   NAND2_X1 i_257_76_9336 (.A1(n_257_76_9251), .A2(n_257_76_9319), .ZN(
      n_257_76_9320));
   NOR2_X1 i_257_76_9337 (.A1(n_257_76_9318), .A2(n_257_76_9320), .ZN(
      n_257_76_9321));
   NAND4_X1 i_257_76_9338 (.A1(n_257_76_9220), .A2(n_257_76_9315), .A3(
      n_257_76_9221), .A4(n_257_76_9321), .ZN(n_257_76_9322));
   INV_X1 i_257_76_9339 (.A(n_257_76_9322), .ZN(n_257_76_9323));
   NAND2_X1 i_257_76_9340 (.A1(n_257_76_18066), .A2(n_257_76_9323), .ZN(
      n_257_76_9324));
   NAND3_X1 i_257_76_9341 (.A1(n_257_76_9285), .A2(n_257_76_9295), .A3(
      n_257_76_9324), .ZN(n_257_76_9325));
   NOR2_X1 i_257_76_9342 (.A1(n_257_76_9277), .A2(n_257_76_9325), .ZN(
      n_257_76_9326));
   NAND3_X1 i_257_76_9343 (.A1(n_257_441), .A2(n_257_979), .A3(n_257_76_9278), 
      .ZN(n_257_76_9327));
   INV_X1 i_257_76_9344 (.A(n_257_76_9327), .ZN(n_257_76_9328));
   NAND3_X1 i_257_76_9345 (.A1(n_257_76_9220), .A2(n_257_76_9221), .A3(
      n_257_76_9328), .ZN(n_257_76_9329));
   INV_X1 i_257_76_9346 (.A(n_257_76_9329), .ZN(n_257_76_9330));
   NAND2_X1 i_257_76_9347 (.A1(n_257_76_18071), .A2(n_257_76_9330), .ZN(
      n_257_76_9331));
   NAND2_X1 i_257_76_9348 (.A1(n_257_76_9242), .A2(n_257_76_9243), .ZN(
      n_257_76_9332));
   NAND3_X1 i_257_76_9349 (.A1(n_257_76_9223), .A2(n_257_717), .A3(
      n_257_76_15655), .ZN(n_257_76_9333));
   NOR2_X1 i_257_76_9350 (.A1(n_257_76_9332), .A2(n_257_76_9333), .ZN(
      n_257_76_9334));
   NAND2_X1 i_257_76_9351 (.A1(n_257_76_9233), .A2(n_257_76_9235), .ZN(
      n_257_76_9335));
   INV_X1 i_257_76_9352 (.A(n_257_76_9335), .ZN(n_257_76_9336));
   NAND4_X1 i_257_76_9353 (.A1(n_257_76_9255), .A2(n_257_76_9334), .A3(
      n_257_76_9336), .A4(n_257_76_9222), .ZN(n_257_76_9337));
   INV_X1 i_257_76_9354 (.A(n_257_76_9337), .ZN(n_257_76_9338));
   NAND3_X1 i_257_76_9355 (.A1(n_257_76_9313), .A2(n_257_76_9338), .A3(
      n_257_76_9252), .ZN(n_257_76_9339));
   INV_X1 i_257_76_9356 (.A(n_257_76_9339), .ZN(n_257_76_9340));
   NAND3_X1 i_257_76_9357 (.A1(n_257_76_9220), .A2(n_257_76_9221), .A3(
      n_257_76_9340), .ZN(n_257_76_9341));
   INV_X1 i_257_76_9358 (.A(n_257_76_9341), .ZN(n_257_76_9342));
   NAND2_X1 i_257_76_9359 (.A1(n_257_76_18078), .A2(n_257_76_9342), .ZN(
      n_257_76_9343));
   NAND2_X1 i_257_76_9360 (.A1(n_257_76_9241), .A2(n_257_76_9242), .ZN(
      n_257_76_9344));
   INV_X1 i_257_76_9361 (.A(n_257_76_9344), .ZN(n_257_76_9345));
   INV_X1 i_257_76_9362 (.A(n_257_76_9297), .ZN(n_257_76_9346));
   NAND3_X1 i_257_76_9363 (.A1(n_257_581), .A2(n_257_428), .A3(n_257_442), 
      .ZN(n_257_76_9347));
   NOR2_X1 i_257_76_9364 (.A1(n_257_76_9346), .A2(n_257_76_9347), .ZN(
      n_257_76_9348));
   NAND3_X1 i_257_76_9365 (.A1(n_257_76_9243), .A2(n_257_76_9223), .A3(
      n_257_76_9348), .ZN(n_257_76_9349));
   INV_X1 i_257_76_9366 (.A(n_257_76_9349), .ZN(n_257_76_9350));
   NAND4_X1 i_257_76_9367 (.A1(n_257_76_9345), .A2(n_257_76_9350), .A3(
      n_257_76_9234), .A4(n_257_76_9235), .ZN(n_257_76_9351));
   NAND3_X1 i_257_76_9368 (.A1(n_257_76_9222), .A2(n_257_76_9238), .A3(
      n_257_76_9233), .ZN(n_257_76_9352));
   NOR2_X1 i_257_76_9369 (.A1(n_257_76_9351), .A2(n_257_76_9352), .ZN(
      n_257_76_9353));
   NAND4_X1 i_257_76_9370 (.A1(n_257_76_9309), .A2(n_257_76_9255), .A3(
      n_257_76_9247), .A4(n_257_76_9248), .ZN(n_257_76_9354));
   INV_X1 i_257_76_9371 (.A(n_257_76_9354), .ZN(n_257_76_9355));
   NAND4_X1 i_257_76_9372 (.A1(n_257_76_9313), .A2(n_257_76_9353), .A3(
      n_257_76_9355), .A4(n_257_76_9317), .ZN(n_257_76_9356));
   NAND3_X1 i_257_76_9373 (.A1(n_257_76_9251), .A2(n_257_76_9316), .A3(
      n_257_76_9252), .ZN(n_257_76_9357));
   NOR2_X1 i_257_76_9374 (.A1(n_257_76_9356), .A2(n_257_76_9357), .ZN(
      n_257_76_9358));
   NAND3_X1 i_257_76_9375 (.A1(n_257_76_9358), .A2(n_257_76_9220), .A3(
      n_257_76_9221), .ZN(n_257_76_9359));
   INV_X1 i_257_76_9376 (.A(n_257_76_9359), .ZN(n_257_76_9360));
   NAND2_X1 i_257_76_9377 (.A1(n_257_76_18074), .A2(n_257_76_9360), .ZN(
      n_257_76_9361));
   NAND3_X1 i_257_76_9378 (.A1(n_257_76_9331), .A2(n_257_76_9343), .A3(
      n_257_76_9361), .ZN(n_257_76_9362));
   NAND2_X1 i_257_76_9379 (.A1(n_257_1075), .A2(n_257_442), .ZN(n_257_76_9363));
   INV_X1 i_257_76_9380 (.A(n_257_76_9363), .ZN(n_257_76_9364));
   NAND2_X1 i_257_76_9381 (.A1(n_257_13), .A2(n_257_76_9364), .ZN(n_257_76_9365));
   NOR2_X1 i_257_76_9382 (.A1(n_257_1075), .A2(n_257_76_17902), .ZN(
      n_257_76_9366));
   NAND3_X1 i_257_76_9383 (.A1(n_257_76_9366), .A2(n_257_76_9242), .A3(
      n_257_76_9243), .ZN(n_257_76_9367));
   INV_X1 i_257_76_9384 (.A(n_257_76_9367), .ZN(n_257_76_9368));
   NAND4_X1 i_257_76_9385 (.A1(n_257_76_9255), .A2(n_257_877), .A3(n_257_76_9368), 
      .A4(n_257_76_9222), .ZN(n_257_76_9369));
   INV_X1 i_257_76_9386 (.A(n_257_76_9369), .ZN(n_257_76_9370));
   NAND3_X1 i_257_76_9387 (.A1(n_257_76_9220), .A2(n_257_76_9221), .A3(
      n_257_76_9370), .ZN(n_257_76_9371));
   INV_X1 i_257_76_9388 (.A(n_257_76_9371), .ZN(n_257_76_9372));
   NAND2_X1 i_257_76_9389 (.A1(n_257_76_18077), .A2(n_257_76_9372), .ZN(
      n_257_76_9373));
   NAND2_X1 i_257_76_9390 (.A1(n_257_76_9365), .A2(n_257_76_9373), .ZN(
      n_257_76_9374));
   NOR2_X1 i_257_76_9391 (.A1(n_257_76_9362), .A2(n_257_76_9374), .ZN(
      n_257_76_9375));
   NAND3_X1 i_257_76_9392 (.A1(n_257_76_9253), .A2(n_257_749), .A3(n_257_76_9254), 
      .ZN(n_257_76_9376));
   NOR2_X1 i_257_76_9393 (.A1(n_257_1075), .A2(n_257_76_17934), .ZN(
      n_257_76_9377));
   NAND3_X1 i_257_76_9394 (.A1(n_257_76_9377), .A2(n_257_76_9242), .A3(
      n_257_76_9243), .ZN(n_257_76_9378));
   INV_X1 i_257_76_9395 (.A(n_257_76_9378), .ZN(n_257_76_9379));
   NAND4_X1 i_257_76_9396 (.A1(n_257_76_9255), .A2(n_257_76_9336), .A3(
      n_257_76_9379), .A4(n_257_76_9222), .ZN(n_257_76_9380));
   NOR2_X1 i_257_76_9397 (.A1(n_257_76_9376), .A2(n_257_76_9380), .ZN(
      n_257_76_9381));
   NAND3_X1 i_257_76_9398 (.A1(n_257_76_9220), .A2(n_257_76_9221), .A3(
      n_257_76_9381), .ZN(n_257_76_9382));
   INV_X1 i_257_76_9399 (.A(n_257_76_9382), .ZN(n_257_76_9383));
   NAND2_X1 i_257_76_9400 (.A1(n_257_76_18069), .A2(n_257_76_9383), .ZN(
      n_257_76_9384));
   NAND2_X1 i_257_76_9401 (.A1(n_257_76_9297), .A2(n_257_426), .ZN(n_257_76_9385));
   NOR2_X1 i_257_76_9402 (.A1(n_257_76_9296), .A2(n_257_76_9385), .ZN(
      n_257_76_9386));
   NAND3_X1 i_257_76_9403 (.A1(n_257_76_9386), .A2(n_257_76_9243), .A3(
      n_257_76_9223), .ZN(n_257_76_9387));
   INV_X1 i_257_76_9404 (.A(n_257_76_9387), .ZN(n_257_76_9388));
   INV_X1 i_257_76_9405 (.A(n_257_76_9302), .ZN(n_257_76_9389));
   NAND4_X1 i_257_76_9406 (.A1(n_257_76_9388), .A2(n_257_76_9389), .A3(
      n_257_76_9234), .A4(n_257_76_9235), .ZN(n_257_76_9390));
   NOR2_X1 i_257_76_9407 (.A1(n_257_76_9390), .A2(n_257_76_9352), .ZN(
      n_257_76_9391));
   NAND4_X1 i_257_76_9408 (.A1(n_257_76_9309), .A2(n_257_76_9255), .A3(
      n_257_76_9248), .A4(n_257_549), .ZN(n_257_76_9392));
   INV_X1 i_257_76_9409 (.A(n_257_76_9392), .ZN(n_257_76_9393));
   NAND3_X1 i_257_76_9410 (.A1(n_257_76_9391), .A2(n_257_76_9313), .A3(
      n_257_76_9393), .ZN(n_257_76_9394));
   INV_X1 i_257_76_9411 (.A(n_257_76_9394), .ZN(n_257_76_9395));
   NAND3_X1 i_257_76_9412 (.A1(n_257_76_9252), .A2(n_257_76_9317), .A3(
      n_257_76_9247), .ZN(n_257_76_9396));
   INV_X1 i_257_76_9413 (.A(n_257_76_9396), .ZN(n_257_76_9397));
   NAND3_X1 i_257_76_9414 (.A1(n_257_76_9397), .A2(n_257_76_9251), .A3(
      n_257_76_9316), .ZN(n_257_76_9398));
   INV_X1 i_257_76_9415 (.A(n_257_76_9398), .ZN(n_257_76_9399));
   NAND4_X1 i_257_76_9416 (.A1(n_257_76_9220), .A2(n_257_76_9395), .A3(
      n_257_76_9221), .A4(n_257_76_9399), .ZN(n_257_76_9400));
   INV_X1 i_257_76_9417 (.A(n_257_76_9400), .ZN(n_257_76_9401));
   NAND2_X1 i_257_76_9418 (.A1(n_257_76_18076), .A2(n_257_76_9401), .ZN(
      n_257_76_9402));
   INV_X1 i_257_76_9419 (.A(n_257_76_9278), .ZN(n_257_76_9403));
   NOR2_X1 i_257_76_9420 (.A1(n_257_76_9403), .A2(n_257_76_15197), .ZN(
      n_257_76_9404));
   NAND2_X1 i_257_76_9421 (.A1(n_257_1043), .A2(n_257_76_9404), .ZN(
      n_257_76_9405));
   INV_X1 i_257_76_9422 (.A(n_257_76_9405), .ZN(n_257_76_9406));
   NAND2_X1 i_257_76_9423 (.A1(n_257_76_18072), .A2(n_257_76_9406), .ZN(
      n_257_76_9407));
   NAND3_X1 i_257_76_9424 (.A1(n_257_76_9384), .A2(n_257_76_9402), .A3(
      n_257_76_9407), .ZN(n_257_76_9408));
   NOR2_X1 i_257_76_9425 (.A1(n_257_1075), .A2(n_257_76_17951), .ZN(
      n_257_76_9409));
   NAND3_X1 i_257_76_9426 (.A1(n_257_76_9409), .A2(n_257_76_9242), .A3(
      n_257_76_9243), .ZN(n_257_76_9410));
   INV_X1 i_257_76_9427 (.A(n_257_76_9233), .ZN(n_257_76_9411));
   NOR2_X1 i_257_76_9428 (.A1(n_257_76_9410), .A2(n_257_76_9411), .ZN(
      n_257_76_9412));
   NAND3_X1 i_257_76_9429 (.A1(n_257_76_9412), .A2(n_257_813), .A3(n_257_76_9222), 
      .ZN(n_257_76_9413));
   NAND2_X1 i_257_76_9430 (.A1(n_257_76_9254), .A2(n_257_76_9255), .ZN(
      n_257_76_9414));
   NOR2_X1 i_257_76_9431 (.A1(n_257_76_9413), .A2(n_257_76_9414), .ZN(
      n_257_76_9415));
   NAND3_X1 i_257_76_9432 (.A1(n_257_76_9220), .A2(n_257_76_9221), .A3(
      n_257_76_9415), .ZN(n_257_76_9416));
   INV_X1 i_257_76_9433 (.A(n_257_76_9416), .ZN(n_257_76_9417));
   NAND2_X1 i_257_76_9434 (.A1(n_257_22), .A2(n_257_76_9417), .ZN(n_257_76_9418));
   NAND2_X1 i_257_76_9435 (.A1(n_257_444), .A2(n_257_76_9278), .ZN(n_257_76_9419));
   INV_X1 i_257_76_9436 (.A(n_257_76_9419), .ZN(n_257_76_9420));
   NAND3_X1 i_257_76_9437 (.A1(n_257_76_9221), .A2(n_257_1011), .A3(
      n_257_76_9420), .ZN(n_257_76_9421));
   INV_X1 i_257_76_9438 (.A(n_257_76_9421), .ZN(n_257_76_9422));
   NAND2_X1 i_257_76_9439 (.A1(n_257_76_18075), .A2(n_257_76_9422), .ZN(
      n_257_76_9423));
   NAND2_X1 i_257_76_9440 (.A1(n_257_76_9418), .A2(n_257_76_9423), .ZN(
      n_257_76_9424));
   NOR2_X1 i_257_76_9441 (.A1(n_257_76_9408), .A2(n_257_76_9424), .ZN(
      n_257_76_9425));
   NAND3_X1 i_257_76_9442 (.A1(n_257_76_9326), .A2(n_257_76_9375), .A3(
      n_257_76_9425), .ZN(n_257_76_9426));
   INV_X1 i_257_76_9443 (.A(n_257_76_9426), .ZN(n_257_76_9427));
   NOR2_X1 i_257_76_9444 (.A1(n_257_1075), .A2(n_257_76_17633), .ZN(
      n_257_76_9428));
   NAND4_X1 i_257_76_9445 (.A1(n_257_76_9428), .A2(n_257_76_9241), .A3(
      n_257_76_9242), .A4(n_257_76_9243), .ZN(n_257_76_9429));
   INV_X1 i_257_76_9446 (.A(n_257_76_9429), .ZN(n_257_76_9430));
   NAND2_X1 i_257_76_9447 (.A1(n_257_76_9233), .A2(n_257_76_9234), .ZN(
      n_257_76_9431));
   INV_X1 i_257_76_9448 (.A(n_257_76_9431), .ZN(n_257_76_9432));
   NAND2_X1 i_257_76_9449 (.A1(n_257_76_9235), .A2(n_257_51), .ZN(n_257_76_9433));
   INV_X1 i_257_76_9450 (.A(n_257_76_9433), .ZN(n_257_76_9434));
   NAND3_X1 i_257_76_9451 (.A1(n_257_76_9430), .A2(n_257_76_9432), .A3(
      n_257_76_9434), .ZN(n_257_76_9435));
   NOR2_X1 i_257_76_9452 (.A1(n_257_76_9435), .A2(n_257_76_9249), .ZN(
      n_257_76_9436));
   NAND4_X1 i_257_76_9453 (.A1(n_257_76_9436), .A2(n_257_76_9251), .A3(
      n_257_76_9252), .A4(n_257_76_9257), .ZN(n_257_76_9437));
   INV_X1 i_257_76_9454 (.A(n_257_76_9437), .ZN(n_257_76_9438));
   NAND3_X1 i_257_76_9455 (.A1(n_257_76_9220), .A2(n_257_76_9438), .A3(
      n_257_76_9221), .ZN(n_257_76_9439));
   INV_X1 i_257_76_9456 (.A(n_257_76_9439), .ZN(n_257_76_9440));
   NAND2_X1 i_257_76_9457 (.A1(n_257_76_18081), .A2(n_257_76_9440), .ZN(
      n_257_76_9441));
   NAND3_X1 i_257_76_9458 (.A1(n_257_76_9243), .A2(n_257_76_18032), .A3(
      n_257_76_9223), .ZN(n_257_76_9442));
   NOR2_X1 i_257_76_9459 (.A1(n_257_76_9344), .A2(n_257_76_9442), .ZN(
      n_257_76_9443));
   NAND4_X1 i_257_76_9460 (.A1(n_257_76_9443), .A2(n_257_76_9237), .A3(
      n_257_76_9222), .A4(n_257_76_9238), .ZN(n_257_76_9444));
   NAND3_X1 i_257_76_9461 (.A1(n_257_76_9255), .A2(n_257_76_9247), .A3(
      n_257_76_9248), .ZN(n_257_76_9445));
   NOR2_X1 i_257_76_9462 (.A1(n_257_76_9444), .A2(n_257_76_9445), .ZN(
      n_257_76_9446));
   NAND3_X1 i_257_76_9463 (.A1(n_257_76_9253), .A2(n_257_91), .A3(n_257_76_9254), 
      .ZN(n_257_76_9447));
   INV_X1 i_257_76_9464 (.A(n_257_76_9447), .ZN(n_257_76_9448));
   NAND4_X1 i_257_76_9465 (.A1(n_257_76_9446), .A2(n_257_76_9251), .A3(
      n_257_76_9252), .A4(n_257_76_9448), .ZN(n_257_76_9449));
   INV_X1 i_257_76_9466 (.A(n_257_76_9449), .ZN(n_257_76_9450));
   NAND3_X1 i_257_76_9467 (.A1(n_257_76_9450), .A2(n_257_76_9220), .A3(
      n_257_76_9221), .ZN(n_257_76_9451));
   INV_X1 i_257_76_9468 (.A(n_257_76_9451), .ZN(n_257_76_9452));
   NAND2_X1 i_257_76_9469 (.A1(n_257_76_18080), .A2(n_257_76_9452), .ZN(
      n_257_76_9453));
   NAND3_X1 i_257_76_9470 (.A1(n_257_76_18033), .A2(n_257_76_9243), .A3(
      n_257_76_9223), .ZN(n_257_76_9454));
   NOR2_X1 i_257_76_9471 (.A1(n_257_76_9454), .A2(n_257_76_9344), .ZN(
      n_257_76_9455));
   NAND4_X1 i_257_76_9472 (.A1(n_257_76_9237), .A2(n_257_76_9455), .A3(
      n_257_76_9222), .A4(n_257_76_9238), .ZN(n_257_76_9456));
   NOR2_X1 i_257_76_9473 (.A1(n_257_76_9456), .A2(n_257_76_9445), .ZN(
      n_257_76_9457));
   NAND3_X1 i_257_76_9474 (.A1(n_257_76_9253), .A2(n_257_76_9254), .A3(
      n_257_76_9309), .ZN(n_257_76_9458));
   INV_X1 i_257_76_9475 (.A(n_257_168), .ZN(n_257_76_9459));
   NOR2_X1 i_257_76_9476 (.A1(n_257_76_9458), .A2(n_257_76_9459), .ZN(
      n_257_76_9460));
   NAND2_X1 i_257_76_9477 (.A1(n_257_76_9252), .A2(n_257_76_9317), .ZN(
      n_257_76_9461));
   INV_X1 i_257_76_9478 (.A(n_257_76_9461), .ZN(n_257_76_9462));
   NAND4_X1 i_257_76_9479 (.A1(n_257_76_9457), .A2(n_257_76_9460), .A3(
      n_257_76_9462), .A4(n_257_76_9251), .ZN(n_257_76_9463));
   INV_X1 i_257_76_9480 (.A(n_257_76_9463), .ZN(n_257_76_9464));
   NAND3_X1 i_257_76_9481 (.A1(n_257_76_9464), .A2(n_257_76_9220), .A3(
      n_257_76_9221), .ZN(n_257_76_9465));
   INV_X1 i_257_76_9482 (.A(n_257_76_9465), .ZN(n_257_76_9466));
   NAND2_X1 i_257_76_9483 (.A1(n_257_76_18061), .A2(n_257_76_9466), .ZN(
      n_257_76_9467));
   NAND3_X1 i_257_76_9484 (.A1(n_257_76_9441), .A2(n_257_76_9453), .A3(
      n_257_76_9467), .ZN(n_257_76_9468));
   INV_X1 i_257_76_9485 (.A(n_257_76_9468), .ZN(n_257_76_9469));
   INV_X1 i_257_76_9486 (.A(n_257_76_9242), .ZN(n_257_76_9470));
   NAND3_X1 i_257_76_9487 (.A1(n_257_76_9278), .A2(n_257_76_9470), .A3(
      n_257_76_9243), .ZN(n_257_76_9471));
   INV_X1 i_257_76_9488 (.A(n_257_76_9471), .ZN(n_257_76_9472));
   NAND3_X1 i_257_76_9489 (.A1(n_257_76_9255), .A2(n_257_76_9222), .A3(
      n_257_76_9472), .ZN(n_257_76_9473));
   INV_X1 i_257_76_9490 (.A(n_257_76_9473), .ZN(n_257_76_9474));
   NAND3_X1 i_257_76_9491 (.A1(n_257_76_9220), .A2(n_257_76_9221), .A3(
      n_257_76_9474), .ZN(n_257_76_9475));
   INV_X1 i_257_76_9492 (.A(n_257_76_9475), .ZN(n_257_76_9476));
   NAND2_X1 i_257_76_9493 (.A1(n_257_76_18067), .A2(n_257_76_9476), .ZN(
      n_257_76_9477));
   NAND2_X1 i_257_76_9494 (.A1(n_257_76_9222), .A2(n_257_76_9238), .ZN(
      n_257_76_9478));
   INV_X1 i_257_76_9495 (.A(n_257_76_9478), .ZN(n_257_76_9479));
   INV_X1 i_257_76_9496 (.A(n_257_76_9305), .ZN(n_257_76_9480));
   NOR2_X1 i_257_76_9497 (.A1(n_257_76_9431), .A2(n_257_76_9480), .ZN(
      n_257_76_9481));
   NAND2_X1 i_257_76_9498 (.A1(n_257_76_9479), .A2(n_257_76_9481), .ZN(
      n_257_76_9482));
   NAND2_X1 i_257_76_9499 (.A1(n_257_326), .A2(n_257_422), .ZN(n_257_76_9483));
   NAND2_X1 i_257_76_9500 (.A1(n_257_76_9235), .A2(n_257_76_9483), .ZN(
      n_257_76_9484));
   NAND2_X1 i_257_76_9501 (.A1(n_257_76_9241), .A2(n_257_76_9301), .ZN(
      n_257_76_9485));
   NOR2_X1 i_257_76_9502 (.A1(n_257_76_9484), .A2(n_257_76_9485), .ZN(
      n_257_76_9486));
   NAND2_X1 i_257_76_9503 (.A1(n_257_442), .A2(n_257_485), .ZN(n_257_76_9487));
   INV_X1 i_257_76_9504 (.A(n_257_76_18034), .ZN(n_257_76_9488));
   NOR2_X1 i_257_76_9505 (.A1(n_257_76_9488), .A2(n_257_1075), .ZN(n_257_76_9489));
   NAND2_X1 i_257_76_9506 (.A1(n_257_420), .A2(n_257_76_9297), .ZN(n_257_76_9490));
   INV_X1 i_257_76_9507 (.A(n_257_76_9490), .ZN(n_257_76_9491));
   NAND2_X1 i_257_76_9508 (.A1(n_257_76_9489), .A2(n_257_76_9491), .ZN(
      n_257_76_9492));
   NOR2_X1 i_257_76_9509 (.A1(n_257_76_9492), .A2(n_257_76_9332), .ZN(
      n_257_76_9493));
   NAND2_X1 i_257_76_9510 (.A1(n_257_76_9486), .A2(n_257_76_9493), .ZN(
      n_257_76_9494));
   NOR2_X1 i_257_76_9511 (.A1(n_257_76_9482), .A2(n_257_76_9494), .ZN(
      n_257_76_9495));
   NAND2_X1 i_257_76_9512 (.A1(n_257_76_9255), .A2(n_257_76_9247), .ZN(
      n_257_76_9496));
   NAND2_X1 i_257_76_9513 (.A1(n_257_288), .A2(n_257_423), .ZN(n_257_76_9497));
   NAND2_X1 i_257_76_9514 (.A1(n_257_76_9248), .A2(n_257_76_9497), .ZN(
      n_257_76_9498));
   NOR2_X1 i_257_76_9515 (.A1(n_257_76_9496), .A2(n_257_76_9498), .ZN(
      n_257_76_9499));
   NAND2_X1 i_257_76_9516 (.A1(n_257_76_9495), .A2(n_257_76_9499), .ZN(
      n_257_76_9500));
   NAND2_X1 i_257_76_9517 (.A1(n_257_76_9317), .A2(n_257_76_9253), .ZN(
      n_257_76_9501));
   INV_X1 i_257_76_9518 (.A(n_257_76_9501), .ZN(n_257_76_9502));
   NAND2_X1 i_257_76_9519 (.A1(n_257_76_9254), .A2(n_257_76_9308), .ZN(
      n_257_76_9503));
   NAND2_X1 i_257_76_9520 (.A1(n_257_365), .A2(n_257_421), .ZN(n_257_76_9504));
   NAND2_X1 i_257_76_9521 (.A1(n_257_76_9309), .A2(n_257_76_9504), .ZN(
      n_257_76_9505));
   NOR2_X1 i_257_76_9522 (.A1(n_257_76_9503), .A2(n_257_76_9505), .ZN(
      n_257_76_9506));
   NAND2_X1 i_257_76_9523 (.A1(n_257_76_9502), .A2(n_257_76_9506), .ZN(
      n_257_76_9507));
   NOR2_X1 i_257_76_9524 (.A1(n_257_76_9500), .A2(n_257_76_9507), .ZN(
      n_257_76_9508));
   NAND2_X1 i_257_76_9525 (.A1(n_257_76_9316), .A2(n_257_76_9252), .ZN(
      n_257_76_9509));
   NOR2_X1 i_257_76_9526 (.A1(n_257_76_9320), .A2(n_257_76_9509), .ZN(
      n_257_76_9510));
   NAND2_X1 i_257_76_9527 (.A1(n_257_76_9508), .A2(n_257_76_9510), .ZN(
      n_257_76_9511));
   NAND2_X1 i_257_76_9528 (.A1(n_257_76_9220), .A2(n_257_76_9221), .ZN(
      n_257_76_9512));
   NOR2_X1 i_257_76_9529 (.A1(n_257_76_9511), .A2(n_257_76_9512), .ZN(
      n_257_76_9513));
   NAND2_X1 i_257_76_9530 (.A1(n_257_76_18073), .A2(n_257_76_9513), .ZN(
      n_257_76_9514));
   NAND4_X1 i_257_76_9531 (.A1(n_257_76_9248), .A2(n_257_76_9222), .A3(
      n_257_76_9238), .A4(n_257_129), .ZN(n_257_76_9515));
   NAND2_X1 i_257_76_9532 (.A1(n_257_76_9235), .A2(n_257_76_9241), .ZN(
      n_257_76_9516));
   INV_X1 i_257_76_9533 (.A(n_257_76_9516), .ZN(n_257_76_9517));
   NAND4_X1 i_257_76_9534 (.A1(n_257_76_9242), .A2(n_257_76_9243), .A3(
      n_257_76_18035), .A4(n_257_76_9223), .ZN(n_257_76_9518));
   INV_X1 i_257_76_9535 (.A(n_257_76_9518), .ZN(n_257_76_9519));
   NAND3_X1 i_257_76_9536 (.A1(n_257_76_9432), .A2(n_257_76_9517), .A3(
      n_257_76_9519), .ZN(n_257_76_9520));
   NOR2_X1 i_257_76_9537 (.A1(n_257_76_9515), .A2(n_257_76_9520), .ZN(
      n_257_76_9521));
   NAND4_X1 i_257_76_9538 (.A1(n_257_76_9253), .A2(n_257_76_9254), .A3(
      n_257_76_9255), .A4(n_257_76_9247), .ZN(n_257_76_9522));
   INV_X1 i_257_76_9539 (.A(n_257_76_9522), .ZN(n_257_76_9523));
   NAND4_X1 i_257_76_9540 (.A1(n_257_76_9462), .A2(n_257_76_9251), .A3(
      n_257_76_9521), .A4(n_257_76_9523), .ZN(n_257_76_9524));
   INV_X1 i_257_76_9541 (.A(n_257_76_9524), .ZN(n_257_76_9525));
   NAND3_X1 i_257_76_9542 (.A1(n_257_76_9220), .A2(n_257_76_9525), .A3(
      n_257_76_9221), .ZN(n_257_76_9526));
   INV_X1 i_257_76_9543 (.A(n_257_76_9526), .ZN(n_257_76_9527));
   NAND2_X1 i_257_76_9544 (.A1(n_257_76_18068), .A2(n_257_76_9527), .ZN(
      n_257_76_9528));
   NAND3_X1 i_257_76_9545 (.A1(n_257_76_9477), .A2(n_257_76_9514), .A3(
      n_257_76_9528), .ZN(n_257_76_9529));
   INV_X1 i_257_76_9546 (.A(n_257_76_9529), .ZN(n_257_76_9530));
   NAND2_X1 i_257_76_9547 (.A1(n_257_76_9233), .A2(n_257_76_9242), .ZN(
      n_257_76_9531));
   INV_X1 i_257_76_9548 (.A(n_257_76_9531), .ZN(n_257_76_9532));
   NAND2_X1 i_257_76_9549 (.A1(n_257_781), .A2(n_257_442), .ZN(n_257_76_9533));
   NOR2_X1 i_257_76_9550 (.A1(n_257_1075), .A2(n_257_76_9533), .ZN(n_257_76_9534));
   NAND3_X1 i_257_76_9551 (.A1(n_257_76_9534), .A2(n_257_447), .A3(n_257_76_9243), 
      .ZN(n_257_76_9535));
   INV_X1 i_257_76_9552 (.A(n_257_76_9535), .ZN(n_257_76_9536));
   NAND4_X1 i_257_76_9553 (.A1(n_257_76_9255), .A2(n_257_76_9532), .A3(
      n_257_76_9536), .A4(n_257_76_9222), .ZN(n_257_76_9537));
   NOR2_X1 i_257_76_9554 (.A1(n_257_76_9312), .A2(n_257_76_9537), .ZN(
      n_257_76_9538));
   NAND3_X1 i_257_76_9555 (.A1(n_257_76_9220), .A2(n_257_76_9221), .A3(
      n_257_76_9538), .ZN(n_257_76_9539));
   INV_X1 i_257_76_9556 (.A(n_257_76_9539), .ZN(n_257_76_9540));
   NAND3_X1 i_257_76_9557 (.A1(n_257_76_9278), .A2(n_257_76_9241), .A3(n_257_449), 
      .ZN(n_257_76_9541));
   NAND3_X1 i_257_76_9558 (.A1(n_257_76_9242), .A2(n_257_76_9243), .A3(
      n_257_1089), .ZN(n_257_76_9542));
   NOR2_X1 i_257_76_9559 (.A1(n_257_76_9541), .A2(n_257_76_9542), .ZN(
      n_257_76_9543));
   NAND4_X1 i_257_76_9560 (.A1(n_257_76_9543), .A2(n_257_76_9255), .A3(
      n_257_76_9336), .A4(n_257_76_9222), .ZN(n_257_76_9544));
   INV_X1 i_257_76_9561 (.A(n_257_76_9544), .ZN(n_257_76_9545));
   NAND3_X1 i_257_76_9562 (.A1(n_257_76_9545), .A2(n_257_76_9313), .A3(
      n_257_76_9252), .ZN(n_257_76_9546));
   INV_X1 i_257_76_9563 (.A(n_257_76_9251), .ZN(n_257_76_9547));
   NOR2_X1 i_257_76_9564 (.A1(n_257_76_9546), .A2(n_257_76_9547), .ZN(
      n_257_76_9548));
   NAND3_X1 i_257_76_9565 (.A1(n_257_76_9548), .A2(n_257_76_9220), .A3(
      n_257_76_9221), .ZN(n_257_76_9549));
   INV_X1 i_257_76_9566 (.A(n_257_76_9549), .ZN(n_257_76_9550));
   AOI22_X1 i_257_76_9567 (.A1(n_257_76_18085), .A2(n_257_76_9540), .B1(
      n_257_76_18083), .B2(n_257_76_9550), .ZN(n_257_76_9551));
   NAND3_X1 i_257_76_9568 (.A1(n_257_76_9469), .A2(n_257_76_9530), .A3(
      n_257_76_9551), .ZN(n_257_76_9552));
   NAND3_X1 i_257_76_9569 (.A1(n_257_76_9242), .A2(n_257_76_9243), .A3(
      n_257_76_9223), .ZN(n_257_76_9553));
   NOR2_X1 i_257_76_9570 (.A1(n_257_435), .A2(n_257_76_17412), .ZN(n_257_76_9554));
   INV_X1 i_257_76_9571 (.A(n_257_717), .ZN(n_257_76_9555));
   AOI21_X1 i_257_76_9572 (.A(n_257_76_9554), .B1(n_257_76_9555), .B2(n_257_442), 
      .ZN(n_257_76_9556));
   NOR2_X1 i_257_76_9573 (.A1(n_257_76_9553), .A2(n_257_76_9556), .ZN(
      n_257_76_9557));
   NAND2_X1 i_257_76_9574 (.A1(n_257_76_9255), .A2(n_257_76_9557), .ZN(
      n_257_76_9558));
   INV_X1 i_257_76_9575 (.A(n_257_76_9558), .ZN(n_257_76_9559));
   NAND3_X1 i_257_76_9576 (.A1(n_257_76_9233), .A2(n_257_76_9235), .A3(n_257_448), 
      .ZN(n_257_76_9560));
   INV_X1 i_257_76_9577 (.A(n_257_76_9222), .ZN(n_257_76_9561));
   NOR2_X1 i_257_76_9578 (.A1(n_257_76_9560), .A2(n_257_76_9561), .ZN(
      n_257_76_9562));
   NAND4_X1 i_257_76_9579 (.A1(n_257_76_9559), .A2(n_257_76_9562), .A3(
      n_257_76_9253), .A4(n_257_76_9254), .ZN(n_257_76_9563));
   NAND2_X1 i_257_76_9580 (.A1(n_257_685), .A2(n_257_76_9252), .ZN(n_257_76_9564));
   NOR2_X1 i_257_76_9581 (.A1(n_257_76_9563), .A2(n_257_76_9564), .ZN(
      n_257_76_9565));
   NAND3_X1 i_257_76_9582 (.A1(n_257_76_9220), .A2(n_257_76_9221), .A3(
      n_257_76_9565), .ZN(n_257_76_9566));
   INV_X1 i_257_76_9583 (.A(n_257_76_9566), .ZN(n_257_76_9567));
   NAND2_X1 i_257_76_9584 (.A1(n_257_76_18079), .A2(n_257_76_9567), .ZN(
      n_257_76_9568));
   NAND3_X1 i_257_76_9585 (.A1(n_257_76_18031), .A2(n_257_76_9297), .A3(
      n_257_425), .ZN(n_257_76_9569));
   NOR2_X1 i_257_76_9586 (.A1(n_257_76_9569), .A2(n_257_1075), .ZN(n_257_76_9570));
   INV_X1 i_257_76_9587 (.A(n_257_76_9485), .ZN(n_257_76_9571));
   INV_X1 i_257_76_9588 (.A(n_257_76_9332), .ZN(n_257_76_9572));
   NAND3_X1 i_257_76_9589 (.A1(n_257_76_9570), .A2(n_257_76_9571), .A3(
      n_257_76_9572), .ZN(n_257_76_9573));
   NOR2_X1 i_257_76_9590 (.A1(n_257_76_9573), .A2(n_257_76_9236), .ZN(
      n_257_76_9574));
   NAND3_X1 i_257_76_9591 (.A1(n_257_76_9248), .A2(n_257_76_9222), .A3(
      n_257_76_9238), .ZN(n_257_76_9575));
   INV_X1 i_257_76_9592 (.A(n_257_76_9575), .ZN(n_257_76_9576));
   INV_X1 i_257_76_9593 (.A(n_257_76_9496), .ZN(n_257_76_9577));
   NAND3_X1 i_257_76_9594 (.A1(n_257_76_9574), .A2(n_257_76_9576), .A3(
      n_257_76_9577), .ZN(n_257_76_9578));
   NAND4_X1 i_257_76_9595 (.A1(n_257_76_9253), .A2(n_257_76_9254), .A3(
      n_257_76_9308), .A4(n_257_76_9309), .ZN(n_257_76_9579));
   NOR2_X1 i_257_76_9596 (.A1(n_257_76_9578), .A2(n_257_76_9579), .ZN(
      n_257_76_9580));
   NAND3_X1 i_257_76_9597 (.A1(n_257_76_9252), .A2(n_257_76_9317), .A3(n_257_248), 
      .ZN(n_257_76_9581));
   INV_X1 i_257_76_9598 (.A(n_257_76_9581), .ZN(n_257_76_9582));
   NAND4_X1 i_257_76_9599 (.A1(n_257_76_9580), .A2(n_257_76_9582), .A3(
      n_257_76_9251), .A4(n_257_76_9316), .ZN(n_257_76_9583));
   NOR2_X1 i_257_76_9600 (.A1(n_257_76_9583), .A2(n_257_76_9512), .ZN(
      n_257_76_9584));
   NAND2_X1 i_257_76_9601 (.A1(n_257_76_18064), .A2(n_257_76_9584), .ZN(
      n_257_76_9585));
   NAND2_X1 i_257_76_9602 (.A1(n_257_76_9297), .A2(n_257_421), .ZN(n_257_76_9586));
   NOR2_X1 i_257_76_9603 (.A1(n_257_76_9296), .A2(n_257_76_9586), .ZN(
      n_257_76_9587));
   NAND4_X1 i_257_76_9604 (.A1(n_257_76_9587), .A2(n_257_76_9242), .A3(
      n_257_76_9243), .A4(n_257_76_9223), .ZN(n_257_76_9588));
   INV_X1 i_257_76_9605 (.A(n_257_76_9588), .ZN(n_257_76_9589));
   NAND2_X1 i_257_76_9606 (.A1(n_257_76_9234), .A2(n_257_76_9235), .ZN(
      n_257_76_9590));
   INV_X1 i_257_76_9607 (.A(n_257_76_9590), .ZN(n_257_76_9591));
   NAND3_X1 i_257_76_9608 (.A1(n_257_76_9483), .A2(n_257_76_9241), .A3(
      n_257_76_9301), .ZN(n_257_76_9592));
   INV_X1 i_257_76_9609 (.A(n_257_76_9592), .ZN(n_257_76_9593));
   NAND3_X1 i_257_76_9610 (.A1(n_257_76_9589), .A2(n_257_76_9591), .A3(
      n_257_76_9593), .ZN(n_257_76_9594));
   NAND4_X1 i_257_76_9611 (.A1(n_257_76_9238), .A2(n_257_365), .A3(n_257_76_9305), 
      .A4(n_257_76_9233), .ZN(n_257_76_9595));
   NOR2_X1 i_257_76_9612 (.A1(n_257_76_9594), .A2(n_257_76_9595), .ZN(
      n_257_76_9596));
   NAND3_X1 i_257_76_9613 (.A1(n_257_76_9253), .A2(n_257_76_9254), .A3(
      n_257_76_9308), .ZN(n_257_76_9597));
   INV_X1 i_257_76_9614 (.A(n_257_76_9597), .ZN(n_257_76_9598));
   NAND3_X1 i_257_76_9615 (.A1(n_257_76_9248), .A2(n_257_76_9497), .A3(
      n_257_76_9222), .ZN(n_257_76_9599));
   NAND2_X1 i_257_76_9616 (.A1(n_257_76_9309), .A2(n_257_76_9255), .ZN(
      n_257_76_9600));
   NOR2_X1 i_257_76_9617 (.A1(n_257_76_9599), .A2(n_257_76_9600), .ZN(
      n_257_76_9601));
   NAND3_X1 i_257_76_9618 (.A1(n_257_76_9596), .A2(n_257_76_9598), .A3(
      n_257_76_9601), .ZN(n_257_76_9602));
   NOR2_X1 i_257_76_9619 (.A1(n_257_76_9602), .A2(n_257_76_9547), .ZN(
      n_257_76_9603));
   NAND2_X1 i_257_76_9620 (.A1(n_257_76_9319), .A2(n_257_76_9316), .ZN(
      n_257_76_9604));
   NOR2_X1 i_257_76_9621 (.A1(n_257_76_9604), .A2(n_257_76_9396), .ZN(
      n_257_76_9605));
   NAND4_X1 i_257_76_9622 (.A1(n_257_76_9603), .A2(n_257_76_9220), .A3(
      n_257_76_9221), .A4(n_257_76_9605), .ZN(n_257_76_9606));
   INV_X1 i_257_76_9623 (.A(n_257_76_9606), .ZN(n_257_76_9607));
   NAND2_X1 i_257_76_9624 (.A1(n_257_76_18082), .A2(n_257_76_9607), .ZN(
      n_257_76_9608));
   NAND3_X1 i_257_76_9625 (.A1(n_257_76_9568), .A2(n_257_76_9585), .A3(
      n_257_76_9608), .ZN(n_257_76_9609));
   INV_X1 i_257_76_9626 (.A(n_257_76_9609), .ZN(n_257_76_9610));
   NAND3_X1 i_257_76_9627 (.A1(n_257_76_9241), .A2(n_257_76_9242), .A3(
      n_257_76_9243), .ZN(n_257_76_9611));
   INV_X1 i_257_76_9628 (.A(n_257_76_9611), .ZN(n_257_76_9612));
   NAND4_X1 i_257_76_9629 (.A1(n_257_76_9612), .A2(n_257_76_9233), .A3(
      n_257_76_9234), .A4(n_257_76_9235), .ZN(n_257_76_9613));
   NAND2_X1 i_257_76_9630 (.A1(n_257_427), .A2(n_257_76_9297), .ZN(n_257_76_9614));
   INV_X1 i_257_76_9631 (.A(n_257_76_9614), .ZN(n_257_76_9615));
   NAND4_X1 i_257_76_9632 (.A1(n_257_76_9615), .A2(n_257_76_9223), .A3(n_257_208), 
      .A4(n_257_76_18031), .ZN(n_257_76_9616));
   INV_X1 i_257_76_9633 (.A(n_257_76_9616), .ZN(n_257_76_9617));
   NAND3_X1 i_257_76_9634 (.A1(n_257_76_9222), .A2(n_257_76_9617), .A3(
      n_257_76_9238), .ZN(n_257_76_9618));
   NOR2_X1 i_257_76_9635 (.A1(n_257_76_9613), .A2(n_257_76_9618), .ZN(
      n_257_76_9619));
   NAND4_X1 i_257_76_9636 (.A1(n_257_76_9313), .A2(n_257_76_9619), .A3(
      n_257_76_9355), .A4(n_257_76_9317), .ZN(n_257_76_9620));
   NOR2_X1 i_257_76_9637 (.A1(n_257_76_9620), .A2(n_257_76_9357), .ZN(
      n_257_76_9621));
   NAND3_X1 i_257_76_9638 (.A1(n_257_76_9621), .A2(n_257_76_9220), .A3(
      n_257_76_9221), .ZN(n_257_76_9622));
   INV_X1 i_257_76_9639 (.A(n_257_76_9622), .ZN(n_257_76_9623));
   NAND2_X1 i_257_76_9640 (.A1(n_257_76_18065), .A2(n_257_76_9623), .ZN(
      n_257_76_9624));
   NAND3_X1 i_257_76_9641 (.A1(n_257_76_9255), .A2(n_257_76_9248), .A3(
      n_257_76_9222), .ZN(n_257_76_9625));
   INV_X1 i_257_76_9642 (.A(n_257_76_9247), .ZN(n_257_76_9626));
   NAND2_X1 i_257_76_9643 (.A1(n_257_76_9626), .A2(n_257_76_9237), .ZN(
      n_257_76_9627));
   NOR2_X1 i_257_76_9644 (.A1(n_257_76_9625), .A2(n_257_76_9627), .ZN(
      n_257_76_9628));
   NAND3_X1 i_257_76_9645 (.A1(n_257_76_9253), .A2(n_257_76_9254), .A3(
      n_257_76_9557), .ZN(n_257_76_9629));
   INV_X1 i_257_76_9646 (.A(n_257_76_9629), .ZN(n_257_76_9630));
   NAND4_X1 i_257_76_9647 (.A1(n_257_76_9251), .A2(n_257_76_9628), .A3(
      n_257_76_9252), .A4(n_257_76_9630), .ZN(n_257_76_9631));
   INV_X1 i_257_76_9648 (.A(n_257_76_9631), .ZN(n_257_76_9632));
   NAND3_X1 i_257_76_9649 (.A1(n_257_76_9220), .A2(n_257_76_9632), .A3(
      n_257_76_9221), .ZN(n_257_76_9633));
   INV_X1 i_257_76_9650 (.A(n_257_76_9633), .ZN(n_257_76_9634));
   NAND2_X1 i_257_76_9651 (.A1(n_257_76_18063), .A2(n_257_76_9634), .ZN(
      n_257_76_9635));
   NAND3_X1 i_257_76_9652 (.A1(n_257_76_9237), .A2(n_257_76_9248), .A3(
      n_257_76_9222), .ZN(n_257_76_9636));
   NAND3_X1 i_257_76_9653 (.A1(n_257_76_9309), .A2(n_257_76_9255), .A3(
      n_257_76_9247), .ZN(n_257_76_9637));
   NOR2_X1 i_257_76_9654 (.A1(n_257_76_9636), .A2(n_257_76_9637), .ZN(
      n_257_76_9638));
   NAND4_X1 i_257_76_9655 (.A1(n_257_76_9638), .A2(n_257_76_9598), .A3(
      n_257_76_9252), .A4(n_257_76_9317), .ZN(n_257_76_9639));
   NAND2_X1 i_257_76_9656 (.A1(n_257_76_9297), .A2(n_257_424), .ZN(n_257_76_9640));
   NOR2_X1 i_257_76_9657 (.A1(n_257_76_9296), .A2(n_257_76_9640), .ZN(
      n_257_76_9641));
   NAND4_X1 i_257_76_9658 (.A1(n_257_76_9641), .A2(n_257_76_9242), .A3(
      n_257_76_9243), .A4(n_257_76_9223), .ZN(n_257_76_9642));
   INV_X1 i_257_76_9659 (.A(n_257_76_9642), .ZN(n_257_76_9643));
   NAND3_X1 i_257_76_9660 (.A1(n_257_517), .A2(n_257_76_9241), .A3(n_257_76_9301), 
      .ZN(n_257_76_9644));
   INV_X1 i_257_76_9661 (.A(n_257_76_9644), .ZN(n_257_76_9645));
   NAND3_X1 i_257_76_9662 (.A1(n_257_76_9643), .A2(n_257_76_9645), .A3(
      n_257_76_9238), .ZN(n_257_76_9646));
   INV_X1 i_257_76_9663 (.A(n_257_76_9646), .ZN(n_257_76_9647));
   NAND4_X1 i_257_76_9664 (.A1(n_257_76_9251), .A2(n_257_76_9319), .A3(
      n_257_76_9316), .A4(n_257_76_9647), .ZN(n_257_76_9648));
   NOR2_X1 i_257_76_9665 (.A1(n_257_76_9639), .A2(n_257_76_9648), .ZN(
      n_257_76_9649));
   NAND3_X1 i_257_76_9666 (.A1(n_257_76_9649), .A2(n_257_76_9220), .A3(
      n_257_76_9221), .ZN(n_257_76_9650));
   INV_X1 i_257_76_9667 (.A(n_257_76_9650), .ZN(n_257_76_9651));
   NAND2_X1 i_257_76_9668 (.A1(n_257_76_18062), .A2(n_257_76_9651), .ZN(
      n_257_76_9652));
   NAND3_X1 i_257_76_9669 (.A1(n_257_76_9624), .A2(n_257_76_9635), .A3(
      n_257_76_9652), .ZN(n_257_76_9653));
   INV_X1 i_257_76_9670 (.A(n_257_76_9653), .ZN(n_257_76_9654));
   NAND4_X1 i_257_76_9671 (.A1(n_257_76_9241), .A2(n_257_76_9301), .A3(
      n_257_76_9242), .A4(n_257_76_9243), .ZN(n_257_76_9655));
   NOR2_X1 i_257_76_9672 (.A1(n_257_76_9655), .A2(n_257_76_9590), .ZN(
      n_257_76_9656));
   NAND2_X1 i_257_76_9673 (.A1(n_257_76_9297), .A2(n_257_422), .ZN(n_257_76_9657));
   INV_X1 i_257_76_9674 (.A(n_257_76_9657), .ZN(n_257_76_9658));
   NAND4_X1 i_257_76_9675 (.A1(n_257_76_9223), .A2(n_257_326), .A3(
      n_257_76_18031), .A4(n_257_76_9658), .ZN(n_257_76_9659));
   INV_X1 i_257_76_9676 (.A(n_257_76_9659), .ZN(n_257_76_9660));
   NAND3_X1 i_257_76_9677 (.A1(n_257_76_9305), .A2(n_257_76_9660), .A3(
      n_257_76_9233), .ZN(n_257_76_9661));
   INV_X1 i_257_76_9678 (.A(n_257_76_9661), .ZN(n_257_76_9662));
   NAND3_X1 i_257_76_9679 (.A1(n_257_76_9656), .A2(n_257_76_9479), .A3(
      n_257_76_9662), .ZN(n_257_76_9663));
   NAND4_X1 i_257_76_9680 (.A1(n_257_76_9255), .A2(n_257_76_9247), .A3(
      n_257_76_9248), .A4(n_257_76_9497), .ZN(n_257_76_9664));
   NOR2_X1 i_257_76_9681 (.A1(n_257_76_9663), .A2(n_257_76_9664), .ZN(
      n_257_76_9665));
   INV_X1 i_257_76_9682 (.A(n_257_76_9579), .ZN(n_257_76_9666));
   NAND3_X1 i_257_76_9683 (.A1(n_257_76_9665), .A2(n_257_76_9462), .A3(
      n_257_76_9666), .ZN(n_257_76_9667));
   NAND3_X1 i_257_76_9684 (.A1(n_257_76_9251), .A2(n_257_76_9319), .A3(
      n_257_76_9316), .ZN(n_257_76_9668));
   NOR2_X1 i_257_76_9685 (.A1(n_257_76_9667), .A2(n_257_76_9668), .ZN(
      n_257_76_9669));
   NAND3_X1 i_257_76_9686 (.A1(n_257_76_9669), .A2(n_257_76_9220), .A3(
      n_257_76_9221), .ZN(n_257_76_9670));
   INV_X1 i_257_76_9687 (.A(n_257_76_9670), .ZN(n_257_76_9671));
   NAND2_X1 i_257_76_9688 (.A1(n_257_342), .A2(n_257_76_9671), .ZN(n_257_76_9672));
   NAND2_X1 i_257_76_9689 (.A1(n_257_749), .A2(n_257_76_17935), .ZN(
      n_257_76_9673));
   NAND2_X1 i_257_76_9690 (.A1(n_257_91), .A2(n_257_76_17932), .ZN(n_257_76_9674));
   NAND3_X1 i_257_76_9691 (.A1(n_257_76_9673), .A2(n_257_76_9674), .A3(
      n_257_76_9646), .ZN(n_257_76_9675));
   NAND2_X1 i_257_76_9692 (.A1(n_257_168), .A2(n_257_76_17331), .ZN(
      n_257_76_9676));
   INV_X1 i_257_76_9693 (.A(n_257_76_9676), .ZN(n_257_76_9677));
   NOR2_X1 i_257_76_9694 (.A1(n_257_76_9675), .A2(n_257_76_9677), .ZN(
      n_257_76_9678));
   NAND2_X1 i_257_76_9695 (.A1(n_257_645), .A2(n_257_76_17928), .ZN(
      n_257_76_9679));
   NAND3_X1 i_257_76_9696 (.A1(n_257_441), .A2(n_257_979), .A3(n_257_442), 
      .ZN(n_257_76_9680));
   NAND2_X1 i_257_76_9697 (.A1(n_257_76_9679), .A2(n_257_76_9680), .ZN(
      n_257_76_9681));
   INV_X1 i_257_76_9698 (.A(n_257_76_9681), .ZN(n_257_76_9682));
   INV_X1 i_257_76_9699 (.A(Small_Packet_Data_Size[16]), .ZN(n_257_76_9683));
   NAND2_X1 i_257_76_9700 (.A1(n_257_581), .A2(n_257_428), .ZN(n_257_76_9684));
   NAND3_X1 i_257_76_9701 (.A1(n_257_76_18036), .A2(n_257_76_9297), .A3(
      n_257_76_9684), .ZN(n_257_76_9685));
   INV_X1 i_257_76_9702 (.A(n_257_76_9685), .ZN(n_257_76_9686));
   NAND2_X1 i_257_76_9703 (.A1(n_257_420), .A2(n_257_485), .ZN(n_257_76_9687));
   NAND3_X1 i_257_76_9704 (.A1(n_257_76_9223), .A2(n_257_76_9686), .A3(
      n_257_76_9687), .ZN(n_257_76_9688));
   NAND2_X1 i_257_76_9705 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[16]), 
      .ZN(n_257_76_9689));
   NAND2_X1 i_257_76_9706 (.A1(n_257_76_9688), .A2(n_257_76_9689), .ZN(
      n_257_76_9690));
   NAND2_X1 i_257_76_9707 (.A1(n_257_51), .A2(n_257_76_17918), .ZN(n_257_76_9691));
   NAND4_X1 i_257_76_9708 (.A1(n_257_76_9690), .A2(n_257_76_9691), .A3(
      n_257_76_9616), .A4(n_257_76_9659), .ZN(n_257_76_9692));
   INV_X1 i_257_76_9709 (.A(n_257_76_9692), .ZN(n_257_76_9693));
   INV_X1 i_257_76_9710 (.A(n_257_76_9286), .ZN(n_257_76_9694));
   NAND2_X1 i_257_76_9711 (.A1(n_257_446), .A2(n_257_76_9694), .ZN(n_257_76_9695));
   NAND2_X1 i_257_76_9712 (.A1(n_257_449), .A2(n_257_76_16992), .ZN(
      n_257_76_9696));
   INV_X1 i_257_76_9713 (.A(n_257_76_9533), .ZN(n_257_76_9697));
   NAND2_X1 i_257_76_9714 (.A1(n_257_447), .A2(n_257_76_9697), .ZN(n_257_76_9698));
   NAND3_X1 i_257_76_9715 (.A1(n_257_76_9695), .A2(n_257_76_9696), .A3(
      n_257_76_9698), .ZN(n_257_76_9699));
   NAND3_X1 i_257_76_9716 (.A1(n_257_1081), .A2(n_257_438), .A3(n_257_442), 
      .ZN(n_257_76_9700));
   NAND2_X1 i_257_76_9717 (.A1(n_257_717), .A2(n_257_76_15655), .ZN(
      n_257_76_9701));
   NAND2_X1 i_257_76_9718 (.A1(n_257_440), .A2(n_257_76_9225), .ZN(n_257_76_9702));
   NAND3_X1 i_257_76_9719 (.A1(n_257_76_9700), .A2(n_257_76_9701), .A3(
      n_257_76_9702), .ZN(n_257_76_9703));
   NOR2_X1 i_257_76_9720 (.A1(n_257_76_9699), .A2(n_257_76_9703), .ZN(
      n_257_76_9704));
   NAND3_X1 i_257_76_9721 (.A1(n_257_76_9682), .A2(n_257_76_9693), .A3(
      n_257_76_9704), .ZN(n_257_76_9705));
   NAND2_X1 i_257_76_9722 (.A1(n_257_813), .A2(n_257_76_17952), .ZN(
      n_257_76_9706));
   NAND2_X1 i_257_76_9723 (.A1(n_257_877), .A2(n_257_76_17903), .ZN(
      n_257_76_9707));
   NAND2_X1 i_257_76_9724 (.A1(n_257_129), .A2(n_257_76_17925), .ZN(
      n_257_76_9708));
   NAND2_X1 i_257_76_9725 (.A1(n_257_915), .A2(n_257_76_17940), .ZN(
      n_257_76_9709));
   NAND4_X1 i_257_76_9726 (.A1(n_257_76_9706), .A2(n_257_76_9707), .A3(
      n_257_76_9708), .A4(n_257_76_9709), .ZN(n_257_76_9710));
   NOR2_X1 i_257_76_9727 (.A1(n_257_76_9705), .A2(n_257_76_9710), .ZN(
      n_257_76_9711));
   INV_X1 i_257_76_9728 (.A(n_257_76_13584), .ZN(n_257_76_9712));
   NAND2_X1 i_257_76_9729 (.A1(n_257_813), .A2(n_257_76_9712), .ZN(n_257_76_9713));
   INV_X1 i_257_76_9730 (.A(n_257_76_9713), .ZN(n_257_76_9714));
   INV_X1 i_257_76_9731 (.A(n_257_877), .ZN(n_257_76_9715));
   NAND2_X1 i_257_76_9732 (.A1(n_257_76_9715), .A2(n_257_442), .ZN(n_257_76_9716));
   INV_X1 i_257_76_9733 (.A(n_257_915), .ZN(n_257_76_9717));
   NAND2_X1 i_257_76_9734 (.A1(n_257_76_9717), .A2(n_257_442), .ZN(n_257_76_9718));
   NAND3_X1 i_257_76_9735 (.A1(n_257_76_9714), .A2(n_257_76_9716), .A3(
      n_257_76_9718), .ZN(n_257_76_9719));
   NOR2_X1 i_257_76_9736 (.A1(n_257_76_13584), .A2(n_257_442), .ZN(n_257_76_9720));
   NAND3_X1 i_257_76_9737 (.A1(n_257_76_9716), .A2(n_257_76_9718), .A3(
      n_257_76_9720), .ZN(n_257_76_9721));
   NAND3_X1 i_257_76_9738 (.A1(n_257_76_9719), .A2(n_257_76_9721), .A3(
      n_257_76_9626), .ZN(n_257_76_9722));
   NAND2_X1 i_257_76_9739 (.A1(n_257_685), .A2(n_257_76_17958), .ZN(
      n_257_76_9723));
   NAND4_X1 i_257_76_9740 (.A1(n_257_76_9678), .A2(n_257_76_9711), .A3(
      n_257_76_9722), .A4(n_257_76_9723), .ZN(n_257_76_9724));
   NAND3_X1 i_257_76_9741 (.A1(n_257_76_9314), .A2(n_257_76_9602), .A3(
      n_257_76_9394), .ZN(n_257_76_9725));
   NOR2_X1 i_257_76_9742 (.A1(n_257_76_9724), .A2(n_257_76_9725), .ZN(
      n_257_76_9726));
   AOI22_X1 i_257_76_9743 (.A1(n_257_1011), .A2(n_257_76_17964), .B1(n_257_1043), 
      .B2(n_257_76_17969), .ZN(n_257_76_9727));
   NAND3_X1 i_257_76_9744 (.A1(n_257_76_9726), .A2(n_257_76_9583), .A3(
      n_257_76_9727), .ZN(n_257_76_9728));
   INV_X1 i_257_76_9745 (.A(n_257_76_9728), .ZN(n_257_76_9729));
   NAND3_X1 i_257_76_9746 (.A1(n_257_404), .A2(n_257_484), .A3(n_257_442), 
      .ZN(n_257_76_9730));
   INV_X1 i_257_76_9747 (.A(n_257_76_9730), .ZN(n_257_76_9731));
   NAND3_X1 i_257_76_9748 (.A1(n_257_76_9297), .A2(n_257_76_9684), .A3(
      n_257_76_9731), .ZN(n_257_76_9732));
   INV_X1 i_257_76_9749 (.A(n_257_76_9732), .ZN(n_257_76_9733));
   NAND3_X1 i_257_76_9750 (.A1(n_257_76_9223), .A2(n_257_76_9733), .A3(
      n_257_76_9687), .ZN(n_257_76_9734));
   NOR2_X1 i_257_76_9751 (.A1(n_257_76_9332), .A2(n_257_76_9734), .ZN(
      n_257_76_9735));
   NAND3_X1 i_257_76_9752 (.A1(n_257_76_9735), .A2(n_257_76_9591), .A3(
      n_257_76_9593), .ZN(n_257_76_9736));
   NAND4_X1 i_257_76_9753 (.A1(n_257_76_9222), .A2(n_257_76_9238), .A3(
      n_257_76_9305), .A4(n_257_76_9233), .ZN(n_257_76_9737));
   NOR2_X1 i_257_76_9754 (.A1(n_257_76_9736), .A2(n_257_76_9737), .ZN(
      n_257_76_9738));
   NAND4_X1 i_257_76_9755 (.A1(n_257_76_9251), .A2(n_257_76_9738), .A3(
      n_257_76_9319), .A4(n_257_76_9316), .ZN(n_257_76_9739));
   NAND3_X1 i_257_76_9756 (.A1(n_257_76_9309), .A2(n_257_76_9504), .A3(
      n_257_76_9255), .ZN(n_257_76_9740));
   NAND3_X1 i_257_76_9757 (.A1(n_257_76_9247), .A2(n_257_76_9248), .A3(
      n_257_76_9497), .ZN(n_257_76_9741));
   NOR2_X1 i_257_76_9758 (.A1(n_257_76_9740), .A2(n_257_76_9741), .ZN(
      n_257_76_9742));
   NAND4_X1 i_257_76_9759 (.A1(n_257_76_9742), .A2(n_257_76_9598), .A3(
      n_257_76_9252), .A4(n_257_76_9317), .ZN(n_257_76_9743));
   NOR2_X1 i_257_76_9760 (.A1(n_257_76_9739), .A2(n_257_76_9743), .ZN(
      n_257_76_9744));
   NAND3_X1 i_257_76_9761 (.A1(n_257_76_9744), .A2(n_257_76_9220), .A3(
      n_257_76_9221), .ZN(n_257_76_9745));
   INV_X1 i_257_76_9762 (.A(n_257_76_9745), .ZN(n_257_76_9746));
   AOI21_X1 i_257_76_9763 (.A(n_257_76_9729), .B1(n_257_76_18060), .B2(
      n_257_76_9746), .ZN(n_257_76_9747));
   NAND2_X1 i_257_76_9764 (.A1(n_257_76_9672), .A2(n_257_76_9747), .ZN(
      n_257_76_9748));
   INV_X1 i_257_76_9765 (.A(n_257_76_9748), .ZN(n_257_76_9749));
   NAND3_X1 i_257_76_9766 (.A1(n_257_76_9610), .A2(n_257_76_9654), .A3(
      n_257_76_9749), .ZN(n_257_76_9750));
   NOR2_X1 i_257_76_9767 (.A1(n_257_76_9552), .A2(n_257_76_9750), .ZN(
      n_257_76_9751));
   NAND2_X1 i_257_76_9768 (.A1(n_257_76_9427), .A2(n_257_76_9751), .ZN(n_16));
   NAND2_X1 i_257_76_9769 (.A1(n_257_1012), .A2(n_257_444), .ZN(n_257_76_9752));
   NAND2_X1 i_257_76_9770 (.A1(n_257_441), .A2(n_257_980), .ZN(n_257_76_9753));
   NAND2_X1 i_257_76_9771 (.A1(n_257_948), .A2(n_257_442), .ZN(n_257_76_9754));
   NOR2_X1 i_257_76_9772 (.A1(n_257_1076), .A2(n_257_76_9754), .ZN(n_257_76_9755));
   NAND2_X1 i_257_76_9773 (.A1(n_257_440), .A2(n_257_76_9755), .ZN(n_257_76_9756));
   INV_X1 i_257_76_9774 (.A(n_257_76_9756), .ZN(n_257_76_9757));
   NAND2_X1 i_257_76_9775 (.A1(n_257_76_9753), .A2(n_257_76_9757), .ZN(
      n_257_76_9758));
   INV_X1 i_257_76_9776 (.A(n_257_76_9758), .ZN(n_257_76_9759));
   NAND2_X1 i_257_76_9777 (.A1(n_257_76_9752), .A2(n_257_76_9759), .ZN(
      n_257_76_9760));
   INV_X1 i_257_76_9778 (.A(n_257_76_9760), .ZN(n_257_76_9761));
   NAND2_X1 i_257_76_9779 (.A1(n_257_1044), .A2(n_257_443), .ZN(n_257_76_9762));
   NAND2_X1 i_257_76_9780 (.A1(n_257_76_9761), .A2(n_257_76_9762), .ZN(
      n_257_76_9763));
   INV_X1 i_257_76_9781 (.A(n_257_76_9763), .ZN(n_257_76_9764));
   NAND2_X1 i_257_76_9782 (.A1(n_257_17), .A2(n_257_76_9764), .ZN(n_257_76_9765));
   NOR2_X1 i_257_76_9783 (.A1(n_257_1076), .A2(n_257_76_17412), .ZN(
      n_257_76_9766));
   INV_X1 i_257_76_9784 (.A(n_257_76_9766), .ZN(n_257_76_9767));
   NOR2_X1 i_257_76_9785 (.A1(n_257_76_9767), .A2(n_257_76_15197), .ZN(
      n_257_76_9768));
   NAND2_X1 i_257_76_9786 (.A1(n_257_1044), .A2(n_257_76_9768), .ZN(
      n_257_76_9769));
   INV_X1 i_257_76_9787 (.A(n_257_76_9769), .ZN(n_257_76_9770));
   NAND2_X1 i_257_76_9788 (.A1(n_257_76_18072), .A2(n_257_76_9770), .ZN(
      n_257_76_9771));
   INV_X1 i_257_76_9789 (.A(n_257_76_9762), .ZN(n_257_76_9772));
   NAND2_X1 i_257_76_9790 (.A1(n_257_750), .A2(n_257_436), .ZN(n_257_76_9773));
   NAND2_X1 i_257_76_9791 (.A1(n_257_916), .A2(n_257_439), .ZN(n_257_76_9774));
   NAND2_X1 i_257_76_9792 (.A1(n_257_814), .A2(n_257_437), .ZN(n_257_76_9775));
   NAND4_X1 i_257_76_9793 (.A1(n_257_76_9773), .A2(n_257_76_9774), .A3(
      n_257_76_9775), .A4(n_257_76_9753), .ZN(n_257_76_9776));
   NAND2_X1 i_257_76_9794 (.A1(n_257_449), .A2(n_257_1090), .ZN(n_257_76_9777));
   NAND2_X1 i_257_76_9795 (.A1(n_257_447), .A2(n_257_782), .ZN(n_257_76_9778));
   NAND3_X1 i_257_76_9796 (.A1(n_257_76_9777), .A2(n_257_76_9778), .A3(n_257_646), 
      .ZN(n_257_76_9779));
   INV_X1 i_257_76_9797 (.A(n_257_76_9779), .ZN(n_257_76_9780));
   NAND2_X1 i_257_76_9798 (.A1(n_257_878), .A2(n_257_445), .ZN(n_257_76_9781));
   NAND2_X1 i_257_76_9799 (.A1(n_257_446), .A2(n_257_846), .ZN(n_257_76_9782));
   NAND2_X1 i_257_76_9800 (.A1(n_257_76_9781), .A2(n_257_76_9782), .ZN(
      n_257_76_9783));
   INV_X1 i_257_76_9801 (.A(n_257_76_9783), .ZN(n_257_76_9784));
   NAND2_X1 i_257_76_9802 (.A1(n_257_438), .A2(n_257_1082), .ZN(n_257_76_9785));
   NAND2_X1 i_257_76_9803 (.A1(n_257_440), .A2(n_257_948), .ZN(n_257_76_9786));
   NAND2_X1 i_257_76_9804 (.A1(n_257_718), .A2(n_257_435), .ZN(n_257_76_9787));
   NOR2_X1 i_257_76_9805 (.A1(n_257_76_17927), .A2(n_257_1076), .ZN(
      n_257_76_9788));
   NAND4_X1 i_257_76_9806 (.A1(n_257_76_9785), .A2(n_257_76_9786), .A3(
      n_257_76_9787), .A4(n_257_76_9788), .ZN(n_257_76_9789));
   INV_X1 i_257_76_9807 (.A(n_257_76_9789), .ZN(n_257_76_9790));
   NAND3_X1 i_257_76_9808 (.A1(n_257_76_9780), .A2(n_257_76_9784), .A3(
      n_257_76_9790), .ZN(n_257_76_9791));
   NOR2_X1 i_257_76_9809 (.A1(n_257_76_9776), .A2(n_257_76_9791), .ZN(
      n_257_76_9792));
   NAND2_X1 i_257_76_9810 (.A1(n_257_686), .A2(n_257_448), .ZN(n_257_76_9793));
   NAND3_X1 i_257_76_9811 (.A1(n_257_76_9752), .A2(n_257_76_9792), .A3(
      n_257_76_9793), .ZN(n_257_76_9794));
   NOR2_X1 i_257_76_9812 (.A1(n_257_76_9772), .A2(n_257_76_9794), .ZN(
      n_257_76_9795));
   NAND2_X1 i_257_76_9813 (.A1(n_257_28), .A2(n_257_76_9795), .ZN(n_257_76_9796));
   NAND3_X1 i_257_76_9814 (.A1(n_257_76_9765), .A2(n_257_76_9771), .A3(
      n_257_76_9796), .ZN(n_257_76_9797));
   NAND2_X1 i_257_76_9815 (.A1(n_257_846), .A2(n_257_442), .ZN(n_257_76_9798));
   NOR2_X1 i_257_76_9816 (.A1(n_257_1076), .A2(n_257_76_9798), .ZN(n_257_76_9799));
   NAND4_X1 i_257_76_9817 (.A1(n_257_446), .A2(n_257_76_9785), .A3(n_257_76_9786), 
      .A4(n_257_76_9799), .ZN(n_257_76_9800));
   INV_X1 i_257_76_9818 (.A(n_257_76_9800), .ZN(n_257_76_9801));
   NAND4_X1 i_257_76_9819 (.A1(n_257_76_9774), .A2(n_257_76_9801), .A3(
      n_257_76_9753), .A4(n_257_76_9781), .ZN(n_257_76_9802));
   INV_X1 i_257_76_9820 (.A(n_257_76_9802), .ZN(n_257_76_9803));
   NAND2_X1 i_257_76_9821 (.A1(n_257_76_9752), .A2(n_257_76_9803), .ZN(
      n_257_76_9804));
   INV_X1 i_257_76_9822 (.A(n_257_76_9804), .ZN(n_257_76_9805));
   NAND2_X1 i_257_76_9823 (.A1(n_257_76_9805), .A2(n_257_76_9762), .ZN(
      n_257_76_9806));
   INV_X1 i_257_76_9824 (.A(n_257_76_9806), .ZN(n_257_76_9807));
   NAND2_X1 i_257_76_9825 (.A1(n_257_76_18070), .A2(n_257_76_9807), .ZN(
      n_257_76_9808));
   INV_X1 i_257_76_9826 (.A(n_257_76_9786), .ZN(n_257_76_9809));
   NAND2_X1 i_257_76_9827 (.A1(n_257_439), .A2(n_257_76_9766), .ZN(n_257_76_9810));
   NOR2_X1 i_257_76_9828 (.A1(n_257_76_9809), .A2(n_257_76_9810), .ZN(
      n_257_76_9811));
   NAND3_X1 i_257_76_9829 (.A1(n_257_76_9753), .A2(n_257_76_9811), .A3(n_257_916), 
      .ZN(n_257_76_9812));
   INV_X1 i_257_76_9830 (.A(n_257_76_9812), .ZN(n_257_76_9813));
   NAND2_X1 i_257_76_9831 (.A1(n_257_76_9752), .A2(n_257_76_9813), .ZN(
      n_257_76_9814));
   INV_X1 i_257_76_9832 (.A(n_257_76_9814), .ZN(n_257_76_9815));
   NAND2_X1 i_257_76_9833 (.A1(n_257_76_9815), .A2(n_257_76_9762), .ZN(
      n_257_76_9816));
   INV_X1 i_257_76_9834 (.A(n_257_76_9816), .ZN(n_257_76_9817));
   NAND2_X1 i_257_76_9835 (.A1(n_257_76_18084), .A2(n_257_76_9817), .ZN(
      n_257_76_9818));
   NAND2_X1 i_257_76_9836 (.A1(n_257_550), .A2(n_257_426), .ZN(n_257_76_9819));
   NAND2_X1 i_257_76_9837 (.A1(n_257_130), .A2(n_257_430), .ZN(n_257_76_9820));
   NAND3_X1 i_257_76_9838 (.A1(n_257_76_9819), .A2(n_257_76_9773), .A3(
      n_257_76_9820), .ZN(n_257_76_9821));
   INV_X1 i_257_76_9839 (.A(n_257_1076), .ZN(n_257_76_9822));
   NAND2_X1 i_257_76_9840 (.A1(n_257_432), .A2(n_257_614), .ZN(n_257_76_9823));
   NAND4_X1 i_257_76_9841 (.A1(n_257_76_18027), .A2(n_257_76_9822), .A3(
      n_257_76_9823), .A4(n_257_423), .ZN(n_257_76_9824));
   INV_X1 i_257_76_9842 (.A(n_257_76_9824), .ZN(n_257_76_9825));
   NAND4_X1 i_257_76_9843 (.A1(n_257_76_9825), .A2(n_257_76_9785), .A3(
      n_257_76_9786), .A4(n_257_76_9787), .ZN(n_257_76_9826));
   INV_X1 i_257_76_9844 (.A(n_257_76_9826), .ZN(n_257_76_9827));
   NAND2_X1 i_257_76_9845 (.A1(n_257_518), .A2(n_257_424), .ZN(n_257_76_9828));
   NAND2_X1 i_257_76_9846 (.A1(n_257_76_9828), .A2(n_257_76_9781), .ZN(
      n_257_76_9829));
   INV_X1 i_257_76_9847 (.A(n_257_76_9829), .ZN(n_257_76_9830));
   NAND2_X1 i_257_76_9848 (.A1(n_257_52), .A2(n_257_433), .ZN(n_257_76_9831));
   NAND2_X1 i_257_76_9849 (.A1(n_257_209), .A2(n_257_427), .ZN(n_257_76_9832));
   NAND3_X1 i_257_76_9850 (.A1(n_257_76_9831), .A2(n_257_289), .A3(n_257_76_9832), 
      .ZN(n_257_76_9833));
   INV_X1 i_257_76_9851 (.A(n_257_76_9833), .ZN(n_257_76_9834));
   NAND3_X1 i_257_76_9852 (.A1(n_257_76_9827), .A2(n_257_76_9830), .A3(
      n_257_76_9834), .ZN(n_257_76_9835));
   NOR2_X1 i_257_76_9853 (.A1(n_257_76_9821), .A2(n_257_76_9835), .ZN(
      n_257_76_9836));
   NAND2_X1 i_257_76_9854 (.A1(n_257_76_9777), .A2(n_257_76_9778), .ZN(
      n_257_76_9837));
   INV_X1 i_257_76_9855 (.A(n_257_76_9837), .ZN(n_257_76_9838));
   NAND2_X1 i_257_76_9856 (.A1(n_257_646), .A2(n_257_450), .ZN(n_257_76_9839));
   NAND4_X1 i_257_76_9857 (.A1(n_257_76_9838), .A2(n_257_76_9753), .A3(
      n_257_76_9839), .A4(n_257_76_9782), .ZN(n_257_76_9840));
   NAND2_X1 i_257_76_9858 (.A1(n_257_451), .A2(n_257_469), .ZN(n_257_76_9841));
   NAND3_X1 i_257_76_9859 (.A1(n_257_76_9774), .A2(n_257_76_9775), .A3(
      n_257_76_9841), .ZN(n_257_76_9842));
   NOR2_X1 i_257_76_9860 (.A1(n_257_76_9840), .A2(n_257_76_9842), .ZN(
      n_257_76_9843));
   NAND2_X1 i_257_76_9861 (.A1(n_257_169), .A2(n_257_429), .ZN(n_257_76_9844));
   NAND2_X1 i_257_76_9862 (.A1(n_257_249), .A2(n_257_425), .ZN(n_257_76_9845));
   NAND4_X1 i_257_76_9863 (.A1(n_257_76_9836), .A2(n_257_76_9843), .A3(
      n_257_76_9844), .A4(n_257_76_9845), .ZN(n_257_76_9846));
   INV_X1 i_257_76_9864 (.A(n_257_76_9846), .ZN(n_257_76_9847));
   NAND2_X1 i_257_76_9865 (.A1(n_257_92), .A2(n_257_431), .ZN(n_257_76_9848));
   NAND3_X1 i_257_76_9866 (.A1(n_257_76_9752), .A2(n_257_76_9793), .A3(
      n_257_76_9848), .ZN(n_257_76_9849));
   INV_X1 i_257_76_9867 (.A(n_257_76_9849), .ZN(n_257_76_9850));
   NAND3_X1 i_257_76_9868 (.A1(n_257_76_9847), .A2(n_257_76_9850), .A3(
      n_257_76_9762), .ZN(n_257_76_9851));
   INV_X1 i_257_76_9869 (.A(n_257_76_9851), .ZN(n_257_76_9852));
   NAND2_X1 i_257_76_9870 (.A1(n_257_76_18066), .A2(n_257_76_9852), .ZN(
      n_257_76_9853));
   NAND3_X1 i_257_76_9871 (.A1(n_257_76_9808), .A2(n_257_76_9818), .A3(
      n_257_76_9853), .ZN(n_257_76_9854));
   NOR2_X1 i_257_76_9872 (.A1(n_257_76_9797), .A2(n_257_76_9854), .ZN(
      n_257_76_9855));
   NAND3_X1 i_257_76_9873 (.A1(n_257_441), .A2(n_257_980), .A3(n_257_76_9766), 
      .ZN(n_257_76_9856));
   INV_X1 i_257_76_9874 (.A(n_257_76_9856), .ZN(n_257_76_9857));
   NAND2_X1 i_257_76_9875 (.A1(n_257_76_9752), .A2(n_257_76_9857), .ZN(
      n_257_76_9858));
   INV_X1 i_257_76_9876 (.A(n_257_76_9858), .ZN(n_257_76_9859));
   NAND2_X1 i_257_76_9877 (.A1(n_257_76_9859), .A2(n_257_76_9762), .ZN(
      n_257_76_9860));
   INV_X1 i_257_76_9878 (.A(n_257_76_9860), .ZN(n_257_76_9861));
   NAND2_X1 i_257_76_9879 (.A1(n_257_76_18071), .A2(n_257_76_9861), .ZN(
      n_257_76_9862));
   NAND2_X1 i_257_76_9880 (.A1(n_257_76_9782), .A2(n_257_76_9778), .ZN(
      n_257_76_9863));
   INV_X1 i_257_76_9881 (.A(n_257_76_9863), .ZN(n_257_76_9864));
   NAND3_X1 i_257_76_9882 (.A1(n_257_718), .A2(n_257_76_15655), .A3(
      n_257_76_9822), .ZN(n_257_76_9865));
   INV_X1 i_257_76_9883 (.A(n_257_76_9865), .ZN(n_257_76_9866));
   NAND3_X1 i_257_76_9884 (.A1(n_257_76_9866), .A2(n_257_76_9785), .A3(
      n_257_76_9786), .ZN(n_257_76_9867));
   INV_X1 i_257_76_9885 (.A(n_257_76_9867), .ZN(n_257_76_9868));
   NAND4_X1 i_257_76_9886 (.A1(n_257_76_9864), .A2(n_257_76_9868), .A3(
      n_257_76_9753), .A4(n_257_76_9781), .ZN(n_257_76_9869));
   NAND3_X1 i_257_76_9887 (.A1(n_257_76_9773), .A2(n_257_76_9774), .A3(
      n_257_76_9775), .ZN(n_257_76_9870));
   NOR2_X1 i_257_76_9888 (.A1(n_257_76_9869), .A2(n_257_76_9870), .ZN(
      n_257_76_9871));
   NAND2_X1 i_257_76_9889 (.A1(n_257_76_9752), .A2(n_257_76_9871), .ZN(
      n_257_76_9872));
   INV_X1 i_257_76_9890 (.A(n_257_76_9872), .ZN(n_257_76_9873));
   NAND2_X1 i_257_76_9891 (.A1(n_257_76_9873), .A2(n_257_76_9762), .ZN(
      n_257_76_9874));
   INV_X1 i_257_76_9892 (.A(n_257_76_9874), .ZN(n_257_76_9875));
   NAND2_X1 i_257_76_9893 (.A1(n_257_76_18078), .A2(n_257_76_9875), .ZN(
      n_257_76_9876));
   NAND4_X1 i_257_76_9894 (.A1(n_257_76_9775), .A2(n_257_76_9841), .A3(
      n_257_76_9753), .A4(n_257_76_9839), .ZN(n_257_76_9877));
   NAND3_X1 i_257_76_9895 (.A1(n_257_76_9773), .A2(n_257_76_9820), .A3(
      n_257_76_9774), .ZN(n_257_76_9878));
   NOR2_X1 i_257_76_9896 (.A1(n_257_76_9877), .A2(n_257_76_9878), .ZN(
      n_257_76_9879));
   NAND2_X1 i_257_76_9897 (.A1(n_257_76_9785), .A2(n_257_76_9786), .ZN(
      n_257_76_9880));
   INV_X1 i_257_76_9898 (.A(n_257_76_9880), .ZN(n_257_76_9881));
   NAND3_X1 i_257_76_9899 (.A1(n_257_582), .A2(n_257_428), .A3(n_257_442), 
      .ZN(n_257_76_9882));
   INV_X1 i_257_76_9900 (.A(n_257_76_9882), .ZN(n_257_76_9883));
   NAND3_X1 i_257_76_9901 (.A1(n_257_76_9883), .A2(n_257_76_9822), .A3(
      n_257_76_9823), .ZN(n_257_76_9884));
   INV_X1 i_257_76_9902 (.A(n_257_76_9884), .ZN(n_257_76_9885));
   NAND2_X1 i_257_76_9903 (.A1(n_257_76_9885), .A2(n_257_76_9787), .ZN(
      n_257_76_9886));
   INV_X1 i_257_76_9904 (.A(n_257_76_9886), .ZN(n_257_76_9887));
   NAND4_X1 i_257_76_9905 (.A1(n_257_76_9881), .A2(n_257_76_9887), .A3(
      n_257_76_9778), .A4(n_257_76_9831), .ZN(n_257_76_9888));
   NAND3_X1 i_257_76_9906 (.A1(n_257_76_9781), .A2(n_257_76_9782), .A3(
      n_257_76_9777), .ZN(n_257_76_9889));
   NOR2_X1 i_257_76_9907 (.A1(n_257_76_9888), .A2(n_257_76_9889), .ZN(
      n_257_76_9890));
   NAND4_X1 i_257_76_9908 (.A1(n_257_76_9879), .A2(n_257_76_9848), .A3(
      n_257_76_9844), .A4(n_257_76_9890), .ZN(n_257_76_9891));
   INV_X1 i_257_76_9909 (.A(n_257_76_9891), .ZN(n_257_76_9892));
   NAND2_X1 i_257_76_9910 (.A1(n_257_76_9752), .A2(n_257_76_9793), .ZN(
      n_257_76_9893));
   INV_X1 i_257_76_9911 (.A(n_257_76_9893), .ZN(n_257_76_9894));
   NAND3_X1 i_257_76_9912 (.A1(n_257_76_9892), .A2(n_257_76_9894), .A3(
      n_257_76_9762), .ZN(n_257_76_9895));
   INV_X1 i_257_76_9913 (.A(n_257_76_9895), .ZN(n_257_76_9896));
   NAND2_X1 i_257_76_9914 (.A1(n_257_76_18074), .A2(n_257_76_9896), .ZN(
      n_257_76_9897));
   NAND3_X1 i_257_76_9915 (.A1(n_257_76_9862), .A2(n_257_76_9876), .A3(
      n_257_76_9897), .ZN(n_257_76_9898));
   NAND2_X1 i_257_76_9916 (.A1(n_257_1076), .A2(n_257_442), .ZN(n_257_76_9899));
   INV_X1 i_257_76_9917 (.A(n_257_76_9899), .ZN(n_257_76_9900));
   NAND2_X1 i_257_76_9918 (.A1(n_257_13), .A2(n_257_76_9900), .ZN(n_257_76_9901));
   NOR2_X1 i_257_76_9919 (.A1(n_257_76_9767), .A2(n_257_76_11918), .ZN(
      n_257_76_9902));
   NAND4_X1 i_257_76_9920 (.A1(n_257_76_9902), .A2(n_257_878), .A3(n_257_76_9785), 
      .A4(n_257_76_9786), .ZN(n_257_76_9903));
   INV_X1 i_257_76_9921 (.A(n_257_76_9903), .ZN(n_257_76_9904));
   NAND3_X1 i_257_76_9922 (.A1(n_257_76_9904), .A2(n_257_76_9774), .A3(
      n_257_76_9753), .ZN(n_257_76_9905));
   INV_X1 i_257_76_9923 (.A(n_257_76_9905), .ZN(n_257_76_9906));
   NAND2_X1 i_257_76_9924 (.A1(n_257_76_9752), .A2(n_257_76_9906), .ZN(
      n_257_76_9907));
   INV_X1 i_257_76_9925 (.A(n_257_76_9907), .ZN(n_257_76_9908));
   NAND2_X1 i_257_76_9926 (.A1(n_257_76_9908), .A2(n_257_76_9762), .ZN(
      n_257_76_9909));
   INV_X1 i_257_76_9927 (.A(n_257_76_9909), .ZN(n_257_76_9910));
   NAND2_X1 i_257_76_9928 (.A1(n_257_76_18077), .A2(n_257_76_9910), .ZN(
      n_257_76_9911));
   NAND2_X1 i_257_76_9929 (.A1(n_257_76_9901), .A2(n_257_76_9911), .ZN(
      n_257_76_9912));
   NOR2_X1 i_257_76_9930 (.A1(n_257_76_9898), .A2(n_257_76_9912), .ZN(
      n_257_76_9913));
   INV_X1 i_257_76_9931 (.A(n_257_76_9752), .ZN(n_257_76_9914));
   NAND4_X1 i_257_76_9932 (.A1(n_257_76_18027), .A2(n_257_76_9822), .A3(
      n_257_76_9823), .A4(n_257_426), .ZN(n_257_76_9915));
   INV_X1 i_257_76_9933 (.A(n_257_76_9787), .ZN(n_257_76_9916));
   NOR2_X1 i_257_76_9934 (.A1(n_257_76_9915), .A2(n_257_76_9916), .ZN(
      n_257_76_9917));
   NAND3_X1 i_257_76_9935 (.A1(n_257_76_9917), .A2(n_257_76_9881), .A3(
      n_257_76_9832), .ZN(n_257_76_9918));
   NAND4_X1 i_257_76_9936 (.A1(n_257_76_9782), .A2(n_257_76_9777), .A3(
      n_257_76_9778), .A4(n_257_76_9831), .ZN(n_257_76_9919));
   NOR2_X1 i_257_76_9937 (.A1(n_257_76_9918), .A2(n_257_76_9919), .ZN(
      n_257_76_9920));
   INV_X1 i_257_76_9938 (.A(n_257_76_9878), .ZN(n_257_76_9921));
   NAND4_X1 i_257_76_9939 (.A1(n_257_76_9775), .A2(n_257_550), .A3(n_257_76_9839), 
      .A4(n_257_76_9781), .ZN(n_257_76_9922));
   INV_X1 i_257_76_9940 (.A(n_257_76_9922), .ZN(n_257_76_9923));
   NAND3_X1 i_257_76_9941 (.A1(n_257_76_9920), .A2(n_257_76_9921), .A3(
      n_257_76_9923), .ZN(n_257_76_9924));
   NOR2_X1 i_257_76_9942 (.A1(n_257_76_9914), .A2(n_257_76_9924), .ZN(
      n_257_76_9925));
   NAND2_X1 i_257_76_9943 (.A1(n_257_76_9841), .A2(n_257_76_9753), .ZN(
      n_257_76_9926));
   INV_X1 i_257_76_9944 (.A(n_257_76_9926), .ZN(n_257_76_9927));
   NAND4_X1 i_257_76_9945 (.A1(n_257_76_9793), .A2(n_257_76_9848), .A3(
      n_257_76_9844), .A4(n_257_76_9927), .ZN(n_257_76_9928));
   INV_X1 i_257_76_9946 (.A(n_257_76_9928), .ZN(n_257_76_9929));
   NAND3_X1 i_257_76_9947 (.A1(n_257_76_9925), .A2(n_257_76_9929), .A3(
      n_257_76_9762), .ZN(n_257_76_9930));
   INV_X1 i_257_76_9948 (.A(n_257_76_9930), .ZN(n_257_76_9931));
   NAND2_X1 i_257_76_9949 (.A1(n_257_76_18076), .A2(n_257_76_9931), .ZN(
      n_257_76_9932));
   INV_X1 i_257_76_9950 (.A(n_257_76_9778), .ZN(n_257_76_9933));
   NOR2_X1 i_257_76_9951 (.A1(n_257_76_17934), .A2(n_257_1076), .ZN(
      n_257_76_9934));
   NAND3_X1 i_257_76_9952 (.A1(n_257_76_9785), .A2(n_257_76_9786), .A3(
      n_257_76_9934), .ZN(n_257_76_9935));
   NOR2_X1 i_257_76_9953 (.A1(n_257_76_9933), .A2(n_257_76_9935), .ZN(
      n_257_76_9936));
   NAND3_X1 i_257_76_9954 (.A1(n_257_76_9936), .A2(n_257_76_9784), .A3(n_257_750), 
      .ZN(n_257_76_9937));
   NAND3_X1 i_257_76_9955 (.A1(n_257_76_9774), .A2(n_257_76_9775), .A3(
      n_257_76_9753), .ZN(n_257_76_9938));
   NOR2_X1 i_257_76_9956 (.A1(n_257_76_9937), .A2(n_257_76_9938), .ZN(
      n_257_76_9939));
   NAND2_X1 i_257_76_9957 (.A1(n_257_76_9752), .A2(n_257_76_9939), .ZN(
      n_257_76_9940));
   NOR2_X1 i_257_76_9958 (.A1(n_257_76_9772), .A2(n_257_76_9940), .ZN(
      n_257_76_9941));
   NAND2_X1 i_257_76_9959 (.A1(n_257_76_18069), .A2(n_257_76_9941), .ZN(
      n_257_76_9942));
   NAND2_X1 i_257_76_9960 (.A1(n_257_76_9778), .A2(n_257_76_9831), .ZN(
      n_257_76_9943));
   NAND3_X1 i_257_76_9961 (.A1(n_257_432), .A2(n_257_614), .A3(n_257_442), 
      .ZN(n_257_76_9944));
   NOR2_X1 i_257_76_9962 (.A1(n_257_76_9944), .A2(n_257_1076), .ZN(n_257_76_9945));
   NAND4_X1 i_257_76_9963 (.A1(n_257_76_9785), .A2(n_257_76_9786), .A3(
      n_257_76_9787), .A4(n_257_76_9945), .ZN(n_257_76_9946));
   NOR2_X1 i_257_76_9964 (.A1(n_257_76_9943), .A2(n_257_76_9946), .ZN(
      n_257_76_9947));
   NAND2_X1 i_257_76_9965 (.A1(n_257_76_9753), .A2(n_257_76_9839), .ZN(
      n_257_76_9948));
   INV_X1 i_257_76_9966 (.A(n_257_76_9948), .ZN(n_257_76_9949));
   INV_X1 i_257_76_9967 (.A(n_257_76_9889), .ZN(n_257_76_9950));
   NAND3_X1 i_257_76_9968 (.A1(n_257_76_9947), .A2(n_257_76_9949), .A3(
      n_257_76_9950), .ZN(n_257_76_9951));
   NAND4_X1 i_257_76_9969 (.A1(n_257_76_9773), .A2(n_257_76_9774), .A3(
      n_257_76_9775), .A4(n_257_76_9841), .ZN(n_257_76_9952));
   NOR2_X1 i_257_76_9970 (.A1(n_257_76_9951), .A2(n_257_76_9952), .ZN(
      n_257_76_9953));
   NAND3_X1 i_257_76_9971 (.A1(n_257_76_9953), .A2(n_257_76_9752), .A3(
      n_257_76_9793), .ZN(n_257_76_9954));
   NOR2_X1 i_257_76_9972 (.A1(n_257_76_9954), .A2(n_257_76_9772), .ZN(
      n_257_76_9955));
   NAND2_X1 i_257_76_9973 (.A1(n_257_68), .A2(n_257_76_9955), .ZN(n_257_76_9956));
   NAND3_X1 i_257_76_9974 (.A1(n_257_76_9932), .A2(n_257_76_9942), .A3(
      n_257_76_9956), .ZN(n_257_76_9957));
   NOR2_X1 i_257_76_9975 (.A1(n_257_76_17951), .A2(n_257_1076), .ZN(
      n_257_76_9958));
   NAND3_X1 i_257_76_9976 (.A1(n_257_76_9785), .A2(n_257_76_9786), .A3(
      n_257_76_9958), .ZN(n_257_76_9959));
   INV_X1 i_257_76_9977 (.A(n_257_76_9959), .ZN(n_257_76_9960));
   NAND4_X1 i_257_76_9978 (.A1(n_257_76_9960), .A2(n_257_814), .A3(n_257_76_9781), 
      .A4(n_257_76_9782), .ZN(n_257_76_9961));
   NAND2_X1 i_257_76_9979 (.A1(n_257_76_9774), .A2(n_257_76_9753), .ZN(
      n_257_76_9962));
   NOR2_X1 i_257_76_9980 (.A1(n_257_76_9961), .A2(n_257_76_9962), .ZN(
      n_257_76_9963));
   NAND2_X1 i_257_76_9981 (.A1(n_257_76_9752), .A2(n_257_76_9963), .ZN(
      n_257_76_9964));
   INV_X1 i_257_76_9982 (.A(n_257_76_9964), .ZN(n_257_76_9965));
   NAND2_X1 i_257_76_9983 (.A1(n_257_76_9965), .A2(n_257_76_9762), .ZN(
      n_257_76_9966));
   INV_X1 i_257_76_9984 (.A(n_257_76_9966), .ZN(n_257_76_9967));
   NAND2_X1 i_257_76_9985 (.A1(n_257_22), .A2(n_257_76_9967), .ZN(n_257_76_9968));
   NAND2_X1 i_257_76_9986 (.A1(n_257_444), .A2(n_257_76_9766), .ZN(n_257_76_9969));
   INV_X1 i_257_76_9987 (.A(n_257_76_9969), .ZN(n_257_76_9970));
   NAND2_X1 i_257_76_9988 (.A1(n_257_1012), .A2(n_257_76_9970), .ZN(
      n_257_76_9971));
   INV_X1 i_257_76_9989 (.A(n_257_76_9971), .ZN(n_257_76_9972));
   NAND2_X1 i_257_76_9990 (.A1(n_257_76_9762), .A2(n_257_76_9972), .ZN(
      n_257_76_9973));
   INV_X1 i_257_76_9991 (.A(n_257_76_9973), .ZN(n_257_76_9974));
   NAND2_X1 i_257_76_9992 (.A1(n_257_76_18075), .A2(n_257_76_9974), .ZN(
      n_257_76_9975));
   NAND2_X1 i_257_76_9993 (.A1(n_257_76_9968), .A2(n_257_76_9975), .ZN(
      n_257_76_9976));
   NOR2_X1 i_257_76_9994 (.A1(n_257_76_9957), .A2(n_257_76_9976), .ZN(
      n_257_76_9977));
   NAND3_X1 i_257_76_9995 (.A1(n_257_76_9855), .A2(n_257_76_9913), .A3(
      n_257_76_9977), .ZN(n_257_76_9978));
   INV_X1 i_257_76_9996 (.A(n_257_76_9978), .ZN(n_257_76_9979));
   NOR2_X1 i_257_76_9997 (.A1(n_257_1076), .A2(n_257_76_17633), .ZN(
      n_257_76_9980));
   NAND3_X1 i_257_76_9998 (.A1(n_257_52), .A2(n_257_76_9787), .A3(n_257_76_9980), 
      .ZN(n_257_76_9981));
   INV_X1 i_257_76_9999 (.A(n_257_76_9981), .ZN(n_257_76_9982));
   NAND3_X1 i_257_76_10000 (.A1(n_257_76_9982), .A2(n_257_76_9881), .A3(
      n_257_76_9778), .ZN(n_257_76_9983));
   INV_X1 i_257_76_10001 (.A(n_257_76_9983), .ZN(n_257_76_9984));
   NAND3_X1 i_257_76_10002 (.A1(n_257_76_9949), .A2(n_257_76_9984), .A3(
      n_257_76_9950), .ZN(n_257_76_9985));
   NOR2_X1 i_257_76_10003 (.A1(n_257_76_9985), .A2(n_257_76_9952), .ZN(
      n_257_76_9986));
   NAND3_X1 i_257_76_10004 (.A1(n_257_76_9986), .A2(n_257_76_9752), .A3(
      n_257_76_9793), .ZN(n_257_76_9987));
   NOR2_X1 i_257_76_10005 (.A1(n_257_76_9772), .A2(n_257_76_9987), .ZN(
      n_257_76_9988));
   NAND2_X1 i_257_76_10006 (.A1(n_257_76_18081), .A2(n_257_76_9988), .ZN(
      n_257_76_9989));
   NAND3_X1 i_257_76_10007 (.A1(n_257_76_9781), .A2(n_257_76_9782), .A3(
      n_257_76_9778), .ZN(n_257_76_9990));
   INV_X1 i_257_76_10008 (.A(n_257_76_9990), .ZN(n_257_76_9991));
   NAND3_X1 i_257_76_10009 (.A1(n_257_449), .A2(n_257_76_9785), .A3(
      n_257_76_9786), .ZN(n_257_76_9992));
   NAND3_X1 i_257_76_10010 (.A1(n_257_76_9787), .A2(n_257_76_9766), .A3(
      n_257_1090), .ZN(n_257_76_9993));
   NOR2_X1 i_257_76_10011 (.A1(n_257_76_9992), .A2(n_257_76_9993), .ZN(
      n_257_76_9994));
   NAND3_X1 i_257_76_10012 (.A1(n_257_76_9991), .A2(n_257_76_9994), .A3(
      n_257_76_9753), .ZN(n_257_76_9995));
   NOR2_X1 i_257_76_10013 (.A1(n_257_76_9995), .A2(n_257_76_9870), .ZN(
      n_257_76_9996));
   NAND3_X1 i_257_76_10014 (.A1(n_257_76_9752), .A2(n_257_76_9996), .A3(
      n_257_76_9793), .ZN(n_257_76_9997));
   NOR2_X1 i_257_76_10015 (.A1(n_257_76_9772), .A2(n_257_76_9997), .ZN(
      n_257_76_9998));
   NAND2_X1 i_257_76_10016 (.A1(n_257_76_18083), .A2(n_257_76_9998), .ZN(
      n_257_76_9999));
   NAND3_X1 i_257_76_10017 (.A1(n_257_76_18028), .A2(n_257_76_9822), .A3(
      n_257_429), .ZN(n_257_76_10000));
   NOR2_X1 i_257_76_10018 (.A1(n_257_76_9916), .A2(n_257_76_10000), .ZN(
      n_257_76_10001));
   NAND4_X1 i_257_76_10019 (.A1(n_257_76_10001), .A2(n_257_76_9881), .A3(
      n_257_76_9778), .A4(n_257_76_9831), .ZN(n_257_76_10002));
   NOR2_X1 i_257_76_10020 (.A1(n_257_76_10002), .A2(n_257_76_9889), .ZN(
      n_257_76_10003));
   INV_X1 i_257_76_10021 (.A(n_257_76_9877), .ZN(n_257_76_10004));
   NAND4_X1 i_257_76_10022 (.A1(n_257_76_10003), .A2(n_257_76_9921), .A3(
      n_257_76_10004), .A4(n_257_169), .ZN(n_257_76_10005));
   INV_X1 i_257_76_10023 (.A(n_257_76_9848), .ZN(n_257_76_10006));
   NOR2_X1 i_257_76_10024 (.A1(n_257_76_10005), .A2(n_257_76_10006), .ZN(
      n_257_76_10007));
   NAND3_X1 i_257_76_10025 (.A1(n_257_76_10007), .A2(n_257_76_9894), .A3(
      n_257_76_9762), .ZN(n_257_76_10008));
   INV_X1 i_257_76_10026 (.A(n_257_76_10008), .ZN(n_257_76_10009));
   NAND2_X1 i_257_76_10027 (.A1(n_257_76_18061), .A2(n_257_76_10009), .ZN(
      n_257_76_10010));
   NAND3_X1 i_257_76_10028 (.A1(n_257_76_9989), .A2(n_257_76_9999), .A3(
      n_257_76_10010), .ZN(n_257_76_10011));
   INV_X1 i_257_76_10029 (.A(n_257_76_10011), .ZN(n_257_76_10012));
   NAND3_X1 i_257_76_10030 (.A1(n_257_76_9766), .A2(n_257_438), .A3(n_257_1082), 
      .ZN(n_257_76_10013));
   NOR2_X1 i_257_76_10031 (.A1(n_257_76_10013), .A2(n_257_76_9809), .ZN(
      n_257_76_10014));
   NAND3_X1 i_257_76_10032 (.A1(n_257_76_9774), .A2(n_257_76_9753), .A3(
      n_257_76_10014), .ZN(n_257_76_10015));
   INV_X1 i_257_76_10033 (.A(n_257_76_10015), .ZN(n_257_76_10016));
   NAND2_X1 i_257_76_10034 (.A1(n_257_76_9752), .A2(n_257_76_10016), .ZN(
      n_257_76_10017));
   INV_X1 i_257_76_10035 (.A(n_257_76_10017), .ZN(n_257_76_10018));
   NAND2_X1 i_257_76_10036 (.A1(n_257_76_10018), .A2(n_257_76_9762), .ZN(
      n_257_76_10019));
   INV_X1 i_257_76_10037 (.A(n_257_76_10019), .ZN(n_257_76_10020));
   NAND2_X1 i_257_76_10038 (.A1(n_257_76_18067), .A2(n_257_76_10020), .ZN(
      n_257_76_10021));
   NAND2_X1 i_257_76_10039 (.A1(n_257_366), .A2(n_257_421), .ZN(n_257_76_10022));
   NAND4_X1 i_257_76_10040 (.A1(n_257_76_9819), .A2(n_257_76_10022), .A3(
      n_257_76_9773), .A4(n_257_76_9820), .ZN(n_257_76_10023));
   INV_X1 i_257_76_10041 (.A(n_257_76_10023), .ZN(n_257_76_10024));
   NAND2_X1 i_257_76_10042 (.A1(n_257_289), .A2(n_257_423), .ZN(n_257_76_10025));
   NAND3_X1 i_257_76_10043 (.A1(n_257_76_9753), .A2(n_257_76_9839), .A3(
      n_257_76_10025), .ZN(n_257_76_10026));
   NOR2_X1 i_257_76_10044 (.A1(n_257_76_9842), .A2(n_257_76_10026), .ZN(
      n_257_76_10027));
   NAND2_X1 i_257_76_10045 (.A1(n_257_442), .A2(n_257_486), .ZN(n_257_76_10028));
   NAND4_X1 i_257_76_10046 (.A1(n_257_76_18029), .A2(n_257_76_9822), .A3(
      n_257_420), .A4(n_257_76_9823), .ZN(n_257_76_10029));
   INV_X1 i_257_76_10047 (.A(n_257_76_10029), .ZN(n_257_76_10030));
   NAND2_X1 i_257_76_10048 (.A1(n_257_327), .A2(n_257_422), .ZN(n_257_76_10031));
   NAND3_X1 i_257_76_10049 (.A1(n_257_76_10030), .A2(n_257_76_10031), .A3(
      n_257_76_9832), .ZN(n_257_76_10032));
   NAND3_X1 i_257_76_10050 (.A1(n_257_76_9785), .A2(n_257_76_9786), .A3(
      n_257_76_9787), .ZN(n_257_76_10033));
   NOR2_X1 i_257_76_10051 (.A1(n_257_76_10032), .A2(n_257_76_10033), .ZN(
      n_257_76_10034));
   NAND3_X1 i_257_76_10052 (.A1(n_257_76_9828), .A2(n_257_76_9781), .A3(
      n_257_76_9782), .ZN(n_257_76_10035));
   INV_X1 i_257_76_10053 (.A(n_257_76_10035), .ZN(n_257_76_10036));
   NAND3_X1 i_257_76_10054 (.A1(n_257_76_9777), .A2(n_257_76_9778), .A3(
      n_257_76_9831), .ZN(n_257_76_10037));
   INV_X1 i_257_76_10055 (.A(n_257_76_10037), .ZN(n_257_76_10038));
   NAND3_X1 i_257_76_10056 (.A1(n_257_76_10034), .A2(n_257_76_10036), .A3(
      n_257_76_10038), .ZN(n_257_76_10039));
   INV_X1 i_257_76_10057 (.A(n_257_76_10039), .ZN(n_257_76_10040));
   NAND3_X1 i_257_76_10058 (.A1(n_257_76_10024), .A2(n_257_76_10027), .A3(
      n_257_76_10040), .ZN(n_257_76_10041));
   NAND2_X1 i_257_76_10059 (.A1(n_257_76_9844), .A2(n_257_76_9845), .ZN(
      n_257_76_10042));
   NOR2_X1 i_257_76_10060 (.A1(n_257_76_10041), .A2(n_257_76_10042), .ZN(
      n_257_76_10043));
   NAND3_X1 i_257_76_10061 (.A1(n_257_76_10043), .A2(n_257_76_9850), .A3(
      n_257_76_9762), .ZN(n_257_76_10044));
   INV_X1 i_257_76_10062 (.A(n_257_76_10044), .ZN(n_257_76_10045));
   NAND2_X1 i_257_76_10063 (.A1(n_257_76_18073), .A2(n_257_76_10045), .ZN(
      n_257_76_10046));
   INV_X1 i_257_76_10064 (.A(n_257_614), .ZN(n_257_76_10047));
   NAND2_X1 i_257_76_10065 (.A1(n_257_76_17925), .A2(n_257_76_10047), .ZN(
      n_257_76_10048));
   AOI21_X1 i_257_76_10066 (.A(n_257_1076), .B1(n_257_76_15482), .B2(
      n_257_76_10048), .ZN(n_257_76_10049));
   NAND4_X1 i_257_76_10067 (.A1(n_257_76_10049), .A2(n_257_76_9785), .A3(
      n_257_76_9786), .A4(n_257_76_9787), .ZN(n_257_76_10050));
   NOR2_X1 i_257_76_10068 (.A1(n_257_76_9943), .A2(n_257_76_10050), .ZN(
      n_257_76_10051));
   NAND4_X1 i_257_76_10069 (.A1(n_257_130), .A2(n_257_76_9781), .A3(
      n_257_76_9782), .A4(n_257_76_9777), .ZN(n_257_76_10052));
   INV_X1 i_257_76_10070 (.A(n_257_76_10052), .ZN(n_257_76_10053));
   NAND3_X1 i_257_76_10071 (.A1(n_257_76_10051), .A2(n_257_76_10053), .A3(
      n_257_76_9949), .ZN(n_257_76_10054));
   NOR2_X1 i_257_76_10072 (.A1(n_257_76_10054), .A2(n_257_76_9952), .ZN(
      n_257_76_10055));
   NAND4_X1 i_257_76_10073 (.A1(n_257_76_10055), .A2(n_257_76_9752), .A3(
      n_257_76_9793), .A4(n_257_76_9848), .ZN(n_257_76_10056));
   NOR2_X1 i_257_76_10074 (.A1(n_257_76_10056), .A2(n_257_76_9772), .ZN(
      n_257_76_10057));
   NAND2_X1 i_257_76_10075 (.A1(n_257_76_18068), .A2(n_257_76_10057), .ZN(
      n_257_76_10058));
   NAND3_X1 i_257_76_10076 (.A1(n_257_76_10021), .A2(n_257_76_10046), .A3(
      n_257_76_10058), .ZN(n_257_76_10059));
   INV_X1 i_257_76_10077 (.A(n_257_76_10059), .ZN(n_257_76_10060));
   NAND2_X1 i_257_76_10078 (.A1(n_257_447), .A2(n_257_76_9785), .ZN(
      n_257_76_10061));
   INV_X1 i_257_76_10079 (.A(n_257_76_10061), .ZN(n_257_76_10062));
   NAND2_X1 i_257_76_10080 (.A1(n_257_782), .A2(n_257_442), .ZN(n_257_76_10063));
   NOR2_X1 i_257_76_10081 (.A1(n_257_1076), .A2(n_257_76_10063), .ZN(
      n_257_76_10064));
   NAND2_X1 i_257_76_10082 (.A1(n_257_76_9786), .A2(n_257_76_10064), .ZN(
      n_257_76_10065));
   INV_X1 i_257_76_10083 (.A(n_257_76_10065), .ZN(n_257_76_10066));
   NAND4_X1 i_257_76_10084 (.A1(n_257_76_10062), .A2(n_257_76_10066), .A3(
      n_257_76_9781), .A4(n_257_76_9782), .ZN(n_257_76_10067));
   NOR2_X1 i_257_76_10085 (.A1(n_257_76_9938), .A2(n_257_76_10067), .ZN(
      n_257_76_10068));
   NAND2_X1 i_257_76_10086 (.A1(n_257_76_9752), .A2(n_257_76_10068), .ZN(
      n_257_76_10069));
   INV_X1 i_257_76_10087 (.A(n_257_76_10069), .ZN(n_257_76_10070));
   NAND2_X1 i_257_76_10088 (.A1(n_257_76_10070), .A2(n_257_76_9762), .ZN(
      n_257_76_10071));
   INV_X1 i_257_76_10089 (.A(n_257_76_10071), .ZN(n_257_76_10072));
   INV_X1 i_257_76_10090 (.A(n_257_76_9870), .ZN(n_257_76_10073));
   NAND2_X1 i_257_76_10091 (.A1(n_257_92), .A2(n_257_76_10073), .ZN(
      n_257_76_10074));
   INV_X1 i_257_76_10092 (.A(n_257_76_10074), .ZN(n_257_76_10075));
   NAND4_X1 i_257_76_10093 (.A1(n_257_76_9841), .A2(n_257_76_9753), .A3(
      n_257_76_9839), .A4(n_257_76_9781), .ZN(n_257_76_10076));
   NAND2_X1 i_257_76_10094 (.A1(n_257_76_9782), .A2(n_257_76_9777), .ZN(
      n_257_76_10077));
   INV_X1 i_257_76_10095 (.A(n_257_76_10077), .ZN(n_257_76_10078));
   INV_X1 i_257_76_10096 (.A(n_257_76_9943), .ZN(n_257_76_10079));
   NAND2_X1 i_257_76_10097 (.A1(n_257_76_17932), .A2(n_257_76_10047), .ZN(
      n_257_76_10080));
   AOI21_X1 i_257_76_10098 (.A(n_257_1076), .B1(n_257_76_15507), .B2(
      n_257_76_10080), .ZN(n_257_76_10081));
   NAND4_X1 i_257_76_10099 (.A1(n_257_76_10081), .A2(n_257_76_9785), .A3(
      n_257_76_9786), .A4(n_257_76_9787), .ZN(n_257_76_10082));
   INV_X1 i_257_76_10100 (.A(n_257_76_10082), .ZN(n_257_76_10083));
   NAND3_X1 i_257_76_10101 (.A1(n_257_76_10078), .A2(n_257_76_10079), .A3(
      n_257_76_10083), .ZN(n_257_76_10084));
   NOR2_X1 i_257_76_10102 (.A1(n_257_76_10076), .A2(n_257_76_10084), .ZN(
      n_257_76_10085));
   NAND4_X1 i_257_76_10103 (.A1(n_257_76_9752), .A2(n_257_76_10075), .A3(
      n_257_76_10085), .A4(n_257_76_9793), .ZN(n_257_76_10086));
   NOR2_X1 i_257_76_10104 (.A1(n_257_76_10086), .A2(n_257_76_9772), .ZN(
      n_257_76_10087));
   AOI22_X1 i_257_76_10105 (.A1(n_257_76_18085), .A2(n_257_76_10072), .B1(
      n_257_76_18080), .B2(n_257_76_10087), .ZN(n_257_76_10088));
   NAND3_X1 i_257_76_10106 (.A1(n_257_76_10012), .A2(n_257_76_10060), .A3(
      n_257_76_10088), .ZN(n_257_76_10089));
   OAI21_X1 i_257_76_10107 (.A(n_257_76_17761), .B1(n_257_718), .B2(
      n_257_76_17412), .ZN(n_257_76_10090));
   NAND4_X1 i_257_76_10108 (.A1(n_257_76_10090), .A2(n_257_76_9785), .A3(
      n_257_76_9786), .A4(n_257_76_9822), .ZN(n_257_76_10091));
   INV_X1 i_257_76_10109 (.A(n_257_76_9781), .ZN(n_257_76_10092));
   NOR2_X1 i_257_76_10110 (.A1(n_257_76_10091), .A2(n_257_76_10092), .ZN(
      n_257_76_10093));
   NAND2_X1 i_257_76_10111 (.A1(n_257_76_9773), .A2(n_257_76_10093), .ZN(
      n_257_76_10094));
   NAND3_X1 i_257_76_10112 (.A1(n_257_76_9782), .A2(n_257_76_9778), .A3(
      n_257_448), .ZN(n_257_76_10095));
   INV_X1 i_257_76_10113 (.A(n_257_76_10095), .ZN(n_257_76_10096));
   NAND4_X1 i_257_76_10114 (.A1(n_257_76_10096), .A2(n_257_76_9774), .A3(
      n_257_76_9775), .A4(n_257_76_9753), .ZN(n_257_76_10097));
   NOR2_X1 i_257_76_10115 (.A1(n_257_76_10094), .A2(n_257_76_10097), .ZN(
      n_257_76_10098));
   NAND3_X1 i_257_76_10116 (.A1(n_257_76_10098), .A2(n_257_76_9752), .A3(
      n_257_686), .ZN(n_257_76_10099));
   NOR2_X1 i_257_76_10117 (.A1(n_257_76_10099), .A2(n_257_76_9772), .ZN(
      n_257_76_10100));
   NAND2_X1 i_257_76_10118 (.A1(n_257_76_18079), .A2(n_257_76_10100), .ZN(
      n_257_76_10101));
   NAND2_X1 i_257_76_10119 (.A1(n_257_76_9832), .A2(n_257_76_9785), .ZN(
      n_257_76_10102));
   INV_X1 i_257_76_10120 (.A(n_257_76_10102), .ZN(n_257_76_10103));
   NAND2_X1 i_257_76_10121 (.A1(n_257_76_9786), .A2(n_257_76_9787), .ZN(
      n_257_76_10104));
   INV_X1 i_257_76_10122 (.A(n_257_76_10104), .ZN(n_257_76_10105));
   NAND4_X1 i_257_76_10123 (.A1(n_257_76_18027), .A2(n_257_76_9822), .A3(
      n_257_76_9823), .A4(n_257_425), .ZN(n_257_76_10106));
   INV_X1 i_257_76_10124 (.A(n_257_76_10106), .ZN(n_257_76_10107));
   NAND4_X1 i_257_76_10125 (.A1(n_257_76_10103), .A2(n_257_76_10105), .A3(
      n_257_76_9831), .A4(n_257_76_10107), .ZN(n_257_76_10108));
   INV_X1 i_257_76_10126 (.A(n_257_76_10108), .ZN(n_257_76_10109));
   NAND4_X1 i_257_76_10127 (.A1(n_257_76_9781), .A2(n_257_76_9782), .A3(
      n_257_76_9777), .A4(n_257_76_9778), .ZN(n_257_76_10110));
   INV_X1 i_257_76_10128 (.A(n_257_76_10110), .ZN(n_257_76_10111));
   NAND2_X1 i_257_76_10129 (.A1(n_257_76_10109), .A2(n_257_76_10111), .ZN(
      n_257_76_10112));
   NOR3_X1 i_257_76_10130 (.A1(n_257_76_10112), .A2(n_257_76_9877), .A3(
      n_257_76_9878), .ZN(n_257_76_10113));
   INV_X1 i_257_76_10131 (.A(n_257_76_9844), .ZN(n_257_76_10114));
   NAND2_X1 i_257_76_10132 (.A1(n_257_249), .A2(n_257_76_9819), .ZN(
      n_257_76_10115));
   NOR2_X1 i_257_76_10133 (.A1(n_257_76_10114), .A2(n_257_76_10115), .ZN(
      n_257_76_10116));
   NAND4_X1 i_257_76_10134 (.A1(n_257_76_10113), .A2(n_257_76_10116), .A3(
      n_257_76_9793), .A4(n_257_76_9848), .ZN(n_257_76_10117));
   NAND2_X1 i_257_76_10135 (.A1(n_257_76_9762), .A2(n_257_76_9752), .ZN(
      n_257_76_10118));
   NOR2_X1 i_257_76_10136 (.A1(n_257_76_10117), .A2(n_257_76_10118), .ZN(
      n_257_76_10119));
   NAND2_X1 i_257_76_10137 (.A1(n_257_76_18064), .A2(n_257_76_10119), .ZN(
      n_257_76_10120));
   NAND3_X1 i_257_76_10138 (.A1(n_257_76_10031), .A2(n_257_76_9832), .A3(
      n_257_76_9785), .ZN(n_257_76_10121));
   INV_X1 i_257_76_10139 (.A(n_257_76_10121), .ZN(n_257_76_10122));
   NAND3_X1 i_257_76_10140 (.A1(n_257_76_9822), .A2(n_257_76_9823), .A3(
      n_257_421), .ZN(n_257_76_10123));
   INV_X1 i_257_76_10141 (.A(n_257_76_10123), .ZN(n_257_76_10124));
   NAND4_X1 i_257_76_10142 (.A1(n_257_76_9786), .A2(n_257_76_10124), .A3(
      n_257_76_9787), .A4(n_257_76_18027), .ZN(n_257_76_10125));
   INV_X1 i_257_76_10143 (.A(n_257_76_10125), .ZN(n_257_76_10126));
   NAND2_X1 i_257_76_10144 (.A1(n_257_76_10122), .A2(n_257_76_10126), .ZN(
      n_257_76_10127));
   NOR3_X1 i_257_76_10145 (.A1(n_257_76_10127), .A2(n_257_76_10035), .A3(
      n_257_76_10037), .ZN(n_257_76_10128));
   INV_X1 i_257_76_10146 (.A(n_257_76_9821), .ZN(n_257_76_10129));
   NAND2_X1 i_257_76_10147 (.A1(n_257_76_9774), .A2(n_257_76_9775), .ZN(
      n_257_76_10130));
   NAND3_X1 i_257_76_10148 (.A1(n_257_76_9839), .A2(n_257_366), .A3(
      n_257_76_10025), .ZN(n_257_76_10131));
   NOR2_X1 i_257_76_10149 (.A1(n_257_76_10130), .A2(n_257_76_10131), .ZN(
      n_257_76_10132));
   NAND3_X1 i_257_76_10150 (.A1(n_257_76_10128), .A2(n_257_76_10129), .A3(
      n_257_76_10132), .ZN(n_257_76_10133));
   INV_X1 i_257_76_10151 (.A(n_257_76_10133), .ZN(n_257_76_10134));
   NAND4_X1 i_257_76_10152 (.A1(n_257_76_9848), .A2(n_257_76_9844), .A3(
      n_257_76_9845), .A4(n_257_76_9927), .ZN(n_257_76_10135));
   INV_X1 i_257_76_10153 (.A(n_257_76_10135), .ZN(n_257_76_10136));
   NAND4_X1 i_257_76_10154 (.A1(n_257_76_10134), .A2(n_257_76_10136), .A3(
      n_257_76_9894), .A4(n_257_76_9762), .ZN(n_257_76_10137));
   INV_X1 i_257_76_10155 (.A(n_257_76_10137), .ZN(n_257_76_10138));
   NAND2_X1 i_257_76_10156 (.A1(n_257_76_18082), .A2(n_257_76_10138), .ZN(
      n_257_76_10139));
   NAND3_X1 i_257_76_10157 (.A1(n_257_76_10101), .A2(n_257_76_10120), .A3(
      n_257_76_10139), .ZN(n_257_76_10140));
   INV_X1 i_257_76_10158 (.A(n_257_76_10140), .ZN(n_257_76_10141));
   NAND4_X1 i_257_76_10159 (.A1(n_257_76_18027), .A2(n_257_427), .A3(
      n_257_76_9822), .A4(n_257_76_9823), .ZN(n_257_76_10142));
   INV_X1 i_257_76_10160 (.A(n_257_209), .ZN(n_257_76_10143));
   NOR2_X1 i_257_76_10161 (.A1(n_257_76_10142), .A2(n_257_76_10143), .ZN(
      n_257_76_10144));
   INV_X1 i_257_76_10162 (.A(n_257_76_10033), .ZN(n_257_76_10145));
   NAND4_X1 i_257_76_10163 (.A1(n_257_76_10144), .A2(n_257_76_10145), .A3(
      n_257_76_9781), .A4(n_257_76_9831), .ZN(n_257_76_10146));
   NOR2_X1 i_257_76_10164 (.A1(n_257_76_9878), .A2(n_257_76_10146), .ZN(
      n_257_76_10147));
   NAND3_X1 i_257_76_10165 (.A1(n_257_76_9775), .A2(n_257_76_9841), .A3(
      n_257_76_9753), .ZN(n_257_76_10148));
   NAND4_X1 i_257_76_10166 (.A1(n_257_76_9839), .A2(n_257_76_9782), .A3(
      n_257_76_9777), .A4(n_257_76_9778), .ZN(n_257_76_10149));
   NOR2_X1 i_257_76_10167 (.A1(n_257_76_10148), .A2(n_257_76_10149), .ZN(
      n_257_76_10150));
   NAND4_X1 i_257_76_10168 (.A1(n_257_76_9848), .A2(n_257_76_10147), .A3(
      n_257_76_10150), .A4(n_257_76_9844), .ZN(n_257_76_10151));
   INV_X1 i_257_76_10169 (.A(n_257_76_10151), .ZN(n_257_76_10152));
   NAND3_X1 i_257_76_10170 (.A1(n_257_76_10152), .A2(n_257_76_9894), .A3(
      n_257_76_9762), .ZN(n_257_76_10153));
   INV_X1 i_257_76_10171 (.A(n_257_76_10153), .ZN(n_257_76_10154));
   NAND2_X1 i_257_76_10172 (.A1(n_257_76_18065), .A2(n_257_76_10154), .ZN(
      n_257_76_10155));
   NAND4_X1 i_257_76_10173 (.A1(n_257_76_10093), .A2(n_257_76_9773), .A3(
      n_257_76_9774), .A4(n_257_76_9775), .ZN(n_257_76_10156));
   NAND3_X1 i_257_76_10174 (.A1(n_257_469), .A2(n_257_76_9777), .A3(
      n_257_76_9778), .ZN(n_257_76_10157));
   INV_X1 i_257_76_10175 (.A(n_257_76_10157), .ZN(n_257_76_10158));
   NAND2_X1 i_257_76_10176 (.A1(n_257_451), .A2(n_257_76_9782), .ZN(
      n_257_76_10159));
   INV_X1 i_257_76_10177 (.A(n_257_76_10159), .ZN(n_257_76_10160));
   NAND4_X1 i_257_76_10178 (.A1(n_257_76_10158), .A2(n_257_76_10160), .A3(
      n_257_76_9753), .A4(n_257_76_9839), .ZN(n_257_76_10161));
   NOR2_X1 i_257_76_10179 (.A1(n_257_76_10156), .A2(n_257_76_10161), .ZN(
      n_257_76_10162));
   NAND3_X1 i_257_76_10180 (.A1(n_257_76_10162), .A2(n_257_76_9752), .A3(
      n_257_76_9793), .ZN(n_257_76_10163));
   NOR2_X1 i_257_76_10181 (.A1(n_257_76_10163), .A2(n_257_76_9772), .ZN(
      n_257_76_10164));
   NAND2_X1 i_257_76_10182 (.A1(n_257_76_18063), .A2(n_257_76_10164), .ZN(
      n_257_76_10165));
   NAND3_X1 i_257_76_10183 (.A1(n_257_518), .A2(n_257_76_9832), .A3(
      n_257_76_9785), .ZN(n_257_76_10166));
   INV_X1 i_257_76_10184 (.A(n_257_76_10166), .ZN(n_257_76_10167));
   NAND3_X1 i_257_76_10185 (.A1(n_257_76_9822), .A2(n_257_76_9823), .A3(
      n_257_424), .ZN(n_257_76_10168));
   INV_X1 i_257_76_10186 (.A(n_257_76_10168), .ZN(n_257_76_10169));
   NAND4_X1 i_257_76_10187 (.A1(n_257_76_9786), .A2(n_257_76_10169), .A3(
      n_257_76_9787), .A4(n_257_76_18027), .ZN(n_257_76_10170));
   INV_X1 i_257_76_10188 (.A(n_257_76_10170), .ZN(n_257_76_10171));
   NAND4_X1 i_257_76_10189 (.A1(n_257_76_10167), .A2(n_257_76_10171), .A3(
      n_257_76_9781), .A4(n_257_76_9831), .ZN(n_257_76_10172));
   NOR2_X1 i_257_76_10190 (.A1(n_257_76_9821), .A2(n_257_76_10172), .ZN(
      n_257_76_10173));
   NAND4_X1 i_257_76_10191 (.A1(n_257_76_10173), .A2(n_257_76_9843), .A3(
      n_257_76_9844), .A4(n_257_76_9845), .ZN(n_257_76_10174));
   INV_X1 i_257_76_10192 (.A(n_257_76_10174), .ZN(n_257_76_10175));
   NAND3_X1 i_257_76_10193 (.A1(n_257_76_10175), .A2(n_257_76_9850), .A3(
      n_257_76_9762), .ZN(n_257_76_10176));
   INV_X1 i_257_76_10194 (.A(n_257_76_10176), .ZN(n_257_76_10177));
   NAND2_X1 i_257_76_10195 (.A1(n_257_76_18062), .A2(n_257_76_10177), .ZN(
      n_257_76_10178));
   NAND3_X1 i_257_76_10196 (.A1(n_257_76_10155), .A2(n_257_76_10165), .A3(
      n_257_76_10178), .ZN(n_257_76_10179));
   INV_X1 i_257_76_10197 (.A(n_257_76_10179), .ZN(n_257_76_10180));
   NAND4_X1 i_257_76_10198 (.A1(n_257_76_9819), .A2(n_257_76_9773), .A3(
      n_257_76_9820), .A4(n_257_76_9774), .ZN(n_257_76_10181));
   INV_X1 i_257_76_10199 (.A(n_257_76_10181), .ZN(n_257_76_10182));
   NAND2_X1 i_257_76_10200 (.A1(n_257_76_10025), .A2(n_257_76_9828), .ZN(
      n_257_76_10183));
   INV_X1 i_257_76_10201 (.A(n_257_76_10183), .ZN(n_257_76_10184));
   NAND3_X1 i_257_76_10202 (.A1(n_257_76_9822), .A2(n_257_76_9823), .A3(
      n_257_422), .ZN(n_257_76_10185));
   INV_X1 i_257_76_10203 (.A(n_257_76_10185), .ZN(n_257_76_10186));
   NAND3_X1 i_257_76_10204 (.A1(n_257_76_10186), .A2(n_257_327), .A3(
      n_257_76_18027), .ZN(n_257_76_10187));
   NOR2_X1 i_257_76_10205 (.A1(n_257_76_10033), .A2(n_257_76_10187), .ZN(
      n_257_76_10188));
   NAND3_X1 i_257_76_10206 (.A1(n_257_76_9781), .A2(n_257_76_9831), .A3(
      n_257_76_9832), .ZN(n_257_76_10189));
   INV_X1 i_257_76_10207 (.A(n_257_76_10189), .ZN(n_257_76_10190));
   NAND3_X1 i_257_76_10208 (.A1(n_257_76_10184), .A2(n_257_76_10188), .A3(
      n_257_76_10190), .ZN(n_257_76_10191));
   INV_X1 i_257_76_10209 (.A(n_257_76_10191), .ZN(n_257_76_10192));
   NAND3_X1 i_257_76_10210 (.A1(n_257_76_10150), .A2(n_257_76_10182), .A3(
      n_257_76_10192), .ZN(n_257_76_10193));
   NOR2_X1 i_257_76_10211 (.A1(n_257_76_10193), .A2(n_257_76_10042), .ZN(
      n_257_76_10194));
   NAND3_X1 i_257_76_10212 (.A1(n_257_76_10194), .A2(n_257_76_9850), .A3(
      n_257_76_9762), .ZN(n_257_76_10195));
   INV_X1 i_257_76_10213 (.A(n_257_76_10195), .ZN(n_257_76_10196));
   NAND2_X1 i_257_76_10214 (.A1(n_257_342), .A2(n_257_76_10196), .ZN(
      n_257_76_10197));
   NAND3_X1 i_257_76_10215 (.A1(n_257_76_9819), .A2(n_257_76_10022), .A3(
      n_257_76_9773), .ZN(n_257_76_10198));
   INV_X1 i_257_76_10216 (.A(n_257_76_10198), .ZN(n_257_76_10199));
   NAND3_X1 i_257_76_10217 (.A1(n_257_76_9820), .A2(n_257_76_9774), .A3(
      n_257_76_9775), .ZN(n_257_76_10200));
   INV_X1 i_257_76_10218 (.A(n_257_76_10200), .ZN(n_257_76_10201));
   NAND4_X1 i_257_76_10219 (.A1(n_257_76_9841), .A2(n_257_76_9753), .A3(
      n_257_76_9839), .A4(n_257_76_10025), .ZN(n_257_76_10202));
   INV_X1 i_257_76_10220 (.A(n_257_76_10202), .ZN(n_257_76_10203));
   NAND3_X1 i_257_76_10221 (.A1(n_257_76_10199), .A2(n_257_76_10201), .A3(
      n_257_76_10203), .ZN(n_257_76_10204));
   NOR2_X1 i_257_76_10222 (.A1(n_257_76_10042), .A2(n_257_76_10204), .ZN(
      n_257_76_10205));
   NAND2_X1 i_257_76_10223 (.A1(n_257_582), .A2(n_257_428), .ZN(n_257_76_10206));
   NAND3_X1 i_257_76_10224 (.A1(n_257_405), .A2(n_257_484), .A3(n_257_442), 
      .ZN(n_257_76_10207));
   INV_X1 i_257_76_10225 (.A(n_257_76_10207), .ZN(n_257_76_10208));
   NAND4_X1 i_257_76_10226 (.A1(n_257_76_9822), .A2(n_257_76_9823), .A3(
      n_257_76_10206), .A4(n_257_76_10208), .ZN(n_257_76_10209));
   INV_X1 i_257_76_10227 (.A(n_257_76_10209), .ZN(n_257_76_10210));
   NAND2_X1 i_257_76_10228 (.A1(n_257_420), .A2(n_257_486), .ZN(n_257_76_10211));
   NAND4_X1 i_257_76_10229 (.A1(n_257_76_9786), .A2(n_257_76_10210), .A3(
      n_257_76_9787), .A4(n_257_76_10211), .ZN(n_257_76_10212));
   INV_X1 i_257_76_10230 (.A(n_257_76_10212), .ZN(n_257_76_10213));
   NAND2_X1 i_257_76_10231 (.A1(n_257_76_10122), .A2(n_257_76_10213), .ZN(
      n_257_76_10214));
   NOR3_X1 i_257_76_10232 (.A1(n_257_76_10214), .A2(n_257_76_10035), .A3(
      n_257_76_10037), .ZN(n_257_76_10215));
   NAND2_X1 i_257_76_10233 (.A1(n_257_76_9752), .A2(n_257_76_10215), .ZN(
      n_257_76_10216));
   INV_X1 i_257_76_10234 (.A(n_257_76_10216), .ZN(n_257_76_10217));
   NAND2_X1 i_257_76_10235 (.A1(n_257_76_9793), .A2(n_257_76_9848), .ZN(
      n_257_76_10218));
   INV_X1 i_257_76_10236 (.A(n_257_76_10218), .ZN(n_257_76_10219));
   NAND4_X1 i_257_76_10237 (.A1(n_257_76_10205), .A2(n_257_76_10217), .A3(
      n_257_76_9762), .A4(n_257_76_10219), .ZN(n_257_76_10220));
   INV_X1 i_257_76_10238 (.A(n_257_76_10220), .ZN(n_257_76_10221));
   NAND2_X1 i_257_76_10239 (.A1(n_257_76_18060), .A2(n_257_76_10221), .ZN(
      n_257_76_10222));
   INV_X1 i_257_76_10240 (.A(n_257_76_9798), .ZN(n_257_76_10223));
   AOI22_X1 i_257_76_10241 (.A1(n_257_446), .A2(n_257_76_10223), .B1(n_257_449), 
      .B2(n_257_76_17546), .ZN(n_257_76_10224));
   INV_X1 i_257_76_10242 (.A(n_257_76_10063), .ZN(n_257_76_10225));
   NAND2_X1 i_257_76_10243 (.A1(n_257_447), .A2(n_257_76_10225), .ZN(
      n_257_76_10226));
   NAND2_X1 i_257_76_10244 (.A1(n_257_52), .A2(n_257_76_17918), .ZN(
      n_257_76_10227));
   INV_X1 i_257_76_10245 (.A(Small_Packet_Data_Size[17]), .ZN(n_257_76_10228));
   NAND4_X1 i_257_76_10246 (.A1(n_257_76_9822), .A2(n_257_76_9823), .A3(
      n_257_76_18030), .A4(n_257_76_10206), .ZN(n_257_76_10229));
   NAND2_X1 i_257_76_10247 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[17]), 
      .ZN(n_257_76_10230));
   NAND2_X1 i_257_76_10248 (.A1(n_257_76_10229), .A2(n_257_76_10230), .ZN(
      n_257_76_10231));
   NAND3_X1 i_257_76_10249 (.A1(n_257_76_10226), .A2(n_257_76_10227), .A3(
      n_257_76_10231), .ZN(n_257_76_10232));
   INV_X1 i_257_76_10250 (.A(n_257_76_10232), .ZN(n_257_76_10233));
   NAND3_X1 i_257_76_10251 (.A1(n_257_438), .A2(n_257_1082), .A3(n_257_442), 
      .ZN(n_257_76_10234));
   INV_X1 i_257_76_10252 (.A(n_257_76_9754), .ZN(n_257_76_10235));
   NAND2_X1 i_257_76_10253 (.A1(n_257_440), .A2(n_257_76_10235), .ZN(
      n_257_76_10236));
   NAND2_X1 i_257_76_10254 (.A1(n_257_718), .A2(n_257_76_15655), .ZN(
      n_257_76_10237));
   NAND4_X1 i_257_76_10255 (.A1(n_257_76_10234), .A2(n_257_76_10236), .A3(
      n_257_76_10029), .A4(n_257_76_10237), .ZN(n_257_76_10238));
   INV_X1 i_257_76_10256 (.A(n_257_76_10238), .ZN(n_257_76_10239));
   NAND3_X1 i_257_76_10257 (.A1(n_257_76_10224), .A2(n_257_76_10233), .A3(
      n_257_76_10239), .ZN(n_257_76_10240));
   NAND2_X1 i_257_76_10258 (.A1(n_257_814), .A2(n_257_76_17952), .ZN(
      n_257_76_10241));
   NAND3_X1 i_257_76_10259 (.A1(n_257_441), .A2(n_257_980), .A3(n_257_442), 
      .ZN(n_257_76_10242));
   NAND2_X1 i_257_76_10260 (.A1(n_257_646), .A2(n_257_76_17928), .ZN(
      n_257_76_10243));
   NAND2_X1 i_257_76_10261 (.A1(n_257_878), .A2(n_257_76_17903), .ZN(
      n_257_76_10244));
   NAND4_X1 i_257_76_10262 (.A1(n_257_76_10241), .A2(n_257_76_10242), .A3(
      n_257_76_10243), .A4(n_257_76_10244), .ZN(n_257_76_10245));
   NOR2_X1 i_257_76_10263 (.A1(n_257_76_10240), .A2(n_257_76_10245), .ZN(
      n_257_76_10246));
   NAND2_X1 i_257_76_10264 (.A1(n_257_76_9835), .A2(n_257_76_10172), .ZN(
      n_257_76_10247));
   INV_X1 i_257_76_10265 (.A(n_257_76_10247), .ZN(n_257_76_10248));
   NAND2_X1 i_257_76_10266 (.A1(n_257_750), .A2(n_257_76_17935), .ZN(
      n_257_76_10249));
   NAND2_X1 i_257_76_10267 (.A1(n_257_130), .A2(n_257_76_17925), .ZN(
      n_257_76_10250));
   NAND2_X1 i_257_76_10268 (.A1(n_257_916), .A2(n_257_76_17940), .ZN(
      n_257_76_10251));
   NAND3_X1 i_257_76_10269 (.A1(n_257_76_10249), .A2(n_257_76_10250), .A3(
      n_257_76_10251), .ZN(n_257_76_10252));
   INV_X1 i_257_76_10270 (.A(n_257_76_10146), .ZN(n_257_76_10253));
   NOR2_X1 i_257_76_10271 (.A1(n_257_76_10252), .A2(n_257_76_10253), .ZN(
      n_257_76_10254));
   NAND3_X1 i_257_76_10272 (.A1(n_257_76_10246), .A2(n_257_76_10248), .A3(
      n_257_76_10254), .ZN(n_257_76_10255));
   NAND2_X1 i_257_76_10273 (.A1(n_257_92), .A2(n_257_76_17932), .ZN(
      n_257_76_10256));
   NAND2_X1 i_257_76_10274 (.A1(n_257_169), .A2(n_257_76_17331), .ZN(
      n_257_76_10257));
   NAND3_X1 i_257_76_10275 (.A1(n_257_76_10256), .A2(n_257_76_10257), .A3(
      n_257_76_10191), .ZN(n_257_76_10258));
   NOR2_X1 i_257_76_10276 (.A1(n_257_76_10255), .A2(n_257_76_10258), .ZN(
      n_257_76_10259));
   INV_X1 i_257_76_10277 (.A(n_257_1044), .ZN(n_257_76_10260));
   OAI21_X1 i_257_76_10278 (.A(n_257_76_10133), .B1(n_257_76_10260), .B2(
      n_257_76_17968), .ZN(n_257_76_10261));
   INV_X1 i_257_76_10279 (.A(n_257_76_10261), .ZN(n_257_76_10262));
   NAND2_X1 i_257_76_10280 (.A1(n_257_1012), .A2(n_257_76_17964), .ZN(
      n_257_76_10263));
   INV_X1 i_257_76_10281 (.A(n_257_750), .ZN(n_257_76_10264));
   NAND2_X1 i_257_76_10282 (.A1(n_257_76_10264), .A2(n_257_442), .ZN(
      n_257_76_10265));
   INV_X1 i_257_76_10283 (.A(n_257_916), .ZN(n_257_76_10266));
   NAND2_X1 i_257_76_10284 (.A1(n_257_76_10266), .A2(n_257_442), .ZN(
      n_257_76_10267));
   INV_X1 i_257_76_10285 (.A(n_257_814), .ZN(n_257_76_10268));
   NAND2_X1 i_257_76_10286 (.A1(n_257_76_10268), .A2(n_257_442), .ZN(
      n_257_76_10269));
   NAND4_X1 i_257_76_10287 (.A1(n_257_76_10265), .A2(n_257_76_10267), .A3(
      n_257_76_10269), .A4(n_257_76_13029), .ZN(n_257_76_10270));
   INV_X1 i_257_76_10288 (.A(n_257_76_9841), .ZN(n_257_76_10271));
   NAND2_X1 i_257_76_10289 (.A1(n_257_76_10270), .A2(n_257_76_10271), .ZN(
      n_257_76_10272));
   NAND2_X1 i_257_76_10290 (.A1(n_257_686), .A2(n_257_76_17958), .ZN(
      n_257_76_10273));
   NAND4_X1 i_257_76_10291 (.A1(n_257_76_10263), .A2(n_257_76_9924), .A3(
      n_257_76_10272), .A4(n_257_76_10273), .ZN(n_257_76_10274));
   INV_X1 i_257_76_10292 (.A(n_257_76_10274), .ZN(n_257_76_10275));
   NAND4_X1 i_257_76_10293 (.A1(n_257_76_10259), .A2(n_257_76_10117), .A3(
      n_257_76_10262), .A4(n_257_76_10275), .ZN(n_257_76_10276));
   NAND3_X1 i_257_76_10294 (.A1(n_257_76_10197), .A2(n_257_76_10222), .A3(
      n_257_76_10276), .ZN(n_257_76_10277));
   INV_X1 i_257_76_10295 (.A(n_257_76_10277), .ZN(n_257_76_10278));
   NAND3_X1 i_257_76_10296 (.A1(n_257_76_10141), .A2(n_257_76_10180), .A3(
      n_257_76_10278), .ZN(n_257_76_10279));
   NOR2_X1 i_257_76_10297 (.A1(n_257_76_10089), .A2(n_257_76_10279), .ZN(
      n_257_76_10280));
   NAND2_X1 i_257_76_10298 (.A1(n_257_76_9979), .A2(n_257_76_10280), .ZN(n_17));
   NAND2_X1 i_257_76_10299 (.A1(n_257_1045), .A2(n_257_443), .ZN(n_257_76_10281));
   INV_X1 i_257_76_10300 (.A(n_257_76_10281), .ZN(n_257_76_10282));
   NAND2_X1 i_257_76_10301 (.A1(n_257_1013), .A2(n_257_444), .ZN(n_257_76_10283));
   NAND2_X1 i_257_76_10302 (.A1(n_257_441), .A2(n_257_981), .ZN(n_257_76_10284));
   NAND2_X1 i_257_76_10303 (.A1(n_257_949), .A2(n_257_442), .ZN(n_257_76_10285));
   NOR2_X1 i_257_76_10304 (.A1(n_257_1077), .A2(n_257_76_10285), .ZN(
      n_257_76_10286));
   NAND2_X1 i_257_76_10305 (.A1(n_257_440), .A2(n_257_76_10286), .ZN(
      n_257_76_10287));
   INV_X1 i_257_76_10306 (.A(n_257_76_10287), .ZN(n_257_76_10288));
   NAND2_X1 i_257_76_10307 (.A1(n_257_76_10284), .A2(n_257_76_10288), .ZN(
      n_257_76_10289));
   INV_X1 i_257_76_10308 (.A(n_257_76_10289), .ZN(n_257_76_10290));
   NAND2_X1 i_257_76_10309 (.A1(n_257_76_10283), .A2(n_257_76_10290), .ZN(
      n_257_76_10291));
   NOR2_X1 i_257_76_10310 (.A1(n_257_76_10282), .A2(n_257_76_10291), .ZN(
      n_257_76_10292));
   NAND2_X1 i_257_76_10311 (.A1(n_257_17), .A2(n_257_76_10292), .ZN(
      n_257_76_10293));
   NOR2_X1 i_257_76_10312 (.A1(n_257_1077), .A2(n_257_76_17412), .ZN(
      n_257_76_10294));
   INV_X1 i_257_76_10313 (.A(n_257_76_10294), .ZN(n_257_76_10295));
   NOR2_X1 i_257_76_10314 (.A1(n_257_76_10295), .A2(n_257_76_15197), .ZN(
      n_257_76_10296));
   NAND2_X1 i_257_76_10315 (.A1(n_257_1045), .A2(n_257_76_10296), .ZN(
      n_257_76_10297));
   INV_X1 i_257_76_10316 (.A(n_257_76_10297), .ZN(n_257_76_10298));
   NAND2_X1 i_257_76_10317 (.A1(n_257_76_18072), .A2(n_257_76_10298), .ZN(
      n_257_76_10299));
   NAND2_X1 i_257_76_10318 (.A1(n_257_719), .A2(n_257_435), .ZN(n_257_76_10300));
   NAND3_X1 i_257_76_10319 (.A1(n_257_76_10294), .A2(n_257_76_10300), .A3(
      n_257_450), .ZN(n_257_76_10301));
   INV_X1 i_257_76_10320 (.A(n_257_76_10301), .ZN(n_257_76_10302));
   NAND2_X1 i_257_76_10321 (.A1(n_257_440), .A2(n_257_949), .ZN(n_257_76_10303));
   NAND2_X1 i_257_76_10322 (.A1(n_257_438), .A2(n_257_1083), .ZN(n_257_76_10304));
   NAND4_X1 i_257_76_10323 (.A1(n_257_76_10302), .A2(n_257_76_10303), .A3(
      n_257_647), .A4(n_257_76_10304), .ZN(n_257_76_10305));
   INV_X1 i_257_76_10324 (.A(n_257_76_10305), .ZN(n_257_76_10306));
   NAND2_X1 i_257_76_10325 (.A1(n_257_446), .A2(n_257_847), .ZN(n_257_76_10307));
   NAND2_X1 i_257_76_10326 (.A1(n_257_449), .A2(n_257_893), .ZN(n_257_76_10308));
   NAND2_X1 i_257_76_10327 (.A1(n_257_76_10307), .A2(n_257_76_10308), .ZN(
      n_257_76_10309));
   INV_X1 i_257_76_10328 (.A(n_257_76_10309), .ZN(n_257_76_10310));
   NAND2_X1 i_257_76_10329 (.A1(n_257_447), .A2(n_257_783), .ZN(n_257_76_10311));
   NAND2_X1 i_257_76_10330 (.A1(n_257_879), .A2(n_257_445), .ZN(n_257_76_10312));
   NAND2_X1 i_257_76_10331 (.A1(n_257_76_10311), .A2(n_257_76_10312), .ZN(
      n_257_76_10313));
   INV_X1 i_257_76_10332 (.A(n_257_76_10313), .ZN(n_257_76_10314));
   NAND3_X1 i_257_76_10333 (.A1(n_257_76_10306), .A2(n_257_76_10310), .A3(
      n_257_76_10314), .ZN(n_257_76_10315));
   NAND2_X1 i_257_76_10334 (.A1(n_257_751), .A2(n_257_436), .ZN(n_257_76_10316));
   NAND2_X1 i_257_76_10335 (.A1(n_257_815), .A2(n_257_437), .ZN(n_257_76_10317));
   NAND2_X1 i_257_76_10336 (.A1(n_257_917), .A2(n_257_439), .ZN(n_257_76_10318));
   NAND4_X1 i_257_76_10337 (.A1(n_257_76_10316), .A2(n_257_76_10284), .A3(
      n_257_76_10317), .A4(n_257_76_10318), .ZN(n_257_76_10319));
   NOR2_X1 i_257_76_10338 (.A1(n_257_76_10315), .A2(n_257_76_10319), .ZN(
      n_257_76_10320));
   NAND2_X1 i_257_76_10339 (.A1(n_257_687), .A2(n_257_448), .ZN(n_257_76_10321));
   NAND3_X1 i_257_76_10340 (.A1(n_257_76_10320), .A2(n_257_76_10283), .A3(
      n_257_76_10321), .ZN(n_257_76_10322));
   NOR2_X1 i_257_76_10341 (.A1(n_257_76_10322), .A2(n_257_76_10282), .ZN(
      n_257_76_10323));
   NAND2_X1 i_257_76_10342 (.A1(n_257_28), .A2(n_257_76_10323), .ZN(
      n_257_76_10324));
   NAND3_X1 i_257_76_10343 (.A1(n_257_76_10293), .A2(n_257_76_10299), .A3(
      n_257_76_10324), .ZN(n_257_76_10325));
   NAND2_X1 i_257_76_10344 (.A1(n_257_847), .A2(n_257_442), .ZN(n_257_76_10326));
   NOR2_X1 i_257_76_10345 (.A1(n_257_1077), .A2(n_257_76_10326), .ZN(
      n_257_76_10327));
   NAND3_X1 i_257_76_10346 (.A1(n_257_76_10303), .A2(n_257_76_10304), .A3(
      n_257_76_10327), .ZN(n_257_76_10328));
   INV_X1 i_257_76_10347 (.A(n_257_76_10328), .ZN(n_257_76_10329));
   NAND2_X1 i_257_76_10348 (.A1(n_257_76_10312), .A2(n_257_446), .ZN(
      n_257_76_10330));
   INV_X1 i_257_76_10349 (.A(n_257_76_10330), .ZN(n_257_76_10331));
   NAND4_X1 i_257_76_10350 (.A1(n_257_76_10284), .A2(n_257_76_10329), .A3(
      n_257_76_10318), .A4(n_257_76_10331), .ZN(n_257_76_10332));
   INV_X1 i_257_76_10351 (.A(n_257_76_10332), .ZN(n_257_76_10333));
   NAND2_X1 i_257_76_10352 (.A1(n_257_76_10283), .A2(n_257_76_10333), .ZN(
      n_257_76_10334));
   NOR2_X1 i_257_76_10353 (.A1(n_257_76_10282), .A2(n_257_76_10334), .ZN(
      n_257_76_10335));
   NAND2_X1 i_257_76_10354 (.A1(n_257_76_18070), .A2(n_257_76_10335), .ZN(
      n_257_76_10336));
   NAND2_X1 i_257_76_10355 (.A1(n_257_439), .A2(n_257_76_10294), .ZN(
      n_257_76_10337));
   INV_X1 i_257_76_10356 (.A(n_257_76_10337), .ZN(n_257_76_10338));
   NAND3_X1 i_257_76_10357 (.A1(n_257_76_10338), .A2(n_257_917), .A3(
      n_257_76_10303), .ZN(n_257_76_10339));
   INV_X1 i_257_76_10358 (.A(n_257_76_10339), .ZN(n_257_76_10340));
   NAND2_X1 i_257_76_10359 (.A1(n_257_76_10340), .A2(n_257_76_10284), .ZN(
      n_257_76_10341));
   INV_X1 i_257_76_10360 (.A(n_257_76_10341), .ZN(n_257_76_10342));
   NAND2_X1 i_257_76_10361 (.A1(n_257_76_10283), .A2(n_257_76_10342), .ZN(
      n_257_76_10343));
   NOR2_X1 i_257_76_10362 (.A1(n_257_76_10282), .A2(n_257_76_10343), .ZN(
      n_257_76_10344));
   NAND2_X1 i_257_76_10363 (.A1(n_257_76_18084), .A2(n_257_76_10344), .ZN(
      n_257_76_10345));
   NAND2_X1 i_257_76_10364 (.A1(n_257_551), .A2(n_257_426), .ZN(n_257_76_10346));
   NAND3_X1 i_257_76_10365 (.A1(n_257_76_10316), .A2(n_257_76_10284), .A3(
      n_257_76_10346), .ZN(n_257_76_10347));
   NAND2_X1 i_257_76_10366 (.A1(n_257_131), .A2(n_257_430), .ZN(n_257_76_10348));
   NAND2_X1 i_257_76_10367 (.A1(n_257_451), .A2(n_257_470), .ZN(n_257_76_10349));
   NAND4_X1 i_257_76_10368 (.A1(n_257_76_10317), .A2(n_257_76_10348), .A3(
      n_257_76_10318), .A4(n_257_76_10349), .ZN(n_257_76_10350));
   NOR2_X1 i_257_76_10369 (.A1(n_257_76_10347), .A2(n_257_76_10350), .ZN(
      n_257_76_10351));
   NAND2_X1 i_257_76_10370 (.A1(n_257_93), .A2(n_257_431), .ZN(n_257_76_10352));
   INV_X1 i_257_76_10371 (.A(n_257_1077), .ZN(n_257_76_10353));
   NAND2_X1 i_257_76_10372 (.A1(n_257_432), .A2(n_257_615), .ZN(n_257_76_10354));
   NAND4_X1 i_257_76_10373 (.A1(n_257_76_10353), .A2(n_257_76_18023), .A3(
      n_257_76_10354), .A4(n_257_423), .ZN(n_257_76_10355));
   INV_X1 i_257_76_10374 (.A(n_257_76_10300), .ZN(n_257_76_10356));
   NOR2_X1 i_257_76_10375 (.A1(n_257_76_10355), .A2(n_257_76_10356), .ZN(
      n_257_76_10357));
   NAND2_X1 i_257_76_10376 (.A1(n_257_519), .A2(n_257_424), .ZN(n_257_76_10358));
   NAND2_X1 i_257_76_10377 (.A1(n_257_53), .A2(n_257_433), .ZN(n_257_76_10359));
   NAND4_X1 i_257_76_10378 (.A1(n_257_76_10357), .A2(n_257_76_10358), .A3(
      n_257_76_10359), .A4(n_257_290), .ZN(n_257_76_10360));
   INV_X1 i_257_76_10379 (.A(n_257_76_10360), .ZN(n_257_76_10361));
   NAND2_X1 i_257_76_10380 (.A1(n_257_76_10352), .A2(n_257_76_10361), .ZN(
      n_257_76_10362));
   INV_X1 i_257_76_10381 (.A(n_257_76_10362), .ZN(n_257_76_10363));
   NAND2_X1 i_257_76_10382 (.A1(n_257_170), .A2(n_257_429), .ZN(n_257_76_10364));
   NAND2_X1 i_257_76_10383 (.A1(n_257_76_10312), .A2(n_257_76_10303), .ZN(
      n_257_76_10365));
   INV_X1 i_257_76_10384 (.A(n_257_76_10365), .ZN(n_257_76_10366));
   NAND2_X1 i_257_76_10385 (.A1(n_257_647), .A2(n_257_450), .ZN(n_257_76_10367));
   NAND2_X1 i_257_76_10386 (.A1(n_257_427), .A2(n_257_210), .ZN(n_257_76_10368));
   NAND2_X1 i_257_76_10387 (.A1(n_257_76_10304), .A2(n_257_76_10368), .ZN(
      n_257_76_10369));
   INV_X1 i_257_76_10388 (.A(n_257_76_10369), .ZN(n_257_76_10370));
   NAND3_X1 i_257_76_10389 (.A1(n_257_76_10366), .A2(n_257_76_10367), .A3(
      n_257_76_10370), .ZN(n_257_76_10371));
   NAND3_X1 i_257_76_10390 (.A1(n_257_76_10307), .A2(n_257_76_10308), .A3(
      n_257_76_10311), .ZN(n_257_76_10372));
   NOR2_X1 i_257_76_10391 (.A1(n_257_76_10371), .A2(n_257_76_10372), .ZN(
      n_257_76_10373));
   NAND4_X1 i_257_76_10392 (.A1(n_257_76_10351), .A2(n_257_76_10363), .A3(
      n_257_76_10364), .A4(n_257_76_10373), .ZN(n_257_76_10374));
   INV_X1 i_257_76_10393 (.A(n_257_76_10374), .ZN(n_257_76_10375));
   NAND2_X1 i_257_76_10394 (.A1(n_257_250), .A2(n_257_425), .ZN(n_257_76_10376));
   NAND2_X1 i_257_76_10395 (.A1(n_257_76_10376), .A2(n_257_76_10321), .ZN(
      n_257_76_10377));
   INV_X1 i_257_76_10396 (.A(n_257_76_10377), .ZN(n_257_76_10378));
   NAND4_X1 i_257_76_10397 (.A1(n_257_76_10375), .A2(n_257_76_10378), .A3(
      n_257_76_10281), .A4(n_257_76_10283), .ZN(n_257_76_10379));
   INV_X1 i_257_76_10398 (.A(n_257_76_10379), .ZN(n_257_76_10380));
   NAND2_X1 i_257_76_10399 (.A1(n_257_76_18066), .A2(n_257_76_10380), .ZN(
      n_257_76_10381));
   NAND3_X1 i_257_76_10400 (.A1(n_257_76_10336), .A2(n_257_76_10345), .A3(
      n_257_76_10381), .ZN(n_257_76_10382));
   NOR2_X1 i_257_76_10401 (.A1(n_257_76_10325), .A2(n_257_76_10382), .ZN(
      n_257_76_10383));
   NAND2_X1 i_257_76_10402 (.A1(n_257_981), .A2(n_257_76_10294), .ZN(
      n_257_76_10384));
   INV_X1 i_257_76_10403 (.A(n_257_76_10384), .ZN(n_257_76_10385));
   NAND2_X1 i_257_76_10404 (.A1(n_257_441), .A2(n_257_76_10385), .ZN(
      n_257_76_10386));
   INV_X1 i_257_76_10405 (.A(n_257_76_10386), .ZN(n_257_76_10387));
   NAND2_X1 i_257_76_10406 (.A1(n_257_76_10283), .A2(n_257_76_10387), .ZN(
      n_257_76_10388));
   NOR2_X1 i_257_76_10407 (.A1(n_257_76_10282), .A2(n_257_76_10388), .ZN(
      n_257_76_10389));
   NAND2_X1 i_257_76_10408 (.A1(n_257_76_18071), .A2(n_257_76_10389), .ZN(
      n_257_76_10390));
   NOR2_X1 i_257_76_10409 (.A1(n_257_76_10295), .A2(n_257_76_10300), .ZN(
      n_257_76_10391));
   NAND4_X1 i_257_76_10410 (.A1(n_257_76_10391), .A2(n_257_76_10312), .A3(
      n_257_76_10303), .A4(n_257_76_10304), .ZN(n_257_76_10392));
   INV_X1 i_257_76_10411 (.A(n_257_76_10392), .ZN(n_257_76_10393));
   NAND2_X1 i_257_76_10412 (.A1(n_257_76_10307), .A2(n_257_76_10311), .ZN(
      n_257_76_10394));
   INV_X1 i_257_76_10413 (.A(n_257_76_10394), .ZN(n_257_76_10395));
   NAND3_X1 i_257_76_10414 (.A1(n_257_76_10393), .A2(n_257_76_10395), .A3(
      n_257_76_10318), .ZN(n_257_76_10396));
   NAND3_X1 i_257_76_10415 (.A1(n_257_76_10316), .A2(n_257_76_10284), .A3(
      n_257_76_10317), .ZN(n_257_76_10397));
   NOR2_X1 i_257_76_10416 (.A1(n_257_76_10396), .A2(n_257_76_10397), .ZN(
      n_257_76_10398));
   NAND2_X1 i_257_76_10417 (.A1(n_257_76_10283), .A2(n_257_76_10398), .ZN(
      n_257_76_10399));
   NOR2_X1 i_257_76_10418 (.A1(n_257_76_10282), .A2(n_257_76_10399), .ZN(
      n_257_76_10400));
   NAND2_X1 i_257_76_10419 (.A1(n_257_76_18078), .A2(n_257_76_10400), .ZN(
      n_257_76_10401));
   NAND3_X1 i_257_76_10420 (.A1(n_257_428), .A2(n_257_583), .A3(n_257_442), 
      .ZN(n_257_76_10402));
   INV_X1 i_257_76_10421 (.A(n_257_76_10402), .ZN(n_257_76_10403));
   NAND3_X1 i_257_76_10422 (.A1(n_257_76_10353), .A2(n_257_76_10354), .A3(
      n_257_76_10403), .ZN(n_257_76_10404));
   NOR2_X1 i_257_76_10423 (.A1(n_257_76_10404), .A2(n_257_76_10356), .ZN(
      n_257_76_10405));
   NAND4_X1 i_257_76_10424 (.A1(n_257_76_10405), .A2(n_257_76_10303), .A3(
      n_257_76_10304), .A4(n_257_76_10359), .ZN(n_257_76_10406));
   NAND2_X1 i_257_76_10425 (.A1(n_257_76_10367), .A2(n_257_76_10312), .ZN(
      n_257_76_10407));
   NOR2_X1 i_257_76_10426 (.A1(n_257_76_10406), .A2(n_257_76_10407), .ZN(
      n_257_76_10408));
   NAND3_X1 i_257_76_10427 (.A1(n_257_76_10348), .A2(n_257_76_10318), .A3(
      n_257_76_10349), .ZN(n_257_76_10409));
   INV_X1 i_257_76_10428 (.A(n_257_76_10409), .ZN(n_257_76_10410));
   INV_X1 i_257_76_10429 (.A(n_257_76_10372), .ZN(n_257_76_10411));
   NAND3_X1 i_257_76_10430 (.A1(n_257_76_10408), .A2(n_257_76_10410), .A3(
      n_257_76_10411), .ZN(n_257_76_10412));
   NAND2_X1 i_257_76_10431 (.A1(n_257_76_10284), .A2(n_257_76_10317), .ZN(
      n_257_76_10413));
   INV_X1 i_257_76_10432 (.A(n_257_76_10413), .ZN(n_257_76_10414));
   NAND3_X1 i_257_76_10433 (.A1(n_257_76_10414), .A2(n_257_76_10352), .A3(
      n_257_76_10316), .ZN(n_257_76_10415));
   NOR2_X1 i_257_76_10434 (.A1(n_257_76_10412), .A2(n_257_76_10415), .ZN(
      n_257_76_10416));
   NAND2_X1 i_257_76_10435 (.A1(n_257_76_10321), .A2(n_257_76_10364), .ZN(
      n_257_76_10417));
   INV_X1 i_257_76_10436 (.A(n_257_76_10417), .ZN(n_257_76_10418));
   NAND4_X1 i_257_76_10437 (.A1(n_257_76_10416), .A2(n_257_76_10281), .A3(
      n_257_76_10283), .A4(n_257_76_10418), .ZN(n_257_76_10419));
   INV_X1 i_257_76_10438 (.A(n_257_76_10419), .ZN(n_257_76_10420));
   NAND2_X1 i_257_76_10439 (.A1(n_257_76_18074), .A2(n_257_76_10420), .ZN(
      n_257_76_10421));
   NAND3_X1 i_257_76_10440 (.A1(n_257_76_10390), .A2(n_257_76_10401), .A3(
      n_257_76_10421), .ZN(n_257_76_10422));
   NAND2_X1 i_257_76_10441 (.A1(n_257_1077), .A2(n_257_442), .ZN(n_257_76_10423));
   INV_X1 i_257_76_10442 (.A(n_257_76_10423), .ZN(n_257_76_10424));
   NAND2_X1 i_257_76_10443 (.A1(n_257_13), .A2(n_257_76_10424), .ZN(
      n_257_76_10425));
   NAND2_X1 i_257_76_10444 (.A1(n_257_76_10303), .A2(n_257_76_10304), .ZN(
      n_257_76_10426));
   NAND3_X1 i_257_76_10445 (.A1(n_257_879), .A2(n_257_76_10294), .A3(n_257_445), 
      .ZN(n_257_76_10427));
   NOR2_X1 i_257_76_10446 (.A1(n_257_76_10426), .A2(n_257_76_10427), .ZN(
      n_257_76_10428));
   NAND3_X1 i_257_76_10447 (.A1(n_257_76_10428), .A2(n_257_76_10284), .A3(
      n_257_76_10318), .ZN(n_257_76_10429));
   INV_X1 i_257_76_10448 (.A(n_257_76_10429), .ZN(n_257_76_10430));
   NAND2_X1 i_257_76_10449 (.A1(n_257_76_10283), .A2(n_257_76_10430), .ZN(
      n_257_76_10431));
   NOR2_X1 i_257_76_10450 (.A1(n_257_76_10282), .A2(n_257_76_10431), .ZN(
      n_257_76_10432));
   NAND2_X1 i_257_76_10451 (.A1(n_257_76_18077), .A2(n_257_76_10432), .ZN(
      n_257_76_10433));
   NAND2_X1 i_257_76_10452 (.A1(n_257_76_10425), .A2(n_257_76_10433), .ZN(
      n_257_76_10434));
   NOR2_X1 i_257_76_10453 (.A1(n_257_76_10422), .A2(n_257_76_10434), .ZN(
      n_257_76_10435));
   INV_X1 i_257_76_10454 (.A(n_257_76_10321), .ZN(n_257_76_10436));
   NAND2_X1 i_257_76_10455 (.A1(n_257_76_10300), .A2(n_257_76_10353), .ZN(
      n_257_76_10437));
   INV_X1 i_257_76_10456 (.A(n_257_76_10437), .ZN(n_257_76_10438));
   NAND3_X1 i_257_76_10457 (.A1(n_257_76_10354), .A2(n_257_76_18023), .A3(
      n_257_426), .ZN(n_257_76_10439));
   INV_X1 i_257_76_10458 (.A(n_257_76_10439), .ZN(n_257_76_10440));
   NAND4_X1 i_257_76_10459 (.A1(n_257_76_10438), .A2(n_257_76_10359), .A3(
      n_257_76_10368), .A4(n_257_76_10440), .ZN(n_257_76_10441));
   NAND3_X1 i_257_76_10460 (.A1(n_257_76_10312), .A2(n_257_76_10303), .A3(
      n_257_76_10304), .ZN(n_257_76_10442));
   NOR2_X1 i_257_76_10461 (.A1(n_257_76_10441), .A2(n_257_76_10442), .ZN(
      n_257_76_10443));
   NAND2_X1 i_257_76_10462 (.A1(n_257_76_10317), .A2(n_257_76_10348), .ZN(
      n_257_76_10444));
   INV_X1 i_257_76_10463 (.A(n_257_76_10444), .ZN(n_257_76_10445));
   NAND3_X1 i_257_76_10464 (.A1(n_257_76_10318), .A2(n_257_551), .A3(
      n_257_76_10367), .ZN(n_257_76_10446));
   INV_X1 i_257_76_10465 (.A(n_257_76_10446), .ZN(n_257_76_10447));
   NAND3_X1 i_257_76_10466 (.A1(n_257_76_10443), .A2(n_257_76_10445), .A3(
      n_257_76_10447), .ZN(n_257_76_10448));
   NOR2_X1 i_257_76_10467 (.A1(n_257_76_10436), .A2(n_257_76_10448), .ZN(
      n_257_76_10449));
   NAND4_X1 i_257_76_10468 (.A1(n_257_76_10349), .A2(n_257_76_10307), .A3(
      n_257_76_10308), .A4(n_257_76_10311), .ZN(n_257_76_10450));
   INV_X1 i_257_76_10469 (.A(n_257_76_10450), .ZN(n_257_76_10451));
   NAND2_X1 i_257_76_10470 (.A1(n_257_76_10316), .A2(n_257_76_10284), .ZN(
      n_257_76_10452));
   INV_X1 i_257_76_10471 (.A(n_257_76_10452), .ZN(n_257_76_10453));
   NAND4_X1 i_257_76_10472 (.A1(n_257_76_10364), .A2(n_257_76_10451), .A3(
      n_257_76_10453), .A4(n_257_76_10352), .ZN(n_257_76_10454));
   INV_X1 i_257_76_10473 (.A(n_257_76_10454), .ZN(n_257_76_10455));
   NAND4_X1 i_257_76_10474 (.A1(n_257_76_10449), .A2(n_257_76_10281), .A3(
      n_257_76_10283), .A4(n_257_76_10455), .ZN(n_257_76_10456));
   INV_X1 i_257_76_10475 (.A(n_257_76_10456), .ZN(n_257_76_10457));
   NAND2_X1 i_257_76_10476 (.A1(n_257_76_18076), .A2(n_257_76_10457), .ZN(
      n_257_76_10458));
   NAND4_X1 i_257_76_10477 (.A1(n_257_76_10284), .A2(n_257_76_10317), .A3(
      n_257_76_10318), .A4(n_257_751), .ZN(n_257_76_10459));
   INV_X1 i_257_76_10478 (.A(n_257_76_10304), .ZN(n_257_76_10460));
   NAND2_X1 i_257_76_10479 (.A1(n_257_76_10294), .A2(n_257_436), .ZN(
      n_257_76_10461));
   NOR2_X1 i_257_76_10480 (.A1(n_257_76_10460), .A2(n_257_76_10461), .ZN(
      n_257_76_10462));
   NAND4_X1 i_257_76_10481 (.A1(n_257_76_10462), .A2(n_257_76_10366), .A3(
      n_257_76_10307), .A4(n_257_76_10311), .ZN(n_257_76_10463));
   NOR2_X1 i_257_76_10482 (.A1(n_257_76_10459), .A2(n_257_76_10463), .ZN(
      n_257_76_10464));
   NAND2_X1 i_257_76_10483 (.A1(n_257_76_10283), .A2(n_257_76_10464), .ZN(
      n_257_76_10465));
   NOR2_X1 i_257_76_10484 (.A1(n_257_76_10282), .A2(n_257_76_10465), .ZN(
      n_257_76_10466));
   NAND2_X1 i_257_76_10485 (.A1(n_257_76_18069), .A2(n_257_76_10466), .ZN(
      n_257_76_10467));
   NAND2_X1 i_257_76_10486 (.A1(n_257_615), .A2(n_257_442), .ZN(n_257_76_10468));
   INV_X1 i_257_76_10487 (.A(n_257_76_10468), .ZN(n_257_76_10469));
   NAND2_X1 i_257_76_10488 (.A1(n_257_432), .A2(n_257_76_10469), .ZN(
      n_257_76_10470));
   NOR2_X1 i_257_76_10489 (.A1(n_257_76_10470), .A2(n_257_1077), .ZN(
      n_257_76_10471));
   NAND3_X1 i_257_76_10490 (.A1(n_257_76_10359), .A2(n_257_76_10300), .A3(
      n_257_76_10471), .ZN(n_257_76_10472));
   NOR2_X1 i_257_76_10491 (.A1(n_257_76_10442), .A2(n_257_76_10472), .ZN(
      n_257_76_10473));
   NAND3_X1 i_257_76_10492 (.A1(n_257_76_10308), .A2(n_257_76_10311), .A3(
      n_257_76_10367), .ZN(n_257_76_10474));
   INV_X1 i_257_76_10493 (.A(n_257_76_10474), .ZN(n_257_76_10475));
   NAND2_X1 i_257_76_10494 (.A1(n_257_76_10349), .A2(n_257_76_10307), .ZN(
      n_257_76_10476));
   INV_X1 i_257_76_10495 (.A(n_257_76_10476), .ZN(n_257_76_10477));
   NAND3_X1 i_257_76_10496 (.A1(n_257_76_10473), .A2(n_257_76_10475), .A3(
      n_257_76_10477), .ZN(n_257_76_10478));
   NOR2_X1 i_257_76_10497 (.A1(n_257_76_10478), .A2(n_257_76_10319), .ZN(
      n_257_76_10479));
   NAND3_X1 i_257_76_10498 (.A1(n_257_76_10479), .A2(n_257_76_10283), .A3(
      n_257_76_10321), .ZN(n_257_76_10480));
   NOR2_X1 i_257_76_10499 (.A1(n_257_76_10480), .A2(n_257_76_10282), .ZN(
      n_257_76_10481));
   NAND2_X1 i_257_76_10500 (.A1(n_257_68), .A2(n_257_76_10481), .ZN(
      n_257_76_10482));
   NAND3_X1 i_257_76_10501 (.A1(n_257_76_10458), .A2(n_257_76_10467), .A3(
      n_257_76_10482), .ZN(n_257_76_10483));
   NAND2_X1 i_257_76_10502 (.A1(n_257_76_10307), .A2(n_257_815), .ZN(
      n_257_76_10484));
   INV_X1 i_257_76_10503 (.A(n_257_76_10484), .ZN(n_257_76_10485));
   NOR2_X1 i_257_76_10504 (.A1(n_257_76_10295), .A2(n_257_76_15924), .ZN(
      n_257_76_10486));
   NAND4_X1 i_257_76_10505 (.A1(n_257_76_10486), .A2(n_257_76_10312), .A3(
      n_257_76_10303), .A4(n_257_76_10304), .ZN(n_257_76_10487));
   INV_X1 i_257_76_10506 (.A(n_257_76_10487), .ZN(n_257_76_10488));
   NAND4_X1 i_257_76_10507 (.A1(n_257_76_10485), .A2(n_257_76_10488), .A3(
      n_257_76_10284), .A4(n_257_76_10318), .ZN(n_257_76_10489));
   INV_X1 i_257_76_10508 (.A(n_257_76_10489), .ZN(n_257_76_10490));
   NAND2_X1 i_257_76_10509 (.A1(n_257_76_10283), .A2(n_257_76_10490), .ZN(
      n_257_76_10491));
   NOR2_X1 i_257_76_10510 (.A1(n_257_76_10282), .A2(n_257_76_10491), .ZN(
      n_257_76_10492));
   NAND2_X1 i_257_76_10511 (.A1(n_257_22), .A2(n_257_76_10492), .ZN(
      n_257_76_10493));
   NAND2_X1 i_257_76_10512 (.A1(n_257_444), .A2(n_257_76_10294), .ZN(
      n_257_76_10494));
   INV_X1 i_257_76_10513 (.A(n_257_76_10494), .ZN(n_257_76_10495));
   NAND2_X1 i_257_76_10514 (.A1(n_257_1013), .A2(n_257_76_10495), .ZN(
      n_257_76_10496));
   INV_X1 i_257_76_10515 (.A(n_257_76_10496), .ZN(n_257_76_10497));
   NAND2_X1 i_257_76_10516 (.A1(n_257_76_10281), .A2(n_257_76_10497), .ZN(
      n_257_76_10498));
   INV_X1 i_257_76_10517 (.A(n_257_76_10498), .ZN(n_257_76_10499));
   NAND2_X1 i_257_76_10518 (.A1(n_257_76_18075), .A2(n_257_76_10499), .ZN(
      n_257_76_10500));
   NAND2_X1 i_257_76_10519 (.A1(n_257_76_10493), .A2(n_257_76_10500), .ZN(
      n_257_76_10501));
   NOR2_X1 i_257_76_10520 (.A1(n_257_76_10483), .A2(n_257_76_10501), .ZN(
      n_257_76_10502));
   NAND3_X1 i_257_76_10521 (.A1(n_257_76_10383), .A2(n_257_76_10435), .A3(
      n_257_76_10502), .ZN(n_257_76_10503));
   INV_X1 i_257_76_10522 (.A(n_257_76_10503), .ZN(n_257_76_10504));
   NOR2_X1 i_257_76_10523 (.A1(n_257_1077), .A2(n_257_76_17633), .ZN(
      n_257_76_10505));
   NAND3_X1 i_257_76_10524 (.A1(n_257_76_10505), .A2(n_257_53), .A3(
      n_257_76_10300), .ZN(n_257_76_10506));
   INV_X1 i_257_76_10525 (.A(n_257_76_10506), .ZN(n_257_76_10507));
   NAND4_X1 i_257_76_10526 (.A1(n_257_76_10507), .A2(n_257_76_10312), .A3(
      n_257_76_10303), .A4(n_257_76_10304), .ZN(n_257_76_10508));
   INV_X1 i_257_76_10527 (.A(n_257_76_10508), .ZN(n_257_76_10509));
   NAND3_X1 i_257_76_10528 (.A1(n_257_76_10475), .A2(n_257_76_10477), .A3(
      n_257_76_10509), .ZN(n_257_76_10510));
   NOR2_X1 i_257_76_10529 (.A1(n_257_76_10510), .A2(n_257_76_10319), .ZN(
      n_257_76_10511));
   NAND3_X1 i_257_76_10530 (.A1(n_257_76_10511), .A2(n_257_76_10283), .A3(
      n_257_76_10321), .ZN(n_257_76_10512));
   NOR2_X1 i_257_76_10531 (.A1(n_257_76_10512), .A2(n_257_76_10282), .ZN(
      n_257_76_10513));
   NAND2_X1 i_257_76_10532 (.A1(n_257_76_18081), .A2(n_257_76_10513), .ZN(
      n_257_76_10514));
   NOR2_X1 i_257_76_10533 (.A1(n_257_1077), .A2(n_257_76_14899), .ZN(
      n_257_76_10515));
   NAND2_X1 i_257_76_10534 (.A1(n_257_76_10300), .A2(n_257_76_10515), .ZN(
      n_257_76_10516));
   INV_X1 i_257_76_10535 (.A(n_257_76_10516), .ZN(n_257_76_10517));
   NAND4_X1 i_257_76_10536 (.A1(n_257_76_10517), .A2(n_257_449), .A3(
      n_257_76_10303), .A4(n_257_76_10304), .ZN(n_257_76_10518));
   NOR2_X1 i_257_76_10537 (.A1(n_257_76_10518), .A2(n_257_76_10313), .ZN(
      n_257_76_10519));
   NAND3_X1 i_257_76_10538 (.A1(n_257_76_10317), .A2(n_257_76_10318), .A3(
      n_257_76_10307), .ZN(n_257_76_10520));
   INV_X1 i_257_76_10539 (.A(n_257_76_10520), .ZN(n_257_76_10521));
   NAND3_X1 i_257_76_10540 (.A1(n_257_76_10519), .A2(n_257_76_10453), .A3(
      n_257_76_10521), .ZN(n_257_76_10522));
   NOR2_X1 i_257_76_10541 (.A1(n_257_76_10522), .A2(n_257_76_10436), .ZN(
      n_257_76_10523));
   NAND3_X1 i_257_76_10542 (.A1(n_257_76_10523), .A2(n_257_76_10281), .A3(
      n_257_76_10283), .ZN(n_257_76_10524));
   INV_X1 i_257_76_10543 (.A(n_257_76_10524), .ZN(n_257_76_10525));
   NAND2_X1 i_257_76_10544 (.A1(n_257_76_18083), .A2(n_257_76_10525), .ZN(
      n_257_76_10526));
   NAND3_X1 i_257_76_10545 (.A1(n_257_76_10318), .A2(n_257_76_10349), .A3(
      n_257_76_10307), .ZN(n_257_76_10527));
   INV_X1 i_257_76_10546 (.A(n_257_76_10527), .ZN(n_257_76_10528));
   NAND3_X1 i_257_76_10547 (.A1(n_257_76_10353), .A2(n_257_76_10354), .A3(
      n_257_76_17331), .ZN(n_257_76_10529));
   INV_X1 i_257_76_10548 (.A(n_257_76_10529), .ZN(n_257_76_10530));
   NAND3_X1 i_257_76_10549 (.A1(n_257_76_10359), .A2(n_257_76_10300), .A3(
      n_257_76_10530), .ZN(n_257_76_10531));
   NOR2_X1 i_257_76_10550 (.A1(n_257_76_10442), .A2(n_257_76_10531), .ZN(
      n_257_76_10532));
   NAND3_X1 i_257_76_10551 (.A1(n_257_76_10528), .A2(n_257_76_10475), .A3(
      n_257_76_10532), .ZN(n_257_76_10533));
   NAND4_X1 i_257_76_10552 (.A1(n_257_76_10316), .A2(n_257_76_10284), .A3(
      n_257_76_10317), .A4(n_257_76_10348), .ZN(n_257_76_10534));
   NOR2_X1 i_257_76_10553 (.A1(n_257_76_10533), .A2(n_257_76_10534), .ZN(
      n_257_76_10535));
   NAND2_X1 i_257_76_10554 (.A1(n_257_76_10352), .A2(n_257_170), .ZN(
      n_257_76_10536));
   INV_X1 i_257_76_10555 (.A(n_257_76_10536), .ZN(n_257_76_10537));
   NAND2_X1 i_257_76_10556 (.A1(n_257_76_10321), .A2(n_257_76_10537), .ZN(
      n_257_76_10538));
   INV_X1 i_257_76_10557 (.A(n_257_76_10538), .ZN(n_257_76_10539));
   NAND4_X1 i_257_76_10558 (.A1(n_257_76_10281), .A2(n_257_76_10535), .A3(
      n_257_76_10539), .A4(n_257_76_10283), .ZN(n_257_76_10540));
   INV_X1 i_257_76_10559 (.A(n_257_76_10540), .ZN(n_257_76_10541));
   NAND2_X1 i_257_76_10560 (.A1(n_257_76_18061), .A2(n_257_76_10541), .ZN(
      n_257_76_10542));
   NAND3_X1 i_257_76_10561 (.A1(n_257_76_10514), .A2(n_257_76_10526), .A3(
      n_257_76_10542), .ZN(n_257_76_10543));
   INV_X1 i_257_76_10562 (.A(n_257_76_10543), .ZN(n_257_76_10544));
   NAND3_X1 i_257_76_10563 (.A1(n_257_76_10294), .A2(n_257_438), .A3(n_257_1083), 
      .ZN(n_257_76_10545));
   INV_X1 i_257_76_10564 (.A(n_257_76_10303), .ZN(n_257_76_10546));
   NOR2_X1 i_257_76_10565 (.A1(n_257_76_10545), .A2(n_257_76_10546), .ZN(
      n_257_76_10547));
   NAND3_X1 i_257_76_10566 (.A1(n_257_76_10284), .A2(n_257_76_10547), .A3(
      n_257_76_10318), .ZN(n_257_76_10548));
   INV_X1 i_257_76_10567 (.A(n_257_76_10548), .ZN(n_257_76_10549));
   NAND2_X1 i_257_76_10568 (.A1(n_257_76_10283), .A2(n_257_76_10549), .ZN(
      n_257_76_10550));
   NOR2_X1 i_257_76_10569 (.A1(n_257_76_10282), .A2(n_257_76_10550), .ZN(
      n_257_76_10551));
   NAND2_X1 i_257_76_10570 (.A1(n_257_76_18067), .A2(n_257_76_10551), .ZN(
      n_257_76_10552));
   NAND2_X1 i_257_76_10571 (.A1(n_257_367), .A2(n_257_421), .ZN(n_257_76_10553));
   NAND2_X1 i_257_76_10572 (.A1(n_257_76_10553), .A2(n_257_76_10352), .ZN(
      n_257_76_10554));
   INV_X1 i_257_76_10573 (.A(n_257_76_10554), .ZN(n_257_76_10555));
   NAND2_X1 i_257_76_10574 (.A1(n_257_76_10555), .A2(n_257_76_10364), .ZN(
      n_257_76_10556));
   NOR2_X1 i_257_76_10575 (.A1(n_257_76_10556), .A2(n_257_76_10436), .ZN(
      n_257_76_10557));
   NAND2_X1 i_257_76_10576 (.A1(n_257_76_10346), .A2(n_257_76_10317), .ZN(
      n_257_76_10558));
   NOR2_X1 i_257_76_10577 (.A1(n_257_76_10452), .A2(n_257_76_10558), .ZN(
      n_257_76_10559));
   NAND2_X1 i_257_76_10578 (.A1(n_257_76_10348), .A2(n_257_76_10318), .ZN(
      n_257_76_10560));
   NOR2_X1 i_257_76_10579 (.A1(n_257_76_10560), .A2(n_257_76_10476), .ZN(
      n_257_76_10561));
   NAND2_X1 i_257_76_10580 (.A1(n_257_76_10559), .A2(n_257_76_10561), .ZN(
      n_257_76_10562));
   NAND2_X1 i_257_76_10581 (.A1(n_257_290), .A2(n_257_423), .ZN(n_257_76_10563));
   NAND2_X1 i_257_76_10582 (.A1(n_257_76_10563), .A2(n_257_76_10358), .ZN(
      n_257_76_10564));
   NOR2_X1 i_257_76_10583 (.A1(n_257_76_10564), .A2(n_257_76_10365), .ZN(
      n_257_76_10565));
   NAND2_X1 i_257_76_10584 (.A1(n_257_76_10368), .A2(n_257_76_10300), .ZN(
      n_257_76_10566));
   INV_X1 i_257_76_10585 (.A(n_257_76_10566), .ZN(n_257_76_10567));
   NAND2_X1 i_257_76_10586 (.A1(n_257_442), .A2(n_257_487), .ZN(n_257_76_10568));
   NAND2_X1 i_257_76_10587 (.A1(n_257_76_10353), .A2(n_257_76_18024), .ZN(
      n_257_76_10569));
   NAND2_X1 i_257_76_10588 (.A1(n_257_76_10354), .A2(n_257_420), .ZN(
      n_257_76_10570));
   NOR2_X1 i_257_76_10589 (.A1(n_257_76_10569), .A2(n_257_76_10570), .ZN(
      n_257_76_10571));
   NAND2_X1 i_257_76_10590 (.A1(n_257_76_10567), .A2(n_257_76_10571), .ZN(
      n_257_76_10572));
   NAND2_X1 i_257_76_10591 (.A1(n_257_76_10304), .A2(n_257_76_10359), .ZN(
      n_257_76_10573));
   NOR2_X1 i_257_76_10592 (.A1(n_257_76_10572), .A2(n_257_76_10573), .ZN(
      n_257_76_10574));
   NAND2_X1 i_257_76_10593 (.A1(n_257_76_10565), .A2(n_257_76_10574), .ZN(
      n_257_76_10575));
   INV_X1 i_257_76_10594 (.A(n_257_76_10575), .ZN(n_257_76_10576));
   NAND2_X1 i_257_76_10595 (.A1(n_257_76_10308), .A2(n_257_76_10311), .ZN(
      n_257_76_10577));
   NAND2_X1 i_257_76_10596 (.A1(n_257_328), .A2(n_257_422), .ZN(n_257_76_10578));
   NAND2_X1 i_257_76_10597 (.A1(n_257_76_10367), .A2(n_257_76_10578), .ZN(
      n_257_76_10579));
   NOR2_X1 i_257_76_10598 (.A1(n_257_76_10577), .A2(n_257_76_10579), .ZN(
      n_257_76_10580));
   NAND2_X1 i_257_76_10599 (.A1(n_257_76_10576), .A2(n_257_76_10580), .ZN(
      n_257_76_10581));
   NOR2_X1 i_257_76_10600 (.A1(n_257_76_10562), .A2(n_257_76_10581), .ZN(
      n_257_76_10582));
   NAND2_X1 i_257_76_10601 (.A1(n_257_76_10557), .A2(n_257_76_10582), .ZN(
      n_257_76_10583));
   NAND2_X1 i_257_76_10602 (.A1(n_257_76_10283), .A2(n_257_76_10376), .ZN(
      n_257_76_10584));
   INV_X1 i_257_76_10603 (.A(n_257_76_10584), .ZN(n_257_76_10585));
   NAND2_X1 i_257_76_10604 (.A1(n_257_76_10585), .A2(n_257_76_10281), .ZN(
      n_257_76_10586));
   NOR2_X1 i_257_76_10605 (.A1(n_257_76_10583), .A2(n_257_76_10586), .ZN(
      n_257_76_10587));
   NAND2_X1 i_257_76_10606 (.A1(n_257_76_18073), .A2(n_257_76_10587), .ZN(
      n_257_76_10588));
   NAND3_X1 i_257_76_10607 (.A1(n_257_131), .A2(n_257_76_10312), .A3(
      n_257_76_10303), .ZN(n_257_76_10589));
   NAND3_X1 i_257_76_10608 (.A1(n_257_76_10353), .A2(n_257_76_10354), .A3(
      n_257_76_17925), .ZN(n_257_76_10590));
   INV_X1 i_257_76_10609 (.A(n_257_76_10590), .ZN(n_257_76_10591));
   NAND4_X1 i_257_76_10610 (.A1(n_257_76_10304), .A2(n_257_76_10359), .A3(
      n_257_76_10300), .A4(n_257_76_10591), .ZN(n_257_76_10592));
   NOR2_X1 i_257_76_10611 (.A1(n_257_76_10589), .A2(n_257_76_10592), .ZN(
      n_257_76_10593));
   NAND3_X1 i_257_76_10612 (.A1(n_257_76_10593), .A2(n_257_76_10528), .A3(
      n_257_76_10475), .ZN(n_257_76_10594));
   INV_X1 i_257_76_10613 (.A(n_257_76_10594), .ZN(n_257_76_10595));
   INV_X1 i_257_76_10614 (.A(n_257_76_10352), .ZN(n_257_76_10596));
   NOR2_X1 i_257_76_10615 (.A1(n_257_76_10397), .A2(n_257_76_10596), .ZN(
      n_257_76_10597));
   NAND3_X1 i_257_76_10616 (.A1(n_257_76_10321), .A2(n_257_76_10595), .A3(
      n_257_76_10597), .ZN(n_257_76_10598));
   INV_X1 i_257_76_10617 (.A(n_257_76_10598), .ZN(n_257_76_10599));
   NAND3_X1 i_257_76_10618 (.A1(n_257_76_10599), .A2(n_257_76_10281), .A3(
      n_257_76_10283), .ZN(n_257_76_10600));
   INV_X1 i_257_76_10619 (.A(n_257_76_10600), .ZN(n_257_76_10601));
   NAND2_X1 i_257_76_10620 (.A1(n_257_76_18068), .A2(n_257_76_10601), .ZN(
      n_257_76_10602));
   NAND3_X1 i_257_76_10621 (.A1(n_257_76_10552), .A2(n_257_76_10588), .A3(
      n_257_76_10602), .ZN(n_257_76_10603));
   INV_X1 i_257_76_10622 (.A(n_257_76_10603), .ZN(n_257_76_10604));
   NAND3_X1 i_257_76_10623 (.A1(n_257_76_10284), .A2(n_257_76_10317), .A3(
      n_257_76_10318), .ZN(n_257_76_10605));
   NAND2_X1 i_257_76_10624 (.A1(n_257_783), .A2(n_257_442), .ZN(n_257_76_10606));
   NOR2_X1 i_257_76_10625 (.A1(n_257_1077), .A2(n_257_76_10606), .ZN(
      n_257_76_10607));
   NAND3_X1 i_257_76_10626 (.A1(n_257_76_10303), .A2(n_257_76_10304), .A3(
      n_257_76_10607), .ZN(n_257_76_10608));
   INV_X1 i_257_76_10627 (.A(n_257_76_10608), .ZN(n_257_76_10609));
   NAND2_X1 i_257_76_10628 (.A1(n_257_76_10312), .A2(n_257_447), .ZN(
      n_257_76_10610));
   INV_X1 i_257_76_10629 (.A(n_257_76_10610), .ZN(n_257_76_10611));
   NAND3_X1 i_257_76_10630 (.A1(n_257_76_10609), .A2(n_257_76_10611), .A3(
      n_257_76_10307), .ZN(n_257_76_10612));
   NOR2_X1 i_257_76_10631 (.A1(n_257_76_10605), .A2(n_257_76_10612), .ZN(
      n_257_76_10613));
   NAND2_X1 i_257_76_10632 (.A1(n_257_76_10283), .A2(n_257_76_10613), .ZN(
      n_257_76_10614));
   NOR2_X1 i_257_76_10633 (.A1(n_257_76_10282), .A2(n_257_76_10614), .ZN(
      n_257_76_10615));
   NAND3_X1 i_257_76_10634 (.A1(n_257_76_10353), .A2(n_257_76_10354), .A3(
      n_257_76_17932), .ZN(n_257_76_10616));
   INV_X1 i_257_76_10635 (.A(n_257_76_10616), .ZN(n_257_76_10617));
   NAND3_X1 i_257_76_10636 (.A1(n_257_76_10359), .A2(n_257_76_10300), .A3(
      n_257_76_10617), .ZN(n_257_76_10618));
   NOR2_X1 i_257_76_10637 (.A1(n_257_76_10442), .A2(n_257_76_10618), .ZN(
      n_257_76_10619));
   NAND3_X1 i_257_76_10638 (.A1(n_257_76_10528), .A2(n_257_76_10475), .A3(
      n_257_76_10619), .ZN(n_257_76_10620));
   NAND4_X1 i_257_76_10639 (.A1(n_257_76_10316), .A2(n_257_93), .A3(
      n_257_76_10284), .A4(n_257_76_10317), .ZN(n_257_76_10621));
   NOR2_X1 i_257_76_10640 (.A1(n_257_76_10620), .A2(n_257_76_10621), .ZN(
      n_257_76_10622));
   NAND3_X1 i_257_76_10641 (.A1(n_257_76_10622), .A2(n_257_76_10283), .A3(
      n_257_76_10321), .ZN(n_257_76_10623));
   NOR2_X1 i_257_76_10642 (.A1(n_257_76_10623), .A2(n_257_76_10282), .ZN(
      n_257_76_10624));
   AOI22_X1 i_257_76_10643 (.A1(n_257_76_18085), .A2(n_257_76_10615), .B1(
      n_257_76_18080), .B2(n_257_76_10624), .ZN(n_257_76_10625));
   NAND3_X1 i_257_76_10644 (.A1(n_257_76_10544), .A2(n_257_76_10604), .A3(
      n_257_76_10625), .ZN(n_257_76_10626));
   NAND3_X1 i_257_76_10645 (.A1(n_257_76_10304), .A2(n_257_76_18025), .A3(
      n_257_76_10353), .ZN(n_257_76_10627));
   INV_X1 i_257_76_10646 (.A(n_257_76_10627), .ZN(n_257_76_10628));
   NAND4_X1 i_257_76_10647 (.A1(n_257_76_10317), .A2(n_257_76_10628), .A3(
      n_257_76_10366), .A4(n_257_76_10318), .ZN(n_257_76_10629));
   INV_X1 i_257_76_10648 (.A(n_257_76_10629), .ZN(n_257_76_10630));
   NAND3_X1 i_257_76_10649 (.A1(n_257_76_10307), .A2(n_257_76_10311), .A3(
      n_257_448), .ZN(n_257_76_10631));
   INV_X1 i_257_76_10650 (.A(n_257_76_10631), .ZN(n_257_76_10632));
   NAND4_X1 i_257_76_10651 (.A1(n_257_76_10630), .A2(n_257_687), .A3(
      n_257_76_10453), .A4(n_257_76_10632), .ZN(n_257_76_10633));
   INV_X1 i_257_76_10652 (.A(n_257_76_10633), .ZN(n_257_76_10634));
   NAND3_X1 i_257_76_10653 (.A1(n_257_76_10281), .A2(n_257_76_10283), .A3(
      n_257_76_10634), .ZN(n_257_76_10635));
   INV_X1 i_257_76_10654 (.A(n_257_76_10635), .ZN(n_257_76_10636));
   NAND2_X1 i_257_76_10655 (.A1(n_257_76_18079), .A2(n_257_76_10636), .ZN(
      n_257_76_10637));
   NAND2_X1 i_257_76_10656 (.A1(n_257_76_10352), .A2(n_257_76_10316), .ZN(
      n_257_76_10638));
   NAND4_X1 i_257_76_10657 (.A1(n_257_76_10284), .A2(n_257_76_10346), .A3(
      n_257_76_10317), .A4(n_257_76_10348), .ZN(n_257_76_10639));
   NOR2_X1 i_257_76_10658 (.A1(n_257_76_10638), .A2(n_257_76_10639), .ZN(
      n_257_76_10640));
   NAND2_X1 i_257_76_10659 (.A1(n_257_250), .A2(n_257_76_10364), .ZN(
      n_257_76_10641));
   INV_X1 i_257_76_10660 (.A(n_257_76_10641), .ZN(n_257_76_10642));
   NAND3_X1 i_257_76_10661 (.A1(n_257_76_10354), .A2(n_257_76_18023), .A3(
      n_257_425), .ZN(n_257_76_10643));
   INV_X1 i_257_76_10662 (.A(n_257_76_10643), .ZN(n_257_76_10644));
   NAND4_X1 i_257_76_10663 (.A1(n_257_76_10438), .A2(n_257_76_10359), .A3(
      n_257_76_10368), .A4(n_257_76_10644), .ZN(n_257_76_10645));
   NOR2_X1 i_257_76_10664 (.A1(n_257_76_10645), .A2(n_257_76_10442), .ZN(
      n_257_76_10646));
   NAND3_X1 i_257_76_10665 (.A1(n_257_76_10646), .A2(n_257_76_10528), .A3(
      n_257_76_10475), .ZN(n_257_76_10647));
   INV_X1 i_257_76_10666 (.A(n_257_76_10647), .ZN(n_257_76_10648));
   NAND4_X1 i_257_76_10667 (.A1(n_257_76_10640), .A2(n_257_76_10642), .A3(
      n_257_76_10321), .A4(n_257_76_10648), .ZN(n_257_76_10649));
   NAND2_X1 i_257_76_10668 (.A1(n_257_76_10281), .A2(n_257_76_10283), .ZN(
      n_257_76_10650));
   NOR2_X1 i_257_76_10669 (.A1(n_257_76_10649), .A2(n_257_76_10650), .ZN(
      n_257_76_10651));
   NAND2_X1 i_257_76_10670 (.A1(n_257_76_18064), .A2(n_257_76_10651), .ZN(
      n_257_76_10652));
   NAND3_X1 i_257_76_10671 (.A1(n_257_76_10284), .A2(n_257_76_10346), .A3(
      n_257_76_10317), .ZN(n_257_76_10653));
   NAND4_X1 i_257_76_10672 (.A1(n_257_76_10348), .A2(n_257_76_10318), .A3(
      n_257_76_10349), .A4(n_257_76_10307), .ZN(n_257_76_10654));
   NOR2_X1 i_257_76_10673 (.A1(n_257_76_10653), .A2(n_257_76_10654), .ZN(
      n_257_76_10655));
   NAND3_X1 i_257_76_10674 (.A1(n_257_76_10303), .A2(n_257_76_10304), .A3(
      n_257_76_10359), .ZN(n_257_76_10656));
   INV_X1 i_257_76_10675 (.A(n_257_76_18023), .ZN(n_257_76_10657));
   NOR2_X1 i_257_76_10676 (.A1(n_257_76_10657), .A2(n_257_1077), .ZN(
      n_257_76_10658));
   NAND2_X1 i_257_76_10677 (.A1(n_257_76_10354), .A2(n_257_421), .ZN(
      n_257_76_10659));
   INV_X1 i_257_76_10678 (.A(n_257_76_10659), .ZN(n_257_76_10660));
   NAND4_X1 i_257_76_10679 (.A1(n_257_76_10658), .A2(n_257_76_10368), .A3(
      n_257_76_10300), .A4(n_257_76_10660), .ZN(n_257_76_10661));
   NOR2_X1 i_257_76_10680 (.A1(n_257_76_10656), .A2(n_257_76_10661), .ZN(
      n_257_76_10662));
   NAND4_X1 i_257_76_10681 (.A1(n_257_76_10578), .A2(n_257_76_10563), .A3(
      n_257_76_10358), .A4(n_257_76_10312), .ZN(n_257_76_10663));
   INV_X1 i_257_76_10682 (.A(n_257_76_10663), .ZN(n_257_76_10664));
   NAND3_X1 i_257_76_10683 (.A1(n_257_76_10662), .A2(n_257_76_10475), .A3(
      n_257_76_10664), .ZN(n_257_76_10665));
   INV_X1 i_257_76_10684 (.A(n_257_76_10665), .ZN(n_257_76_10666));
   NAND2_X1 i_257_76_10685 (.A1(n_257_367), .A2(n_257_76_10316), .ZN(
      n_257_76_10667));
   NOR2_X1 i_257_76_10686 (.A1(n_257_76_10596), .A2(n_257_76_10667), .ZN(
      n_257_76_10668));
   NAND3_X1 i_257_76_10687 (.A1(n_257_76_10655), .A2(n_257_76_10666), .A3(
      n_257_76_10668), .ZN(n_257_76_10669));
   INV_X1 i_257_76_10688 (.A(n_257_76_10669), .ZN(n_257_76_10670));
   NAND2_X1 i_257_76_10689 (.A1(n_257_76_10281), .A2(n_257_76_10670), .ZN(
      n_257_76_10671));
   NAND4_X1 i_257_76_10690 (.A1(n_257_76_10283), .A2(n_257_76_10376), .A3(
      n_257_76_10321), .A4(n_257_76_10364), .ZN(n_257_76_10672));
   NOR2_X1 i_257_76_10691 (.A1(n_257_76_10671), .A2(n_257_76_10672), .ZN(
      n_257_76_10673));
   NAND2_X1 i_257_76_10692 (.A1(n_257_76_18082), .A2(n_257_76_10673), .ZN(
      n_257_76_10674));
   NAND3_X1 i_257_76_10693 (.A1(n_257_76_10637), .A2(n_257_76_10652), .A3(
      n_257_76_10674), .ZN(n_257_76_10675));
   INV_X1 i_257_76_10694 (.A(n_257_76_10675), .ZN(n_257_76_10676));
   NOR2_X1 i_257_76_10695 (.A1(n_257_76_10444), .A2(n_257_76_10527), .ZN(
      n_257_76_10677));
   NAND4_X1 i_257_76_10696 (.A1(n_257_210), .A2(n_257_76_10353), .A3(
      n_257_76_18023), .A4(n_257_76_10354), .ZN(n_257_76_10678));
   INV_X1 i_257_76_10697 (.A(n_257_76_10678), .ZN(n_257_76_10679));
   NAND2_X1 i_257_76_10698 (.A1(n_257_76_10300), .A2(n_257_427), .ZN(
      n_257_76_10680));
   INV_X1 i_257_76_10699 (.A(n_257_76_10680), .ZN(n_257_76_10681));
   NAND3_X1 i_257_76_10700 (.A1(n_257_76_10679), .A2(n_257_76_10681), .A3(
      n_257_76_10359), .ZN(n_257_76_10682));
   INV_X1 i_257_76_10701 (.A(n_257_76_10682), .ZN(n_257_76_10683));
   NAND3_X1 i_257_76_10702 (.A1(n_257_76_10316), .A2(n_257_76_10284), .A3(
      n_257_76_10683), .ZN(n_257_76_10684));
   INV_X1 i_257_76_10703 (.A(n_257_76_10684), .ZN(n_257_76_10685));
   NOR2_X1 i_257_76_10704 (.A1(n_257_76_10474), .A2(n_257_76_10442), .ZN(
      n_257_76_10686));
   NAND4_X1 i_257_76_10705 (.A1(n_257_76_10677), .A2(n_257_76_10685), .A3(
      n_257_76_10352), .A4(n_257_76_10686), .ZN(n_257_76_10687));
   INV_X1 i_257_76_10706 (.A(n_257_76_10687), .ZN(n_257_76_10688));
   NAND4_X1 i_257_76_10707 (.A1(n_257_76_10688), .A2(n_257_76_10281), .A3(
      n_257_76_10283), .A4(n_257_76_10418), .ZN(n_257_76_10689));
   INV_X1 i_257_76_10708 (.A(n_257_76_10689), .ZN(n_257_76_10690));
   NAND2_X1 i_257_76_10709 (.A1(n_257_76_18065), .A2(n_257_76_10690), .ZN(
      n_257_76_10691));
   NOR2_X1 i_257_76_10710 (.A1(n_257_76_10629), .A2(n_257_76_10452), .ZN(
      n_257_76_10692));
   NAND3_X1 i_257_76_10711 (.A1(n_257_76_10367), .A2(n_257_451), .A3(n_257_470), 
      .ZN(n_257_76_10693));
   NOR2_X1 i_257_76_10712 (.A1(n_257_76_10372), .A2(n_257_76_10693), .ZN(
      n_257_76_10694));
   NAND3_X1 i_257_76_10713 (.A1(n_257_76_10692), .A2(n_257_76_10321), .A3(
      n_257_76_10694), .ZN(n_257_76_10695));
   INV_X1 i_257_76_10714 (.A(n_257_76_10695), .ZN(n_257_76_10696));
   NAND3_X1 i_257_76_10715 (.A1(n_257_76_10696), .A2(n_257_76_10281), .A3(
      n_257_76_10283), .ZN(n_257_76_10697));
   INV_X1 i_257_76_10716 (.A(n_257_76_10697), .ZN(n_257_76_10698));
   NAND2_X1 i_257_76_10717 (.A1(n_257_76_18063), .A2(n_257_76_10698), .ZN(
      n_257_76_10699));
   NAND3_X1 i_257_76_10718 (.A1(n_257_76_10354), .A2(n_257_76_18023), .A3(
      n_257_424), .ZN(n_257_76_10700));
   INV_X1 i_257_76_10719 (.A(n_257_76_10700), .ZN(n_257_76_10701));
   NAND4_X1 i_257_76_10720 (.A1(n_257_76_10438), .A2(n_257_76_10359), .A3(
      n_257_519), .A4(n_257_76_10701), .ZN(n_257_76_10702));
   INV_X1 i_257_76_10721 (.A(n_257_76_10702), .ZN(n_257_76_10703));
   NAND3_X1 i_257_76_10722 (.A1(n_257_76_10316), .A2(n_257_76_10703), .A3(
      n_257_76_10284), .ZN(n_257_76_10704));
   INV_X1 i_257_76_10723 (.A(n_257_76_10704), .ZN(n_257_76_10705));
   NAND3_X1 i_257_76_10724 (.A1(n_257_76_10364), .A2(n_257_76_10705), .A3(
      n_257_76_10352), .ZN(n_257_76_10706));
   INV_X1 i_257_76_10725 (.A(n_257_76_10706), .ZN(n_257_76_10707));
   NAND2_X1 i_257_76_10726 (.A1(n_257_76_10311), .A2(n_257_76_10367), .ZN(
      n_257_76_10708));
   NAND4_X1 i_257_76_10727 (.A1(n_257_76_10312), .A2(n_257_76_10303), .A3(
      n_257_76_10304), .A4(n_257_76_10368), .ZN(n_257_76_10709));
   NOR2_X1 i_257_76_10728 (.A1(n_257_76_10708), .A2(n_257_76_10709), .ZN(
      n_257_76_10710));
   NAND3_X1 i_257_76_10729 (.A1(n_257_76_10346), .A2(n_257_76_10317), .A3(
      n_257_76_10348), .ZN(n_257_76_10711));
   INV_X1 i_257_76_10730 (.A(n_257_76_10711), .ZN(n_257_76_10712));
   NAND4_X1 i_257_76_10731 (.A1(n_257_76_10318), .A2(n_257_76_10349), .A3(
      n_257_76_10307), .A4(n_257_76_10308), .ZN(n_257_76_10713));
   INV_X1 i_257_76_10732 (.A(n_257_76_10713), .ZN(n_257_76_10714));
   NAND3_X1 i_257_76_10733 (.A1(n_257_76_10710), .A2(n_257_76_10712), .A3(
      n_257_76_10714), .ZN(n_257_76_10715));
   INV_X1 i_257_76_10734 (.A(n_257_76_10715), .ZN(n_257_76_10716));
   NAND4_X1 i_257_76_10735 (.A1(n_257_76_10707), .A2(n_257_76_10716), .A3(
      n_257_76_10376), .A4(n_257_76_10321), .ZN(n_257_76_10717));
   NOR2_X1 i_257_76_10736 (.A1(n_257_76_10717), .A2(n_257_76_10650), .ZN(
      n_257_76_10718));
   NAND2_X1 i_257_76_10737 (.A1(n_257_76_18062), .A2(n_257_76_10718), .ZN(
      n_257_76_10719));
   NAND3_X1 i_257_76_10738 (.A1(n_257_76_10691), .A2(n_257_76_10699), .A3(
      n_257_76_10719), .ZN(n_257_76_10720));
   INV_X1 i_257_76_10739 (.A(n_257_76_10720), .ZN(n_257_76_10721));
   NAND4_X1 i_257_76_10740 (.A1(n_257_76_10455), .A2(n_257_76_10283), .A3(
      n_257_76_10376), .A4(n_257_76_10321), .ZN(n_257_76_10722));
   NAND4_X1 i_257_76_10741 (.A1(n_257_76_10353), .A2(n_257_76_18023), .A3(
      n_257_76_10354), .A4(n_257_422), .ZN(n_257_76_10723));
   INV_X1 i_257_76_10742 (.A(n_257_76_10723), .ZN(n_257_76_10724));
   NAND4_X1 i_257_76_10743 (.A1(n_257_76_10567), .A2(n_257_76_10724), .A3(
      n_257_76_10359), .A4(n_257_328), .ZN(n_257_76_10725));
   NAND4_X1 i_257_76_10744 (.A1(n_257_76_10358), .A2(n_257_76_10312), .A3(
      n_257_76_10303), .A4(n_257_76_10304), .ZN(n_257_76_10726));
   NOR2_X1 i_257_76_10745 (.A1(n_257_76_10725), .A2(n_257_76_10726), .ZN(
      n_257_76_10727));
   NAND4_X1 i_257_76_10746 (.A1(n_257_76_10348), .A2(n_257_76_10318), .A3(
      n_257_76_10367), .A4(n_257_76_10563), .ZN(n_257_76_10728));
   INV_X1 i_257_76_10747 (.A(n_257_76_10728), .ZN(n_257_76_10729));
   INV_X1 i_257_76_10748 (.A(n_257_76_10558), .ZN(n_257_76_10730));
   NAND3_X1 i_257_76_10749 (.A1(n_257_76_10727), .A2(n_257_76_10729), .A3(
      n_257_76_10730), .ZN(n_257_76_10731));
   INV_X1 i_257_76_10750 (.A(n_257_76_10731), .ZN(n_257_76_10732));
   NAND2_X1 i_257_76_10751 (.A1(n_257_76_10281), .A2(n_257_76_10732), .ZN(
      n_257_76_10733));
   NOR2_X1 i_257_76_10752 (.A1(n_257_76_10722), .A2(n_257_76_10733), .ZN(
      n_257_76_10734));
   NAND2_X1 i_257_76_10753 (.A1(n_257_342), .A2(n_257_76_10734), .ZN(
      n_257_76_10735));
   NAND2_X1 i_257_76_10754 (.A1(n_257_76_10358), .A2(n_257_76_10312), .ZN(
      n_257_76_10736));
   INV_X1 i_257_76_10755 (.A(n_257_76_10736), .ZN(n_257_76_10737));
   INV_X1 i_257_76_10756 (.A(n_257_76_10656), .ZN(n_257_76_10738));
   NAND2_X1 i_257_76_10757 (.A1(n_257_428), .A2(n_257_583), .ZN(n_257_76_10739));
   NAND3_X1 i_257_76_10758 (.A1(n_257_484), .A2(n_257_406), .A3(n_257_442), 
      .ZN(n_257_76_10740));
   INV_X1 i_257_76_10759 (.A(n_257_76_10740), .ZN(n_257_76_10741));
   NAND2_X1 i_257_76_10760 (.A1(n_257_76_10739), .A2(n_257_76_10741), .ZN(
      n_257_76_10742));
   INV_X1 i_257_76_10761 (.A(n_257_76_10742), .ZN(n_257_76_10743));
   NAND2_X1 i_257_76_10762 (.A1(n_257_420), .A2(n_257_487), .ZN(n_257_76_10744));
   NAND4_X1 i_257_76_10763 (.A1(n_257_76_10353), .A2(n_257_76_10743), .A3(
      n_257_76_10744), .A4(n_257_76_10354), .ZN(n_257_76_10745));
   NOR2_X1 i_257_76_10764 (.A1(n_257_76_10566), .A2(n_257_76_10745), .ZN(
      n_257_76_10746));
   NAND3_X1 i_257_76_10765 (.A1(n_257_76_10737), .A2(n_257_76_10738), .A3(
      n_257_76_10746), .ZN(n_257_76_10747));
   NAND4_X1 i_257_76_10766 (.A1(n_257_76_10311), .A2(n_257_76_10367), .A3(
      n_257_76_10578), .A4(n_257_76_10563), .ZN(n_257_76_10748));
   NOR2_X1 i_257_76_10767 (.A1(n_257_76_10747), .A2(n_257_76_10748), .ZN(
      n_257_76_10749));
   NAND3_X1 i_257_76_10768 (.A1(n_257_76_10321), .A2(n_257_76_10749), .A3(
      n_257_76_10364), .ZN(n_257_76_10750));
   INV_X1 i_257_76_10769 (.A(n_257_76_10750), .ZN(n_257_76_10751));
   NAND2_X1 i_257_76_10770 (.A1(n_257_76_10284), .A2(n_257_76_10346), .ZN(
      n_257_76_10752));
   INV_X1 i_257_76_10771 (.A(n_257_76_10752), .ZN(n_257_76_10753));
   NAND3_X1 i_257_76_10772 (.A1(n_257_76_10317), .A2(n_257_76_10348), .A3(
      n_257_76_10318), .ZN(n_257_76_10754));
   INV_X1 i_257_76_10773 (.A(n_257_76_10754), .ZN(n_257_76_10755));
   NAND3_X1 i_257_76_10774 (.A1(n_257_76_10349), .A2(n_257_76_10307), .A3(
      n_257_76_10308), .ZN(n_257_76_10756));
   INV_X1 i_257_76_10775 (.A(n_257_76_10756), .ZN(n_257_76_10757));
   NAND3_X1 i_257_76_10776 (.A1(n_257_76_10753), .A2(n_257_76_10755), .A3(
      n_257_76_10757), .ZN(n_257_76_10758));
   NAND3_X1 i_257_76_10777 (.A1(n_257_76_10553), .A2(n_257_76_10352), .A3(
      n_257_76_10316), .ZN(n_257_76_10759));
   NOR2_X1 i_257_76_10778 (.A1(n_257_76_10758), .A2(n_257_76_10759), .ZN(
      n_257_76_10760));
   NAND4_X1 i_257_76_10779 (.A1(n_257_76_10585), .A2(n_257_76_10751), .A3(
      n_257_76_10281), .A4(n_257_76_10760), .ZN(n_257_76_10761));
   INV_X1 i_257_76_10780 (.A(n_257_76_10761), .ZN(n_257_76_10762));
   NAND2_X1 i_257_76_10781 (.A1(n_257_76_18060), .A2(n_257_76_10762), .ZN(
      n_257_76_10763));
   INV_X1 i_257_76_10782 (.A(n_257_76_10326), .ZN(n_257_76_10764));
   NAND2_X1 i_257_76_10783 (.A1(n_257_446), .A2(n_257_76_10764), .ZN(
      n_257_76_10765));
   NAND2_X1 i_257_76_10784 (.A1(n_257_449), .A2(n_257_76_15108), .ZN(
      n_257_76_10766));
   INV_X1 i_257_76_10785 (.A(n_257_76_10606), .ZN(n_257_76_10767));
   NAND2_X1 i_257_76_10786 (.A1(n_257_447), .A2(n_257_76_10767), .ZN(
      n_257_76_10768));
   NAND3_X1 i_257_76_10787 (.A1(n_257_76_10765), .A2(n_257_76_10766), .A3(
      n_257_76_10768), .ZN(n_257_76_10769));
   NAND2_X1 i_257_76_10788 (.A1(n_257_647), .A2(n_257_76_17928), .ZN(
      n_257_76_10770));
   INV_X1 i_257_76_10789 (.A(Small_Packet_Data_Size[18]), .ZN(n_257_76_10771));
   NAND2_X1 i_257_76_10790 (.A1(n_257_76_10739), .A2(n_257_76_18026), .ZN(
      n_257_76_10772));
   INV_X1 i_257_76_10791 (.A(n_257_76_10772), .ZN(n_257_76_10773));
   NAND3_X1 i_257_76_10792 (.A1(n_257_76_10773), .A2(n_257_76_10353), .A3(
      n_257_76_10744), .ZN(n_257_76_10774));
   NAND2_X1 i_257_76_10793 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[18]), 
      .ZN(n_257_76_10775));
   NAND2_X1 i_257_76_10794 (.A1(n_257_76_10774), .A2(n_257_76_10775), .ZN(
      n_257_76_10776));
   NAND2_X1 i_257_76_10795 (.A1(n_257_879), .A2(n_257_76_17903), .ZN(
      n_257_76_10777));
   NAND3_X1 i_257_76_10796 (.A1(n_257_76_10770), .A2(n_257_76_10776), .A3(
      n_257_76_10777), .ZN(n_257_76_10778));
   NAND3_X1 i_257_76_10797 (.A1(n_257_719), .A2(n_257_435), .A3(n_257_442), 
      .ZN(n_257_76_10779));
   NAND2_X1 i_257_76_10798 (.A1(n_257_76_10779), .A2(n_257_76_10470), .ZN(
      n_257_76_10780));
   INV_X1 i_257_76_10799 (.A(n_257_76_10780), .ZN(n_257_76_10781));
   INV_X1 i_257_76_10800 (.A(n_257_76_10285), .ZN(n_257_76_10782));
   NAND2_X1 i_257_76_10801 (.A1(n_257_440), .A2(n_257_76_10782), .ZN(
      n_257_76_10783));
   NAND2_X1 i_257_76_10802 (.A1(n_257_438), .A2(n_257_76_13741), .ZN(
      n_257_76_10784));
   NAND2_X1 i_257_76_10803 (.A1(n_257_53), .A2(n_257_76_17918), .ZN(
      n_257_76_10785));
   NAND4_X1 i_257_76_10804 (.A1(n_257_76_10781), .A2(n_257_76_10783), .A3(
      n_257_76_10784), .A4(n_257_76_10785), .ZN(n_257_76_10786));
   NOR3_X1 i_257_76_10805 (.A1(n_257_76_10769), .A2(n_257_76_10778), .A3(
      n_257_76_10786), .ZN(n_257_76_10787));
   NAND2_X1 i_257_76_10806 (.A1(n_257_93), .A2(n_257_76_17932), .ZN(
      n_257_76_10788));
   NAND2_X1 i_257_76_10807 (.A1(n_257_751), .A2(n_257_76_17935), .ZN(
      n_257_76_10789));
   NAND3_X1 i_257_76_10808 (.A1(n_257_76_10788), .A2(n_257_76_10360), .A3(
      n_257_76_10789), .ZN(n_257_76_10790));
   INV_X1 i_257_76_10809 (.A(n_257_76_10790), .ZN(n_257_76_10791));
   NAND2_X1 i_257_76_10810 (.A1(n_257_170), .A2(n_257_76_17331), .ZN(
      n_257_76_10792));
   NAND2_X1 i_257_76_10811 (.A1(n_257_981), .A2(n_257_442), .ZN(n_257_76_10793));
   INV_X1 i_257_76_10812 (.A(n_257_76_10793), .ZN(n_257_76_10794));
   NAND2_X1 i_257_76_10813 (.A1(n_257_441), .A2(n_257_76_10794), .ZN(
      n_257_76_10795));
   NAND2_X1 i_257_76_10814 (.A1(n_257_815), .A2(n_257_76_17952), .ZN(
      n_257_76_10796));
   NAND3_X1 i_257_76_10815 (.A1(n_257_76_10795), .A2(n_257_76_10702), .A3(
      n_257_76_10796), .ZN(n_257_76_10797));
   NAND2_X1 i_257_76_10816 (.A1(n_257_131), .A2(n_257_76_17925), .ZN(
      n_257_76_10798));
   NAND2_X1 i_257_76_10817 (.A1(n_257_917), .A2(n_257_76_17940), .ZN(
      n_257_76_10799));
   NAND3_X1 i_257_76_10818 (.A1(n_257_76_10682), .A2(n_257_76_10798), .A3(
      n_257_76_10799), .ZN(n_257_76_10800));
   NOR2_X1 i_257_76_10819 (.A1(n_257_76_10797), .A2(n_257_76_10800), .ZN(
      n_257_76_10801));
   NAND4_X1 i_257_76_10820 (.A1(n_257_76_10787), .A2(n_257_76_10791), .A3(
      n_257_76_10792), .A4(n_257_76_10801), .ZN(n_257_76_10802));
   NAND2_X1 i_257_76_10821 (.A1(n_257_687), .A2(n_257_76_17958), .ZN(
      n_257_76_10803));
   INV_X1 i_257_76_10822 (.A(n_257_815), .ZN(n_257_76_10804));
   NAND2_X1 i_257_76_10823 (.A1(n_257_76_10804), .A2(n_257_442), .ZN(
      n_257_76_10805));
   INV_X1 i_257_76_10824 (.A(n_257_917), .ZN(n_257_76_10806));
   NAND2_X1 i_257_76_10825 (.A1(n_257_76_10806), .A2(n_257_442), .ZN(
      n_257_76_10807));
   NAND3_X1 i_257_76_10826 (.A1(n_257_76_10805), .A2(n_257_76_10807), .A3(
      n_257_76_13029), .ZN(n_257_76_10808));
   INV_X1 i_257_76_10827 (.A(n_257_76_10349), .ZN(n_257_76_10809));
   NAND2_X1 i_257_76_10828 (.A1(n_257_76_10808), .A2(n_257_76_10809), .ZN(
      n_257_76_10810));
   NAND4_X1 i_257_76_10829 (.A1(n_257_76_10731), .A2(n_257_76_10803), .A3(
      n_257_76_10448), .A4(n_257_76_10810), .ZN(n_257_76_10811));
   NOR2_X1 i_257_76_10830 (.A1(n_257_76_10802), .A2(n_257_76_10811), .ZN(
      n_257_76_10812));
   NAND2_X1 i_257_76_10831 (.A1(n_257_1045), .A2(n_257_76_17969), .ZN(
      n_257_76_10813));
   NAND2_X1 i_257_76_10832 (.A1(n_257_1013), .A2(n_257_76_17964), .ZN(
      n_257_76_10814));
   NAND3_X1 i_257_76_10833 (.A1(n_257_76_10813), .A2(n_257_76_10669), .A3(
      n_257_76_10814), .ZN(n_257_76_10815));
   INV_X1 i_257_76_10834 (.A(n_257_76_10815), .ZN(n_257_76_10816));
   NAND3_X1 i_257_76_10835 (.A1(n_257_76_10812), .A2(n_257_76_10816), .A3(
      n_257_76_10649), .ZN(n_257_76_10817));
   NAND3_X1 i_257_76_10836 (.A1(n_257_76_10735), .A2(n_257_76_10763), .A3(
      n_257_76_10817), .ZN(n_257_76_10818));
   INV_X1 i_257_76_10837 (.A(n_257_76_10818), .ZN(n_257_76_10819));
   NAND3_X1 i_257_76_10838 (.A1(n_257_76_10676), .A2(n_257_76_10721), .A3(
      n_257_76_10819), .ZN(n_257_76_10820));
   NOR2_X1 i_257_76_10839 (.A1(n_257_76_10626), .A2(n_257_76_10820), .ZN(
      n_257_76_10821));
   NAND2_X1 i_257_76_10840 (.A1(n_257_76_10504), .A2(n_257_76_10821), .ZN(n_18));
   NAND2_X1 i_257_76_10841 (.A1(n_257_1046), .A2(n_257_443), .ZN(n_257_76_10822));
   NAND2_X1 i_257_76_10842 (.A1(n_257_1014), .A2(n_257_444), .ZN(n_257_76_10823));
   NAND2_X1 i_257_76_10843 (.A1(n_257_441), .A2(n_257_982), .ZN(n_257_76_10824));
   INV_X1 i_257_76_10844 (.A(n_257_1078), .ZN(n_257_76_10825));
   NAND2_X1 i_257_76_10845 (.A1(n_257_950), .A2(n_257_442), .ZN(n_257_76_10826));
   INV_X1 i_257_76_10846 (.A(n_257_76_10826), .ZN(n_257_76_10827));
   NAND3_X1 i_257_76_10847 (.A1(n_257_440), .A2(n_257_76_10825), .A3(
      n_257_76_10827), .ZN(n_257_76_10828));
   INV_X1 i_257_76_10848 (.A(n_257_76_10828), .ZN(n_257_76_10829));
   NAND2_X1 i_257_76_10849 (.A1(n_257_76_10824), .A2(n_257_76_10829), .ZN(
      n_257_76_10830));
   INV_X1 i_257_76_10850 (.A(n_257_76_10830), .ZN(n_257_76_10831));
   NAND2_X1 i_257_76_10851 (.A1(n_257_76_10823), .A2(n_257_76_10831), .ZN(
      n_257_76_10832));
   INV_X1 i_257_76_10852 (.A(n_257_76_10832), .ZN(n_257_76_10833));
   NAND2_X1 i_257_76_10853 (.A1(n_257_76_10822), .A2(n_257_76_10833), .ZN(
      n_257_76_10834));
   INV_X1 i_257_76_10854 (.A(n_257_76_10834), .ZN(n_257_76_10835));
   NAND2_X1 i_257_76_10855 (.A1(n_257_17), .A2(n_257_76_10835), .ZN(
      n_257_76_10836));
   NOR2_X1 i_257_76_10856 (.A1(n_257_1078), .A2(n_257_76_17412), .ZN(
      n_257_76_10837));
   INV_X1 i_257_76_10857 (.A(n_257_76_10837), .ZN(n_257_76_10838));
   NOR2_X1 i_257_76_10858 (.A1(n_257_76_10838), .A2(n_257_76_15197), .ZN(
      n_257_76_10839));
   NAND2_X1 i_257_76_10859 (.A1(n_257_1046), .A2(n_257_76_10839), .ZN(
      n_257_76_10840));
   INV_X1 i_257_76_10860 (.A(n_257_76_10840), .ZN(n_257_76_10841));
   NAND2_X1 i_257_76_10861 (.A1(n_257_76_18072), .A2(n_257_76_10841), .ZN(
      n_257_76_10842));
   NAND2_X1 i_257_76_10862 (.A1(n_257_447), .A2(n_257_784), .ZN(n_257_76_10843));
   NAND2_X1 i_257_76_10863 (.A1(n_257_880), .A2(n_257_445), .ZN(n_257_76_10844));
   NAND3_X1 i_257_76_10864 (.A1(n_257_76_10843), .A2(n_257_648), .A3(
      n_257_76_10844), .ZN(n_257_76_10845));
   INV_X1 i_257_76_10865 (.A(n_257_76_10845), .ZN(n_257_76_10846));
   NAND2_X1 i_257_76_10866 (.A1(n_257_446), .A2(n_257_848), .ZN(n_257_76_10847));
   NAND2_X1 i_257_76_10867 (.A1(n_257_449), .A2(n_257_894), .ZN(n_257_76_10848));
   NAND2_X1 i_257_76_10868 (.A1(n_257_76_10847), .A2(n_257_76_10848), .ZN(
      n_257_76_10849));
   INV_X1 i_257_76_10869 (.A(n_257_76_10849), .ZN(n_257_76_10850));
   OAI21_X1 i_257_76_10870 (.A(n_257_76_17761), .B1(n_257_720), .B2(
      n_257_76_17412), .ZN(n_257_76_10851));
   NAND2_X1 i_257_76_10871 (.A1(n_257_440), .A2(n_257_950), .ZN(n_257_76_10852));
   NAND2_X1 i_257_76_10872 (.A1(n_257_438), .A2(n_257_1084), .ZN(n_257_76_10853));
   NOR2_X1 i_257_76_10873 (.A1(n_257_1078), .A2(n_257_76_14694), .ZN(
      n_257_76_10854));
   NAND4_X1 i_257_76_10874 (.A1(n_257_76_10851), .A2(n_257_76_10852), .A3(
      n_257_76_10853), .A4(n_257_76_10854), .ZN(n_257_76_10855));
   INV_X1 i_257_76_10875 (.A(n_257_76_10855), .ZN(n_257_76_10856));
   NAND3_X1 i_257_76_10876 (.A1(n_257_76_10846), .A2(n_257_76_10850), .A3(
      n_257_76_10856), .ZN(n_257_76_10857));
   NAND2_X1 i_257_76_10877 (.A1(n_257_816), .A2(n_257_437), .ZN(n_257_76_10858));
   NAND2_X1 i_257_76_10878 (.A1(n_257_752), .A2(n_257_436), .ZN(n_257_76_10859));
   NAND2_X1 i_257_76_10879 (.A1(n_257_918), .A2(n_257_439), .ZN(n_257_76_10860));
   NAND4_X1 i_257_76_10880 (.A1(n_257_76_10858), .A2(n_257_76_10859), .A3(
      n_257_76_10824), .A4(n_257_76_10860), .ZN(n_257_76_10861));
   NOR2_X1 i_257_76_10881 (.A1(n_257_76_10857), .A2(n_257_76_10861), .ZN(
      n_257_76_10862));
   NAND2_X1 i_257_76_10882 (.A1(n_257_688), .A2(n_257_448), .ZN(n_257_76_10863));
   NAND3_X1 i_257_76_10883 (.A1(n_257_76_10862), .A2(n_257_76_10823), .A3(
      n_257_76_10863), .ZN(n_257_76_10864));
   INV_X1 i_257_76_10884 (.A(n_257_76_10864), .ZN(n_257_76_10865));
   NAND2_X1 i_257_76_10885 (.A1(n_257_76_10822), .A2(n_257_76_10865), .ZN(
      n_257_76_10866));
   INV_X1 i_257_76_10886 (.A(n_257_76_10866), .ZN(n_257_76_10867));
   NAND2_X1 i_257_76_10887 (.A1(n_257_28), .A2(n_257_76_10867), .ZN(
      n_257_76_10868));
   NAND3_X1 i_257_76_10888 (.A1(n_257_76_10836), .A2(n_257_76_10842), .A3(
      n_257_76_10868), .ZN(n_257_76_10869));
   NAND2_X1 i_257_76_10889 (.A1(n_257_76_10844), .A2(n_257_446), .ZN(
      n_257_76_10870));
   INV_X1 i_257_76_10890 (.A(n_257_76_10870), .ZN(n_257_76_10871));
   NAND2_X1 i_257_76_10891 (.A1(n_257_848), .A2(n_257_442), .ZN(n_257_76_10872));
   NOR2_X1 i_257_76_10892 (.A1(n_257_1078), .A2(n_257_76_10872), .ZN(
      n_257_76_10873));
   NAND3_X1 i_257_76_10893 (.A1(n_257_76_10852), .A2(n_257_76_10853), .A3(
      n_257_76_10873), .ZN(n_257_76_10874));
   INV_X1 i_257_76_10894 (.A(n_257_76_10874), .ZN(n_257_76_10875));
   NAND4_X1 i_257_76_10895 (.A1(n_257_76_10824), .A2(n_257_76_10871), .A3(
      n_257_76_10860), .A4(n_257_76_10875), .ZN(n_257_76_10876));
   INV_X1 i_257_76_10896 (.A(n_257_76_10876), .ZN(n_257_76_10877));
   NAND2_X1 i_257_76_10897 (.A1(n_257_76_10823), .A2(n_257_76_10877), .ZN(
      n_257_76_10878));
   INV_X1 i_257_76_10898 (.A(n_257_76_10878), .ZN(n_257_76_10879));
   NAND2_X1 i_257_76_10899 (.A1(n_257_76_10822), .A2(n_257_76_10879), .ZN(
      n_257_76_10880));
   INV_X1 i_257_76_10900 (.A(n_257_76_10880), .ZN(n_257_76_10881));
   NAND2_X1 i_257_76_10901 (.A1(n_257_76_18070), .A2(n_257_76_10881), .ZN(
      n_257_76_10882));
   NOR2_X1 i_257_76_10902 (.A1(n_257_76_10838), .A2(n_257_76_13028), .ZN(
      n_257_76_10883));
   NAND3_X1 i_257_76_10903 (.A1(n_257_76_10883), .A2(n_257_918), .A3(
      n_257_76_10852), .ZN(n_257_76_10884));
   INV_X1 i_257_76_10904 (.A(n_257_76_10824), .ZN(n_257_76_10885));
   NOR2_X1 i_257_76_10905 (.A1(n_257_76_10884), .A2(n_257_76_10885), .ZN(
      n_257_76_10886));
   NAND2_X1 i_257_76_10906 (.A1(n_257_76_10823), .A2(n_257_76_10886), .ZN(
      n_257_76_10887));
   INV_X1 i_257_76_10907 (.A(n_257_76_10887), .ZN(n_257_76_10888));
   NAND2_X1 i_257_76_10908 (.A1(n_257_76_10822), .A2(n_257_76_10888), .ZN(
      n_257_76_10889));
   INV_X1 i_257_76_10909 (.A(n_257_76_10889), .ZN(n_257_76_10890));
   NAND2_X1 i_257_76_10910 (.A1(n_257_76_18084), .A2(n_257_76_10890), .ZN(
      n_257_76_10891));
   INV_X1 i_257_76_10911 (.A(n_257_76_18020), .ZN(n_257_76_10892));
   NOR2_X1 i_257_76_10912 (.A1(n_257_76_10892), .A2(n_257_1078), .ZN(
      n_257_76_10893));
   NAND2_X1 i_257_76_10913 (.A1(n_257_211), .A2(n_257_427), .ZN(n_257_76_10894));
   NAND2_X1 i_257_76_10914 (.A1(n_257_720), .A2(n_257_435), .ZN(n_257_76_10895));
   NAND2_X1 i_257_76_10915 (.A1(n_257_432), .A2(n_257_616), .ZN(n_257_76_10896));
   NAND2_X1 i_257_76_10916 (.A1(n_257_76_10896), .A2(n_257_423), .ZN(
      n_257_76_10897));
   INV_X1 i_257_76_10917 (.A(n_257_76_10897), .ZN(n_257_76_10898));
   NAND4_X1 i_257_76_10918 (.A1(n_257_76_10893), .A2(n_257_76_10894), .A3(
      n_257_76_10895), .A4(n_257_76_10898), .ZN(n_257_76_10899));
   NAND2_X1 i_257_76_10919 (.A1(n_257_76_10852), .A2(n_257_76_10853), .ZN(
      n_257_76_10900));
   NOR2_X1 i_257_76_10920 (.A1(n_257_76_10899), .A2(n_257_76_10900), .ZN(
      n_257_76_10901));
   NAND2_X1 i_257_76_10921 (.A1(n_257_76_10848), .A2(n_257_76_10843), .ZN(
      n_257_76_10902));
   INV_X1 i_257_76_10922 (.A(n_257_76_10902), .ZN(n_257_76_10903));
   NAND2_X1 i_257_76_10923 (.A1(n_257_54), .A2(n_257_433), .ZN(n_257_76_10904));
   NAND2_X1 i_257_76_10924 (.A1(n_257_76_10904), .A2(n_257_76_10844), .ZN(
      n_257_76_10905));
   INV_X1 i_257_76_10925 (.A(n_257_76_10905), .ZN(n_257_76_10906));
   NAND3_X1 i_257_76_10926 (.A1(n_257_76_10901), .A2(n_257_76_10903), .A3(
      n_257_76_10906), .ZN(n_257_76_10907));
   NAND2_X1 i_257_76_10927 (.A1(n_257_451), .A2(n_257_471), .ZN(n_257_76_10908));
   NAND2_X1 i_257_76_10928 (.A1(n_257_648), .A2(n_257_450), .ZN(n_257_76_10909));
   NAND4_X1 i_257_76_10929 (.A1(n_257_76_10908), .A2(n_257_76_10909), .A3(
      n_257_291), .A4(n_257_76_10847), .ZN(n_257_76_10910));
   NOR2_X1 i_257_76_10930 (.A1(n_257_76_10907), .A2(n_257_76_10910), .ZN(
      n_257_76_10911));
   NAND2_X1 i_257_76_10931 (.A1(n_257_94), .A2(n_257_431), .ZN(n_257_76_10912));
   NAND2_X1 i_257_76_10932 (.A1(n_257_552), .A2(n_257_426), .ZN(n_257_76_10913));
   NAND2_X1 i_257_76_10933 (.A1(n_257_76_10912), .A2(n_257_76_10913), .ZN(
      n_257_76_10914));
   INV_X1 i_257_76_10934 (.A(n_257_76_10914), .ZN(n_257_76_10915));
   NAND2_X1 i_257_76_10935 (.A1(n_257_520), .A2(n_257_424), .ZN(n_257_76_10916));
   NAND3_X1 i_257_76_10936 (.A1(n_257_76_10916), .A2(n_257_76_10858), .A3(
      n_257_76_10859), .ZN(n_257_76_10917));
   NAND2_X1 i_257_76_10937 (.A1(n_257_132), .A2(n_257_430), .ZN(n_257_76_10918));
   NAND3_X1 i_257_76_10938 (.A1(n_257_76_10824), .A2(n_257_76_10918), .A3(
      n_257_76_10860), .ZN(n_257_76_10919));
   NOR2_X1 i_257_76_10939 (.A1(n_257_76_10917), .A2(n_257_76_10919), .ZN(
      n_257_76_10920));
   NAND3_X1 i_257_76_10940 (.A1(n_257_76_10911), .A2(n_257_76_10915), .A3(
      n_257_76_10920), .ZN(n_257_76_10921));
   NAND2_X1 i_257_76_10941 (.A1(n_257_171), .A2(n_257_429), .ZN(n_257_76_10922));
   NAND2_X1 i_257_76_10942 (.A1(n_257_251), .A2(n_257_425), .ZN(n_257_76_10923));
   NAND2_X1 i_257_76_10943 (.A1(n_257_76_10922), .A2(n_257_76_10923), .ZN(
      n_257_76_10924));
   INV_X1 i_257_76_10944 (.A(n_257_76_10924), .ZN(n_257_76_10925));
   NAND3_X1 i_257_76_10945 (.A1(n_257_76_10925), .A2(n_257_76_10823), .A3(
      n_257_76_10863), .ZN(n_257_76_10926));
   NOR2_X1 i_257_76_10946 (.A1(n_257_76_10921), .A2(n_257_76_10926), .ZN(
      n_257_76_10927));
   NAND2_X1 i_257_76_10947 (.A1(n_257_76_10822), .A2(n_257_76_10927), .ZN(
      n_257_76_10928));
   INV_X1 i_257_76_10948 (.A(n_257_76_10928), .ZN(n_257_76_10929));
   NAND2_X1 i_257_76_10949 (.A1(n_257_76_18066), .A2(n_257_76_10929), .ZN(
      n_257_76_10930));
   NAND3_X1 i_257_76_10950 (.A1(n_257_76_10882), .A2(n_257_76_10891), .A3(
      n_257_76_10930), .ZN(n_257_76_10931));
   NOR2_X1 i_257_76_10951 (.A1(n_257_76_10869), .A2(n_257_76_10931), .ZN(
      n_257_76_10932));
   NAND2_X1 i_257_76_10952 (.A1(n_257_982), .A2(n_257_76_10837), .ZN(
      n_257_76_10933));
   NOR2_X1 i_257_76_10953 (.A1(n_257_76_13147), .A2(n_257_76_10933), .ZN(
      n_257_76_10934));
   NAND2_X1 i_257_76_10954 (.A1(n_257_76_10823), .A2(n_257_76_10934), .ZN(
      n_257_76_10935));
   INV_X1 i_257_76_10955 (.A(n_257_76_10935), .ZN(n_257_76_10936));
   NAND2_X1 i_257_76_10956 (.A1(n_257_76_10822), .A2(n_257_76_10936), .ZN(
      n_257_76_10937));
   INV_X1 i_257_76_10957 (.A(n_257_76_10937), .ZN(n_257_76_10938));
   NAND2_X1 i_257_76_10958 (.A1(n_257_76_18071), .A2(n_257_76_10938), .ZN(
      n_257_76_10939));
   NAND3_X1 i_257_76_10959 (.A1(n_257_76_10825), .A2(n_257_720), .A3(
      n_257_76_15655), .ZN(n_257_76_10940));
   INV_X1 i_257_76_10960 (.A(n_257_76_10940), .ZN(n_257_76_10941));
   NAND4_X1 i_257_76_10961 (.A1(n_257_76_10844), .A2(n_257_76_10941), .A3(
      n_257_76_10852), .A4(n_257_76_10853), .ZN(n_257_76_10942));
   INV_X1 i_257_76_10962 (.A(n_257_76_10942), .ZN(n_257_76_10943));
   NAND2_X1 i_257_76_10963 (.A1(n_257_76_10847), .A2(n_257_76_10843), .ZN(
      n_257_76_10944));
   INV_X1 i_257_76_10964 (.A(n_257_76_10944), .ZN(n_257_76_10945));
   NAND3_X1 i_257_76_10965 (.A1(n_257_76_10943), .A2(n_257_76_10945), .A3(
      n_257_76_10860), .ZN(n_257_76_10946));
   NAND3_X1 i_257_76_10966 (.A1(n_257_76_10858), .A2(n_257_76_10859), .A3(
      n_257_76_10824), .ZN(n_257_76_10947));
   NOR2_X1 i_257_76_10967 (.A1(n_257_76_10946), .A2(n_257_76_10947), .ZN(
      n_257_76_10948));
   NAND2_X1 i_257_76_10968 (.A1(n_257_76_10823), .A2(n_257_76_10948), .ZN(
      n_257_76_10949));
   INV_X1 i_257_76_10969 (.A(n_257_76_10949), .ZN(n_257_76_10950));
   NAND2_X1 i_257_76_10970 (.A1(n_257_76_10822), .A2(n_257_76_10950), .ZN(
      n_257_76_10951));
   INV_X1 i_257_76_10971 (.A(n_257_76_10951), .ZN(n_257_76_10952));
   NAND2_X1 i_257_76_10972 (.A1(n_257_76_18078), .A2(n_257_76_10952), .ZN(
      n_257_76_10953));
   NAND3_X1 i_257_76_10973 (.A1(n_257_76_10918), .A2(n_257_76_10860), .A3(
      n_257_76_10908), .ZN(n_257_76_10954));
   NOR2_X1 i_257_76_10974 (.A1(n_257_76_10947), .A2(n_257_76_10954), .ZN(
      n_257_76_10955));
   NAND4_X1 i_257_76_10975 (.A1(n_257_76_10909), .A2(n_257_76_10847), .A3(
      n_257_76_10848), .A4(n_257_76_10843), .ZN(n_257_76_10956));
   INV_X1 i_257_76_10976 (.A(n_257_76_10900), .ZN(n_257_76_10957));
   NAND3_X1 i_257_76_10977 (.A1(n_257_584), .A2(n_257_428), .A3(n_257_442), 
      .ZN(n_257_76_10958));
   INV_X1 i_257_76_10978 (.A(n_257_76_10958), .ZN(n_257_76_10959));
   NAND2_X1 i_257_76_10979 (.A1(n_257_76_10896), .A2(n_257_76_10959), .ZN(
      n_257_76_10960));
   INV_X1 i_257_76_10980 (.A(n_257_76_10960), .ZN(n_257_76_10961));
   NAND3_X1 i_257_76_10981 (.A1(n_257_76_10895), .A2(n_257_76_10961), .A3(
      n_257_76_10825), .ZN(n_257_76_10962));
   INV_X1 i_257_76_10982 (.A(n_257_76_10962), .ZN(n_257_76_10963));
   NAND4_X1 i_257_76_10983 (.A1(n_257_76_10957), .A2(n_257_76_10963), .A3(
      n_257_76_10904), .A4(n_257_76_10844), .ZN(n_257_76_10964));
   NOR2_X1 i_257_76_10984 (.A1(n_257_76_10956), .A2(n_257_76_10964), .ZN(
      n_257_76_10965));
   NAND4_X1 i_257_76_10985 (.A1(n_257_76_10922), .A2(n_257_76_10955), .A3(
      n_257_76_10912), .A4(n_257_76_10965), .ZN(n_257_76_10966));
   NAND2_X1 i_257_76_10986 (.A1(n_257_76_10823), .A2(n_257_76_10863), .ZN(
      n_257_76_10967));
   NOR2_X1 i_257_76_10987 (.A1(n_257_76_10966), .A2(n_257_76_10967), .ZN(
      n_257_76_10968));
   NAND2_X1 i_257_76_10988 (.A1(n_257_76_10822), .A2(n_257_76_10968), .ZN(
      n_257_76_10969));
   INV_X1 i_257_76_10989 (.A(n_257_76_10969), .ZN(n_257_76_10970));
   NAND2_X1 i_257_76_10990 (.A1(n_257_76_18074), .A2(n_257_76_10970), .ZN(
      n_257_76_10971));
   NAND3_X1 i_257_76_10991 (.A1(n_257_76_10939), .A2(n_257_76_10953), .A3(
      n_257_76_10971), .ZN(n_257_76_10972));
   NAND2_X1 i_257_76_10992 (.A1(n_257_1078), .A2(n_257_442), .ZN(n_257_76_10973));
   INV_X1 i_257_76_10993 (.A(n_257_76_10973), .ZN(n_257_76_10974));
   NAND2_X1 i_257_76_10994 (.A1(n_257_13), .A2(n_257_76_10974), .ZN(
      n_257_76_10975));
   NOR2_X1 i_257_76_10995 (.A1(n_257_76_17902), .A2(n_257_1078), .ZN(
      n_257_76_10976));
   NAND4_X1 i_257_76_10996 (.A1(n_257_76_10976), .A2(n_257_76_10852), .A3(
      n_257_76_10853), .A4(n_257_880), .ZN(n_257_76_10977));
   INV_X1 i_257_76_10997 (.A(n_257_76_10977), .ZN(n_257_76_10978));
   NAND3_X1 i_257_76_10998 (.A1(n_257_76_10978), .A2(n_257_76_10824), .A3(
      n_257_76_10860), .ZN(n_257_76_10979));
   INV_X1 i_257_76_10999 (.A(n_257_76_10979), .ZN(n_257_76_10980));
   NAND2_X1 i_257_76_11000 (.A1(n_257_76_10823), .A2(n_257_76_10980), .ZN(
      n_257_76_10981));
   INV_X1 i_257_76_11001 (.A(n_257_76_10981), .ZN(n_257_76_10982));
   NAND2_X1 i_257_76_11002 (.A1(n_257_76_10822), .A2(n_257_76_10982), .ZN(
      n_257_76_10983));
   INV_X1 i_257_76_11003 (.A(n_257_76_10983), .ZN(n_257_76_10984));
   NAND2_X1 i_257_76_11004 (.A1(n_257_76_18077), .A2(n_257_76_10984), .ZN(
      n_257_76_10985));
   NAND2_X1 i_257_76_11005 (.A1(n_257_76_10975), .A2(n_257_76_10985), .ZN(
      n_257_76_10986));
   NOR2_X1 i_257_76_11006 (.A1(n_257_76_10972), .A2(n_257_76_10986), .ZN(
      n_257_76_10987));
   NAND3_X1 i_257_76_11007 (.A1(n_257_76_10823), .A2(n_257_76_10863), .A3(
      n_257_76_10922), .ZN(n_257_76_10988));
   NAND4_X1 i_257_76_11008 (.A1(n_257_76_10847), .A2(n_257_76_10848), .A3(
      n_257_76_10843), .A4(n_257_76_10904), .ZN(n_257_76_10989));
   NAND3_X1 i_257_76_11009 (.A1(n_257_76_18020), .A2(n_257_76_10896), .A3(
      n_257_426), .ZN(n_257_76_10990));
   NOR2_X1 i_257_76_11010 (.A1(n_257_76_10990), .A2(n_257_1078), .ZN(
      n_257_76_10991));
   NAND2_X1 i_257_76_11011 (.A1(n_257_76_10894), .A2(n_257_76_10895), .ZN(
      n_257_76_10992));
   INV_X1 i_257_76_11012 (.A(n_257_76_10992), .ZN(n_257_76_10993));
   NAND4_X1 i_257_76_11013 (.A1(n_257_76_10957), .A2(n_257_76_10991), .A3(
      n_257_76_10844), .A4(n_257_76_10993), .ZN(n_257_76_10994));
   NOR2_X1 i_257_76_11014 (.A1(n_257_76_10989), .A2(n_257_76_10994), .ZN(
      n_257_76_10995));
   NAND4_X1 i_257_76_11015 (.A1(n_257_76_10858), .A2(n_257_76_10859), .A3(
      n_257_76_10824), .A4(n_257_76_10918), .ZN(n_257_76_10996));
   INV_X1 i_257_76_11016 (.A(n_257_76_10996), .ZN(n_257_76_10997));
   NAND4_X1 i_257_76_11017 (.A1(n_257_552), .A2(n_257_76_10860), .A3(
      n_257_76_10908), .A4(n_257_76_10909), .ZN(n_257_76_10998));
   INV_X1 i_257_76_11018 (.A(n_257_76_10998), .ZN(n_257_76_10999));
   NAND4_X1 i_257_76_11019 (.A1(n_257_76_10995), .A2(n_257_76_10997), .A3(
      n_257_76_10912), .A4(n_257_76_10999), .ZN(n_257_76_11000));
   NOR2_X1 i_257_76_11020 (.A1(n_257_76_10988), .A2(n_257_76_11000), .ZN(
      n_257_76_11001));
   NAND2_X1 i_257_76_11021 (.A1(n_257_76_10822), .A2(n_257_76_11001), .ZN(
      n_257_76_11002));
   INV_X1 i_257_76_11022 (.A(n_257_76_11002), .ZN(n_257_76_11003));
   NAND2_X1 i_257_76_11023 (.A1(n_257_76_18076), .A2(n_257_76_11003), .ZN(
      n_257_76_11004));
   NAND2_X1 i_257_76_11024 (.A1(n_257_752), .A2(n_257_76_10847), .ZN(
      n_257_76_11005));
   INV_X1 i_257_76_11025 (.A(n_257_76_11005), .ZN(n_257_76_11006));
   NAND2_X1 i_257_76_11026 (.A1(n_257_76_10843), .A2(n_257_76_10844), .ZN(
      n_257_76_11007));
   INV_X1 i_257_76_11027 (.A(n_257_76_11007), .ZN(n_257_76_11008));
   NOR2_X1 i_257_76_11028 (.A1(n_257_1078), .A2(n_257_76_17934), .ZN(
      n_257_76_11009));
   NAND3_X1 i_257_76_11029 (.A1(n_257_76_10852), .A2(n_257_76_10853), .A3(
      n_257_76_11009), .ZN(n_257_76_11010));
   INV_X1 i_257_76_11030 (.A(n_257_76_11010), .ZN(n_257_76_11011));
   NAND3_X1 i_257_76_11031 (.A1(n_257_76_11006), .A2(n_257_76_11008), .A3(
      n_257_76_11011), .ZN(n_257_76_11012));
   NAND3_X1 i_257_76_11032 (.A1(n_257_76_10858), .A2(n_257_76_10824), .A3(
      n_257_76_10860), .ZN(n_257_76_11013));
   NOR2_X1 i_257_76_11033 (.A1(n_257_76_11012), .A2(n_257_76_11013), .ZN(
      n_257_76_11014));
   NAND2_X1 i_257_76_11034 (.A1(n_257_76_10823), .A2(n_257_76_11014), .ZN(
      n_257_76_11015));
   INV_X1 i_257_76_11035 (.A(n_257_76_11015), .ZN(n_257_76_11016));
   NAND2_X1 i_257_76_11036 (.A1(n_257_76_10822), .A2(n_257_76_11016), .ZN(
      n_257_76_11017));
   INV_X1 i_257_76_11037 (.A(n_257_76_11017), .ZN(n_257_76_11018));
   NAND2_X1 i_257_76_11038 (.A1(n_257_76_18069), .A2(n_257_76_11018), .ZN(
      n_257_76_11019));
   NAND2_X1 i_257_76_11039 (.A1(n_257_616), .A2(n_257_442), .ZN(n_257_76_11020));
   INV_X1 i_257_76_11040 (.A(n_257_76_11020), .ZN(n_257_76_11021));
   NAND2_X1 i_257_76_11041 (.A1(n_257_432), .A2(n_257_76_11021), .ZN(
      n_257_76_11022));
   NOR2_X1 i_257_76_11042 (.A1(n_257_1078), .A2(n_257_76_11022), .ZN(
      n_257_76_11023));
   NAND4_X1 i_257_76_11043 (.A1(n_257_76_10852), .A2(n_257_76_10853), .A3(
      n_257_76_11023), .A4(n_257_76_10895), .ZN(n_257_76_11024));
   NOR2_X1 i_257_76_11044 (.A1(n_257_76_11024), .A2(n_257_76_10905), .ZN(
      n_257_76_11025));
   NAND2_X1 i_257_76_11045 (.A1(n_257_76_10908), .A2(n_257_76_10909), .ZN(
      n_257_76_11026));
   INV_X1 i_257_76_11046 (.A(n_257_76_11026), .ZN(n_257_76_11027));
   NAND3_X1 i_257_76_11047 (.A1(n_257_76_10847), .A2(n_257_76_10848), .A3(
      n_257_76_10843), .ZN(n_257_76_11028));
   INV_X1 i_257_76_11048 (.A(n_257_76_11028), .ZN(n_257_76_11029));
   NAND3_X1 i_257_76_11049 (.A1(n_257_76_11025), .A2(n_257_76_11027), .A3(
      n_257_76_11029), .ZN(n_257_76_11030));
   NOR2_X1 i_257_76_11050 (.A1(n_257_76_11030), .A2(n_257_76_10861), .ZN(
      n_257_76_11031));
   NAND3_X1 i_257_76_11051 (.A1(n_257_76_11031), .A2(n_257_76_10823), .A3(
      n_257_76_10863), .ZN(n_257_76_11032));
   INV_X1 i_257_76_11052 (.A(n_257_76_11032), .ZN(n_257_76_11033));
   NAND2_X1 i_257_76_11053 (.A1(n_257_76_10822), .A2(n_257_76_11033), .ZN(
      n_257_76_11034));
   INV_X1 i_257_76_11054 (.A(n_257_76_11034), .ZN(n_257_76_11035));
   NAND2_X1 i_257_76_11055 (.A1(n_257_68), .A2(n_257_76_11035), .ZN(
      n_257_76_11036));
   NAND3_X1 i_257_76_11056 (.A1(n_257_76_11004), .A2(n_257_76_11019), .A3(
      n_257_76_11036), .ZN(n_257_76_11037));
   NOR2_X1 i_257_76_11057 (.A1(n_257_1078), .A2(n_257_76_17951), .ZN(
      n_257_76_11038));
   NAND3_X1 i_257_76_11058 (.A1(n_257_76_10852), .A2(n_257_76_10853), .A3(
      n_257_76_11038), .ZN(n_257_76_11039));
   INV_X1 i_257_76_11059 (.A(n_257_76_11039), .ZN(n_257_76_11040));
   NAND4_X1 i_257_76_11060 (.A1(n_257_76_11040), .A2(n_257_816), .A3(
      n_257_76_10847), .A4(n_257_76_10844), .ZN(n_257_76_11041));
   NAND2_X1 i_257_76_11061 (.A1(n_257_76_10824), .A2(n_257_76_10860), .ZN(
      n_257_76_11042));
   NOR2_X1 i_257_76_11062 (.A1(n_257_76_11041), .A2(n_257_76_11042), .ZN(
      n_257_76_11043));
   NAND2_X1 i_257_76_11063 (.A1(n_257_76_10823), .A2(n_257_76_11043), .ZN(
      n_257_76_11044));
   INV_X1 i_257_76_11064 (.A(n_257_76_11044), .ZN(n_257_76_11045));
   NAND2_X1 i_257_76_11065 (.A1(n_257_76_10822), .A2(n_257_76_11045), .ZN(
      n_257_76_11046));
   INV_X1 i_257_76_11066 (.A(n_257_76_11046), .ZN(n_257_76_11047));
   NAND2_X1 i_257_76_11067 (.A1(n_257_22), .A2(n_257_76_11047), .ZN(
      n_257_76_11048));
   NAND2_X1 i_257_76_11068 (.A1(n_257_444), .A2(n_257_76_10837), .ZN(
      n_257_76_11049));
   INV_X1 i_257_76_11069 (.A(n_257_76_11049), .ZN(n_257_76_11050));
   NAND2_X1 i_257_76_11070 (.A1(n_257_1014), .A2(n_257_76_11050), .ZN(
      n_257_76_11051));
   INV_X1 i_257_76_11071 (.A(n_257_76_11051), .ZN(n_257_76_11052));
   NAND2_X1 i_257_76_11072 (.A1(n_257_76_10822), .A2(n_257_76_11052), .ZN(
      n_257_76_11053));
   INV_X1 i_257_76_11073 (.A(n_257_76_11053), .ZN(n_257_76_11054));
   NAND2_X1 i_257_76_11074 (.A1(n_257_76_18075), .A2(n_257_76_11054), .ZN(
      n_257_76_11055));
   NAND2_X1 i_257_76_11075 (.A1(n_257_76_11048), .A2(n_257_76_11055), .ZN(
      n_257_76_11056));
   NOR2_X1 i_257_76_11076 (.A1(n_257_76_11037), .A2(n_257_76_11056), .ZN(
      n_257_76_11057));
   NAND3_X1 i_257_76_11077 (.A1(n_257_76_10932), .A2(n_257_76_10987), .A3(
      n_257_76_11057), .ZN(n_257_76_11058));
   INV_X1 i_257_76_11078 (.A(n_257_76_11058), .ZN(n_257_76_11059));
   NAND3_X1 i_257_76_11079 (.A1(n_257_76_10853), .A2(n_257_54), .A3(
      n_257_76_10825), .ZN(n_257_76_11060));
   INV_X1 i_257_76_11080 (.A(n_257_76_11060), .ZN(n_257_76_11061));
   NAND2_X1 i_257_76_11081 (.A1(n_257_76_17760), .A2(n_257_76_17918), .ZN(
      n_257_76_11062));
   OAI21_X1 i_257_76_11082 (.A(n_257_76_11062), .B1(n_257_720), .B2(
      n_257_76_17633), .ZN(n_257_76_11063));
   NAND2_X1 i_257_76_11083 (.A1(n_257_76_10852), .A2(n_257_76_11063), .ZN(
      n_257_76_11064));
   INV_X1 i_257_76_11084 (.A(n_257_76_11064), .ZN(n_257_76_11065));
   NAND3_X1 i_257_76_11085 (.A1(n_257_76_11061), .A2(n_257_76_11065), .A3(
      n_257_76_10844), .ZN(n_257_76_11066));
   NOR2_X1 i_257_76_11086 (.A1(n_257_76_11066), .A2(n_257_76_11028), .ZN(
      n_257_76_11067));
   INV_X1 i_257_76_11087 (.A(n_257_76_10947), .ZN(n_257_76_11068));
   NAND3_X1 i_257_76_11088 (.A1(n_257_76_10860), .A2(n_257_76_10908), .A3(
      n_257_76_10909), .ZN(n_257_76_11069));
   INV_X1 i_257_76_11089 (.A(n_257_76_11069), .ZN(n_257_76_11070));
   NAND3_X1 i_257_76_11090 (.A1(n_257_76_11067), .A2(n_257_76_11068), .A3(
      n_257_76_11070), .ZN(n_257_76_11071));
   INV_X1 i_257_76_11091 (.A(n_257_76_11071), .ZN(n_257_76_11072));
   NAND3_X1 i_257_76_11092 (.A1(n_257_76_11072), .A2(n_257_76_10823), .A3(
      n_257_76_10863), .ZN(n_257_76_11073));
   INV_X1 i_257_76_11093 (.A(n_257_76_11073), .ZN(n_257_76_11074));
   NAND2_X1 i_257_76_11094 (.A1(n_257_76_10822), .A2(n_257_76_11074), .ZN(
      n_257_76_11075));
   INV_X1 i_257_76_11095 (.A(n_257_76_11075), .ZN(n_257_76_11076));
   NAND2_X1 i_257_76_11096 (.A1(n_257_76_18081), .A2(n_257_76_11076), .ZN(
      n_257_76_11077));
   NAND2_X1 i_257_76_11097 (.A1(n_257_76_17760), .A2(n_257_76_15658), .ZN(
      n_257_76_11078));
   OAI21_X1 i_257_76_11098 (.A(n_257_76_11078), .B1(n_257_720), .B2(
      n_257_76_15434), .ZN(n_257_76_11079));
   NAND3_X1 i_257_76_11099 (.A1(n_257_76_10844), .A2(n_257_76_11079), .A3(
      n_257_449), .ZN(n_257_76_11080));
   INV_X1 i_257_76_11100 (.A(n_257_76_11080), .ZN(n_257_76_11081));
   NAND3_X1 i_257_76_11101 (.A1(n_257_76_10852), .A2(n_257_76_10853), .A3(
      n_257_76_10825), .ZN(n_257_76_11082));
   INV_X1 i_257_76_11102 (.A(n_257_76_11082), .ZN(n_257_76_11083));
   NAND3_X1 i_257_76_11103 (.A1(n_257_76_10945), .A2(n_257_76_11081), .A3(
      n_257_76_11083), .ZN(n_257_76_11084));
   NOR2_X1 i_257_76_11104 (.A1(n_257_76_10861), .A2(n_257_76_11084), .ZN(
      n_257_76_11085));
   NAND3_X1 i_257_76_11105 (.A1(n_257_76_10823), .A2(n_257_76_11085), .A3(
      n_257_76_10863), .ZN(n_257_76_11086));
   INV_X1 i_257_76_11106 (.A(n_257_76_11086), .ZN(n_257_76_11087));
   NAND2_X1 i_257_76_11107 (.A1(n_257_76_10822), .A2(n_257_76_11087), .ZN(
      n_257_76_11088));
   INV_X1 i_257_76_11108 (.A(n_257_76_11088), .ZN(n_257_76_11089));
   NAND2_X1 i_257_76_11109 (.A1(n_257_76_18083), .A2(n_257_76_11089), .ZN(
      n_257_76_11090));
   NAND3_X1 i_257_76_11110 (.A1(n_257_76_10843), .A2(n_257_76_10904), .A3(
      n_257_76_10844), .ZN(n_257_76_11091));
   INV_X1 i_257_76_11111 (.A(n_257_76_11091), .ZN(n_257_76_11092));
   INV_X1 i_257_76_11112 (.A(n_257_616), .ZN(n_257_76_11093));
   NAND2_X1 i_257_76_11113 (.A1(n_257_76_11093), .A2(n_257_442), .ZN(
      n_257_76_11094));
   OAI21_X1 i_257_76_11114 (.A(n_257_76_11094), .B1(n_257_432), .B2(
      n_257_76_17412), .ZN(n_257_76_11095));
   NAND4_X1 i_257_76_11115 (.A1(n_257_76_10895), .A2(n_257_76_10825), .A3(
      n_257_76_11095), .A4(n_257_429), .ZN(n_257_76_11096));
   NOR2_X1 i_257_76_11116 (.A1(n_257_76_10900), .A2(n_257_76_11096), .ZN(
      n_257_76_11097));
   NAND3_X1 i_257_76_11117 (.A1(n_257_76_11092), .A2(n_257_76_10850), .A3(
      n_257_76_11097), .ZN(n_257_76_11098));
   NAND4_X1 i_257_76_11118 (.A1(n_257_76_10918), .A2(n_257_76_10860), .A3(
      n_257_76_10908), .A4(n_257_76_10909), .ZN(n_257_76_11099));
   NOR2_X1 i_257_76_11119 (.A1(n_257_76_11098), .A2(n_257_76_11099), .ZN(
      n_257_76_11100));
   NAND3_X1 i_257_76_11120 (.A1(n_257_76_11068), .A2(n_257_76_10912), .A3(
      n_257_171), .ZN(n_257_76_11101));
   INV_X1 i_257_76_11121 (.A(n_257_76_11101), .ZN(n_257_76_11102));
   NAND4_X1 i_257_76_11122 (.A1(n_257_76_10823), .A2(n_257_76_11100), .A3(
      n_257_76_10863), .A4(n_257_76_11102), .ZN(n_257_76_11103));
   INV_X1 i_257_76_11123 (.A(n_257_76_11103), .ZN(n_257_76_11104));
   NAND2_X1 i_257_76_11124 (.A1(n_257_76_10822), .A2(n_257_76_11104), .ZN(
      n_257_76_11105));
   INV_X1 i_257_76_11125 (.A(n_257_76_11105), .ZN(n_257_76_11106));
   NAND2_X1 i_257_76_11126 (.A1(n_257_76_18061), .A2(n_257_76_11106), .ZN(
      n_257_76_11107));
   NAND3_X1 i_257_76_11127 (.A1(n_257_76_11077), .A2(n_257_76_11090), .A3(
      n_257_76_11107), .ZN(n_257_76_11108));
   INV_X1 i_257_76_11128 (.A(n_257_76_11108), .ZN(n_257_76_11109));
   NAND2_X1 i_257_76_11129 (.A1(n_257_438), .A2(n_257_76_10825), .ZN(
      n_257_76_11110));
   INV_X1 i_257_76_11130 (.A(n_257_76_11110), .ZN(n_257_76_11111));
   NAND3_X1 i_257_76_11131 (.A1(n_257_76_11111), .A2(n_257_76_10852), .A3(
      n_257_76_14266), .ZN(n_257_76_11112));
   INV_X1 i_257_76_11132 (.A(n_257_76_11112), .ZN(n_257_76_11113));
   NAND3_X1 i_257_76_11133 (.A1(n_257_76_10824), .A2(n_257_76_10860), .A3(
      n_257_76_11113), .ZN(n_257_76_11114));
   INV_X1 i_257_76_11134 (.A(n_257_76_11114), .ZN(n_257_76_11115));
   NAND2_X1 i_257_76_11135 (.A1(n_257_76_10823), .A2(n_257_76_11115), .ZN(
      n_257_76_11116));
   INV_X1 i_257_76_11136 (.A(n_257_76_11116), .ZN(n_257_76_11117));
   NAND2_X1 i_257_76_11137 (.A1(n_257_76_10822), .A2(n_257_76_11117), .ZN(
      n_257_76_11118));
   INV_X1 i_257_76_11138 (.A(n_257_76_11118), .ZN(n_257_76_11119));
   NAND2_X1 i_257_76_11139 (.A1(n_257_76_18067), .A2(n_257_76_11119), .ZN(
      n_257_76_11120));
   NAND2_X1 i_257_76_11140 (.A1(n_257_76_10858), .A2(n_257_76_10859), .ZN(
      n_257_76_11121));
   INV_X1 i_257_76_11141 (.A(n_257_76_10916), .ZN(n_257_76_11122));
   NOR2_X1 i_257_76_11142 (.A1(n_257_76_11121), .A2(n_257_76_11122), .ZN(
      n_257_76_11123));
   NAND2_X1 i_257_76_11143 (.A1(n_257_76_10824), .A2(n_257_76_10918), .ZN(
      n_257_76_11124));
   NAND2_X1 i_257_76_11144 (.A1(n_257_76_10860), .A2(n_257_76_10908), .ZN(
      n_257_76_11125));
   NOR2_X1 i_257_76_11145 (.A1(n_257_76_11124), .A2(n_257_76_11125), .ZN(
      n_257_76_11126));
   NAND2_X1 i_257_76_11146 (.A1(n_257_76_11123), .A2(n_257_76_11126), .ZN(
      n_257_76_11127));
   INV_X1 i_257_76_11147 (.A(n_257_76_11127), .ZN(n_257_76_11128));
   NAND2_X1 i_257_76_11148 (.A1(n_257_442), .A2(n_257_488), .ZN(n_257_76_11129));
   NAND2_X1 i_257_76_11149 (.A1(n_257_76_10825), .A2(n_257_76_18021), .ZN(
      n_257_76_11130));
   NAND2_X1 i_257_76_11150 (.A1(n_257_76_10896), .A2(n_257_420), .ZN(
      n_257_76_11131));
   NOR2_X1 i_257_76_11151 (.A1(n_257_76_11130), .A2(n_257_76_11131), .ZN(
      n_257_76_11132));
   NAND2_X1 i_257_76_11152 (.A1(n_257_76_10993), .A2(n_257_76_11132), .ZN(
      n_257_76_11133));
   NOR2_X1 i_257_76_11153 (.A1(n_257_76_11133), .A2(n_257_76_10900), .ZN(
      n_257_76_11134));
   INV_X1 i_257_76_11154 (.A(n_257_76_10843), .ZN(n_257_76_11135));
   NOR2_X1 i_257_76_11155 (.A1(n_257_76_10905), .A2(n_257_76_11135), .ZN(
      n_257_76_11136));
   NAND2_X1 i_257_76_11156 (.A1(n_257_76_11134), .A2(n_257_76_11136), .ZN(
      n_257_76_11137));
   NAND2_X1 i_257_76_11157 (.A1(n_257_329), .A2(n_257_422), .ZN(n_257_76_11138));
   NAND2_X1 i_257_76_11158 (.A1(n_257_76_10909), .A2(n_257_76_11138), .ZN(
      n_257_76_11139));
   INV_X1 i_257_76_11159 (.A(n_257_76_11139), .ZN(n_257_76_11140));
   NAND2_X1 i_257_76_11160 (.A1(n_257_76_11140), .A2(n_257_76_10850), .ZN(
      n_257_76_11141));
   NOR2_X1 i_257_76_11161 (.A1(n_257_76_11137), .A2(n_257_76_11141), .ZN(
      n_257_76_11142));
   NAND2_X1 i_257_76_11162 (.A1(n_257_76_11128), .A2(n_257_76_11142), .ZN(
      n_257_76_11143));
   NAND2_X1 i_257_76_11163 (.A1(n_257_368), .A2(n_257_421), .ZN(n_257_76_11144));
   NAND2_X1 i_257_76_11164 (.A1(n_257_76_10923), .A2(n_257_76_11144), .ZN(
      n_257_76_11145));
   INV_X1 i_257_76_11165 (.A(n_257_76_11145), .ZN(n_257_76_11146));
   INV_X1 i_257_76_11166 (.A(n_257_76_10912), .ZN(n_257_76_11147));
   NAND2_X1 i_257_76_11167 (.A1(n_257_291), .A2(n_257_423), .ZN(n_257_76_11148));
   NAND2_X1 i_257_76_11168 (.A1(n_257_76_10913), .A2(n_257_76_11148), .ZN(
      n_257_76_11149));
   NOR2_X1 i_257_76_11169 (.A1(n_257_76_11147), .A2(n_257_76_11149), .ZN(
      n_257_76_11150));
   NAND2_X1 i_257_76_11170 (.A1(n_257_76_11146), .A2(n_257_76_11150), .ZN(
      n_257_76_11151));
   NOR2_X1 i_257_76_11171 (.A1(n_257_76_11143), .A2(n_257_76_11151), .ZN(
      n_257_76_11152));
   INV_X1 i_257_76_11172 (.A(n_257_76_10823), .ZN(n_257_76_11153));
   NAND2_X1 i_257_76_11173 (.A1(n_257_76_10863), .A2(n_257_76_10922), .ZN(
      n_257_76_11154));
   NOR2_X1 i_257_76_11174 (.A1(n_257_76_11153), .A2(n_257_76_11154), .ZN(
      n_257_76_11155));
   NAND2_X1 i_257_76_11175 (.A1(n_257_76_11152), .A2(n_257_76_11155), .ZN(
      n_257_76_11156));
   INV_X1 i_257_76_11176 (.A(n_257_76_10822), .ZN(n_257_76_11157));
   NOR2_X1 i_257_76_11177 (.A1(n_257_76_11156), .A2(n_257_76_11157), .ZN(
      n_257_76_11158));
   NAND2_X1 i_257_76_11178 (.A1(n_257_76_18073), .A2(n_257_76_11158), .ZN(
      n_257_76_11159));
   NAND4_X1 i_257_76_11179 (.A1(n_257_76_10895), .A2(n_257_76_10825), .A3(
      n_257_76_11095), .A4(n_257_430), .ZN(n_257_76_11160));
   NOR2_X1 i_257_76_11180 (.A1(n_257_76_10900), .A2(n_257_76_11160), .ZN(
      n_257_76_11161));
   NAND3_X1 i_257_76_11181 (.A1(n_257_76_11161), .A2(n_257_76_10906), .A3(
      n_257_132), .ZN(n_257_76_11162));
   NOR2_X1 i_257_76_11182 (.A1(n_257_76_11162), .A2(n_257_76_10956), .ZN(
      n_257_76_11163));
   NAND3_X1 i_257_76_11183 (.A1(n_257_76_10824), .A2(n_257_76_10860), .A3(
      n_257_76_10908), .ZN(n_257_76_11164));
   INV_X1 i_257_76_11184 (.A(n_257_76_11164), .ZN(n_257_76_11165));
   INV_X1 i_257_76_11185 (.A(n_257_76_11121), .ZN(n_257_76_11166));
   NAND3_X1 i_257_76_11186 (.A1(n_257_76_11165), .A2(n_257_76_10912), .A3(
      n_257_76_11166), .ZN(n_257_76_11167));
   INV_X1 i_257_76_11187 (.A(n_257_76_11167), .ZN(n_257_76_11168));
   NAND4_X1 i_257_76_11188 (.A1(n_257_76_10823), .A2(n_257_76_11163), .A3(
      n_257_76_11168), .A4(n_257_76_10863), .ZN(n_257_76_11169));
   INV_X1 i_257_76_11189 (.A(n_257_76_11169), .ZN(n_257_76_11170));
   NAND2_X1 i_257_76_11190 (.A1(n_257_76_10822), .A2(n_257_76_11170), .ZN(
      n_257_76_11171));
   INV_X1 i_257_76_11191 (.A(n_257_76_11171), .ZN(n_257_76_11172));
   NAND2_X1 i_257_76_11192 (.A1(n_257_76_18068), .A2(n_257_76_11172), .ZN(
      n_257_76_11173));
   NAND3_X1 i_257_76_11193 (.A1(n_257_76_11120), .A2(n_257_76_11159), .A3(
      n_257_76_11173), .ZN(n_257_76_11174));
   INV_X1 i_257_76_11194 (.A(n_257_76_11174), .ZN(n_257_76_11175));
   NAND2_X1 i_257_76_11195 (.A1(n_257_447), .A2(n_257_76_10852), .ZN(
      n_257_76_11176));
   INV_X1 i_257_76_11196 (.A(n_257_76_11176), .ZN(n_257_76_11177));
   NAND2_X1 i_257_76_11197 (.A1(n_257_784), .A2(n_257_442), .ZN(n_257_76_11178));
   NOR2_X1 i_257_76_11198 (.A1(n_257_1078), .A2(n_257_76_11178), .ZN(
      n_257_76_11179));
   NAND2_X1 i_257_76_11199 (.A1(n_257_76_10853), .A2(n_257_76_11179), .ZN(
      n_257_76_11180));
   INV_X1 i_257_76_11200 (.A(n_257_76_11180), .ZN(n_257_76_11181));
   NAND4_X1 i_257_76_11201 (.A1(n_257_76_11177), .A2(n_257_76_11181), .A3(
      n_257_76_10847), .A4(n_257_76_10844), .ZN(n_257_76_11182));
   NOR2_X1 i_257_76_11202 (.A1(n_257_76_11013), .A2(n_257_76_11182), .ZN(
      n_257_76_11183));
   NAND2_X1 i_257_76_11203 (.A1(n_257_76_10823), .A2(n_257_76_11183), .ZN(
      n_257_76_11184));
   INV_X1 i_257_76_11204 (.A(n_257_76_11184), .ZN(n_257_76_11185));
   NAND2_X1 i_257_76_11205 (.A1(n_257_76_10822), .A2(n_257_76_11185), .ZN(
      n_257_76_11186));
   INV_X1 i_257_76_11206 (.A(n_257_76_11186), .ZN(n_257_76_11187));
   NAND3_X1 i_257_76_11207 (.A1(n_257_76_10908), .A2(n_257_76_10909), .A3(
      n_257_76_10847), .ZN(n_257_76_11188));
   NAND4_X1 i_257_76_11208 (.A1(n_257_76_10895), .A2(n_257_76_10825), .A3(
      n_257_76_11095), .A4(n_257_431), .ZN(n_257_76_11189));
   INV_X1 i_257_76_11209 (.A(n_257_76_11189), .ZN(n_257_76_11190));
   NAND3_X1 i_257_76_11210 (.A1(n_257_76_10957), .A2(n_257_76_11190), .A3(
      n_257_76_10844), .ZN(n_257_76_11191));
   NAND3_X1 i_257_76_11211 (.A1(n_257_76_10848), .A2(n_257_76_10843), .A3(
      n_257_76_10904), .ZN(n_257_76_11192));
   NOR3_X1 i_257_76_11212 (.A1(n_257_76_11188), .A2(n_257_76_11191), .A3(
      n_257_76_11192), .ZN(n_257_76_11193));
   NAND2_X1 i_257_76_11213 (.A1(n_257_94), .A2(n_257_76_10858), .ZN(
      n_257_76_11194));
   NAND3_X1 i_257_76_11214 (.A1(n_257_76_10859), .A2(n_257_76_10824), .A3(
      n_257_76_10860), .ZN(n_257_76_11195));
   NOR2_X1 i_257_76_11215 (.A1(n_257_76_11194), .A2(n_257_76_11195), .ZN(
      n_257_76_11196));
   NAND3_X1 i_257_76_11216 (.A1(n_257_76_11193), .A2(n_257_76_10863), .A3(
      n_257_76_11196), .ZN(n_257_76_11197));
   NOR2_X1 i_257_76_11217 (.A1(n_257_76_11197), .A2(n_257_76_11153), .ZN(
      n_257_76_11198));
   NAND2_X1 i_257_76_11218 (.A1(n_257_76_10822), .A2(n_257_76_11198), .ZN(
      n_257_76_11199));
   INV_X1 i_257_76_11219 (.A(n_257_76_11199), .ZN(n_257_76_11200));
   AOI22_X1 i_257_76_11220 (.A1(n_257_76_18085), .A2(n_257_76_11187), .B1(
      n_257_76_18080), .B2(n_257_76_11200), .ZN(n_257_76_11201));
   NAND3_X1 i_257_76_11221 (.A1(n_257_76_11109), .A2(n_257_76_11175), .A3(
      n_257_76_11201), .ZN(n_257_76_11202));
   NAND4_X1 i_257_76_11222 (.A1(n_257_76_10844), .A2(n_257_76_10852), .A3(
      n_257_76_10853), .A4(n_257_448), .ZN(n_257_76_11203));
   NOR2_X1 i_257_76_11223 (.A1(n_257_76_11203), .A2(n_257_76_10944), .ZN(
      n_257_76_11204));
   NAND2_X1 i_257_76_11224 (.A1(n_257_76_10851), .A2(n_257_76_10825), .ZN(
      n_257_76_11205));
   INV_X1 i_257_76_11225 (.A(n_257_76_11205), .ZN(n_257_76_11206));
   NAND3_X1 i_257_76_11226 (.A1(n_257_76_10824), .A2(n_257_76_10860), .A3(
      n_257_76_11206), .ZN(n_257_76_11207));
   INV_X1 i_257_76_11227 (.A(n_257_76_11207), .ZN(n_257_76_11208));
   NAND4_X1 i_257_76_11228 (.A1(n_257_688), .A2(n_257_76_11204), .A3(
      n_257_76_11166), .A4(n_257_76_11208), .ZN(n_257_76_11209));
   NOR2_X1 i_257_76_11229 (.A1(n_257_76_11153), .A2(n_257_76_11209), .ZN(
      n_257_76_11210));
   NAND2_X1 i_257_76_11230 (.A1(n_257_76_10822), .A2(n_257_76_11210), .ZN(
      n_257_76_11211));
   INV_X1 i_257_76_11231 (.A(n_257_76_11211), .ZN(n_257_76_11212));
   NAND2_X1 i_257_76_11232 (.A1(n_257_76_18079), .A2(n_257_76_11212), .ZN(
      n_257_76_11213));
   NAND3_X1 i_257_76_11233 (.A1(n_257_76_18020), .A2(n_257_76_10896), .A3(
      n_257_425), .ZN(n_257_76_11214));
   NOR2_X1 i_257_76_11234 (.A1(n_257_76_11214), .A2(n_257_1078), .ZN(
      n_257_76_11215));
   NAND4_X1 i_257_76_11235 (.A1(n_257_76_11215), .A2(n_257_76_10993), .A3(
      n_257_76_10852), .A4(n_257_76_10853), .ZN(n_257_76_11216));
   NOR2_X1 i_257_76_11236 (.A1(n_257_76_11216), .A2(n_257_76_11091), .ZN(
      n_257_76_11217));
   INV_X1 i_257_76_11237 (.A(n_257_76_10919), .ZN(n_257_76_11218));
   NAND4_X1 i_257_76_11238 (.A1(n_257_76_10908), .A2(n_257_76_10909), .A3(
      n_257_76_10847), .A4(n_257_76_10848), .ZN(n_257_76_11219));
   INV_X1 i_257_76_11239 (.A(n_257_76_11219), .ZN(n_257_76_11220));
   NAND3_X1 i_257_76_11240 (.A1(n_257_76_11217), .A2(n_257_76_11218), .A3(
      n_257_76_11220), .ZN(n_257_76_11221));
   INV_X1 i_257_76_11241 (.A(n_257_76_11221), .ZN(n_257_76_11222));
   NAND4_X1 i_257_76_11242 (.A1(n_257_76_10912), .A2(n_257_76_11166), .A3(
      n_257_251), .A4(n_257_76_10913), .ZN(n_257_76_11223));
   INV_X1 i_257_76_11243 (.A(n_257_76_11223), .ZN(n_257_76_11224));
   NAND4_X1 i_257_76_11244 (.A1(n_257_76_11222), .A2(n_257_76_11224), .A3(
      n_257_76_10863), .A4(n_257_76_10922), .ZN(n_257_76_11225));
   INV_X1 i_257_76_11245 (.A(n_257_76_11225), .ZN(n_257_76_11226));
   NAND2_X1 i_257_76_11246 (.A1(n_257_76_11226), .A2(n_257_76_10823), .ZN(
      n_257_76_11227));
   NOR2_X1 i_257_76_11247 (.A1(n_257_76_11227), .A2(n_257_76_11157), .ZN(
      n_257_76_11228));
   NAND2_X1 i_257_76_11248 (.A1(n_257_76_18064), .A2(n_257_76_11228), .ZN(
      n_257_76_11229));
   NAND2_X1 i_257_76_11249 (.A1(n_257_76_10896), .A2(n_257_421), .ZN(
      n_257_76_11230));
   INV_X1 i_257_76_11250 (.A(n_257_76_11230), .ZN(n_257_76_11231));
   NAND4_X1 i_257_76_11251 (.A1(n_257_76_10893), .A2(n_257_76_10894), .A3(
      n_257_76_10895), .A4(n_257_76_11231), .ZN(n_257_76_11232));
   NOR2_X1 i_257_76_11252 (.A1(n_257_76_11232), .A2(n_257_76_10900), .ZN(
      n_257_76_11233));
   NAND3_X1 i_257_76_11253 (.A1(n_257_76_11233), .A2(n_257_76_11092), .A3(
      n_257_76_10850), .ZN(n_257_76_11234));
   NAND4_X1 i_257_76_11254 (.A1(n_257_76_10860), .A2(n_257_76_10908), .A3(
      n_257_76_10909), .A4(n_257_76_11138), .ZN(n_257_76_11235));
   NOR2_X1 i_257_76_11255 (.A1(n_257_76_11234), .A2(n_257_76_11235), .ZN(
      n_257_76_11236));
   NAND2_X1 i_257_76_11256 (.A1(n_257_76_10913), .A2(n_257_368), .ZN(
      n_257_76_11237));
   NOR2_X1 i_257_76_11257 (.A1(n_257_76_11147), .A2(n_257_76_11237), .ZN(
      n_257_76_11238));
   NAND3_X1 i_257_76_11258 (.A1(n_257_76_11148), .A2(n_257_76_10916), .A3(
      n_257_76_10858), .ZN(n_257_76_11239));
   NAND3_X1 i_257_76_11259 (.A1(n_257_76_10859), .A2(n_257_76_10824), .A3(
      n_257_76_10918), .ZN(n_257_76_11240));
   NOR2_X1 i_257_76_11260 (.A1(n_257_76_11239), .A2(n_257_76_11240), .ZN(
      n_257_76_11241));
   NAND3_X1 i_257_76_11261 (.A1(n_257_76_11236), .A2(n_257_76_11238), .A3(
      n_257_76_11241), .ZN(n_257_76_11242));
   NOR2_X1 i_257_76_11262 (.A1(n_257_76_11242), .A2(n_257_76_10926), .ZN(
      n_257_76_11243));
   NAND2_X1 i_257_76_11263 (.A1(n_257_76_10822), .A2(n_257_76_11243), .ZN(
      n_257_76_11244));
   INV_X1 i_257_76_11264 (.A(n_257_76_11244), .ZN(n_257_76_11245));
   NAND2_X1 i_257_76_11265 (.A1(n_257_76_18082), .A2(n_257_76_11245), .ZN(
      n_257_76_11246));
   NAND3_X1 i_257_76_11266 (.A1(n_257_76_11213), .A2(n_257_76_11229), .A3(
      n_257_76_11246), .ZN(n_257_76_11247));
   INV_X1 i_257_76_11267 (.A(n_257_76_11247), .ZN(n_257_76_11248));
   INV_X1 i_257_76_11268 (.A(n_257_76_10895), .ZN(n_257_76_11249));
   NAND2_X1 i_257_76_11269 (.A1(n_257_76_18020), .A2(n_257_76_10896), .ZN(
      n_257_76_11250));
   NOR2_X1 i_257_76_11270 (.A1(n_257_76_11249), .A2(n_257_76_11250), .ZN(
      n_257_76_11251));
   NAND3_X1 i_257_76_11271 (.A1(n_257_76_10825), .A2(n_257_211), .A3(n_257_427), 
      .ZN(n_257_76_11252));
   INV_X1 i_257_76_11272 (.A(n_257_76_11252), .ZN(n_257_76_11253));
   NAND3_X1 i_257_76_11273 (.A1(n_257_76_11251), .A2(n_257_76_10904), .A3(
      n_257_76_11253), .ZN(n_257_76_11254));
   INV_X1 i_257_76_11274 (.A(n_257_76_11254), .ZN(n_257_76_11255));
   NAND2_X1 i_257_76_11275 (.A1(n_257_76_10912), .A2(n_257_76_11255), .ZN(
      n_257_76_11256));
   INV_X1 i_257_76_11276 (.A(n_257_76_11256), .ZN(n_257_76_11257));
   NAND4_X1 i_257_76_11277 (.A1(n_257_76_10957), .A2(n_257_76_10848), .A3(
      n_257_76_10843), .A4(n_257_76_10844), .ZN(n_257_76_11258));
   NAND2_X1 i_257_76_11278 (.A1(n_257_76_10909), .A2(n_257_76_10847), .ZN(
      n_257_76_11259));
   NOR2_X1 i_257_76_11279 (.A1(n_257_76_11258), .A2(n_257_76_11259), .ZN(
      n_257_76_11260));
   NAND4_X1 i_257_76_11280 (.A1(n_257_76_10955), .A2(n_257_76_11257), .A3(
      n_257_76_10922), .A4(n_257_76_11260), .ZN(n_257_76_11261));
   NOR2_X1 i_257_76_11281 (.A1(n_257_76_11261), .A2(n_257_76_10967), .ZN(
      n_257_76_11262));
   NAND2_X1 i_257_76_11282 (.A1(n_257_76_10822), .A2(n_257_76_11262), .ZN(
      n_257_76_11263));
   INV_X1 i_257_76_11283 (.A(n_257_76_11263), .ZN(n_257_76_11264));
   NAND2_X1 i_257_76_11284 (.A1(n_257_76_18065), .A2(n_257_76_11264), .ZN(
      n_257_76_11265));
   NAND3_X1 i_257_76_11285 (.A1(n_257_471), .A2(n_257_76_10852), .A3(
      n_257_76_10853), .ZN(n_257_76_11266));
   NAND2_X1 i_257_76_11286 (.A1(n_257_451), .A2(n_257_76_10844), .ZN(
      n_257_76_11267));
   NOR2_X1 i_257_76_11287 (.A1(n_257_76_11266), .A2(n_257_76_11267), .ZN(
      n_257_76_11268));
   NAND2_X1 i_257_76_11288 (.A1(n_257_76_10909), .A2(n_257_76_11206), .ZN(
      n_257_76_11269));
   INV_X1 i_257_76_11289 (.A(n_257_76_11269), .ZN(n_257_76_11270));
   NAND3_X1 i_257_76_11290 (.A1(n_257_76_11268), .A2(n_257_76_11270), .A3(
      n_257_76_11029), .ZN(n_257_76_11271));
   NOR2_X1 i_257_76_11291 (.A1(n_257_76_11271), .A2(n_257_76_10861), .ZN(
      n_257_76_11272));
   NAND3_X1 i_257_76_11292 (.A1(n_257_76_11272), .A2(n_257_76_10823), .A3(
      n_257_76_10863), .ZN(n_257_76_11273));
   INV_X1 i_257_76_11293 (.A(n_257_76_11273), .ZN(n_257_76_11274));
   NAND2_X1 i_257_76_11294 (.A1(n_257_76_10822), .A2(n_257_76_11274), .ZN(
      n_257_76_11275));
   INV_X1 i_257_76_11295 (.A(n_257_76_11275), .ZN(n_257_76_11276));
   NAND2_X1 i_257_76_11296 (.A1(n_257_76_18063), .A2(n_257_76_11276), .ZN(
      n_257_76_11277));
   NAND2_X1 i_257_76_11297 (.A1(n_257_76_10923), .A2(n_257_76_10912), .ZN(
      n_257_76_11278));
   INV_X1 i_257_76_11298 (.A(n_257_76_11278), .ZN(n_257_76_11279));
   NAND2_X1 i_257_76_11299 (.A1(n_257_76_10824), .A2(n_257_76_10908), .ZN(
      n_257_76_11280));
   INV_X1 i_257_76_11300 (.A(n_257_76_11280), .ZN(n_257_76_11281));
   NAND3_X1 i_257_76_11301 (.A1(n_257_76_11281), .A2(n_257_76_10913), .A3(
      n_257_76_11029), .ZN(n_257_76_11282));
   INV_X1 i_257_76_11302 (.A(n_257_76_11282), .ZN(n_257_76_11283));
   NAND4_X1 i_257_76_11303 (.A1(n_257_76_11279), .A2(n_257_76_10863), .A3(
      n_257_76_11283), .A4(n_257_76_10922), .ZN(n_257_76_11284));
   INV_X1 i_257_76_11304 (.A(n_257_76_11284), .ZN(n_257_76_11285));
   NAND3_X1 i_257_76_11305 (.A1(n_257_76_18020), .A2(n_257_76_10896), .A3(
      n_257_424), .ZN(n_257_76_11286));
   NOR2_X1 i_257_76_11306 (.A1(n_257_76_11286), .A2(n_257_1078), .ZN(
      n_257_76_11287));
   NAND4_X1 i_257_76_11307 (.A1(n_257_76_11287), .A2(n_257_76_10993), .A3(
      n_257_76_10852), .A4(n_257_76_10853), .ZN(n_257_76_11288));
   NAND3_X1 i_257_76_11308 (.A1(n_257_520), .A2(n_257_76_10904), .A3(
      n_257_76_10844), .ZN(n_257_76_11289));
   NOR2_X1 i_257_76_11309 (.A1(n_257_76_11288), .A2(n_257_76_11289), .ZN(
      n_257_76_11290));
   NAND3_X1 i_257_76_11310 (.A1(n_257_76_10918), .A2(n_257_76_10860), .A3(
      n_257_76_10909), .ZN(n_257_76_11291));
   INV_X1 i_257_76_11311 (.A(n_257_76_11291), .ZN(n_257_76_11292));
   NAND3_X1 i_257_76_11312 (.A1(n_257_76_11290), .A2(n_257_76_11292), .A3(
      n_257_76_11166), .ZN(n_257_76_11293));
   NOR2_X1 i_257_76_11313 (.A1(n_257_76_11153), .A2(n_257_76_11293), .ZN(
      n_257_76_11294));
   NAND2_X1 i_257_76_11314 (.A1(n_257_76_11285), .A2(n_257_76_11294), .ZN(
      n_257_76_11295));
   NOR2_X1 i_257_76_11315 (.A1(n_257_76_11157), .A2(n_257_76_11295), .ZN(
      n_257_76_11296));
   NAND2_X1 i_257_76_11316 (.A1(n_257_76_18062), .A2(n_257_76_11296), .ZN(
      n_257_76_11297));
   NAND3_X1 i_257_76_11317 (.A1(n_257_76_11265), .A2(n_257_76_11277), .A3(
      n_257_76_11297), .ZN(n_257_76_11298));
   INV_X1 i_257_76_11318 (.A(n_257_76_11298), .ZN(n_257_76_11299));
   NAND4_X1 i_257_76_11319 (.A1(n_257_76_10903), .A2(n_257_76_10824), .A3(
      n_257_76_10908), .A4(n_257_76_10847), .ZN(n_257_76_11300));
   NOR2_X1 i_257_76_11320 (.A1(n_257_76_11300), .A2(n_257_76_11149), .ZN(
      n_257_76_11301));
   NAND4_X1 i_257_76_11321 (.A1(n_257_76_11301), .A2(n_257_76_11279), .A3(
      n_257_76_10863), .A4(n_257_76_10922), .ZN(n_257_76_11302));
   NAND4_X1 i_257_76_11322 (.A1(n_257_76_10904), .A2(n_257_76_10844), .A3(
      n_257_329), .A4(n_257_76_10852), .ZN(n_257_76_11303));
   INV_X1 i_257_76_11323 (.A(n_257_76_11250), .ZN(n_257_76_11304));
   NAND2_X1 i_257_76_11324 (.A1(n_257_76_10894), .A2(n_257_76_11304), .ZN(
      n_257_76_11305));
   INV_X1 i_257_76_11325 (.A(n_257_76_11305), .ZN(n_257_76_11306));
   NAND3_X1 i_257_76_11326 (.A1(n_257_76_10895), .A2(n_257_76_10825), .A3(
      n_257_422), .ZN(n_257_76_11307));
   INV_X1 i_257_76_11327 (.A(n_257_76_11307), .ZN(n_257_76_11308));
   NAND3_X1 i_257_76_11328 (.A1(n_257_76_11306), .A2(n_257_76_11308), .A3(
      n_257_76_10853), .ZN(n_257_76_11309));
   NOR2_X1 i_257_76_11329 (.A1(n_257_76_11303), .A2(n_257_76_11309), .ZN(
      n_257_76_11310));
   INV_X1 i_257_76_11330 (.A(n_257_76_10917), .ZN(n_257_76_11311));
   NAND3_X1 i_257_76_11331 (.A1(n_257_76_11310), .A2(n_257_76_11311), .A3(
      n_257_76_11292), .ZN(n_257_76_11312));
   INV_X1 i_257_76_11332 (.A(n_257_76_11312), .ZN(n_257_76_11313));
   NAND2_X1 i_257_76_11333 (.A1(n_257_76_10823), .A2(n_257_76_11313), .ZN(
      n_257_76_11314));
   NOR2_X1 i_257_76_11334 (.A1(n_257_76_11302), .A2(n_257_76_11314), .ZN(
      n_257_76_11315));
   NAND2_X1 i_257_76_11335 (.A1(n_257_76_10822), .A2(n_257_76_11315), .ZN(
      n_257_76_11316));
   INV_X1 i_257_76_11336 (.A(n_257_76_11316), .ZN(n_257_76_11317));
   NAND2_X1 i_257_76_11337 (.A1(n_257_342), .A2(n_257_76_11317), .ZN(
      n_257_76_11318));
   NAND4_X1 i_257_76_11338 (.A1(n_257_76_10824), .A2(n_257_76_10918), .A3(
      n_257_76_10860), .A4(n_257_76_10908), .ZN(n_257_76_11319));
   NOR2_X1 i_257_76_11339 (.A1(n_257_76_11319), .A2(n_257_76_10917), .ZN(
      n_257_76_11320));
   NAND4_X1 i_257_76_11340 (.A1(n_257_76_11146), .A2(n_257_76_11150), .A3(
      n_257_76_11320), .A4(n_257_76_10922), .ZN(n_257_76_11321));
   NAND3_X1 i_257_76_11341 (.A1(n_257_76_10852), .A2(n_257_76_10853), .A3(
      n_257_76_10894), .ZN(n_257_76_11322));
   NAND2_X1 i_257_76_11342 (.A1(n_257_584), .A2(n_257_428), .ZN(n_257_76_11323));
   NAND3_X1 i_257_76_11343 (.A1(n_257_484), .A2(n_257_407), .A3(n_257_442), 
      .ZN(n_257_76_11324));
   INV_X1 i_257_76_11344 (.A(n_257_76_11324), .ZN(n_257_76_11325));
   NAND3_X1 i_257_76_11345 (.A1(n_257_76_10896), .A2(n_257_76_11323), .A3(
      n_257_76_11325), .ZN(n_257_76_11326));
   INV_X1 i_257_76_11346 (.A(n_257_76_11326), .ZN(n_257_76_11327));
   NAND2_X1 i_257_76_11347 (.A1(n_257_420), .A2(n_257_488), .ZN(n_257_76_11328));
   NAND4_X1 i_257_76_11348 (.A1(n_257_76_11327), .A2(n_257_76_10895), .A3(
      n_257_76_10825), .A4(n_257_76_11328), .ZN(n_257_76_11329));
   NOR2_X1 i_257_76_11349 (.A1(n_257_76_11322), .A2(n_257_76_11329), .ZN(
      n_257_76_11330));
   NAND2_X1 i_257_76_11350 (.A1(n_257_76_11092), .A2(n_257_76_11330), .ZN(
      n_257_76_11331));
   NAND4_X1 i_257_76_11351 (.A1(n_257_76_10909), .A2(n_257_76_11138), .A3(
      n_257_76_10847), .A4(n_257_76_10848), .ZN(n_257_76_11332));
   NOR2_X1 i_257_76_11352 (.A1(n_257_76_11331), .A2(n_257_76_11332), .ZN(
      n_257_76_11333));
   NAND3_X1 i_257_76_11353 (.A1(n_257_76_10823), .A2(n_257_76_11333), .A3(
      n_257_76_10863), .ZN(n_257_76_11334));
   NOR2_X1 i_257_76_11354 (.A1(n_257_76_11321), .A2(n_257_76_11334), .ZN(
      n_257_76_11335));
   NAND2_X1 i_257_76_11355 (.A1(n_257_76_10822), .A2(n_257_76_11335), .ZN(
      n_257_76_11336));
   INV_X1 i_257_76_11356 (.A(n_257_76_11336), .ZN(n_257_76_11337));
   NAND2_X1 i_257_76_11357 (.A1(n_257_76_18060), .A2(n_257_76_11337), .ZN(
      n_257_76_11338));
   NAND2_X1 i_257_76_11358 (.A1(n_257_171), .A2(n_257_76_17331), .ZN(
      n_257_76_11339));
   AOI21_X1 i_257_76_11359 (.A(n_257_76_11255), .B1(n_257_94), .B2(
      n_257_76_17932), .ZN(n_257_76_11340));
   NAND2_X1 i_257_76_11360 (.A1(n_257_76_11339), .A2(n_257_76_11340), .ZN(
      n_257_76_11341));
   INV_X1 i_257_76_11361 (.A(n_257_76_11341), .ZN(n_257_76_11342));
   INV_X1 i_257_76_11362 (.A(n_257_76_11178), .ZN(n_257_76_11343));
   NAND2_X1 i_257_76_11363 (.A1(n_257_447), .A2(n_257_76_11343), .ZN(
      n_257_76_11344));
   NAND2_X1 i_257_76_11364 (.A1(n_257_880), .A2(n_257_76_17903), .ZN(
      n_257_76_11345));
   NAND2_X1 i_257_76_11365 (.A1(n_257_76_14266), .A2(n_257_438), .ZN(
      n_257_76_11346));
   NAND2_X1 i_257_76_11366 (.A1(n_257_440), .A2(n_257_76_10827), .ZN(
      n_257_76_11347));
   NAND4_X1 i_257_76_11367 (.A1(n_257_76_11344), .A2(n_257_76_11345), .A3(
      n_257_76_11346), .A4(n_257_76_11347), .ZN(n_257_76_11348));
   INV_X1 i_257_76_11368 (.A(n_257_76_10872), .ZN(n_257_76_11349));
   NAND2_X1 i_257_76_11369 (.A1(n_257_446), .A2(n_257_76_11349), .ZN(
      n_257_76_11350));
   NAND2_X1 i_257_76_11370 (.A1(n_257_54), .A2(n_257_76_11063), .ZN(
      n_257_76_11351));
   NAND2_X1 i_257_76_11371 (.A1(n_257_449), .A2(n_257_76_15658), .ZN(
      n_257_76_11352));
   NAND3_X1 i_257_76_11372 (.A1(n_257_76_11350), .A2(n_257_76_11351), .A3(
      n_257_76_11352), .ZN(n_257_76_11353));
   NOR2_X1 i_257_76_11373 (.A1(n_257_76_11348), .A2(n_257_76_11353), .ZN(
      n_257_76_11354));
   NAND2_X1 i_257_76_11374 (.A1(n_257_752), .A2(n_257_76_17935), .ZN(
      n_257_76_11355));
   NAND2_X1 i_257_76_11375 (.A1(n_257_132), .A2(n_257_76_17925), .ZN(
      n_257_76_11356));
   NAND2_X1 i_257_76_11376 (.A1(n_257_918), .A2(n_257_76_17940), .ZN(
      n_257_76_11357));
   NAND2_X1 i_257_76_11377 (.A1(n_257_648), .A2(n_257_76_17928), .ZN(
      n_257_76_11358));
   NAND4_X1 i_257_76_11378 (.A1(n_257_76_11355), .A2(n_257_76_11356), .A3(
      n_257_76_11357), .A4(n_257_76_11358), .ZN(n_257_76_11359));
   INV_X1 i_257_76_11379 (.A(n_257_76_11359), .ZN(n_257_76_11360));
   NAND2_X1 i_257_76_11380 (.A1(n_257_982), .A2(n_257_442), .ZN(n_257_76_11361));
   INV_X1 i_257_76_11381 (.A(n_257_76_11361), .ZN(n_257_76_11362));
   NAND2_X1 i_257_76_11382 (.A1(n_257_76_11362), .A2(n_257_441), .ZN(
      n_257_76_11363));
   NAND2_X1 i_257_76_11383 (.A1(n_257_816), .A2(n_257_76_17952), .ZN(
      n_257_76_11364));
   INV_X1 i_257_76_11384 (.A(Small_Packet_Data_Size[19]), .ZN(n_257_76_11365));
   NAND3_X1 i_257_76_11385 (.A1(n_257_76_10896), .A2(n_257_76_11323), .A3(
      n_257_76_18022), .ZN(n_257_76_11366));
   INV_X1 i_257_76_11386 (.A(n_257_76_11366), .ZN(n_257_76_11367));
   NAND4_X1 i_257_76_11387 (.A1(n_257_76_11367), .A2(n_257_76_10895), .A3(
      n_257_76_10825), .A4(n_257_76_11328), .ZN(n_257_76_11368));
   NAND2_X1 i_257_76_11388 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[19]), 
      .ZN(n_257_76_11369));
   NAND2_X1 i_257_76_11389 (.A1(n_257_76_11368), .A2(n_257_76_11369), .ZN(
      n_257_76_11370));
   NAND3_X1 i_257_76_11390 (.A1(n_257_76_11363), .A2(n_257_76_11364), .A3(
      n_257_76_11370), .ZN(n_257_76_11371));
   INV_X1 i_257_76_11391 (.A(n_257_76_11371), .ZN(n_257_76_11372));
   NAND3_X1 i_257_76_11392 (.A1(n_257_76_11354), .A2(n_257_76_11360), .A3(
      n_257_76_11372), .ZN(n_257_76_11373));
   INV_X1 i_257_76_11393 (.A(n_257_76_11373), .ZN(n_257_76_11374));
   INV_X1 i_257_76_11394 (.A(n_257_816), .ZN(n_257_76_11375));
   NAND2_X1 i_257_76_11395 (.A1(n_257_76_11375), .A2(n_257_442), .ZN(
      n_257_76_11376));
   INV_X1 i_257_76_11396 (.A(n_257_752), .ZN(n_257_76_11377));
   NAND2_X1 i_257_76_11397 (.A1(n_257_76_11377), .A2(n_257_442), .ZN(
      n_257_76_11378));
   INV_X1 i_257_76_11398 (.A(n_257_918), .ZN(n_257_76_11379));
   NAND2_X1 i_257_76_11399 (.A1(n_257_76_11379), .A2(n_257_442), .ZN(
      n_257_76_11380));
   NAND4_X1 i_257_76_11400 (.A1(n_257_76_11376), .A2(n_257_76_11378), .A3(
      n_257_76_11380), .A4(n_257_76_13029), .ZN(n_257_76_11381));
   INV_X1 i_257_76_11401 (.A(n_257_76_10908), .ZN(n_257_76_11382));
   NAND2_X1 i_257_76_11402 (.A1(n_257_76_11381), .A2(n_257_76_11382), .ZN(
      n_257_76_11383));
   NAND2_X1 i_257_76_11403 (.A1(n_257_688), .A2(n_257_76_17958), .ZN(
      n_257_76_11384));
   NAND4_X1 i_257_76_11404 (.A1(n_257_76_11342), .A2(n_257_76_11374), .A3(
      n_257_76_11383), .A4(n_257_76_11384), .ZN(n_257_76_11385));
   NAND2_X1 i_257_76_11405 (.A1(n_257_1014), .A2(n_257_76_17964), .ZN(
      n_257_76_11386));
   NAND4_X1 i_257_76_11406 (.A1(n_257_76_11000), .A2(n_257_76_11386), .A3(
      n_257_76_11293), .A4(n_257_76_11312), .ZN(n_257_76_11387));
   NOR2_X1 i_257_76_11407 (.A1(n_257_76_11385), .A2(n_257_76_11387), .ZN(
      n_257_76_11388));
   NAND3_X1 i_257_76_11408 (.A1(n_257_76_11225), .A2(n_257_76_10921), .A3(
      n_257_76_11242), .ZN(n_257_76_11389));
   INV_X1 i_257_76_11409 (.A(n_257_76_11389), .ZN(n_257_76_11390));
   NAND2_X1 i_257_76_11410 (.A1(n_257_1046), .A2(n_257_76_17969), .ZN(
      n_257_76_11391));
   NAND3_X1 i_257_76_11411 (.A1(n_257_76_11388), .A2(n_257_76_11390), .A3(
      n_257_76_11391), .ZN(n_257_76_11392));
   NAND3_X1 i_257_76_11412 (.A1(n_257_76_11318), .A2(n_257_76_11338), .A3(
      n_257_76_11392), .ZN(n_257_76_11393));
   INV_X1 i_257_76_11413 (.A(n_257_76_11393), .ZN(n_257_76_11394));
   NAND3_X1 i_257_76_11414 (.A1(n_257_76_11248), .A2(n_257_76_11299), .A3(
      n_257_76_11394), .ZN(n_257_76_11395));
   NOR2_X1 i_257_76_11415 (.A1(n_257_76_11202), .A2(n_257_76_11395), .ZN(
      n_257_76_11396));
   NAND2_X1 i_257_76_11416 (.A1(n_257_76_11059), .A2(n_257_76_11396), .ZN(n_19));
   NAND2_X1 i_257_76_11417 (.A1(n_257_1047), .A2(n_257_443), .ZN(n_257_76_11397));
   NAND2_X1 i_257_76_11418 (.A1(n_257_1015), .A2(n_257_444), .ZN(n_257_76_11398));
   NAND2_X1 i_257_76_11419 (.A1(n_257_441), .A2(n_257_983), .ZN(n_257_76_11399));
   INV_X1 i_257_76_11420 (.A(n_257_1079), .ZN(n_257_76_11400));
   NAND2_X1 i_257_76_11421 (.A1(n_257_951), .A2(n_257_442), .ZN(n_257_76_11401));
   INV_X1 i_257_76_11422 (.A(n_257_76_11401), .ZN(n_257_76_11402));
   NAND3_X1 i_257_76_11423 (.A1(n_257_76_11400), .A2(n_257_440), .A3(
      n_257_76_11402), .ZN(n_257_76_11403));
   INV_X1 i_257_76_11424 (.A(n_257_76_11403), .ZN(n_257_76_11404));
   NAND2_X1 i_257_76_11425 (.A1(n_257_76_11399), .A2(n_257_76_11404), .ZN(
      n_257_76_11405));
   INV_X1 i_257_76_11426 (.A(n_257_76_11405), .ZN(n_257_76_11406));
   NAND2_X1 i_257_76_11427 (.A1(n_257_76_11398), .A2(n_257_76_11406), .ZN(
      n_257_76_11407));
   INV_X1 i_257_76_11428 (.A(n_257_76_11407), .ZN(n_257_76_11408));
   NAND2_X1 i_257_76_11429 (.A1(n_257_76_11397), .A2(n_257_76_11408), .ZN(
      n_257_76_11409));
   INV_X1 i_257_76_11430 (.A(n_257_76_11409), .ZN(n_257_76_11410));
   NAND2_X1 i_257_76_11431 (.A1(n_257_17), .A2(n_257_76_11410), .ZN(
      n_257_76_11411));
   NOR2_X1 i_257_76_11432 (.A1(n_257_1079), .A2(n_257_76_17412), .ZN(
      n_257_76_11412));
   INV_X1 i_257_76_11433 (.A(n_257_76_11412), .ZN(n_257_76_11413));
   NOR2_X1 i_257_76_11434 (.A1(n_257_76_11413), .A2(n_257_76_15197), .ZN(
      n_257_76_11414));
   NAND2_X1 i_257_76_11435 (.A1(n_257_1047), .A2(n_257_76_11414), .ZN(
      n_257_76_11415));
   INV_X1 i_257_76_11436 (.A(n_257_76_11415), .ZN(n_257_76_11416));
   NAND2_X1 i_257_76_11437 (.A1(n_257_76_18072), .A2(n_257_76_11416), .ZN(
      n_257_76_11417));
   INV_X1 i_257_76_11438 (.A(n_257_76_11397), .ZN(n_257_76_11418));
   NAND2_X1 i_257_76_11439 (.A1(n_257_919), .A2(n_257_439), .ZN(n_257_76_11419));
   NAND2_X1 i_257_76_11440 (.A1(n_257_753), .A2(n_257_436), .ZN(n_257_76_11420));
   NAND2_X1 i_257_76_11441 (.A1(n_257_817), .A2(n_257_437), .ZN(n_257_76_11421));
   NAND4_X1 i_257_76_11442 (.A1(n_257_76_11419), .A2(n_257_76_11420), .A3(
      n_257_76_11421), .A4(n_257_76_11399), .ZN(n_257_76_11422));
   NAND2_X1 i_257_76_11443 (.A1(n_257_449), .A2(n_257_895), .ZN(n_257_76_11423));
   NAND2_X1 i_257_76_11444 (.A1(n_257_447), .A2(n_257_785), .ZN(n_257_76_11424));
   NAND3_X1 i_257_76_11445 (.A1(n_257_76_11423), .A2(n_257_76_11424), .A3(
      n_257_649), .ZN(n_257_76_11425));
   INV_X1 i_257_76_11446 (.A(n_257_76_11425), .ZN(n_257_76_11426));
   NAND2_X1 i_257_76_11447 (.A1(n_257_881), .A2(n_257_445), .ZN(n_257_76_11427));
   NAND2_X1 i_257_76_11448 (.A1(n_257_446), .A2(n_257_849), .ZN(n_257_76_11428));
   NAND2_X1 i_257_76_11449 (.A1(n_257_76_11427), .A2(n_257_76_11428), .ZN(
      n_257_76_11429));
   INV_X1 i_257_76_11450 (.A(n_257_76_11429), .ZN(n_257_76_11430));
   NOR2_X1 i_257_76_11451 (.A1(n_257_1079), .A2(n_257_76_17927), .ZN(
      n_257_76_11431));
   NAND2_X1 i_257_76_11452 (.A1(n_257_440), .A2(n_257_951), .ZN(n_257_76_11432));
   NAND2_X1 i_257_76_11453 (.A1(n_257_438), .A2(n_257_1085), .ZN(n_257_76_11433));
   NAND2_X1 i_257_76_11454 (.A1(n_257_721), .A2(n_257_435), .ZN(n_257_76_11434));
   NAND4_X1 i_257_76_11455 (.A1(n_257_76_11431), .A2(n_257_76_11432), .A3(
      n_257_76_11433), .A4(n_257_76_11434), .ZN(n_257_76_11435));
   INV_X1 i_257_76_11456 (.A(n_257_76_11435), .ZN(n_257_76_11436));
   NAND3_X1 i_257_76_11457 (.A1(n_257_76_11426), .A2(n_257_76_11430), .A3(
      n_257_76_11436), .ZN(n_257_76_11437));
   NOR2_X1 i_257_76_11458 (.A1(n_257_76_11422), .A2(n_257_76_11437), .ZN(
      n_257_76_11438));
   NAND2_X1 i_257_76_11459 (.A1(n_257_689), .A2(n_257_448), .ZN(n_257_76_11439));
   NAND3_X1 i_257_76_11460 (.A1(n_257_76_11398), .A2(n_257_76_11438), .A3(
      n_257_76_11439), .ZN(n_257_76_11440));
   NOR2_X1 i_257_76_11461 (.A1(n_257_76_11418), .A2(n_257_76_11440), .ZN(
      n_257_76_11441));
   NAND2_X1 i_257_76_11462 (.A1(n_257_28), .A2(n_257_76_11441), .ZN(
      n_257_76_11442));
   NAND3_X1 i_257_76_11463 (.A1(n_257_76_11411), .A2(n_257_76_11417), .A3(
      n_257_76_11442), .ZN(n_257_76_11443));
   NAND2_X1 i_257_76_11464 (.A1(n_257_76_11427), .A2(n_257_446), .ZN(
      n_257_76_11444));
   INV_X1 i_257_76_11465 (.A(n_257_76_11444), .ZN(n_257_76_11445));
   NAND2_X1 i_257_76_11466 (.A1(n_257_849), .A2(n_257_442), .ZN(n_257_76_11446));
   NOR2_X1 i_257_76_11467 (.A1(n_257_1079), .A2(n_257_76_11446), .ZN(
      n_257_76_11447));
   NAND3_X1 i_257_76_11468 (.A1(n_257_76_11447), .A2(n_257_76_11432), .A3(
      n_257_76_11433), .ZN(n_257_76_11448));
   INV_X1 i_257_76_11469 (.A(n_257_76_11448), .ZN(n_257_76_11449));
   NAND4_X1 i_257_76_11470 (.A1(n_257_76_11419), .A2(n_257_76_11445), .A3(
      n_257_76_11399), .A4(n_257_76_11449), .ZN(n_257_76_11450));
   INV_X1 i_257_76_11471 (.A(n_257_76_11450), .ZN(n_257_76_11451));
   NAND2_X1 i_257_76_11472 (.A1(n_257_76_11398), .A2(n_257_76_11451), .ZN(
      n_257_76_11452));
   INV_X1 i_257_76_11473 (.A(n_257_76_11452), .ZN(n_257_76_11453));
   NAND2_X1 i_257_76_11474 (.A1(n_257_76_11397), .A2(n_257_76_11453), .ZN(
      n_257_76_11454));
   INV_X1 i_257_76_11475 (.A(n_257_76_11454), .ZN(n_257_76_11455));
   NAND2_X1 i_257_76_11476 (.A1(n_257_76_18070), .A2(n_257_76_11455), .ZN(
      n_257_76_11456));
   NAND3_X1 i_257_76_11477 (.A1(n_257_76_11412), .A2(n_257_76_11432), .A3(
      n_257_439), .ZN(n_257_76_11457));
   INV_X1 i_257_76_11478 (.A(n_257_76_11457), .ZN(n_257_76_11458));
   NAND3_X1 i_257_76_11479 (.A1(n_257_76_11458), .A2(n_257_76_11399), .A3(
      n_257_919), .ZN(n_257_76_11459));
   INV_X1 i_257_76_11480 (.A(n_257_76_11459), .ZN(n_257_76_11460));
   NAND2_X1 i_257_76_11481 (.A1(n_257_76_11398), .A2(n_257_76_11460), .ZN(
      n_257_76_11461));
   INV_X1 i_257_76_11482 (.A(n_257_76_11461), .ZN(n_257_76_11462));
   NAND2_X1 i_257_76_11483 (.A1(n_257_76_11397), .A2(n_257_76_11462), .ZN(
      n_257_76_11463));
   INV_X1 i_257_76_11484 (.A(n_257_76_11463), .ZN(n_257_76_11464));
   NAND2_X1 i_257_76_11485 (.A1(n_257_76_18084), .A2(n_257_76_11464), .ZN(
      n_257_76_11465));
   NAND2_X1 i_257_76_11486 (.A1(n_257_432), .A2(n_257_617), .ZN(n_257_76_11466));
   NAND3_X1 i_257_76_11487 (.A1(n_257_76_18016), .A2(n_257_76_11466), .A3(
      n_257_423), .ZN(n_257_76_11467));
   INV_X1 i_257_76_11488 (.A(n_257_76_11467), .ZN(n_257_76_11468));
   NAND3_X1 i_257_76_11489 (.A1(n_257_76_11468), .A2(n_257_76_11434), .A3(
      n_257_76_11400), .ZN(n_257_76_11469));
   NAND2_X1 i_257_76_11490 (.A1(n_257_212), .A2(n_257_427), .ZN(n_257_76_11470));
   NAND2_X1 i_257_76_11491 (.A1(n_257_76_11470), .A2(n_257_76_11433), .ZN(
      n_257_76_11471));
   NOR2_X1 i_257_76_11492 (.A1(n_257_76_11469), .A2(n_257_76_11471), .ZN(
      n_257_76_11472));
   NAND2_X1 i_257_76_11493 (.A1(n_257_521), .A2(n_257_424), .ZN(n_257_76_11473));
   NAND2_X1 i_257_76_11494 (.A1(n_257_76_11473), .A2(n_257_76_11427), .ZN(
      n_257_76_11474));
   INV_X1 i_257_76_11495 (.A(n_257_76_11474), .ZN(n_257_76_11475));
   NAND2_X1 i_257_76_11496 (.A1(n_257_649), .A2(n_257_450), .ZN(n_257_76_11476));
   NAND2_X1 i_257_76_11497 (.A1(n_257_55), .A2(n_257_433), .ZN(n_257_76_11477));
   NAND3_X1 i_257_76_11498 (.A1(n_257_76_11477), .A2(n_257_292), .A3(
      n_257_76_11432), .ZN(n_257_76_11478));
   INV_X1 i_257_76_11499 (.A(n_257_76_11478), .ZN(n_257_76_11479));
   NAND4_X1 i_257_76_11500 (.A1(n_257_76_11472), .A2(n_257_76_11475), .A3(
      n_257_76_11476), .A4(n_257_76_11479), .ZN(n_257_76_11480));
   INV_X1 i_257_76_11501 (.A(n_257_76_11480), .ZN(n_257_76_11481));
   NAND2_X1 i_257_76_11502 (.A1(n_257_172), .A2(n_257_429), .ZN(n_257_76_11482));
   NAND2_X1 i_257_76_11503 (.A1(n_257_252), .A2(n_257_425), .ZN(n_257_76_11483));
   NAND3_X1 i_257_76_11504 (.A1(n_257_76_11481), .A2(n_257_76_11482), .A3(
      n_257_76_11483), .ZN(n_257_76_11484));
   NAND2_X1 i_257_76_11505 (.A1(n_257_76_11423), .A2(n_257_76_11424), .ZN(
      n_257_76_11485));
   INV_X1 i_257_76_11506 (.A(n_257_76_11485), .ZN(n_257_76_11486));
   NAND2_X1 i_257_76_11507 (.A1(n_257_451), .A2(n_257_472), .ZN(n_257_76_11487));
   NAND4_X1 i_257_76_11508 (.A1(n_257_76_11486), .A2(n_257_76_11487), .A3(
      n_257_76_11399), .A4(n_257_76_11428), .ZN(n_257_76_11488));
   INV_X1 i_257_76_11509 (.A(n_257_76_11488), .ZN(n_257_76_11489));
   NAND2_X1 i_257_76_11510 (.A1(n_257_553), .A2(n_257_426), .ZN(n_257_76_11490));
   NAND2_X1 i_257_76_11511 (.A1(n_257_76_11490), .A2(n_257_76_11419), .ZN(
      n_257_76_11491));
   INV_X1 i_257_76_11512 (.A(n_257_76_11491), .ZN(n_257_76_11492));
   NAND2_X1 i_257_76_11513 (.A1(n_257_133), .A2(n_257_430), .ZN(n_257_76_11493));
   NAND3_X1 i_257_76_11514 (.A1(n_257_76_11420), .A2(n_257_76_11493), .A3(
      n_257_76_11421), .ZN(n_257_76_11494));
   INV_X1 i_257_76_11515 (.A(n_257_76_11494), .ZN(n_257_76_11495));
   NAND2_X1 i_257_76_11516 (.A1(n_257_95), .A2(n_257_431), .ZN(n_257_76_11496));
   NAND4_X1 i_257_76_11517 (.A1(n_257_76_11489), .A2(n_257_76_11492), .A3(
      n_257_76_11495), .A4(n_257_76_11496), .ZN(n_257_76_11497));
   NOR2_X1 i_257_76_11518 (.A1(n_257_76_11484), .A2(n_257_76_11497), .ZN(
      n_257_76_11498));
   NAND2_X1 i_257_76_11519 (.A1(n_257_76_11398), .A2(n_257_76_11439), .ZN(
      n_257_76_11499));
   INV_X1 i_257_76_11520 (.A(n_257_76_11499), .ZN(n_257_76_11500));
   NAND3_X1 i_257_76_11521 (.A1(n_257_76_11498), .A2(n_257_76_11397), .A3(
      n_257_76_11500), .ZN(n_257_76_11501));
   INV_X1 i_257_76_11522 (.A(n_257_76_11501), .ZN(n_257_76_11502));
   NAND2_X1 i_257_76_11523 (.A1(n_257_76_18066), .A2(n_257_76_11502), .ZN(
      n_257_76_11503));
   NAND3_X1 i_257_76_11524 (.A1(n_257_76_11456), .A2(n_257_76_11465), .A3(
      n_257_76_11503), .ZN(n_257_76_11504));
   NOR2_X1 i_257_76_11525 (.A1(n_257_76_11443), .A2(n_257_76_11504), .ZN(
      n_257_76_11505));
   NAND3_X1 i_257_76_11526 (.A1(n_257_441), .A2(n_257_983), .A3(n_257_76_11412), 
      .ZN(n_257_76_11506));
   INV_X1 i_257_76_11527 (.A(n_257_76_11506), .ZN(n_257_76_11507));
   NAND2_X1 i_257_76_11528 (.A1(n_257_76_11398), .A2(n_257_76_11507), .ZN(
      n_257_76_11508));
   INV_X1 i_257_76_11529 (.A(n_257_76_11508), .ZN(n_257_76_11509));
   NAND2_X1 i_257_76_11530 (.A1(n_257_76_11397), .A2(n_257_76_11509), .ZN(
      n_257_76_11510));
   INV_X1 i_257_76_11531 (.A(n_257_76_11510), .ZN(n_257_76_11511));
   NAND2_X1 i_257_76_11532 (.A1(n_257_76_18071), .A2(n_257_76_11511), .ZN(
      n_257_76_11512));
   NAND2_X1 i_257_76_11533 (.A1(n_257_76_11428), .A2(n_257_76_11424), .ZN(
      n_257_76_11513));
   INV_X1 i_257_76_11534 (.A(n_257_76_11513), .ZN(n_257_76_11514));
   NAND2_X1 i_257_76_11535 (.A1(n_257_76_11432), .A2(n_257_76_11433), .ZN(
      n_257_76_11515));
   NAND3_X1 i_257_76_11536 (.A1(n_257_76_11400), .A2(n_257_721), .A3(
      n_257_76_15655), .ZN(n_257_76_11516));
   NOR2_X1 i_257_76_11537 (.A1(n_257_76_11515), .A2(n_257_76_11516), .ZN(
      n_257_76_11517));
   NAND4_X1 i_257_76_11538 (.A1(n_257_76_11514), .A2(n_257_76_11517), .A3(
      n_257_76_11399), .A4(n_257_76_11427), .ZN(n_257_76_11518));
   NAND3_X1 i_257_76_11539 (.A1(n_257_76_11419), .A2(n_257_76_11420), .A3(
      n_257_76_11421), .ZN(n_257_76_11519));
   NOR2_X1 i_257_76_11540 (.A1(n_257_76_11518), .A2(n_257_76_11519), .ZN(
      n_257_76_11520));
   NAND2_X1 i_257_76_11541 (.A1(n_257_76_11398), .A2(n_257_76_11520), .ZN(
      n_257_76_11521));
   INV_X1 i_257_76_11542 (.A(n_257_76_11521), .ZN(n_257_76_11522));
   NAND2_X1 i_257_76_11543 (.A1(n_257_76_11397), .A2(n_257_76_11522), .ZN(
      n_257_76_11523));
   INV_X1 i_257_76_11544 (.A(n_257_76_11523), .ZN(n_257_76_11524));
   NAND2_X1 i_257_76_11545 (.A1(n_257_76_18078), .A2(n_257_76_11524), .ZN(
      n_257_76_11525));
   NAND3_X1 i_257_76_11546 (.A1(n_257_76_11419), .A2(n_257_76_11420), .A3(
      n_257_76_11493), .ZN(n_257_76_11526));
   NAND3_X1 i_257_76_11547 (.A1(n_257_76_11421), .A2(n_257_76_11487), .A3(
      n_257_76_11399), .ZN(n_257_76_11527));
   NOR2_X1 i_257_76_11548 (.A1(n_257_76_11526), .A2(n_257_76_11527), .ZN(
      n_257_76_11528));
   NAND4_X1 i_257_76_11549 (.A1(n_257_76_11476), .A2(n_257_76_11427), .A3(
      n_257_76_11428), .A4(n_257_76_11423), .ZN(n_257_76_11529));
   NAND3_X1 i_257_76_11550 (.A1(n_257_585), .A2(n_257_428), .A3(n_257_442), 
      .ZN(n_257_76_11530));
   INV_X1 i_257_76_11551 (.A(n_257_76_11530), .ZN(n_257_76_11531));
   NAND2_X1 i_257_76_11552 (.A1(n_257_76_11531), .A2(n_257_76_11466), .ZN(
      n_257_76_11532));
   INV_X1 i_257_76_11553 (.A(n_257_76_11532), .ZN(n_257_76_11533));
   NAND3_X1 i_257_76_11554 (.A1(n_257_76_11434), .A2(n_257_76_11400), .A3(
      n_257_76_11533), .ZN(n_257_76_11534));
   INV_X1 i_257_76_11555 (.A(n_257_76_11534), .ZN(n_257_76_11535));
   INV_X1 i_257_76_11556 (.A(n_257_76_11515), .ZN(n_257_76_11536));
   NAND4_X1 i_257_76_11557 (.A1(n_257_76_11535), .A2(n_257_76_11536), .A3(
      n_257_76_11424), .A4(n_257_76_11477), .ZN(n_257_76_11537));
   NOR2_X1 i_257_76_11558 (.A1(n_257_76_11529), .A2(n_257_76_11537), .ZN(
      n_257_76_11538));
   NAND4_X1 i_257_76_11559 (.A1(n_257_76_11528), .A2(n_257_76_11482), .A3(
      n_257_76_11538), .A4(n_257_76_11496), .ZN(n_257_76_11539));
   INV_X1 i_257_76_11560 (.A(n_257_76_11539), .ZN(n_257_76_11540));
   NAND3_X1 i_257_76_11561 (.A1(n_257_76_11397), .A2(n_257_76_11540), .A3(
      n_257_76_11500), .ZN(n_257_76_11541));
   INV_X1 i_257_76_11562 (.A(n_257_76_11541), .ZN(n_257_76_11542));
   NAND2_X1 i_257_76_11563 (.A1(n_257_76_18074), .A2(n_257_76_11542), .ZN(
      n_257_76_11543));
   NAND3_X1 i_257_76_11564 (.A1(n_257_76_11512), .A2(n_257_76_11525), .A3(
      n_257_76_11543), .ZN(n_257_76_11544));
   NAND2_X1 i_257_76_11565 (.A1(n_257_1079), .A2(n_257_442), .ZN(n_257_76_11545));
   INV_X1 i_257_76_11566 (.A(n_257_76_11545), .ZN(n_257_76_11546));
   NAND2_X1 i_257_76_11567 (.A1(n_257_13), .A2(n_257_76_11546), .ZN(
      n_257_76_11547));
   NAND2_X1 i_257_76_11568 (.A1(n_257_881), .A2(n_257_76_11412), .ZN(
      n_257_76_11548));
   NAND3_X1 i_257_76_11569 (.A1(n_257_76_11432), .A2(n_257_76_11433), .A3(
      n_257_445), .ZN(n_257_76_11549));
   NOR2_X1 i_257_76_11570 (.A1(n_257_76_11548), .A2(n_257_76_11549), .ZN(
      n_257_76_11550));
   NAND3_X1 i_257_76_11571 (.A1(n_257_76_11550), .A2(n_257_76_11419), .A3(
      n_257_76_11399), .ZN(n_257_76_11551));
   INV_X1 i_257_76_11572 (.A(n_257_76_11551), .ZN(n_257_76_11552));
   NAND2_X1 i_257_76_11573 (.A1(n_257_76_11398), .A2(n_257_76_11552), .ZN(
      n_257_76_11553));
   INV_X1 i_257_76_11574 (.A(n_257_76_11553), .ZN(n_257_76_11554));
   NAND2_X1 i_257_76_11575 (.A1(n_257_76_11397), .A2(n_257_76_11554), .ZN(
      n_257_76_11555));
   INV_X1 i_257_76_11576 (.A(n_257_76_11555), .ZN(n_257_76_11556));
   NAND2_X1 i_257_76_11577 (.A1(n_257_76_18077), .A2(n_257_76_11556), .ZN(
      n_257_76_11557));
   NAND2_X1 i_257_76_11578 (.A1(n_257_76_11547), .A2(n_257_76_11557), .ZN(
      n_257_76_11558));
   NOR2_X1 i_257_76_11579 (.A1(n_257_76_11544), .A2(n_257_76_11558), .ZN(
      n_257_76_11559));
   NAND3_X1 i_257_76_11580 (.A1(n_257_76_11399), .A2(n_257_553), .A3(
      n_257_76_11476), .ZN(n_257_76_11560));
   NAND2_X1 i_257_76_11581 (.A1(n_257_76_11421), .A2(n_257_76_11487), .ZN(
      n_257_76_11561));
   NOR2_X1 i_257_76_11582 (.A1(n_257_76_11560), .A2(n_257_76_11561), .ZN(
      n_257_76_11562));
   NAND3_X1 i_257_76_11583 (.A1(n_257_76_18016), .A2(n_257_76_11466), .A3(
      n_257_426), .ZN(n_257_76_11563));
   INV_X1 i_257_76_11584 (.A(n_257_76_11563), .ZN(n_257_76_11564));
   NAND3_X1 i_257_76_11585 (.A1(n_257_76_11564), .A2(n_257_76_11434), .A3(
      n_257_76_11400), .ZN(n_257_76_11565));
   INV_X1 i_257_76_11586 (.A(n_257_76_11565), .ZN(n_257_76_11566));
   NAND3_X1 i_257_76_11587 (.A1(n_257_76_11432), .A2(n_257_76_11470), .A3(
      n_257_76_11433), .ZN(n_257_76_11567));
   INV_X1 i_257_76_11588 (.A(n_257_76_11567), .ZN(n_257_76_11568));
   NAND3_X1 i_257_76_11589 (.A1(n_257_76_11566), .A2(n_257_76_11568), .A3(
      n_257_76_11477), .ZN(n_257_76_11569));
   NAND4_X1 i_257_76_11590 (.A1(n_257_76_11427), .A2(n_257_76_11428), .A3(
      n_257_76_11423), .A4(n_257_76_11424), .ZN(n_257_76_11570));
   NOR2_X1 i_257_76_11591 (.A1(n_257_76_11569), .A2(n_257_76_11570), .ZN(
      n_257_76_11571));
   INV_X1 i_257_76_11592 (.A(n_257_76_11526), .ZN(n_257_76_11572));
   NAND4_X1 i_257_76_11593 (.A1(n_257_76_11562), .A2(n_257_76_11571), .A3(
      n_257_76_11572), .A4(n_257_76_11496), .ZN(n_257_76_11573));
   INV_X1 i_257_76_11594 (.A(n_257_76_11573), .ZN(n_257_76_11574));
   NAND2_X1 i_257_76_11595 (.A1(n_257_76_11439), .A2(n_257_76_11482), .ZN(
      n_257_76_11575));
   INV_X1 i_257_76_11596 (.A(n_257_76_11575), .ZN(n_257_76_11576));
   NAND3_X1 i_257_76_11597 (.A1(n_257_76_11574), .A2(n_257_76_11576), .A3(
      n_257_76_11398), .ZN(n_257_76_11577));
   NOR2_X1 i_257_76_11598 (.A1(n_257_76_11577), .A2(n_257_76_11418), .ZN(
      n_257_76_11578));
   NAND2_X1 i_257_76_11599 (.A1(n_257_76_18076), .A2(n_257_76_11578), .ZN(
      n_257_76_11579));
   NOR2_X1 i_257_76_11600 (.A1(n_257_1079), .A2(n_257_76_17934), .ZN(
      n_257_76_11580));
   NAND3_X1 i_257_76_11601 (.A1(n_257_76_11580), .A2(n_257_76_11432), .A3(
      n_257_76_11433), .ZN(n_257_76_11581));
   INV_X1 i_257_76_11602 (.A(n_257_76_11581), .ZN(n_257_76_11582));
   NAND4_X1 i_257_76_11603 (.A1(n_257_76_11514), .A2(n_257_76_11582), .A3(
      n_257_753), .A4(n_257_76_11427), .ZN(n_257_76_11583));
   NAND3_X1 i_257_76_11604 (.A1(n_257_76_11419), .A2(n_257_76_11421), .A3(
      n_257_76_11399), .ZN(n_257_76_11584));
   NOR2_X1 i_257_76_11605 (.A1(n_257_76_11583), .A2(n_257_76_11584), .ZN(
      n_257_76_11585));
   NAND2_X1 i_257_76_11606 (.A1(n_257_76_11398), .A2(n_257_76_11585), .ZN(
      n_257_76_11586));
   INV_X1 i_257_76_11607 (.A(n_257_76_11586), .ZN(n_257_76_11587));
   NAND2_X1 i_257_76_11608 (.A1(n_257_76_11397), .A2(n_257_76_11587), .ZN(
      n_257_76_11588));
   INV_X1 i_257_76_11609 (.A(n_257_76_11588), .ZN(n_257_76_11589));
   NAND2_X1 i_257_76_11610 (.A1(n_257_76_18069), .A2(n_257_76_11589), .ZN(
      n_257_76_11590));
   NAND3_X1 i_257_76_11611 (.A1(n_257_432), .A2(n_257_617), .A3(n_257_442), 
      .ZN(n_257_76_11591));
   NOR2_X1 i_257_76_11612 (.A1(n_257_1079), .A2(n_257_76_11591), .ZN(
      n_257_76_11592));
   NAND4_X1 i_257_76_11613 (.A1(n_257_76_11592), .A2(n_257_76_11432), .A3(
      n_257_76_11433), .A4(n_257_76_11434), .ZN(n_257_76_11593));
   NAND2_X1 i_257_76_11614 (.A1(n_257_76_11424), .A2(n_257_76_11477), .ZN(
      n_257_76_11594));
   NOR2_X1 i_257_76_11615 (.A1(n_257_76_11593), .A2(n_257_76_11594), .ZN(
      n_257_76_11595));
   NAND2_X1 i_257_76_11616 (.A1(n_257_76_11399), .A2(n_257_76_11476), .ZN(
      n_257_76_11596));
   INV_X1 i_257_76_11617 (.A(n_257_76_11596), .ZN(n_257_76_11597));
   NAND3_X1 i_257_76_11618 (.A1(n_257_76_11427), .A2(n_257_76_11428), .A3(
      n_257_76_11423), .ZN(n_257_76_11598));
   INV_X1 i_257_76_11619 (.A(n_257_76_11598), .ZN(n_257_76_11599));
   NAND3_X1 i_257_76_11620 (.A1(n_257_76_11595), .A2(n_257_76_11597), .A3(
      n_257_76_11599), .ZN(n_257_76_11600));
   NAND4_X1 i_257_76_11621 (.A1(n_257_76_11419), .A2(n_257_76_11420), .A3(
      n_257_76_11421), .A4(n_257_76_11487), .ZN(n_257_76_11601));
   NOR2_X1 i_257_76_11622 (.A1(n_257_76_11600), .A2(n_257_76_11601), .ZN(
      n_257_76_11602));
   NAND3_X1 i_257_76_11623 (.A1(n_257_76_11602), .A2(n_257_76_11398), .A3(
      n_257_76_11439), .ZN(n_257_76_11603));
   NOR2_X1 i_257_76_11624 (.A1(n_257_76_11603), .A2(n_257_76_11418), .ZN(
      n_257_76_11604));
   NAND2_X1 i_257_76_11625 (.A1(n_257_68), .A2(n_257_76_11604), .ZN(
      n_257_76_11605));
   NAND3_X1 i_257_76_11626 (.A1(n_257_76_11579), .A2(n_257_76_11590), .A3(
      n_257_76_11605), .ZN(n_257_76_11606));
   NOR2_X1 i_257_76_11627 (.A1(n_257_1079), .A2(n_257_76_17951), .ZN(
      n_257_76_11607));
   NAND3_X1 i_257_76_11628 (.A1(n_257_76_11607), .A2(n_257_76_11432), .A3(
      n_257_76_11433), .ZN(n_257_76_11608));
   INV_X1 i_257_76_11629 (.A(n_257_76_11608), .ZN(n_257_76_11609));
   NAND4_X1 i_257_76_11630 (.A1(n_257_76_11609), .A2(n_257_817), .A3(
      n_257_76_11427), .A4(n_257_76_11428), .ZN(n_257_76_11610));
   NAND2_X1 i_257_76_11631 (.A1(n_257_76_11419), .A2(n_257_76_11399), .ZN(
      n_257_76_11611));
   NOR2_X1 i_257_76_11632 (.A1(n_257_76_11610), .A2(n_257_76_11611), .ZN(
      n_257_76_11612));
   NAND2_X1 i_257_76_11633 (.A1(n_257_76_11398), .A2(n_257_76_11612), .ZN(
      n_257_76_11613));
   INV_X1 i_257_76_11634 (.A(n_257_76_11613), .ZN(n_257_76_11614));
   NAND2_X1 i_257_76_11635 (.A1(n_257_76_11397), .A2(n_257_76_11614), .ZN(
      n_257_76_11615));
   INV_X1 i_257_76_11636 (.A(n_257_76_11615), .ZN(n_257_76_11616));
   NAND2_X1 i_257_76_11637 (.A1(n_257_22), .A2(n_257_76_11616), .ZN(
      n_257_76_11617));
   NAND2_X1 i_257_76_11638 (.A1(n_257_444), .A2(n_257_76_11412), .ZN(
      n_257_76_11618));
   INV_X1 i_257_76_11639 (.A(n_257_76_11618), .ZN(n_257_76_11619));
   NAND2_X1 i_257_76_11640 (.A1(n_257_1015), .A2(n_257_76_11619), .ZN(
      n_257_76_11620));
   INV_X1 i_257_76_11641 (.A(n_257_76_11620), .ZN(n_257_76_11621));
   NAND2_X1 i_257_76_11642 (.A1(n_257_76_11397), .A2(n_257_76_11621), .ZN(
      n_257_76_11622));
   INV_X1 i_257_76_11643 (.A(n_257_76_11622), .ZN(n_257_76_11623));
   NAND2_X1 i_257_76_11644 (.A1(n_257_76_18075), .A2(n_257_76_11623), .ZN(
      n_257_76_11624));
   NAND2_X1 i_257_76_11645 (.A1(n_257_76_11617), .A2(n_257_76_11624), .ZN(
      n_257_76_11625));
   NOR2_X1 i_257_76_11646 (.A1(n_257_76_11606), .A2(n_257_76_11625), .ZN(
      n_257_76_11626));
   NAND3_X1 i_257_76_11647 (.A1(n_257_76_11505), .A2(n_257_76_11559), .A3(
      n_257_76_11626), .ZN(n_257_76_11627));
   INV_X1 i_257_76_11648 (.A(n_257_76_11627), .ZN(n_257_76_11628));
   NOR2_X1 i_257_76_11649 (.A1(n_257_1079), .A2(n_257_76_17633), .ZN(
      n_257_76_11629));
   NAND4_X1 i_257_76_11650 (.A1(n_257_76_11629), .A2(n_257_55), .A3(
      n_257_76_11433), .A4(n_257_76_11434), .ZN(n_257_76_11630));
   NAND2_X1 i_257_76_11651 (.A1(n_257_76_11424), .A2(n_257_76_11432), .ZN(
      n_257_76_11631));
   NOR2_X1 i_257_76_11652 (.A1(n_257_76_11630), .A2(n_257_76_11631), .ZN(
      n_257_76_11632));
   NAND3_X1 i_257_76_11653 (.A1(n_257_76_11632), .A2(n_257_76_11597), .A3(
      n_257_76_11599), .ZN(n_257_76_11633));
   NOR2_X1 i_257_76_11654 (.A1(n_257_76_11633), .A2(n_257_76_11601), .ZN(
      n_257_76_11634));
   NAND3_X1 i_257_76_11655 (.A1(n_257_76_11634), .A2(n_257_76_11398), .A3(
      n_257_76_11439), .ZN(n_257_76_11635));
   NOR2_X1 i_257_76_11656 (.A1(n_257_76_11635), .A2(n_257_76_11418), .ZN(
      n_257_76_11636));
   NAND2_X1 i_257_76_11657 (.A1(n_257_76_18081), .A2(n_257_76_11636), .ZN(
      n_257_76_11637));
   NAND3_X1 i_257_76_11658 (.A1(n_257_76_11427), .A2(n_257_76_11428), .A3(
      n_257_76_11424), .ZN(n_257_76_11638));
   INV_X1 i_257_76_11659 (.A(n_257_76_11638), .ZN(n_257_76_11639));
   NAND3_X1 i_257_76_11660 (.A1(n_257_449), .A2(n_257_76_11432), .A3(
      n_257_76_11433), .ZN(n_257_76_11640));
   NAND3_X1 i_257_76_11661 (.A1(n_257_76_11434), .A2(n_257_76_11400), .A3(
      n_257_76_16220), .ZN(n_257_76_11641));
   NOR2_X1 i_257_76_11662 (.A1(n_257_76_11640), .A2(n_257_76_11641), .ZN(
      n_257_76_11642));
   NAND3_X1 i_257_76_11663 (.A1(n_257_76_11639), .A2(n_257_76_11642), .A3(
      n_257_76_11399), .ZN(n_257_76_11643));
   NOR2_X1 i_257_76_11664 (.A1(n_257_76_11643), .A2(n_257_76_11519), .ZN(
      n_257_76_11644));
   NAND3_X1 i_257_76_11665 (.A1(n_257_76_11398), .A2(n_257_76_11644), .A3(
      n_257_76_11439), .ZN(n_257_76_11645));
   NOR2_X1 i_257_76_11666 (.A1(n_257_76_11418), .A2(n_257_76_11645), .ZN(
      n_257_76_11646));
   NAND2_X1 i_257_76_11667 (.A1(n_257_76_18083), .A2(n_257_76_11646), .ZN(
      n_257_76_11647));
   NAND3_X1 i_257_76_11668 (.A1(n_257_76_11423), .A2(n_257_76_11424), .A3(
      n_257_76_11477), .ZN(n_257_76_11648));
   INV_X1 i_257_76_11669 (.A(n_257_76_11648), .ZN(n_257_76_11649));
   INV_X1 i_257_76_11670 (.A(n_257_617), .ZN(n_257_76_11650));
   NAND2_X1 i_257_76_11671 (.A1(n_257_76_11650), .A2(n_257_442), .ZN(
      n_257_76_11651));
   AOI21_X1 i_257_76_11672 (.A(n_257_76_17101), .B1(n_257_76_12179), .B2(
      n_257_76_11651), .ZN(n_257_76_11652));
   NAND3_X1 i_257_76_11673 (.A1(n_257_76_11434), .A2(n_257_76_11652), .A3(
      n_257_76_11400), .ZN(n_257_76_11653));
   NOR2_X1 i_257_76_11674 (.A1(n_257_76_11653), .A2(n_257_76_11515), .ZN(
      n_257_76_11654));
   NAND3_X1 i_257_76_11675 (.A1(n_257_76_11649), .A2(n_257_76_11430), .A3(
      n_257_76_11654), .ZN(n_257_76_11655));
   NAND4_X1 i_257_76_11676 (.A1(n_257_76_11421), .A2(n_257_76_11487), .A3(
      n_257_76_11399), .A4(n_257_76_11476), .ZN(n_257_76_11656));
   NOR2_X1 i_257_76_11677 (.A1(n_257_76_11655), .A2(n_257_76_11656), .ZN(
      n_257_76_11657));
   NAND3_X1 i_257_76_11678 (.A1(n_257_76_11572), .A2(n_257_172), .A3(
      n_257_76_11496), .ZN(n_257_76_11658));
   INV_X1 i_257_76_11679 (.A(n_257_76_11658), .ZN(n_257_76_11659));
   NAND4_X1 i_257_76_11680 (.A1(n_257_76_11398), .A2(n_257_76_11657), .A3(
      n_257_76_11659), .A4(n_257_76_11439), .ZN(n_257_76_11660));
   NOR2_X1 i_257_76_11681 (.A1(n_257_76_11660), .A2(n_257_76_11418), .ZN(
      n_257_76_11661));
   NAND2_X1 i_257_76_11682 (.A1(n_257_76_18061), .A2(n_257_76_11661), .ZN(
      n_257_76_11662));
   NAND3_X1 i_257_76_11683 (.A1(n_257_76_11637), .A2(n_257_76_11647), .A3(
      n_257_76_11662), .ZN(n_257_76_11663));
   INV_X1 i_257_76_11684 (.A(n_257_76_11663), .ZN(n_257_76_11664));
   INV_X1 i_257_76_11685 (.A(n_257_76_11433), .ZN(n_257_76_11665));
   NAND3_X1 i_257_76_11686 (.A1(n_257_76_11412), .A2(n_257_76_11665), .A3(
      n_257_76_11432), .ZN(n_257_76_11666));
   INV_X1 i_257_76_11687 (.A(n_257_76_11666), .ZN(n_257_76_11667));
   NAND3_X1 i_257_76_11688 (.A1(n_257_76_11419), .A2(n_257_76_11399), .A3(
      n_257_76_11667), .ZN(n_257_76_11668));
   INV_X1 i_257_76_11689 (.A(n_257_76_11668), .ZN(n_257_76_11669));
   NAND2_X1 i_257_76_11690 (.A1(n_257_76_11398), .A2(n_257_76_11669), .ZN(
      n_257_76_11670));
   INV_X1 i_257_76_11691 (.A(n_257_76_11670), .ZN(n_257_76_11671));
   NAND2_X1 i_257_76_11692 (.A1(n_257_76_11397), .A2(n_257_76_11671), .ZN(
      n_257_76_11672));
   INV_X1 i_257_76_11693 (.A(n_257_76_11672), .ZN(n_257_76_11673));
   NAND2_X1 i_257_76_11694 (.A1(n_257_76_18067), .A2(n_257_76_11673), .ZN(
      n_257_76_11674));
   NAND2_X1 i_257_76_11695 (.A1(n_257_369), .A2(n_257_421), .ZN(n_257_76_11675));
   NAND3_X1 i_257_76_11696 (.A1(n_257_76_11675), .A2(n_257_76_11419), .A3(
      n_257_76_11420), .ZN(n_257_76_11676));
   INV_X1 i_257_76_11697 (.A(n_257_76_11676), .ZN(n_257_76_11677));
   NAND2_X1 i_257_76_11698 (.A1(n_257_330), .A2(n_257_422), .ZN(n_257_76_11678));
   NAND2_X1 i_257_76_11699 (.A1(n_257_442), .A2(n_257_489), .ZN(n_257_76_11679));
   NOR2_X1 i_257_76_11700 (.A1(n_257_585), .A2(n_257_76_11679), .ZN(
      n_257_76_11680));
   NOR2_X1 i_257_76_11701 (.A1(n_257_428), .A2(n_257_76_11679), .ZN(
      n_257_76_11681));
   OAI211_X1 i_257_76_11702 (.A(n_257_420), .B(n_257_76_11466), .C1(
      n_257_76_11680), .C2(n_257_76_11681), .ZN(n_257_76_11682));
   INV_X1 i_257_76_11703 (.A(n_257_76_11682), .ZN(n_257_76_11683));
   NAND3_X1 i_257_76_11704 (.A1(n_257_76_11678), .A2(n_257_76_11683), .A3(
      n_257_76_11400), .ZN(n_257_76_11684));
   INV_X1 i_257_76_11705 (.A(n_257_76_11684), .ZN(n_257_76_11685));
   NAND2_X1 i_257_76_11706 (.A1(n_257_292), .A2(n_257_423), .ZN(n_257_76_11686));
   NAND3_X1 i_257_76_11707 (.A1(n_257_76_11685), .A2(n_257_76_11686), .A3(
      n_257_76_11473), .ZN(n_257_76_11687));
   NOR2_X1 i_257_76_11708 (.A1(n_257_76_11687), .A2(n_257_76_11596), .ZN(
      n_257_76_11688));
   NAND2_X1 i_257_76_11709 (.A1(n_257_76_11432), .A2(n_257_76_11470), .ZN(
      n_257_76_11689));
   INV_X1 i_257_76_11710 (.A(n_257_76_11689), .ZN(n_257_76_11690));
   NAND2_X1 i_257_76_11711 (.A1(n_257_76_11433), .A2(n_257_76_11434), .ZN(
      n_257_76_11691));
   INV_X1 i_257_76_11712 (.A(n_257_76_11691), .ZN(n_257_76_11692));
   NAND4_X1 i_257_76_11713 (.A1(n_257_76_11690), .A2(n_257_76_11692), .A3(
      n_257_76_11424), .A4(n_257_76_11477), .ZN(n_257_76_11693));
   NOR2_X1 i_257_76_11714 (.A1(n_257_76_11693), .A2(n_257_76_11598), .ZN(
      n_257_76_11694));
   NAND3_X1 i_257_76_11715 (.A1(n_257_76_11493), .A2(n_257_76_11421), .A3(
      n_257_76_11487), .ZN(n_257_76_11695));
   INV_X1 i_257_76_11716 (.A(n_257_76_11695), .ZN(n_257_76_11696));
   NAND4_X1 i_257_76_11717 (.A1(n_257_76_11677), .A2(n_257_76_11688), .A3(
      n_257_76_11694), .A4(n_257_76_11696), .ZN(n_257_76_11697));
   NAND2_X1 i_257_76_11718 (.A1(n_257_76_11496), .A2(n_257_76_11490), .ZN(
      n_257_76_11698));
   INV_X1 i_257_76_11719 (.A(n_257_76_11698), .ZN(n_257_76_11699));
   NAND3_X1 i_257_76_11720 (.A1(n_257_76_11699), .A2(n_257_76_11482), .A3(
      n_257_76_11483), .ZN(n_257_76_11700));
   NOR2_X1 i_257_76_11721 (.A1(n_257_76_11697), .A2(n_257_76_11700), .ZN(
      n_257_76_11701));
   NAND3_X1 i_257_76_11722 (.A1(n_257_76_11701), .A2(n_257_76_11397), .A3(
      n_257_76_11500), .ZN(n_257_76_11702));
   INV_X1 i_257_76_11723 (.A(n_257_76_11702), .ZN(n_257_76_11703));
   NAND2_X1 i_257_76_11724 (.A1(n_257_76_18073), .A2(n_257_76_11703), .ZN(
      n_257_76_11704));
   NAND3_X1 i_257_76_11725 (.A1(n_257_76_11434), .A2(n_257_76_18017), .A3(
      n_257_76_11400), .ZN(n_257_76_11705));
   INV_X1 i_257_76_11726 (.A(n_257_76_11705), .ZN(n_257_76_11706));
   NAND3_X1 i_257_76_11727 (.A1(n_257_76_11706), .A2(n_257_76_11536), .A3(
      n_257_76_11477), .ZN(n_257_76_11707));
   NOR2_X1 i_257_76_11728 (.A1(n_257_76_11570), .A2(n_257_76_11707), .ZN(
      n_257_76_11708));
   INV_X1 i_257_76_11729 (.A(n_257_76_11519), .ZN(n_257_76_11709));
   NAND4_X1 i_257_76_11730 (.A1(n_257_76_11487), .A2(n_257_76_11399), .A3(
      n_257_76_11476), .A4(n_257_133), .ZN(n_257_76_11710));
   INV_X1 i_257_76_11731 (.A(n_257_76_11710), .ZN(n_257_76_11711));
   NAND4_X1 i_257_76_11732 (.A1(n_257_76_11708), .A2(n_257_76_11709), .A3(
      n_257_76_11711), .A4(n_257_76_11496), .ZN(n_257_76_11712));
   INV_X1 i_257_76_11733 (.A(n_257_76_11712), .ZN(n_257_76_11713));
   NAND3_X1 i_257_76_11734 (.A1(n_257_76_11713), .A2(n_257_76_11398), .A3(
      n_257_76_11439), .ZN(n_257_76_11714));
   NOR2_X1 i_257_76_11735 (.A1(n_257_76_11714), .A2(n_257_76_11418), .ZN(
      n_257_76_11715));
   NAND2_X1 i_257_76_11736 (.A1(n_257_76_18068), .A2(n_257_76_11715), .ZN(
      n_257_76_11716));
   NAND3_X1 i_257_76_11737 (.A1(n_257_76_11674), .A2(n_257_76_11704), .A3(
      n_257_76_11716), .ZN(n_257_76_11717));
   INV_X1 i_257_76_11738 (.A(n_257_76_11717), .ZN(n_257_76_11718));
   NAND2_X1 i_257_76_11739 (.A1(n_257_785), .A2(n_257_442), .ZN(n_257_76_11719));
   NOR2_X1 i_257_76_11740 (.A1(n_257_1079), .A2(n_257_76_11719), .ZN(
      n_257_76_11720));
   NAND4_X1 i_257_76_11741 (.A1(n_257_76_11720), .A2(n_257_447), .A3(
      n_257_76_11432), .A4(n_257_76_11433), .ZN(n_257_76_11721));
   INV_X1 i_257_76_11742 (.A(n_257_76_11721), .ZN(n_257_76_11722));
   NAND3_X1 i_257_76_11743 (.A1(n_257_76_11430), .A2(n_257_76_11722), .A3(
      n_257_76_11399), .ZN(n_257_76_11723));
   NAND2_X1 i_257_76_11744 (.A1(n_257_76_11419), .A2(n_257_76_11421), .ZN(
      n_257_76_11724));
   NOR2_X1 i_257_76_11745 (.A1(n_257_76_11723), .A2(n_257_76_11724), .ZN(
      n_257_76_11725));
   NAND2_X1 i_257_76_11746 (.A1(n_257_76_11398), .A2(n_257_76_11725), .ZN(
      n_257_76_11726));
   INV_X1 i_257_76_11747 (.A(n_257_76_11726), .ZN(n_257_76_11727));
   NAND2_X1 i_257_76_11748 (.A1(n_257_76_11397), .A2(n_257_76_11727), .ZN(
      n_257_76_11728));
   INV_X1 i_257_76_11749 (.A(n_257_76_11728), .ZN(n_257_76_11729));
   NAND3_X1 i_257_76_11750 (.A1(n_257_76_11434), .A2(n_257_76_18018), .A3(
      n_257_76_11400), .ZN(n_257_76_11730));
   NOR2_X1 i_257_76_11751 (.A1(n_257_76_11730), .A2(n_257_76_11515), .ZN(
      n_257_76_11731));
   NAND2_X1 i_257_76_11752 (.A1(n_257_76_11428), .A2(n_257_76_11423), .ZN(
      n_257_76_11732));
   INV_X1 i_257_76_11753 (.A(n_257_76_11732), .ZN(n_257_76_11733));
   INV_X1 i_257_76_11754 (.A(n_257_76_11594), .ZN(n_257_76_11734));
   NAND3_X1 i_257_76_11755 (.A1(n_257_76_11731), .A2(n_257_76_11733), .A3(
      n_257_76_11734), .ZN(n_257_76_11735));
   NAND3_X1 i_257_76_11756 (.A1(n_257_76_11399), .A2(n_257_76_11476), .A3(
      n_257_76_11427), .ZN(n_257_76_11736));
   NOR2_X1 i_257_76_11757 (.A1(n_257_76_11735), .A2(n_257_76_11736), .ZN(
      n_257_76_11737));
   NAND3_X1 i_257_76_11758 (.A1(n_257_76_11420), .A2(n_257_76_11421), .A3(
      n_257_76_11487), .ZN(n_257_76_11738));
   NAND2_X1 i_257_76_11759 (.A1(n_257_95), .A2(n_257_76_11419), .ZN(
      n_257_76_11739));
   NOR2_X1 i_257_76_11760 (.A1(n_257_76_11738), .A2(n_257_76_11739), .ZN(
      n_257_76_11740));
   NAND3_X1 i_257_76_11761 (.A1(n_257_76_11439), .A2(n_257_76_11737), .A3(
      n_257_76_11740), .ZN(n_257_76_11741));
   INV_X1 i_257_76_11762 (.A(n_257_76_11741), .ZN(n_257_76_11742));
   NAND2_X1 i_257_76_11763 (.A1(n_257_76_11742), .A2(n_257_76_11398), .ZN(
      n_257_76_11743));
   NOR2_X1 i_257_76_11764 (.A1(n_257_76_11743), .A2(n_257_76_11418), .ZN(
      n_257_76_11744));
   AOI22_X1 i_257_76_11765 (.A1(n_257_76_18085), .A2(n_257_76_11729), .B1(
      n_257_76_18080), .B2(n_257_76_11744), .ZN(n_257_76_11745));
   NAND3_X1 i_257_76_11766 (.A1(n_257_76_11664), .A2(n_257_76_11718), .A3(
      n_257_76_11745), .ZN(n_257_76_11746));
   OAI21_X1 i_257_76_11767 (.A(n_257_76_17761), .B1(n_257_721), .B2(
      n_257_76_17412), .ZN(n_257_76_11747));
   NAND4_X1 i_257_76_11768 (.A1(n_257_76_11747), .A2(n_257_76_11432), .A3(
      n_257_76_11433), .A4(n_257_76_11400), .ZN(n_257_76_11748));
   INV_X1 i_257_76_11769 (.A(n_257_76_11427), .ZN(n_257_76_11749));
   NOR2_X1 i_257_76_11770 (.A1(n_257_76_11748), .A2(n_257_76_11749), .ZN(
      n_257_76_11750));
   INV_X1 i_257_76_11771 (.A(n_257_76_11750), .ZN(n_257_76_11751));
   INV_X1 i_257_76_11772 (.A(n_257_76_11419), .ZN(n_257_76_11752));
   NOR2_X1 i_257_76_11773 (.A1(n_257_76_11751), .A2(n_257_76_11752), .ZN(
      n_257_76_11753));
   NAND3_X1 i_257_76_11774 (.A1(n_257_76_11428), .A2(n_257_76_11424), .A3(
      n_257_448), .ZN(n_257_76_11754));
   INV_X1 i_257_76_11775 (.A(n_257_76_11754), .ZN(n_257_76_11755));
   NAND4_X1 i_257_76_11776 (.A1(n_257_76_11755), .A2(n_257_76_11420), .A3(
      n_257_76_11421), .A4(n_257_76_11399), .ZN(n_257_76_11756));
   INV_X1 i_257_76_11777 (.A(n_257_76_11756), .ZN(n_257_76_11757));
   NAND3_X1 i_257_76_11778 (.A1(n_257_76_11753), .A2(n_257_689), .A3(
      n_257_76_11757), .ZN(n_257_76_11758));
   INV_X1 i_257_76_11779 (.A(n_257_76_11758), .ZN(n_257_76_11759));
   NAND2_X1 i_257_76_11780 (.A1(n_257_76_11759), .A2(n_257_76_11398), .ZN(
      n_257_76_11760));
   NOR2_X1 i_257_76_11781 (.A1(n_257_76_11418), .A2(n_257_76_11760), .ZN(
      n_257_76_11761));
   NAND2_X1 i_257_76_11782 (.A1(n_257_76_18079), .A2(n_257_76_11761), .ZN(
      n_257_76_11762));
   INV_X1 i_257_76_11783 (.A(n_257_76_18016), .ZN(n_257_76_11763));
   NOR2_X1 i_257_76_11784 (.A1(n_257_1079), .A2(n_257_76_11763), .ZN(
      n_257_76_11764));
   NAND2_X1 i_257_76_11785 (.A1(n_257_76_11466), .A2(n_257_425), .ZN(
      n_257_76_11765));
   INV_X1 i_257_76_11786 (.A(n_257_76_11765), .ZN(n_257_76_11766));
   NAND4_X1 i_257_76_11787 (.A1(n_257_76_11764), .A2(n_257_76_11433), .A3(
      n_257_76_11434), .A4(n_257_76_11766), .ZN(n_257_76_11767));
   NAND3_X1 i_257_76_11788 (.A1(n_257_76_11477), .A2(n_257_76_11432), .A3(
      n_257_76_11470), .ZN(n_257_76_11768));
   NOR2_X1 i_257_76_11789 (.A1(n_257_76_11767), .A2(n_257_76_11768), .ZN(
      n_257_76_11769));
   INV_X1 i_257_76_11790 (.A(n_257_76_11570), .ZN(n_257_76_11770));
   NAND3_X1 i_257_76_11791 (.A1(n_257_76_11769), .A2(n_257_76_11597), .A3(
      n_257_76_11770), .ZN(n_257_76_11771));
   NAND4_X1 i_257_76_11792 (.A1(n_257_76_11420), .A2(n_257_76_11493), .A3(
      n_257_76_11421), .A4(n_257_76_11487), .ZN(n_257_76_11772));
   NOR2_X1 i_257_76_11793 (.A1(n_257_76_11771), .A2(n_257_76_11772), .ZN(
      n_257_76_11773));
   NAND3_X1 i_257_76_11794 (.A1(n_257_76_11492), .A2(n_257_252), .A3(
      n_257_76_11496), .ZN(n_257_76_11774));
   INV_X1 i_257_76_11795 (.A(n_257_76_11774), .ZN(n_257_76_11775));
   NAND4_X1 i_257_76_11796 (.A1(n_257_76_11773), .A2(n_257_76_11775), .A3(
      n_257_76_11439), .A4(n_257_76_11482), .ZN(n_257_76_11776));
   NAND2_X1 i_257_76_11797 (.A1(n_257_76_11397), .A2(n_257_76_11398), .ZN(
      n_257_76_11777));
   NOR2_X1 i_257_76_11798 (.A1(n_257_76_11776), .A2(n_257_76_11777), .ZN(
      n_257_76_11778));
   NAND2_X1 i_257_76_11799 (.A1(n_257_76_18064), .A2(n_257_76_11778), .ZN(
      n_257_76_11779));
   NAND4_X1 i_257_76_11800 (.A1(n_257_369), .A2(n_257_76_11686), .A3(
      n_257_76_11473), .A4(n_257_76_11427), .ZN(n_257_76_11780));
   NAND3_X1 i_257_76_11801 (.A1(n_257_76_18016), .A2(n_257_76_11466), .A3(
      n_257_421), .ZN(n_257_76_11781));
   INV_X1 i_257_76_11802 (.A(n_257_76_11781), .ZN(n_257_76_11782));
   NAND3_X1 i_257_76_11803 (.A1(n_257_76_11782), .A2(n_257_76_11434), .A3(
      n_257_76_11400), .ZN(n_257_76_11783));
   INV_X1 i_257_76_11804 (.A(n_257_76_11783), .ZN(n_257_76_11784));
   NAND2_X1 i_257_76_11805 (.A1(n_257_76_11678), .A2(n_257_76_11432), .ZN(
      n_257_76_11785));
   INV_X1 i_257_76_11806 (.A(n_257_76_11785), .ZN(n_257_76_11786));
   INV_X1 i_257_76_11807 (.A(n_257_76_11471), .ZN(n_257_76_11787));
   NAND3_X1 i_257_76_11808 (.A1(n_257_76_11784), .A2(n_257_76_11786), .A3(
      n_257_76_11787), .ZN(n_257_76_11788));
   NAND4_X1 i_257_76_11809 (.A1(n_257_76_11428), .A2(n_257_76_11423), .A3(
      n_257_76_11424), .A4(n_257_76_11477), .ZN(n_257_76_11789));
   NOR3_X1 i_257_76_11810 (.A1(n_257_76_11780), .A2(n_257_76_11788), .A3(
      n_257_76_11789), .ZN(n_257_76_11790));
   INV_X1 i_257_76_11811 (.A(n_257_76_11496), .ZN(n_257_76_11791));
   NOR2_X1 i_257_76_11812 (.A1(n_257_76_11791), .A2(n_257_76_11491), .ZN(
      n_257_76_11792));
   NAND3_X1 i_257_76_11813 (.A1(n_257_76_11487), .A2(n_257_76_11399), .A3(
      n_257_76_11476), .ZN(n_257_76_11793));
   NOR2_X1 i_257_76_11814 (.A1(n_257_76_11494), .A2(n_257_76_11793), .ZN(
      n_257_76_11794));
   NAND3_X1 i_257_76_11815 (.A1(n_257_76_11790), .A2(n_257_76_11792), .A3(
      n_257_76_11794), .ZN(n_257_76_11795));
   INV_X1 i_257_76_11816 (.A(n_257_76_11795), .ZN(n_257_76_11796));
   NAND3_X1 i_257_76_11817 (.A1(n_257_76_11439), .A2(n_257_76_11482), .A3(
      n_257_76_11483), .ZN(n_257_76_11797));
   INV_X1 i_257_76_11818 (.A(n_257_76_11398), .ZN(n_257_76_11798));
   NOR2_X1 i_257_76_11819 (.A1(n_257_76_11797), .A2(n_257_76_11798), .ZN(
      n_257_76_11799));
   NAND3_X1 i_257_76_11820 (.A1(n_257_76_11397), .A2(n_257_76_11796), .A3(
      n_257_76_11799), .ZN(n_257_76_11800));
   INV_X1 i_257_76_11821 (.A(n_257_76_11800), .ZN(n_257_76_11801));
   NAND2_X1 i_257_76_11822 (.A1(n_257_76_18082), .A2(n_257_76_11801), .ZN(
      n_257_76_11802));
   NAND3_X1 i_257_76_11823 (.A1(n_257_76_11762), .A2(n_257_76_11779), .A3(
      n_257_76_11802), .ZN(n_257_76_11803));
   INV_X1 i_257_76_11824 (.A(n_257_76_11803), .ZN(n_257_76_11804));
   NAND2_X1 i_257_76_11825 (.A1(n_257_427), .A2(n_257_76_11466), .ZN(
      n_257_76_11805));
   INV_X1 i_257_76_11826 (.A(n_257_76_11805), .ZN(n_257_76_11806));
   NAND4_X1 i_257_76_11827 (.A1(n_257_76_11806), .A2(n_257_76_11400), .A3(
      n_257_212), .A4(n_257_76_18016), .ZN(n_257_76_11807));
   INV_X1 i_257_76_11828 (.A(n_257_76_11807), .ZN(n_257_76_11808));
   NAND4_X1 i_257_76_11829 (.A1(n_257_76_11476), .A2(n_257_76_11808), .A3(
      n_257_76_11427), .A4(n_257_76_11428), .ZN(n_257_76_11809));
   NAND3_X1 i_257_76_11830 (.A1(n_257_76_11432), .A2(n_257_76_11433), .A3(
      n_257_76_11434), .ZN(n_257_76_11810));
   INV_X1 i_257_76_11831 (.A(n_257_76_11810), .ZN(n_257_76_11811));
   NAND4_X1 i_257_76_11832 (.A1(n_257_76_11811), .A2(n_257_76_11423), .A3(
      n_257_76_11424), .A4(n_257_76_11477), .ZN(n_257_76_11812));
   NOR2_X1 i_257_76_11833 (.A1(n_257_76_11809), .A2(n_257_76_11812), .ZN(
      n_257_76_11813));
   NAND4_X1 i_257_76_11834 (.A1(n_257_76_11528), .A2(n_257_76_11813), .A3(
      n_257_76_11482), .A4(n_257_76_11496), .ZN(n_257_76_11814));
   INV_X1 i_257_76_11835 (.A(n_257_76_11814), .ZN(n_257_76_11815));
   NAND3_X1 i_257_76_11836 (.A1(n_257_76_11397), .A2(n_257_76_11815), .A3(
      n_257_76_11500), .ZN(n_257_76_11816));
   INV_X1 i_257_76_11837 (.A(n_257_76_11816), .ZN(n_257_76_11817));
   NAND2_X1 i_257_76_11838 (.A1(n_257_76_18065), .A2(n_257_76_11817), .ZN(
      n_257_76_11818));
   NAND4_X1 i_257_76_11839 (.A1(n_257_76_11750), .A2(n_257_76_11419), .A3(
      n_257_76_11420), .A4(n_257_76_11421), .ZN(n_257_76_11819));
   NAND3_X1 i_257_76_11840 (.A1(n_257_76_11423), .A2(n_257_472), .A3(
      n_257_76_11424), .ZN(n_257_76_11820));
   INV_X1 i_257_76_11841 (.A(n_257_76_11820), .ZN(n_257_76_11821));
   NAND2_X1 i_257_76_11842 (.A1(n_257_451), .A2(n_257_76_11428), .ZN(
      n_257_76_11822));
   INV_X1 i_257_76_11843 (.A(n_257_76_11822), .ZN(n_257_76_11823));
   NAND4_X1 i_257_76_11844 (.A1(n_257_76_11821), .A2(n_257_76_11823), .A3(
      n_257_76_11399), .A4(n_257_76_11476), .ZN(n_257_76_11824));
   NOR2_X1 i_257_76_11845 (.A1(n_257_76_11819), .A2(n_257_76_11824), .ZN(
      n_257_76_11825));
   NAND3_X1 i_257_76_11846 (.A1(n_257_76_11825), .A2(n_257_76_11398), .A3(
      n_257_76_11439), .ZN(n_257_76_11826));
   NOR2_X1 i_257_76_11847 (.A1(n_257_76_11826), .A2(n_257_76_11418), .ZN(
      n_257_76_11827));
   NAND2_X1 i_257_76_11848 (.A1(n_257_76_18063), .A2(n_257_76_11827), .ZN(
      n_257_76_11828));
   NAND2_X1 i_257_76_11849 (.A1(n_257_76_11427), .A2(n_257_76_11477), .ZN(
      n_257_76_11829));
   INV_X1 i_257_76_11850 (.A(n_257_76_11829), .ZN(n_257_76_11830));
   NAND2_X1 i_257_76_11851 (.A1(n_257_76_11466), .A2(n_257_424), .ZN(
      n_257_76_11831));
   INV_X1 i_257_76_11852 (.A(n_257_76_11831), .ZN(n_257_76_11832));
   NAND3_X1 i_257_76_11853 (.A1(n_257_76_11400), .A2(n_257_76_18016), .A3(
      n_257_76_11832), .ZN(n_257_76_11833));
   NOR2_X1 i_257_76_11854 (.A1(n_257_76_11691), .A2(n_257_76_11833), .ZN(
      n_257_76_11834));
   NAND3_X1 i_257_76_11855 (.A1(n_257_521), .A2(n_257_76_11432), .A3(
      n_257_76_11470), .ZN(n_257_76_11835));
   INV_X1 i_257_76_11856 (.A(n_257_76_11835), .ZN(n_257_76_11836));
   NAND4_X1 i_257_76_11857 (.A1(n_257_76_11830), .A2(n_257_76_11834), .A3(
      n_257_76_11476), .A4(n_257_76_11836), .ZN(n_257_76_11837));
   INV_X1 i_257_76_11858 (.A(n_257_76_11837), .ZN(n_257_76_11838));
   NAND3_X1 i_257_76_11859 (.A1(n_257_76_11482), .A2(n_257_76_11483), .A3(
      n_257_76_11838), .ZN(n_257_76_11839));
   NOR2_X1 i_257_76_11860 (.A1(n_257_76_11839), .A2(n_257_76_11497), .ZN(
      n_257_76_11840));
   NAND3_X1 i_257_76_11861 (.A1(n_257_76_11840), .A2(n_257_76_11397), .A3(
      n_257_76_11500), .ZN(n_257_76_11841));
   INV_X1 i_257_76_11862 (.A(n_257_76_11841), .ZN(n_257_76_11842));
   NAND2_X1 i_257_76_11863 (.A1(n_257_76_18062), .A2(n_257_76_11842), .ZN(
      n_257_76_11843));
   NAND3_X1 i_257_76_11864 (.A1(n_257_76_11818), .A2(n_257_76_11828), .A3(
      n_257_76_11843), .ZN(n_257_76_11844));
   INV_X1 i_257_76_11865 (.A(n_257_76_11844), .ZN(n_257_76_11845));
   NAND3_X1 i_257_76_11866 (.A1(n_257_76_11490), .A2(n_257_76_11419), .A3(
      n_257_76_11420), .ZN(n_257_76_11846));
   INV_X1 i_257_76_11867 (.A(n_257_76_11846), .ZN(n_257_76_11847));
   NAND2_X1 i_257_76_11868 (.A1(n_257_76_11466), .A2(n_257_422), .ZN(
      n_257_76_11848));
   INV_X1 i_257_76_11869 (.A(n_257_76_11848), .ZN(n_257_76_11849));
   NAND4_X1 i_257_76_11870 (.A1(n_257_76_11400), .A2(n_257_76_11849), .A3(
      n_257_330), .A4(n_257_76_18016), .ZN(n_257_76_11850));
   INV_X1 i_257_76_11871 (.A(n_257_76_11850), .ZN(n_257_76_11851));
   NAND3_X1 i_257_76_11872 (.A1(n_257_76_11686), .A2(n_257_76_11851), .A3(
      n_257_76_11473), .ZN(n_257_76_11852));
   NOR2_X1 i_257_76_11873 (.A1(n_257_76_11596), .A2(n_257_76_11852), .ZN(
      n_257_76_11853));
   NAND4_X1 i_257_76_11874 (.A1(n_257_76_11847), .A2(n_257_76_11853), .A3(
      n_257_76_11694), .A4(n_257_76_11696), .ZN(n_257_76_11854));
   NAND3_X1 i_257_76_11875 (.A1(n_257_76_11482), .A2(n_257_76_11483), .A3(
      n_257_76_11496), .ZN(n_257_76_11855));
   NOR2_X1 i_257_76_11876 (.A1(n_257_76_11854), .A2(n_257_76_11855), .ZN(
      n_257_76_11856));
   NAND3_X1 i_257_76_11877 (.A1(n_257_76_11856), .A2(n_257_76_11397), .A3(
      n_257_76_11500), .ZN(n_257_76_11857));
   INV_X1 i_257_76_11878 (.A(n_257_76_11857), .ZN(n_257_76_11858));
   NAND2_X1 i_257_76_11879 (.A1(n_257_342), .A2(n_257_76_11858), .ZN(
      n_257_76_11859));
   NAND2_X1 i_257_76_11880 (.A1(n_257_420), .A2(n_257_489), .ZN(n_257_76_11860));
   NAND2_X1 i_257_76_11881 (.A1(n_257_585), .A2(n_257_428), .ZN(n_257_76_11861));
   NAND3_X1 i_257_76_11882 (.A1(n_257_408), .A2(n_257_484), .A3(n_257_442), 
      .ZN(n_257_76_11862));
   INV_X1 i_257_76_11883 (.A(n_257_76_11862), .ZN(n_257_76_11863));
   NAND2_X1 i_257_76_11884 (.A1(n_257_76_11861), .A2(n_257_76_11863), .ZN(
      n_257_76_11864));
   INV_X1 i_257_76_11885 (.A(n_257_76_11864), .ZN(n_257_76_11865));
   NAND3_X1 i_257_76_11886 (.A1(n_257_76_11860), .A2(n_257_76_11865), .A3(
      n_257_76_11466), .ZN(n_257_76_11866));
   INV_X1 i_257_76_11887 (.A(n_257_76_11866), .ZN(n_257_76_11867));
   NAND4_X1 i_257_76_11888 (.A1(n_257_76_11867), .A2(n_257_76_11433), .A3(
      n_257_76_11434), .A4(n_257_76_11400), .ZN(n_257_76_11868));
   INV_X1 i_257_76_11889 (.A(n_257_76_11868), .ZN(n_257_76_11869));
   NAND3_X1 i_257_76_11890 (.A1(n_257_76_11678), .A2(n_257_76_11432), .A3(
      n_257_76_11470), .ZN(n_257_76_11870));
   INV_X1 i_257_76_11891 (.A(n_257_76_11870), .ZN(n_257_76_11871));
   NAND2_X1 i_257_76_11892 (.A1(n_257_76_11869), .A2(n_257_76_11871), .ZN(
      n_257_76_11872));
   NAND3_X1 i_257_76_11893 (.A1(n_257_76_11473), .A2(n_257_76_11427), .A3(
      n_257_76_11428), .ZN(n_257_76_11873));
   NOR3_X1 i_257_76_11894 (.A1(n_257_76_11872), .A2(n_257_76_11873), .A3(
      n_257_76_11648), .ZN(n_257_76_11874));
   NAND2_X1 i_257_76_11895 (.A1(n_257_76_11439), .A2(n_257_76_11874), .ZN(
      n_257_76_11875));
   NOR2_X1 i_257_76_11896 (.A1(n_257_76_11875), .A2(n_257_76_11798), .ZN(
      n_257_76_11876));
   NAND3_X1 i_257_76_11897 (.A1(n_257_76_11490), .A2(n_257_76_11675), .A3(
      n_257_76_11419), .ZN(n_257_76_11877));
   INV_X1 i_257_76_11898 (.A(n_257_76_11877), .ZN(n_257_76_11878));
   NAND4_X1 i_257_76_11899 (.A1(n_257_76_11487), .A2(n_257_76_11399), .A3(
      n_257_76_11476), .A4(n_257_76_11686), .ZN(n_257_76_11879));
   INV_X1 i_257_76_11900 (.A(n_257_76_11879), .ZN(n_257_76_11880));
   NAND4_X1 i_257_76_11901 (.A1(n_257_76_11878), .A2(n_257_76_11880), .A3(
      n_257_76_11495), .A4(n_257_76_11496), .ZN(n_257_76_11881));
   NAND2_X1 i_257_76_11902 (.A1(n_257_76_11482), .A2(n_257_76_11483), .ZN(
      n_257_76_11882));
   NOR2_X1 i_257_76_11903 (.A1(n_257_76_11881), .A2(n_257_76_11882), .ZN(
      n_257_76_11883));
   NAND3_X1 i_257_76_11904 (.A1(n_257_76_11876), .A2(n_257_76_11397), .A3(
      n_257_76_11883), .ZN(n_257_76_11884));
   INV_X1 i_257_76_11905 (.A(n_257_76_11884), .ZN(n_257_76_11885));
   NAND2_X1 i_257_76_11906 (.A1(n_257_76_18060), .A2(n_257_76_11885), .ZN(
      n_257_76_11886));
   NAND2_X1 i_257_76_11907 (.A1(n_257_817), .A2(n_257_76_17952), .ZN(
      n_257_76_11887));
   NAND3_X1 i_257_76_11908 (.A1(n_257_441), .A2(n_257_983), .A3(n_257_442), 
      .ZN(n_257_76_11888));
   NAND2_X1 i_257_76_11909 (.A1(n_257_649), .A2(n_257_76_17928), .ZN(
      n_257_76_11889));
   NAND3_X1 i_257_76_11910 (.A1(n_257_76_11887), .A2(n_257_76_11888), .A3(
      n_257_76_11889), .ZN(n_257_76_11890));
   INV_X1 i_257_76_11911 (.A(n_257_76_11890), .ZN(n_257_76_11891));
   NAND2_X1 i_257_76_11912 (.A1(n_257_449), .A2(n_257_76_16220), .ZN(
      n_257_76_11892));
   INV_X1 i_257_76_11913 (.A(n_257_76_11719), .ZN(n_257_76_11893));
   NAND2_X1 i_257_76_11914 (.A1(n_257_447), .A2(n_257_76_11893), .ZN(
      n_257_76_11894));
   NAND3_X1 i_257_76_11915 (.A1(n_257_76_11892), .A2(n_257_76_11850), .A3(
      n_257_76_11894), .ZN(n_257_76_11895));
   NAND2_X1 i_257_76_11916 (.A1(n_257_55), .A2(n_257_76_17918), .ZN(
      n_257_76_11896));
   NAND3_X1 i_257_76_11917 (.A1(n_257_438), .A2(n_257_1085), .A3(n_257_442), 
      .ZN(n_257_76_11897));
   NAND2_X1 i_257_76_11918 (.A1(n_257_440), .A2(n_257_76_11402), .ZN(
      n_257_76_11898));
   NAND2_X1 i_257_76_11919 (.A1(n_257_721), .A2(n_257_76_15655), .ZN(
      n_257_76_11899));
   NAND4_X1 i_257_76_11920 (.A1(n_257_76_11896), .A2(n_257_76_11897), .A3(
      n_257_76_11898), .A4(n_257_76_11899), .ZN(n_257_76_11900));
   NOR2_X1 i_257_76_11921 (.A1(n_257_76_11895), .A2(n_257_76_11900), .ZN(
      n_257_76_11901));
   AOI22_X1 i_257_76_11922 (.A1(n_257_753), .A2(n_257_76_17935), .B1(n_257_133), 
      .B2(n_257_76_17925), .ZN(n_257_76_11902));
   NAND2_X1 i_257_76_11923 (.A1(n_257_881), .A2(n_257_76_17903), .ZN(
      n_257_76_11903));
   INV_X1 i_257_76_11924 (.A(n_257_76_11446), .ZN(n_257_76_11904));
   NAND2_X1 i_257_76_11925 (.A1(n_257_446), .A2(n_257_76_11904), .ZN(
      n_257_76_11905));
   NAND2_X1 i_257_76_11926 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[20]), 
      .ZN(n_257_76_11906));
   INV_X1 i_257_76_11927 (.A(Small_Packet_Data_Size[20]), .ZN(n_257_76_11907));
   NAND3_X1 i_257_76_11928 (.A1(n_257_76_11466), .A2(n_257_76_18019), .A3(
      n_257_76_11861), .ZN(n_257_76_11908));
   OAI21_X1 i_257_76_11929 (.A(n_257_76_11906), .B1(n_257_1079), .B2(
      n_257_76_11908), .ZN(n_257_76_11909));
   NAND3_X1 i_257_76_11930 (.A1(n_257_76_11903), .A2(n_257_76_11905), .A3(
      n_257_76_11909), .ZN(n_257_76_11910));
   NAND2_X1 i_257_76_11931 (.A1(n_257_76_11684), .A2(n_257_76_11807), .ZN(
      n_257_76_11911));
   NOR2_X1 i_257_76_11932 (.A1(n_257_76_11910), .A2(n_257_76_11911), .ZN(
      n_257_76_11912));
   NAND4_X1 i_257_76_11933 (.A1(n_257_76_11891), .A2(n_257_76_11901), .A3(
      n_257_76_11902), .A4(n_257_76_11912), .ZN(n_257_76_11913));
   INV_X1 i_257_76_11934 (.A(n_257_76_11913), .ZN(n_257_76_11914));
   INV_X1 i_257_76_11935 (.A(n_257_172), .ZN(n_257_76_11915));
   OAI21_X1 i_257_76_11936 (.A(n_257_76_11480), .B1(n_257_76_11915), .B2(
      n_257_76_17660), .ZN(n_257_76_11916));
   INV_X1 i_257_76_11937 (.A(n_257_76_11916), .ZN(n_257_76_11917));
   INV_X1 i_257_76_11938 (.A(n_257_445), .ZN(n_257_76_11918));
   NAND2_X1 i_257_76_11939 (.A1(n_257_76_11918), .A2(n_257_442), .ZN(
      n_257_76_11919));
   OAI21_X1 i_257_76_11940 (.A(n_257_76_11919), .B1(n_257_881), .B2(
      n_257_76_17412), .ZN(n_257_76_11920));
   NAND3_X1 i_257_76_11941 (.A1(n_257_76_11920), .A2(n_257_451), .A3(n_257_472), 
      .ZN(n_257_76_11921));
   NAND2_X1 i_257_76_11942 (.A1(n_257_919), .A2(n_257_76_17940), .ZN(
      n_257_76_11922));
   NAND2_X1 i_257_76_11943 (.A1(n_257_76_11921), .A2(n_257_76_11922), .ZN(
      n_257_76_11923));
   INV_X1 i_257_76_11944 (.A(n_257_76_11923), .ZN(n_257_76_11924));
   NAND2_X1 i_257_76_11945 (.A1(n_257_95), .A2(n_257_76_17932), .ZN(
      n_257_76_11925));
   NAND3_X1 i_257_76_11946 (.A1(n_257_76_11924), .A2(n_257_76_11837), .A3(
      n_257_76_11925), .ZN(n_257_76_11926));
   INV_X1 i_257_76_11947 (.A(n_257_76_11926), .ZN(n_257_76_11927));
   NAND3_X1 i_257_76_11948 (.A1(n_257_76_11914), .A2(n_257_76_11917), .A3(
      n_257_76_11927), .ZN(n_257_76_11928));
   NAND2_X1 i_257_76_11949 (.A1(n_257_1015), .A2(n_257_76_17964), .ZN(
      n_257_76_11929));
   NAND2_X1 i_257_76_11950 (.A1(n_257_689), .A2(n_257_76_17958), .ZN(
      n_257_76_11930));
   NAND3_X1 i_257_76_11951 (.A1(n_257_76_11929), .A2(n_257_76_11573), .A3(
      n_257_76_11930), .ZN(n_257_76_11931));
   NOR2_X1 i_257_76_11952 (.A1(n_257_76_11928), .A2(n_257_76_11931), .ZN(
      n_257_76_11932));
   INV_X1 i_257_76_11953 (.A(n_257_1047), .ZN(n_257_76_11933));
   OAI21_X1 i_257_76_11954 (.A(n_257_76_11795), .B1(n_257_76_11933), .B2(
      n_257_76_17968), .ZN(n_257_76_11934));
   INV_X1 i_257_76_11955 (.A(n_257_76_11934), .ZN(n_257_76_11935));
   NAND3_X1 i_257_76_11956 (.A1(n_257_76_11932), .A2(n_257_76_11935), .A3(
      n_257_76_11776), .ZN(n_257_76_11936));
   NAND3_X1 i_257_76_11957 (.A1(n_257_76_11859), .A2(n_257_76_11886), .A3(
      n_257_76_11936), .ZN(n_257_76_11937));
   INV_X1 i_257_76_11958 (.A(n_257_76_11937), .ZN(n_257_76_11938));
   NAND3_X1 i_257_76_11959 (.A1(n_257_76_11804), .A2(n_257_76_11845), .A3(
      n_257_76_11938), .ZN(n_257_76_11939));
   NOR2_X1 i_257_76_11960 (.A1(n_257_76_11746), .A2(n_257_76_11939), .ZN(
      n_257_76_11940));
   NAND2_X1 i_257_76_11961 (.A1(n_257_76_11628), .A2(n_257_76_11940), .ZN(n_20));
   NAND2_X1 i_257_76_11962 (.A1(n_257_1048), .A2(n_257_443), .ZN(n_257_76_11941));
   INV_X1 i_257_76_11963 (.A(n_257_76_11941), .ZN(n_257_76_11942));
   NAND2_X1 i_257_76_11964 (.A1(n_257_1016), .A2(n_257_444), .ZN(n_257_76_11943));
   NAND2_X1 i_257_76_11965 (.A1(n_257_441), .A2(n_257_984), .ZN(n_257_76_11944));
   NAND2_X1 i_257_76_11966 (.A1(n_257_952), .A2(n_257_442), .ZN(n_257_76_11945));
   INV_X1 i_257_76_11967 (.A(n_257_76_11945), .ZN(n_257_76_11946));
   NAND2_X1 i_257_76_11968 (.A1(n_257_440), .A2(n_257_76_11946), .ZN(
      n_257_76_11947));
   NOR2_X1 i_257_76_11969 (.A1(n_257_76_11947), .A2(n_257_1080), .ZN(
      n_257_76_11948));
   NAND2_X1 i_257_76_11970 (.A1(n_257_76_11944), .A2(n_257_76_11948), .ZN(
      n_257_76_11949));
   INV_X1 i_257_76_11971 (.A(n_257_76_11949), .ZN(n_257_76_11950));
   NAND2_X1 i_257_76_11972 (.A1(n_257_76_11943), .A2(n_257_76_11950), .ZN(
      n_257_76_11951));
   NOR2_X1 i_257_76_11973 (.A1(n_257_76_11942), .A2(n_257_76_11951), .ZN(
      n_257_76_11952));
   NAND2_X1 i_257_76_11974 (.A1(n_257_17), .A2(n_257_76_11952), .ZN(
      n_257_76_11953));
   NOR2_X1 i_257_76_11975 (.A1(n_257_1080), .A2(n_257_76_17412), .ZN(
      n_257_76_11954));
   INV_X1 i_257_76_11976 (.A(n_257_76_11954), .ZN(n_257_76_11955));
   NOR2_X1 i_257_76_11977 (.A1(n_257_76_11955), .A2(n_257_76_15197), .ZN(
      n_257_76_11956));
   NAND2_X1 i_257_76_11978 (.A1(n_257_1048), .A2(n_257_76_11956), .ZN(
      n_257_76_11957));
   INV_X1 i_257_76_11979 (.A(n_257_76_11957), .ZN(n_257_76_11958));
   NAND2_X1 i_257_76_11980 (.A1(n_257_76_18072), .A2(n_257_76_11958), .ZN(
      n_257_76_11959));
   NAND2_X1 i_257_76_11981 (.A1(n_257_690), .A2(n_257_448), .ZN(n_257_76_11960));
   NAND2_X1 i_257_76_11982 (.A1(n_257_882), .A2(n_257_445), .ZN(n_257_76_11961));
   NAND2_X1 i_257_76_11983 (.A1(n_257_650), .A2(n_257_76_11961), .ZN(
      n_257_76_11962));
   INV_X1 i_257_76_11984 (.A(n_257_76_11962), .ZN(n_257_76_11963));
   NAND2_X1 i_257_76_11985 (.A1(n_257_446), .A2(n_257_850), .ZN(n_257_76_11964));
   NAND2_X1 i_257_76_11986 (.A1(n_257_449), .A2(n_257_896), .ZN(n_257_76_11965));
   NAND2_X1 i_257_76_11987 (.A1(n_257_447), .A2(n_257_786), .ZN(n_257_76_11966));
   NAND3_X1 i_257_76_11988 (.A1(n_257_76_11964), .A2(n_257_76_11965), .A3(
      n_257_76_11966), .ZN(n_257_76_11967));
   INV_X1 i_257_76_11989 (.A(n_257_76_11967), .ZN(n_257_76_11968));
   NOR2_X1 i_257_76_11990 (.A1(n_257_1080), .A2(n_257_76_17927), .ZN(
      n_257_76_11969));
   NAND2_X1 i_257_76_11991 (.A1(n_257_722), .A2(n_257_435), .ZN(n_257_76_11970));
   NAND2_X1 i_257_76_11992 (.A1(n_257_438), .A2(n_257_1086), .ZN(n_257_76_11971));
   NAND2_X1 i_257_76_11993 (.A1(n_257_440), .A2(n_257_952), .ZN(n_257_76_11972));
   NAND4_X1 i_257_76_11994 (.A1(n_257_76_11969), .A2(n_257_76_11970), .A3(
      n_257_76_11971), .A4(n_257_76_11972), .ZN(n_257_76_11973));
   INV_X1 i_257_76_11995 (.A(n_257_76_11973), .ZN(n_257_76_11974));
   NAND4_X1 i_257_76_11996 (.A1(n_257_76_11963), .A2(n_257_76_11968), .A3(
      n_257_76_11974), .A4(n_257_76_11944), .ZN(n_257_76_11975));
   NAND2_X1 i_257_76_11997 (.A1(n_257_754), .A2(n_257_436), .ZN(n_257_76_11976));
   NAND2_X1 i_257_76_11998 (.A1(n_257_818), .A2(n_257_437), .ZN(n_257_76_11977));
   NAND2_X1 i_257_76_11999 (.A1(n_257_920), .A2(n_257_439), .ZN(n_257_76_11978));
   NAND3_X1 i_257_76_12000 (.A1(n_257_76_11976), .A2(n_257_76_11977), .A3(
      n_257_76_11978), .ZN(n_257_76_11979));
   NOR2_X1 i_257_76_12001 (.A1(n_257_76_11975), .A2(n_257_76_11979), .ZN(
      n_257_76_11980));
   NAND2_X1 i_257_76_12002 (.A1(n_257_76_11960), .A2(n_257_76_11980), .ZN(
      n_257_76_11981));
   INV_X1 i_257_76_12003 (.A(n_257_76_11981), .ZN(n_257_76_11982));
   NAND3_X1 i_257_76_12004 (.A1(n_257_76_11982), .A2(n_257_76_11941), .A3(
      n_257_76_11943), .ZN(n_257_76_11983));
   INV_X1 i_257_76_12005 (.A(n_257_76_11983), .ZN(n_257_76_11984));
   NAND2_X1 i_257_76_12006 (.A1(n_257_28), .A2(n_257_76_11984), .ZN(
      n_257_76_11985));
   NAND3_X1 i_257_76_12007 (.A1(n_257_76_11953), .A2(n_257_76_11959), .A3(
      n_257_76_11985), .ZN(n_257_76_11986));
   NAND2_X1 i_257_76_12008 (.A1(n_257_850), .A2(n_257_442), .ZN(n_257_76_11987));
   NOR2_X1 i_257_76_12009 (.A1(n_257_1080), .A2(n_257_76_11987), .ZN(
      n_257_76_11988));
   NAND4_X1 i_257_76_12010 (.A1(n_257_76_11988), .A2(n_257_446), .A3(
      n_257_76_11971), .A4(n_257_76_11972), .ZN(n_257_76_11989));
   INV_X1 i_257_76_12011 (.A(n_257_76_11989), .ZN(n_257_76_11990));
   NAND3_X1 i_257_76_12012 (.A1(n_257_76_11990), .A2(n_257_76_11944), .A3(
      n_257_76_11961), .ZN(n_257_76_11991));
   INV_X1 i_257_76_12013 (.A(n_257_76_11978), .ZN(n_257_76_11992));
   NOR2_X1 i_257_76_12014 (.A1(n_257_76_11991), .A2(n_257_76_11992), .ZN(
      n_257_76_11993));
   NAND2_X1 i_257_76_12015 (.A1(n_257_76_11943), .A2(n_257_76_11993), .ZN(
      n_257_76_11994));
   NOR2_X1 i_257_76_12016 (.A1(n_257_76_11942), .A2(n_257_76_11994), .ZN(
      n_257_76_11995));
   NAND2_X1 i_257_76_12017 (.A1(n_257_76_18070), .A2(n_257_76_11995), .ZN(
      n_257_76_11996));
   NAND3_X1 i_257_76_12018 (.A1(n_257_76_11954), .A2(n_257_76_11972), .A3(
      n_257_439), .ZN(n_257_76_11997));
   INV_X1 i_257_76_12019 (.A(n_257_76_11997), .ZN(n_257_76_11998));
   NAND3_X1 i_257_76_12020 (.A1(n_257_76_11998), .A2(n_257_76_11944), .A3(
      n_257_920), .ZN(n_257_76_11999));
   INV_X1 i_257_76_12021 (.A(n_257_76_11999), .ZN(n_257_76_12000));
   NAND2_X1 i_257_76_12022 (.A1(n_257_76_11943), .A2(n_257_76_12000), .ZN(
      n_257_76_12001));
   NOR2_X1 i_257_76_12023 (.A1(n_257_76_11942), .A2(n_257_76_12001), .ZN(
      n_257_76_12002));
   NAND2_X1 i_257_76_12024 (.A1(n_257_76_18084), .A2(n_257_76_12002), .ZN(
      n_257_76_12003));
   NAND2_X1 i_257_76_12025 (.A1(n_257_554), .A2(n_257_426), .ZN(n_257_76_12004));
   NAND2_X1 i_257_76_12026 (.A1(n_257_134), .A2(n_257_430), .ZN(n_257_76_12005));
   NAND4_X1 i_257_76_12027 (.A1(n_257_76_12004), .A2(n_257_76_11976), .A3(
      n_257_76_11977), .A4(n_257_76_12005), .ZN(n_257_76_12006));
   INV_X1 i_257_76_12028 (.A(n_257_76_12006), .ZN(n_257_76_12007));
   NAND2_X1 i_257_76_12029 (.A1(n_257_650), .A2(n_257_450), .ZN(n_257_76_12008));
   NAND3_X1 i_257_76_12030 (.A1(n_257_76_11968), .A2(n_257_76_12008), .A3(
      n_257_76_11944), .ZN(n_257_76_12009));
   NAND2_X1 i_257_76_12031 (.A1(n_257_451), .A2(n_257_473), .ZN(n_257_76_12010));
   NAND2_X1 i_257_76_12032 (.A1(n_257_76_11978), .A2(n_257_76_12010), .ZN(
      n_257_76_12011));
   NOR2_X1 i_257_76_12033 (.A1(n_257_76_12009), .A2(n_257_76_12011), .ZN(
      n_257_76_12012));
   NAND2_X1 i_257_76_12034 (.A1(n_257_253), .A2(n_257_425), .ZN(n_257_76_12013));
   NAND2_X1 i_257_76_12035 (.A1(n_257_173), .A2(n_257_429), .ZN(n_257_76_12014));
   NAND4_X1 i_257_76_12036 (.A1(n_257_76_12007), .A2(n_257_76_12012), .A3(
      n_257_76_12013), .A4(n_257_76_12014), .ZN(n_257_76_12015));
   INV_X1 i_257_76_12037 (.A(n_257_76_12015), .ZN(n_257_76_12016));
   NAND2_X1 i_257_76_12038 (.A1(n_257_96), .A2(n_257_431), .ZN(n_257_76_12017));
   NAND2_X1 i_257_76_12039 (.A1(n_257_213), .A2(n_257_427), .ZN(n_257_76_12018));
   NAND3_X1 i_257_76_12040 (.A1(n_257_76_12018), .A2(n_257_76_11970), .A3(
      n_257_76_11971), .ZN(n_257_76_12019));
   INV_X1 i_257_76_12041 (.A(n_257_1080), .ZN(n_257_76_12020));
   NAND2_X1 i_257_76_12042 (.A1(n_257_432), .A2(n_257_618), .ZN(n_257_76_12021));
   NAND2_X1 i_257_76_12043 (.A1(n_257_76_12021), .A2(n_257_423), .ZN(
      n_257_76_12022));
   INV_X1 i_257_76_12044 (.A(n_257_76_12022), .ZN(n_257_76_12023));
   NAND4_X1 i_257_76_12045 (.A1(n_257_76_11972), .A2(n_257_76_12020), .A3(
      n_257_76_18011), .A4(n_257_76_12023), .ZN(n_257_76_12024));
   NOR2_X1 i_257_76_12046 (.A1(n_257_76_12019), .A2(n_257_76_12024), .ZN(
      n_257_76_12025));
   NAND2_X1 i_257_76_12047 (.A1(n_257_56), .A2(n_257_433), .ZN(n_257_76_12026));
   NAND2_X1 i_257_76_12048 (.A1(n_257_76_12026), .A2(n_257_76_11961), .ZN(
      n_257_76_12027));
   INV_X1 i_257_76_12049 (.A(n_257_76_12027), .ZN(n_257_76_12028));
   NAND2_X1 i_257_76_12050 (.A1(n_257_522), .A2(n_257_424), .ZN(n_257_76_12029));
   NAND2_X1 i_257_76_12051 (.A1(n_257_76_12029), .A2(n_257_293), .ZN(
      n_257_76_12030));
   INV_X1 i_257_76_12052 (.A(n_257_76_12030), .ZN(n_257_76_12031));
   NAND3_X1 i_257_76_12053 (.A1(n_257_76_12025), .A2(n_257_76_12028), .A3(
      n_257_76_12031), .ZN(n_257_76_12032));
   INV_X1 i_257_76_12054 (.A(n_257_76_12032), .ZN(n_257_76_12033));
   NAND3_X1 i_257_76_12055 (.A1(n_257_76_11960), .A2(n_257_76_12017), .A3(
      n_257_76_12033), .ZN(n_257_76_12034));
   INV_X1 i_257_76_12056 (.A(n_257_76_12034), .ZN(n_257_76_12035));
   NAND4_X1 i_257_76_12057 (.A1(n_257_76_12016), .A2(n_257_76_12035), .A3(
      n_257_76_11941), .A4(n_257_76_11943), .ZN(n_257_76_12036));
   INV_X1 i_257_76_12058 (.A(n_257_76_12036), .ZN(n_257_76_12037));
   NAND2_X1 i_257_76_12059 (.A1(n_257_76_18066), .A2(n_257_76_12037), .ZN(
      n_257_76_12038));
   NAND3_X1 i_257_76_12060 (.A1(n_257_76_11996), .A2(n_257_76_12003), .A3(
      n_257_76_12038), .ZN(n_257_76_12039));
   NOR2_X1 i_257_76_12061 (.A1(n_257_76_11986), .A2(n_257_76_12039), .ZN(
      n_257_76_12040));
   NAND3_X1 i_257_76_12062 (.A1(n_257_441), .A2(n_257_984), .A3(n_257_76_11954), 
      .ZN(n_257_76_12041));
   INV_X1 i_257_76_12063 (.A(n_257_76_12041), .ZN(n_257_76_12042));
   NAND2_X1 i_257_76_12064 (.A1(n_257_76_11943), .A2(n_257_76_12042), .ZN(
      n_257_76_12043));
   NOR2_X1 i_257_76_12065 (.A1(n_257_76_11942), .A2(n_257_76_12043), .ZN(
      n_257_76_12044));
   NAND2_X1 i_257_76_12066 (.A1(n_257_76_18071), .A2(n_257_76_12044), .ZN(
      n_257_76_12045));
   NAND2_X1 i_257_76_12067 (.A1(n_257_76_11972), .A2(n_257_76_11971), .ZN(
      n_257_76_12046));
   NAND3_X1 i_257_76_12068 (.A1(n_257_76_12020), .A2(n_257_722), .A3(
      n_257_76_15655), .ZN(n_257_76_12047));
   NOR2_X1 i_257_76_12069 (.A1(n_257_76_12046), .A2(n_257_76_12047), .ZN(
      n_257_76_12048));
   NAND2_X1 i_257_76_12070 (.A1(n_257_76_11964), .A2(n_257_76_11966), .ZN(
      n_257_76_12049));
   INV_X1 i_257_76_12071 (.A(n_257_76_12049), .ZN(n_257_76_12050));
   NAND4_X1 i_257_76_12072 (.A1(n_257_76_12048), .A2(n_257_76_12050), .A3(
      n_257_76_11944), .A4(n_257_76_11961), .ZN(n_257_76_12051));
   NOR2_X1 i_257_76_12073 (.A1(n_257_76_11979), .A2(n_257_76_12051), .ZN(
      n_257_76_12052));
   NAND2_X1 i_257_76_12074 (.A1(n_257_76_11943), .A2(n_257_76_12052), .ZN(
      n_257_76_12053));
   NOR2_X1 i_257_76_12075 (.A1(n_257_76_11942), .A2(n_257_76_12053), .ZN(
      n_257_76_12054));
   NAND2_X1 i_257_76_12076 (.A1(n_257_76_18078), .A2(n_257_76_12054), .ZN(
      n_257_76_12055));
   NAND3_X1 i_257_76_12077 (.A1(n_257_586), .A2(n_257_428), .A3(n_257_442), 
      .ZN(n_257_76_12056));
   INV_X1 i_257_76_12078 (.A(n_257_76_12021), .ZN(n_257_76_12057));
   NOR2_X1 i_257_76_12079 (.A1(n_257_76_12056), .A2(n_257_76_12057), .ZN(
      n_257_76_12058));
   NAND3_X1 i_257_76_12080 (.A1(n_257_76_11972), .A2(n_257_76_12058), .A3(
      n_257_76_12020), .ZN(n_257_76_12059));
   NAND2_X1 i_257_76_12081 (.A1(n_257_76_11970), .A2(n_257_76_11971), .ZN(
      n_257_76_12060));
   NOR2_X1 i_257_76_12082 (.A1(n_257_76_12059), .A2(n_257_76_12060), .ZN(
      n_257_76_12061));
   NAND3_X1 i_257_76_12083 (.A1(n_257_76_12028), .A2(n_257_76_12061), .A3(
      n_257_76_11968), .ZN(n_257_76_12062));
   NAND3_X1 i_257_76_12084 (.A1(n_257_76_12010), .A2(n_257_76_12008), .A3(
      n_257_76_11944), .ZN(n_257_76_12063));
   NOR2_X1 i_257_76_12085 (.A1(n_257_76_12062), .A2(n_257_76_12063), .ZN(
      n_257_76_12064));
   NAND4_X1 i_257_76_12086 (.A1(n_257_76_11976), .A2(n_257_76_11977), .A3(
      n_257_76_12005), .A4(n_257_76_11978), .ZN(n_257_76_12065));
   INV_X1 i_257_76_12087 (.A(n_257_76_12065), .ZN(n_257_76_12066));
   NAND3_X1 i_257_76_12088 (.A1(n_257_76_12064), .A2(n_257_76_12066), .A3(
      n_257_76_12014), .ZN(n_257_76_12067));
   INV_X1 i_257_76_12089 (.A(n_257_76_12067), .ZN(n_257_76_12068));
   NAND2_X1 i_257_76_12090 (.A1(n_257_76_11960), .A2(n_257_76_12017), .ZN(
      n_257_76_12069));
   INV_X1 i_257_76_12091 (.A(n_257_76_12069), .ZN(n_257_76_12070));
   NAND4_X1 i_257_76_12092 (.A1(n_257_76_11941), .A2(n_257_76_12068), .A3(
      n_257_76_12070), .A4(n_257_76_11943), .ZN(n_257_76_12071));
   INV_X1 i_257_76_12093 (.A(n_257_76_12071), .ZN(n_257_76_12072));
   NAND2_X1 i_257_76_12094 (.A1(n_257_76_18074), .A2(n_257_76_12072), .ZN(
      n_257_76_12073));
   NAND3_X1 i_257_76_12095 (.A1(n_257_76_12045), .A2(n_257_76_12055), .A3(
      n_257_76_12073), .ZN(n_257_76_12074));
   NAND2_X1 i_257_76_12096 (.A1(n_257_1080), .A2(n_257_442), .ZN(n_257_76_12075));
   INV_X1 i_257_76_12097 (.A(n_257_76_12075), .ZN(n_257_76_12076));
   NAND2_X1 i_257_76_12098 (.A1(n_257_13), .A2(n_257_76_12076), .ZN(
      n_257_76_12077));
   NOR2_X1 i_257_76_12099 (.A1(n_257_1080), .A2(n_257_76_17902), .ZN(
      n_257_76_12078));
   NAND4_X1 i_257_76_12100 (.A1(n_257_882), .A2(n_257_76_12078), .A3(
      n_257_76_11971), .A4(n_257_76_11972), .ZN(n_257_76_12079));
   INV_X1 i_257_76_12101 (.A(n_257_76_12079), .ZN(n_257_76_12080));
   NAND3_X1 i_257_76_12102 (.A1(n_257_76_12080), .A2(n_257_76_11978), .A3(
      n_257_76_11944), .ZN(n_257_76_12081));
   INV_X1 i_257_76_12103 (.A(n_257_76_12081), .ZN(n_257_76_12082));
   NAND2_X1 i_257_76_12104 (.A1(n_257_76_11943), .A2(n_257_76_12082), .ZN(
      n_257_76_12083));
   NOR2_X1 i_257_76_12105 (.A1(n_257_76_11942), .A2(n_257_76_12083), .ZN(
      n_257_76_12084));
   NAND2_X1 i_257_76_12106 (.A1(n_257_76_18077), .A2(n_257_76_12084), .ZN(
      n_257_76_12085));
   NAND2_X1 i_257_76_12107 (.A1(n_257_76_12077), .A2(n_257_76_12085), .ZN(
      n_257_76_12086));
   NOR2_X1 i_257_76_12108 (.A1(n_257_76_12074), .A2(n_257_76_12086), .ZN(
      n_257_76_12087));
   INV_X1 i_257_76_12109 (.A(n_257_76_12019), .ZN(n_257_76_12088));
   NAND2_X1 i_257_76_12110 (.A1(n_257_76_12021), .A2(n_257_426), .ZN(
      n_257_76_12089));
   INV_X1 i_257_76_12111 (.A(n_257_76_12089), .ZN(n_257_76_12090));
   NAND4_X1 i_257_76_12112 (.A1(n_257_76_11972), .A2(n_257_76_12020), .A3(
      n_257_76_18011), .A4(n_257_76_12090), .ZN(n_257_76_12091));
   INV_X1 i_257_76_12113 (.A(n_257_76_12091), .ZN(n_257_76_12092));
   NAND4_X1 i_257_76_12114 (.A1(n_257_76_12088), .A2(n_257_76_12092), .A3(
      n_257_76_11965), .A4(n_257_76_11966), .ZN(n_257_76_12093));
   NAND4_X1 i_257_76_12115 (.A1(n_257_76_11944), .A2(n_257_76_12026), .A3(
      n_257_76_11961), .A4(n_257_76_11964), .ZN(n_257_76_12094));
   NOR2_X1 i_257_76_12116 (.A1(n_257_76_12093), .A2(n_257_76_12094), .ZN(
      n_257_76_12095));
   NAND3_X1 i_257_76_12117 (.A1(n_257_76_11976), .A2(n_257_76_11977), .A3(
      n_257_76_12005), .ZN(n_257_76_12096));
   INV_X1 i_257_76_12118 (.A(n_257_76_12096), .ZN(n_257_76_12097));
   NAND3_X1 i_257_76_12119 (.A1(n_257_76_11978), .A2(n_257_554), .A3(
      n_257_76_12008), .ZN(n_257_76_12098));
   INV_X1 i_257_76_12120 (.A(n_257_76_12098), .ZN(n_257_76_12099));
   NAND3_X1 i_257_76_12121 (.A1(n_257_76_12095), .A2(n_257_76_12097), .A3(
      n_257_76_12099), .ZN(n_257_76_12100));
   INV_X1 i_257_76_12122 (.A(n_257_76_12100), .ZN(n_257_76_12101));
   NAND2_X1 i_257_76_12123 (.A1(n_257_76_11941), .A2(n_257_76_12101), .ZN(
      n_257_76_12102));
   NAND2_X1 i_257_76_12124 (.A1(n_257_76_12014), .A2(n_257_76_12010), .ZN(
      n_257_76_12103));
   INV_X1 i_257_76_12125 (.A(n_257_76_12103), .ZN(n_257_76_12104));
   NAND4_X1 i_257_76_12126 (.A1(n_257_76_11943), .A2(n_257_76_11960), .A3(
      n_257_76_12017), .A4(n_257_76_12104), .ZN(n_257_76_12105));
   NOR2_X1 i_257_76_12127 (.A1(n_257_76_12102), .A2(n_257_76_12105), .ZN(
      n_257_76_12106));
   NAND2_X1 i_257_76_12128 (.A1(n_257_76_18076), .A2(n_257_76_12106), .ZN(
      n_257_76_12107));
   NAND3_X1 i_257_76_12129 (.A1(n_257_76_11977), .A2(n_257_76_11978), .A3(
      n_257_754), .ZN(n_257_76_12108));
   NOR2_X1 i_257_76_12130 (.A1(n_257_1080), .A2(n_257_76_17934), .ZN(
      n_257_76_12109));
   NAND3_X1 i_257_76_12131 (.A1(n_257_76_12109), .A2(n_257_76_11972), .A3(
      n_257_76_11971), .ZN(n_257_76_12110));
   INV_X1 i_257_76_12132 (.A(n_257_76_12110), .ZN(n_257_76_12111));
   NAND4_X1 i_257_76_12133 (.A1(n_257_76_12050), .A2(n_257_76_12111), .A3(
      n_257_76_11944), .A4(n_257_76_11961), .ZN(n_257_76_12112));
   NOR2_X1 i_257_76_12134 (.A1(n_257_76_12108), .A2(n_257_76_12112), .ZN(
      n_257_76_12113));
   NAND2_X1 i_257_76_12135 (.A1(n_257_76_11943), .A2(n_257_76_12113), .ZN(
      n_257_76_12114));
   NOR2_X1 i_257_76_12136 (.A1(n_257_76_11942), .A2(n_257_76_12114), .ZN(
      n_257_76_12115));
   NAND2_X1 i_257_76_12137 (.A1(n_257_76_18069), .A2(n_257_76_12115), .ZN(
      n_257_76_12116));
   NAND3_X1 i_257_76_12138 (.A1(n_257_432), .A2(n_257_618), .A3(n_257_442), 
      .ZN(n_257_76_12117));
   NOR2_X1 i_257_76_12139 (.A1(n_257_1080), .A2(n_257_76_12117), .ZN(
      n_257_76_12118));
   NAND4_X1 i_257_76_12140 (.A1(n_257_76_12118), .A2(n_257_76_11970), .A3(
      n_257_76_11971), .A4(n_257_76_11972), .ZN(n_257_76_12119));
   NOR2_X1 i_257_76_12141 (.A1(n_257_76_11967), .A2(n_257_76_12119), .ZN(
      n_257_76_12120));
   NAND3_X1 i_257_76_12142 (.A1(n_257_76_11944), .A2(n_257_76_12026), .A3(
      n_257_76_11961), .ZN(n_257_76_12121));
   INV_X1 i_257_76_12143 (.A(n_257_76_12121), .ZN(n_257_76_12122));
   NAND3_X1 i_257_76_12144 (.A1(n_257_76_12120), .A2(n_257_76_12122), .A3(
      n_257_76_12008), .ZN(n_257_76_12123));
   INV_X1 i_257_76_12145 (.A(n_257_76_12123), .ZN(n_257_76_12124));
   NAND4_X1 i_257_76_12146 (.A1(n_257_76_11976), .A2(n_257_76_11977), .A3(
      n_257_76_11978), .A4(n_257_76_12010), .ZN(n_257_76_12125));
   INV_X1 i_257_76_12147 (.A(n_257_76_12125), .ZN(n_257_76_12126));
   NAND2_X1 i_257_76_12148 (.A1(n_257_76_12124), .A2(n_257_76_12126), .ZN(
      n_257_76_12127));
   INV_X1 i_257_76_12149 (.A(n_257_76_11960), .ZN(n_257_76_12128));
   NOR2_X1 i_257_76_12150 (.A1(n_257_76_12127), .A2(n_257_76_12128), .ZN(
      n_257_76_12129));
   NAND3_X1 i_257_76_12151 (.A1(n_257_76_12129), .A2(n_257_76_11941), .A3(
      n_257_76_11943), .ZN(n_257_76_12130));
   INV_X1 i_257_76_12152 (.A(n_257_76_12130), .ZN(n_257_76_12131));
   NAND2_X1 i_257_76_12153 (.A1(n_257_68), .A2(n_257_76_12131), .ZN(
      n_257_76_12132));
   NAND3_X1 i_257_76_12154 (.A1(n_257_76_12107), .A2(n_257_76_12116), .A3(
      n_257_76_12132), .ZN(n_257_76_12133));
   NOR2_X1 i_257_76_12155 (.A1(n_257_1080), .A2(n_257_76_17951), .ZN(
      n_257_76_12134));
   NAND3_X1 i_257_76_12156 (.A1(n_257_76_12134), .A2(n_257_76_11972), .A3(
      n_257_76_11971), .ZN(n_257_76_12135));
   INV_X1 i_257_76_12157 (.A(n_257_76_12135), .ZN(n_257_76_12136));
   NAND4_X1 i_257_76_12158 (.A1(n_257_76_12136), .A2(n_257_76_11944), .A3(
      n_257_76_11961), .A4(n_257_76_11964), .ZN(n_257_76_12137));
   NAND2_X1 i_257_76_12159 (.A1(n_257_76_11978), .A2(n_257_818), .ZN(
      n_257_76_12138));
   NOR2_X1 i_257_76_12160 (.A1(n_257_76_12137), .A2(n_257_76_12138), .ZN(
      n_257_76_12139));
   NAND2_X1 i_257_76_12161 (.A1(n_257_76_11943), .A2(n_257_76_12139), .ZN(
      n_257_76_12140));
   NOR2_X1 i_257_76_12162 (.A1(n_257_76_11942), .A2(n_257_76_12140), .ZN(
      n_257_76_12141));
   NAND2_X1 i_257_76_12163 (.A1(n_257_22), .A2(n_257_76_12141), .ZN(
      n_257_76_12142));
   NAND2_X1 i_257_76_12164 (.A1(n_257_444), .A2(n_257_76_11954), .ZN(
      n_257_76_12143));
   INV_X1 i_257_76_12165 (.A(n_257_76_12143), .ZN(n_257_76_12144));
   NAND2_X1 i_257_76_12166 (.A1(n_257_1016), .A2(n_257_76_12144), .ZN(
      n_257_76_12145));
   INV_X1 i_257_76_12167 (.A(n_257_76_12145), .ZN(n_257_76_12146));
   NAND2_X1 i_257_76_12168 (.A1(n_257_76_11941), .A2(n_257_76_12146), .ZN(
      n_257_76_12147));
   INV_X1 i_257_76_12169 (.A(n_257_76_12147), .ZN(n_257_76_12148));
   NAND2_X1 i_257_76_12170 (.A1(n_257_76_18075), .A2(n_257_76_12148), .ZN(
      n_257_76_12149));
   NAND2_X1 i_257_76_12171 (.A1(n_257_76_12142), .A2(n_257_76_12149), .ZN(
      n_257_76_12150));
   NOR2_X1 i_257_76_12172 (.A1(n_257_76_12133), .A2(n_257_76_12150), .ZN(
      n_257_76_12151));
   NAND3_X1 i_257_76_12173 (.A1(n_257_76_12040), .A2(n_257_76_12087), .A3(
      n_257_76_12151), .ZN(n_257_76_12152));
   INV_X1 i_257_76_12174 (.A(n_257_76_12152), .ZN(n_257_76_12153));
   NOR2_X1 i_257_76_12175 (.A1(n_257_1080), .A2(n_257_76_17633), .ZN(
      n_257_76_12154));
   NAND3_X1 i_257_76_12176 (.A1(n_257_76_12154), .A2(n_257_76_11972), .A3(
      n_257_76_11971), .ZN(n_257_76_12155));
   NAND2_X1 i_257_76_12177 (.A1(n_257_56), .A2(n_257_76_11970), .ZN(
      n_257_76_12156));
   NOR2_X1 i_257_76_12178 (.A1(n_257_76_12155), .A2(n_257_76_12156), .ZN(
      n_257_76_12157));
   NAND2_X1 i_257_76_12179 (.A1(n_257_76_11944), .A2(n_257_76_11961), .ZN(
      n_257_76_12158));
   INV_X1 i_257_76_12180 (.A(n_257_76_12158), .ZN(n_257_76_12159));
   NAND4_X1 i_257_76_12181 (.A1(n_257_76_12157), .A2(n_257_76_12159), .A3(
      n_257_76_12008), .A4(n_257_76_11968), .ZN(n_257_76_12160));
   INV_X1 i_257_76_12182 (.A(n_257_76_12160), .ZN(n_257_76_12161));
   NAND2_X1 i_257_76_12183 (.A1(n_257_76_12161), .A2(n_257_76_12126), .ZN(
      n_257_76_12162));
   NOR2_X1 i_257_76_12184 (.A1(n_257_76_12162), .A2(n_257_76_12128), .ZN(
      n_257_76_12163));
   NAND3_X1 i_257_76_12185 (.A1(n_257_76_12163), .A2(n_257_76_11941), .A3(
      n_257_76_11943), .ZN(n_257_76_12164));
   INV_X1 i_257_76_12186 (.A(n_257_76_12164), .ZN(n_257_76_12165));
   NAND2_X1 i_257_76_12187 (.A1(n_257_76_18081), .A2(n_257_76_12165), .ZN(
      n_257_76_12166));
   INV_X1 i_257_76_12188 (.A(n_257_76_11979), .ZN(n_257_76_12167));
   NAND3_X1 i_257_76_12189 (.A1(n_257_76_11970), .A2(n_257_449), .A3(
      n_257_76_11971), .ZN(n_257_76_12168));
   INV_X1 i_257_76_12190 (.A(n_257_76_16553), .ZN(n_257_76_12169));
   NAND3_X1 i_257_76_12191 (.A1(n_257_76_11972), .A2(n_257_76_12020), .A3(
      n_257_76_12169), .ZN(n_257_76_12170));
   NOR2_X1 i_257_76_12192 (.A1(n_257_76_12168), .A2(n_257_76_12170), .ZN(
      n_257_76_12171));
   NAND4_X1 i_257_76_12193 (.A1(n_257_76_12171), .A2(n_257_76_12050), .A3(
      n_257_76_11944), .A4(n_257_76_11961), .ZN(n_257_76_12172));
   INV_X1 i_257_76_12194 (.A(n_257_76_12172), .ZN(n_257_76_12173));
   NAND2_X1 i_257_76_12195 (.A1(n_257_76_12167), .A2(n_257_76_12173), .ZN(
      n_257_76_12174));
   NOR2_X1 i_257_76_12196 (.A1(n_257_76_12128), .A2(n_257_76_12174), .ZN(
      n_257_76_12175));
   NAND3_X1 i_257_76_12197 (.A1(n_257_76_12175), .A2(n_257_76_11941), .A3(
      n_257_76_11943), .ZN(n_257_76_12176));
   INV_X1 i_257_76_12198 (.A(n_257_76_12176), .ZN(n_257_76_12177));
   NAND2_X1 i_257_76_12199 (.A1(n_257_76_18083), .A2(n_257_76_12177), .ZN(
      n_257_76_12178));
   NAND2_X1 i_257_76_12200 (.A1(n_257_76_15481), .A2(n_257_442), .ZN(
      n_257_76_12179));
   INV_X1 i_257_76_12201 (.A(n_257_618), .ZN(n_257_76_12180));
   NAND2_X1 i_257_76_12202 (.A1(n_257_76_12180), .A2(n_257_442), .ZN(
      n_257_76_12181));
   AOI21_X1 i_257_76_12203 (.A(n_257_76_17101), .B1(n_257_76_12179), .B2(
      n_257_76_12181), .ZN(n_257_76_12182));
   NAND3_X1 i_257_76_12204 (.A1(n_257_76_11972), .A2(n_257_76_12182), .A3(
      n_257_76_12020), .ZN(n_257_76_12183));
   INV_X1 i_257_76_12205 (.A(n_257_76_12183), .ZN(n_257_76_12184));
   INV_X1 i_257_76_12206 (.A(n_257_76_12060), .ZN(n_257_76_12185));
   NAND4_X1 i_257_76_12207 (.A1(n_257_76_12184), .A2(n_257_76_12185), .A3(
      n_257_76_11965), .A4(n_257_76_11966), .ZN(n_257_76_12186));
   NOR2_X1 i_257_76_12208 (.A1(n_257_76_12094), .A2(n_257_76_12186), .ZN(
      n_257_76_12187));
   NAND3_X1 i_257_76_12209 (.A1(n_257_76_11978), .A2(n_257_76_12010), .A3(
      n_257_76_12008), .ZN(n_257_76_12188));
   INV_X1 i_257_76_12210 (.A(n_257_76_12188), .ZN(n_257_76_12189));
   NAND4_X1 i_257_76_12211 (.A1(n_257_76_12187), .A2(n_257_76_12097), .A3(
      n_257_173), .A4(n_257_76_12189), .ZN(n_257_76_12190));
   INV_X1 i_257_76_12212 (.A(n_257_76_12190), .ZN(n_257_76_12191));
   NAND4_X1 i_257_76_12213 (.A1(n_257_76_11941), .A2(n_257_76_12070), .A3(
      n_257_76_12191), .A4(n_257_76_11943), .ZN(n_257_76_12192));
   INV_X1 i_257_76_12214 (.A(n_257_76_12192), .ZN(n_257_76_12193));
   NAND2_X1 i_257_76_12215 (.A1(n_257_76_18061), .A2(n_257_76_12193), .ZN(
      n_257_76_12194));
   NAND3_X1 i_257_76_12216 (.A1(n_257_76_12166), .A2(n_257_76_12178), .A3(
      n_257_76_12194), .ZN(n_257_76_12195));
   NAND2_X1 i_257_76_12217 (.A1(n_257_786), .A2(n_257_442), .ZN(n_257_76_12196));
   NOR2_X1 i_257_76_12218 (.A1(n_257_1080), .A2(n_257_76_12196), .ZN(
      n_257_76_12197));
   NAND4_X1 i_257_76_12219 (.A1(n_257_76_12197), .A2(n_257_447), .A3(
      n_257_76_11972), .A4(n_257_76_11971), .ZN(n_257_76_12198));
   INV_X1 i_257_76_12220 (.A(n_257_76_12198), .ZN(n_257_76_12199));
   NAND4_X1 i_257_76_12221 (.A1(n_257_76_12199), .A2(n_257_76_11944), .A3(
      n_257_76_11961), .A4(n_257_76_11964), .ZN(n_257_76_12200));
   NAND2_X1 i_257_76_12222 (.A1(n_257_76_11977), .A2(n_257_76_11978), .ZN(
      n_257_76_12201));
   NOR2_X1 i_257_76_12223 (.A1(n_257_76_12200), .A2(n_257_76_12201), .ZN(
      n_257_76_12202));
   NAND2_X1 i_257_76_12224 (.A1(n_257_76_11943), .A2(n_257_76_12202), .ZN(
      n_257_76_12203));
   NOR2_X1 i_257_76_12225 (.A1(n_257_76_11942), .A2(n_257_76_12203), .ZN(
      n_257_76_12204));
   NAND2_X1 i_257_76_12226 (.A1(n_257_76_18085), .A2(n_257_76_12204), .ZN(
      n_257_76_12205));
   NAND3_X1 i_257_76_12227 (.A1(n_257_76_11972), .A2(n_257_76_18012), .A3(
      n_257_76_12020), .ZN(n_257_76_12206));
   INV_X1 i_257_76_12228 (.A(n_257_76_12206), .ZN(n_257_76_12207));
   NAND4_X1 i_257_76_12229 (.A1(n_257_76_12207), .A2(n_257_76_12185), .A3(
      n_257_76_11965), .A4(n_257_76_11966), .ZN(n_257_76_12208));
   NOR2_X1 i_257_76_12230 (.A1(n_257_76_12094), .A2(n_257_76_12208), .ZN(
      n_257_76_12209));
   NAND2_X1 i_257_76_12231 (.A1(n_257_76_11976), .A2(n_257_76_11977), .ZN(
      n_257_76_12210));
   INV_X1 i_257_76_12232 (.A(n_257_76_12210), .ZN(n_257_76_12211));
   NAND4_X1 i_257_76_12233 (.A1(n_257_76_12209), .A2(n_257_96), .A3(
      n_257_76_12211), .A4(n_257_76_12189), .ZN(n_257_76_12212));
   INV_X1 i_257_76_12234 (.A(n_257_76_12212), .ZN(n_257_76_12213));
   NAND3_X1 i_257_76_12235 (.A1(n_257_76_12213), .A2(n_257_76_11943), .A3(
      n_257_76_11960), .ZN(n_257_76_12214));
   NOR2_X1 i_257_76_12236 (.A1(n_257_76_12214), .A2(n_257_76_11942), .ZN(
      n_257_76_12215));
   NAND2_X1 i_257_76_12237 (.A1(n_257_76_18080), .A2(n_257_76_12215), .ZN(
      n_257_76_12216));
   NAND2_X1 i_257_76_12238 (.A1(n_257_76_12205), .A2(n_257_76_12216), .ZN(
      n_257_76_12217));
   NOR2_X1 i_257_76_12239 (.A1(n_257_76_12195), .A2(n_257_76_12217), .ZN(
      n_257_76_12218));
   NAND2_X1 i_257_76_12240 (.A1(n_257_76_11971), .A2(n_257_76_18013), .ZN(
      n_257_76_12219));
   INV_X1 i_257_76_12241 (.A(n_257_76_12219), .ZN(n_257_76_12220));
   NAND2_X1 i_257_76_12242 (.A1(n_257_76_11972), .A2(n_257_76_12020), .ZN(
      n_257_76_12221));
   INV_X1 i_257_76_12243 (.A(n_257_76_12221), .ZN(n_257_76_12222));
   NAND3_X1 i_257_76_12244 (.A1(n_257_76_12220), .A2(n_257_76_12222), .A3(
      n_257_76_11970), .ZN(n_257_76_12223));
   NOR2_X1 i_257_76_12245 (.A1(n_257_76_12223), .A2(n_257_76_11967), .ZN(
      n_257_76_12224));
   NAND2_X1 i_257_76_12246 (.A1(n_257_76_12008), .A2(n_257_76_11944), .ZN(
      n_257_76_12225));
   INV_X1 i_257_76_12247 (.A(n_257_76_12225), .ZN(n_257_76_12226));
   NAND3_X1 i_257_76_12248 (.A1(n_257_134), .A2(n_257_76_12026), .A3(
      n_257_76_11961), .ZN(n_257_76_12227));
   INV_X1 i_257_76_12249 (.A(n_257_76_12227), .ZN(n_257_76_12228));
   NAND3_X1 i_257_76_12250 (.A1(n_257_76_12224), .A2(n_257_76_12226), .A3(
      n_257_76_12228), .ZN(n_257_76_12229));
   NOR2_X1 i_257_76_12251 (.A1(n_257_76_12229), .A2(n_257_76_12125), .ZN(
      n_257_76_12230));
   NAND3_X1 i_257_76_12252 (.A1(n_257_76_12230), .A2(n_257_76_11960), .A3(
      n_257_76_12017), .ZN(n_257_76_12231));
   INV_X1 i_257_76_12253 (.A(n_257_76_12231), .ZN(n_257_76_12232));
   NAND3_X1 i_257_76_12254 (.A1(n_257_76_12232), .A2(n_257_76_11941), .A3(
      n_257_76_11943), .ZN(n_257_76_12233));
   INV_X1 i_257_76_12255 (.A(n_257_76_12233), .ZN(n_257_76_12234));
   NAND2_X1 i_257_76_12256 (.A1(n_257_76_18068), .A2(n_257_76_12234), .ZN(
      n_257_76_12235));
   NAND3_X1 i_257_76_12257 (.A1(n_257_76_11964), .A2(n_257_76_11966), .A3(
      n_257_448), .ZN(n_257_76_12236));
   INV_X1 i_257_76_12258 (.A(n_257_76_12236), .ZN(n_257_76_12237));
   NAND4_X1 i_257_76_12259 (.A1(n_257_76_11977), .A2(n_257_76_12237), .A3(
      n_257_76_11978), .A4(n_257_76_11944), .ZN(n_257_76_12238));
   INV_X1 i_257_76_12260 (.A(n_257_76_12238), .ZN(n_257_76_12239));
   NAND3_X1 i_257_76_12261 (.A1(n_257_76_11972), .A2(n_257_76_11971), .A3(
      n_257_76_12020), .ZN(n_257_76_12240));
   INV_X1 i_257_76_12262 (.A(n_257_76_12240), .ZN(n_257_76_12241));
   OAI21_X1 i_257_76_12263 (.A(n_257_76_17761), .B1(n_257_722), .B2(
      n_257_76_17412), .ZN(n_257_76_12242));
   NAND3_X1 i_257_76_12264 (.A1(n_257_76_11961), .A2(n_257_76_12241), .A3(
      n_257_76_12242), .ZN(n_257_76_12243));
   INV_X1 i_257_76_12265 (.A(n_257_76_12243), .ZN(n_257_76_12244));
   NAND2_X1 i_257_76_12266 (.A1(n_257_76_11976), .A2(n_257_76_12244), .ZN(
      n_257_76_12245));
   INV_X1 i_257_76_12267 (.A(n_257_76_12245), .ZN(n_257_76_12246));
   NAND3_X1 i_257_76_12268 (.A1(n_257_76_12239), .A2(n_257_690), .A3(
      n_257_76_12246), .ZN(n_257_76_12247));
   INV_X1 i_257_76_12269 (.A(n_257_76_12247), .ZN(n_257_76_12248));
   NAND2_X1 i_257_76_12270 (.A1(n_257_76_12248), .A2(n_257_76_11943), .ZN(
      n_257_76_12249));
   NOR2_X1 i_257_76_12271 (.A1(n_257_76_11942), .A2(n_257_76_12249), .ZN(
      n_257_76_12250));
   NAND2_X1 i_257_76_12272 (.A1(n_257_76_18079), .A2(n_257_76_12250), .ZN(
      n_257_76_12251));
   NAND3_X1 i_257_76_12273 (.A1(n_257_76_11941), .A2(n_257_76_11943), .A3(
      n_257_76_11960), .ZN(n_257_76_12252));
   INV_X1 i_257_76_12274 (.A(n_257_76_18011), .ZN(n_257_76_12253));
   NAND2_X1 i_257_76_12275 (.A1(n_257_76_12021), .A2(n_257_425), .ZN(
      n_257_76_12254));
   NOR2_X1 i_257_76_12276 (.A1(n_257_76_12253), .A2(n_257_76_12254), .ZN(
      n_257_76_12255));
   NAND4_X1 i_257_76_12277 (.A1(n_257_76_12255), .A2(n_257_76_11972), .A3(
      n_257_76_11971), .A4(n_257_76_12020), .ZN(n_257_76_12256));
   NAND3_X1 i_257_76_12278 (.A1(n_257_76_11966), .A2(n_257_76_12018), .A3(
      n_257_76_11970), .ZN(n_257_76_12257));
   NOR2_X1 i_257_76_12279 (.A1(n_257_76_12256), .A2(n_257_76_12257), .ZN(
      n_257_76_12258));
   NAND2_X1 i_257_76_12280 (.A1(n_257_76_11944), .A2(n_257_76_12026), .ZN(
      n_257_76_12259));
   INV_X1 i_257_76_12281 (.A(n_257_76_12259), .ZN(n_257_76_12260));
   NAND3_X1 i_257_76_12282 (.A1(n_257_76_11961), .A2(n_257_76_11964), .A3(
      n_257_76_11965), .ZN(n_257_76_12261));
   INV_X1 i_257_76_12283 (.A(n_257_76_12261), .ZN(n_257_76_12262));
   NAND3_X1 i_257_76_12284 (.A1(n_257_76_12258), .A2(n_257_76_12260), .A3(
      n_257_76_12262), .ZN(n_257_76_12263));
   NAND4_X1 i_257_76_12285 (.A1(n_257_76_12005), .A2(n_257_76_11978), .A3(
      n_257_76_12010), .A4(n_257_76_12008), .ZN(n_257_76_12264));
   NOR2_X1 i_257_76_12286 (.A1(n_257_76_12263), .A2(n_257_76_12264), .ZN(
      n_257_76_12265));
   NAND3_X1 i_257_76_12287 (.A1(n_257_76_12004), .A2(n_257_76_11976), .A3(
      n_257_76_11977), .ZN(n_257_76_12266));
   INV_X1 i_257_76_12288 (.A(n_257_253), .ZN(n_257_76_12267));
   NOR2_X1 i_257_76_12289 (.A1(n_257_76_12266), .A2(n_257_76_12267), .ZN(
      n_257_76_12268));
   NAND4_X1 i_257_76_12290 (.A1(n_257_76_12265), .A2(n_257_76_12017), .A3(
      n_257_76_12014), .A4(n_257_76_12268), .ZN(n_257_76_12269));
   NOR2_X1 i_257_76_12291 (.A1(n_257_76_12252), .A2(n_257_76_12269), .ZN(
      n_257_76_12270));
   NAND2_X1 i_257_76_12292 (.A1(n_257_76_18064), .A2(n_257_76_12270), .ZN(
      n_257_76_12271));
   NAND3_X1 i_257_76_12293 (.A1(n_257_76_12235), .A2(n_257_76_12251), .A3(
      n_257_76_12271), .ZN(n_257_76_12272));
   INV_X1 i_257_76_12294 (.A(n_257_76_11971), .ZN(n_257_76_12273));
   NAND3_X1 i_257_76_12295 (.A1(n_257_76_11954), .A2(n_257_76_12273), .A3(
      n_257_76_11972), .ZN(n_257_76_12274));
   INV_X1 i_257_76_12296 (.A(n_257_76_12274), .ZN(n_257_76_12275));
   NAND2_X1 i_257_76_12297 (.A1(n_257_76_12275), .A2(n_257_76_11944), .ZN(
      n_257_76_12276));
   NOR2_X1 i_257_76_12298 (.A1(n_257_76_12276), .A2(n_257_76_11992), .ZN(
      n_257_76_12277));
   NAND2_X1 i_257_76_12299 (.A1(n_257_76_11943), .A2(n_257_76_12277), .ZN(
      n_257_76_12278));
   NOR2_X1 i_257_76_12300 (.A1(n_257_76_11942), .A2(n_257_76_12278), .ZN(
      n_257_76_12279));
   NAND2_X1 i_257_76_12301 (.A1(n_257_76_18067), .A2(n_257_76_12279), .ZN(
      n_257_76_12280));
   NAND2_X1 i_257_76_12302 (.A1(n_257_76_11964), .A2(n_257_76_11965), .ZN(
      n_257_76_12281));
   INV_X1 i_257_76_12303 (.A(n_257_76_12281), .ZN(n_257_76_12282));
   NAND2_X1 i_257_76_12304 (.A1(n_257_76_11966), .A2(n_257_76_12018), .ZN(
      n_257_76_12283));
   INV_X1 i_257_76_12305 (.A(n_257_76_12283), .ZN(n_257_76_12284));
   NAND3_X1 i_257_76_12306 (.A1(n_257_76_11970), .A2(n_257_76_11972), .A3(
      n_257_76_11971), .ZN(n_257_76_12285));
   INV_X1 i_257_76_12307 (.A(n_257_76_12285), .ZN(n_257_76_12286));
   NAND3_X1 i_257_76_12308 (.A1(n_257_76_12282), .A2(n_257_76_12284), .A3(
      n_257_76_12286), .ZN(n_257_76_12287));
   NAND4_X1 i_257_76_12309 (.A1(n_257_76_11944), .A2(n_257_76_12026), .A3(
      n_257_76_11961), .A4(n_257_76_12029), .ZN(n_257_76_12288));
   NOR2_X1 i_257_76_12310 (.A1(n_257_76_12287), .A2(n_257_76_12288), .ZN(
      n_257_76_12289));
   NAND3_X1 i_257_76_12311 (.A1(n_257_76_11977), .A2(n_257_76_12005), .A3(
      n_257_76_11978), .ZN(n_257_76_12290));
   INV_X1 i_257_76_12312 (.A(n_257_76_12290), .ZN(n_257_76_12291));
   NAND2_X1 i_257_76_12313 (.A1(n_257_442), .A2(n_257_490), .ZN(n_257_76_12292));
   INV_X1 i_257_76_12314 (.A(n_257_76_18014), .ZN(n_257_76_12293));
   NOR2_X1 i_257_76_12315 (.A1(n_257_76_12293), .A2(n_257_1080), .ZN(
      n_257_76_12294));
   NAND2_X1 i_257_76_12316 (.A1(n_257_331), .A2(n_257_422), .ZN(n_257_76_12295));
   NAND2_X1 i_257_76_12317 (.A1(n_257_420), .A2(n_257_76_12021), .ZN(
      n_257_76_12296));
   INV_X1 i_257_76_12318 (.A(n_257_76_12296), .ZN(n_257_76_12297));
   NAND3_X1 i_257_76_12319 (.A1(n_257_76_12294), .A2(n_257_76_12295), .A3(
      n_257_76_12297), .ZN(n_257_76_12298));
   INV_X1 i_257_76_12320 (.A(n_257_76_12298), .ZN(n_257_76_12299));
   NAND2_X1 i_257_76_12321 (.A1(n_257_293), .A2(n_257_423), .ZN(n_257_76_12300));
   NAND4_X1 i_257_76_12322 (.A1(n_257_76_12010), .A2(n_257_76_12008), .A3(
      n_257_76_12299), .A4(n_257_76_12300), .ZN(n_257_76_12301));
   INV_X1 i_257_76_12323 (.A(n_257_76_12301), .ZN(n_257_76_12302));
   NAND3_X1 i_257_76_12324 (.A1(n_257_76_12289), .A2(n_257_76_12291), .A3(
      n_257_76_12302), .ZN(n_257_76_12303));
   NAND2_X1 i_257_76_12325 (.A1(n_257_76_12004), .A2(n_257_76_11976), .ZN(
      n_257_76_12304));
   INV_X1 i_257_76_12326 (.A(n_257_76_12304), .ZN(n_257_76_12305));
   NAND2_X1 i_257_76_12327 (.A1(n_257_370), .A2(n_257_421), .ZN(n_257_76_12306));
   NAND3_X1 i_257_76_12328 (.A1(n_257_76_12014), .A2(n_257_76_12305), .A3(
      n_257_76_12306), .ZN(n_257_76_12307));
   NOR2_X1 i_257_76_12329 (.A1(n_257_76_12303), .A2(n_257_76_12307), .ZN(
      n_257_76_12308));
   NAND3_X1 i_257_76_12330 (.A1(n_257_76_11960), .A2(n_257_76_12017), .A3(
      n_257_76_12013), .ZN(n_257_76_12309));
   INV_X1 i_257_76_12331 (.A(n_257_76_12309), .ZN(n_257_76_12310));
   NAND4_X1 i_257_76_12332 (.A1(n_257_76_12308), .A2(n_257_76_11941), .A3(
      n_257_76_12310), .A4(n_257_76_11943), .ZN(n_257_76_12311));
   INV_X1 i_257_76_12333 (.A(n_257_76_12311), .ZN(n_257_76_12312));
   NAND2_X1 i_257_76_12334 (.A1(n_257_76_18073), .A2(n_257_76_12312), .ZN(
      n_257_76_12313));
   NAND2_X1 i_257_76_12335 (.A1(n_257_76_12280), .A2(n_257_76_12313), .ZN(
      n_257_76_12314));
   NOR2_X1 i_257_76_12336 (.A1(n_257_76_12272), .A2(n_257_76_12314), .ZN(
      n_257_76_12315));
   NAND2_X1 i_257_76_12337 (.A1(n_257_76_12021), .A2(n_257_421), .ZN(
      n_257_76_12316));
   NOR2_X1 i_257_76_12338 (.A1(n_257_76_12253), .A2(n_257_76_12316), .ZN(
      n_257_76_12317));
   NAND4_X1 i_257_76_12339 (.A1(n_257_76_12317), .A2(n_257_76_11972), .A3(
      n_257_76_11971), .A4(n_257_76_12020), .ZN(n_257_76_12318));
   NAND3_X1 i_257_76_12340 (.A1(n_257_76_12295), .A2(n_257_76_12018), .A3(
      n_257_76_11970), .ZN(n_257_76_12319));
   NOR2_X1 i_257_76_12341 (.A1(n_257_76_12318), .A2(n_257_76_12319), .ZN(
      n_257_76_12320));
   NAND2_X1 i_257_76_12342 (.A1(n_257_76_11961), .A2(n_257_76_12029), .ZN(
      n_257_76_12321));
   INV_X1 i_257_76_12343 (.A(n_257_76_12321), .ZN(n_257_76_12322));
   NAND3_X1 i_257_76_12344 (.A1(n_257_76_12320), .A2(n_257_76_12322), .A3(
      n_257_76_11968), .ZN(n_257_76_12323));
   NAND4_X1 i_257_76_12345 (.A1(n_257_76_12008), .A2(n_257_76_12300), .A3(
      n_257_76_11944), .A4(n_257_76_12026), .ZN(n_257_76_12324));
   NOR2_X1 i_257_76_12346 (.A1(n_257_76_12323), .A2(n_257_76_12324), .ZN(
      n_257_76_12325));
   NAND2_X1 i_257_76_12347 (.A1(n_257_76_12013), .A2(n_257_76_12014), .ZN(
      n_257_76_12326));
   INV_X1 i_257_76_12348 (.A(n_257_76_12326), .ZN(n_257_76_12327));
   NAND3_X1 i_257_76_12349 (.A1(n_257_76_12004), .A2(n_257_370), .A3(
      n_257_76_11976), .ZN(n_257_76_12328));
   NAND4_X1 i_257_76_12350 (.A1(n_257_76_11977), .A2(n_257_76_12005), .A3(
      n_257_76_11978), .A4(n_257_76_12010), .ZN(n_257_76_12329));
   NOR2_X1 i_257_76_12351 (.A1(n_257_76_12328), .A2(n_257_76_12329), .ZN(
      n_257_76_12330));
   NAND4_X1 i_257_76_12352 (.A1(n_257_76_12325), .A2(n_257_76_12327), .A3(
      n_257_76_12330), .A4(n_257_76_12017), .ZN(n_257_76_12331));
   NOR2_X1 i_257_76_12353 (.A1(n_257_76_12252), .A2(n_257_76_12331), .ZN(
      n_257_76_12332));
   NAND2_X1 i_257_76_12354 (.A1(n_257_76_18082), .A2(n_257_76_12332), .ZN(
      n_257_76_12333));
   NAND2_X1 i_257_76_12355 (.A1(n_257_427), .A2(n_257_76_12021), .ZN(
      n_257_76_12334));
   INV_X1 i_257_76_12356 (.A(n_257_76_12334), .ZN(n_257_76_12335));
   NAND4_X1 i_257_76_12357 (.A1(n_257_76_12020), .A2(n_257_76_12335), .A3(
      n_257_213), .A4(n_257_76_18011), .ZN(n_257_76_12336));
   INV_X1 i_257_76_12358 (.A(n_257_76_12336), .ZN(n_257_76_12337));
   NAND4_X1 i_257_76_12359 (.A1(n_257_76_11944), .A2(n_257_76_12337), .A3(
      n_257_76_12026), .A4(n_257_76_11961), .ZN(n_257_76_12338));
   NAND4_X1 i_257_76_12360 (.A1(n_257_76_12286), .A2(n_257_76_11964), .A3(
      n_257_76_11965), .A4(n_257_76_11966), .ZN(n_257_76_12339));
   NOR2_X1 i_257_76_12361 (.A1(n_257_76_12338), .A2(n_257_76_12339), .ZN(
      n_257_76_12340));
   NAND4_X1 i_257_76_12362 (.A1(n_257_76_12340), .A2(n_257_76_12014), .A3(
      n_257_76_12097), .A4(n_257_76_12189), .ZN(n_257_76_12341));
   INV_X1 i_257_76_12363 (.A(n_257_76_12341), .ZN(n_257_76_12342));
   NAND4_X1 i_257_76_12364 (.A1(n_257_76_11941), .A2(n_257_76_12342), .A3(
      n_257_76_12070), .A4(n_257_76_11943), .ZN(n_257_76_12343));
   INV_X1 i_257_76_12365 (.A(n_257_76_12343), .ZN(n_257_76_12344));
   NAND2_X1 i_257_76_12366 (.A1(n_257_76_18065), .A2(n_257_76_12344), .ZN(
      n_257_76_12345));
   NAND4_X1 i_257_76_12367 (.A1(n_257_473), .A2(n_257_76_11964), .A3(
      n_257_76_11965), .A4(n_257_76_11966), .ZN(n_257_76_12346));
   INV_X1 i_257_76_12368 (.A(n_257_76_12346), .ZN(n_257_76_12347));
   NAND2_X1 i_257_76_12369 (.A1(n_257_76_11944), .A2(n_257_451), .ZN(
      n_257_76_12348));
   INV_X1 i_257_76_12370 (.A(n_257_76_12348), .ZN(n_257_76_12349));
   NAND4_X1 i_257_76_12371 (.A1(n_257_76_12347), .A2(n_257_76_12349), .A3(
      n_257_76_11978), .A4(n_257_76_12008), .ZN(n_257_76_12350));
   NAND3_X1 i_257_76_12372 (.A1(n_257_76_12244), .A2(n_257_76_11976), .A3(
      n_257_76_11977), .ZN(n_257_76_12351));
   NOR2_X1 i_257_76_12373 (.A1(n_257_76_12350), .A2(n_257_76_12351), .ZN(
      n_257_76_12352));
   NAND2_X1 i_257_76_12374 (.A1(n_257_76_11960), .A2(n_257_76_12352), .ZN(
      n_257_76_12353));
   INV_X1 i_257_76_12375 (.A(n_257_76_12353), .ZN(n_257_76_12354));
   NAND3_X1 i_257_76_12376 (.A1(n_257_76_12354), .A2(n_257_76_11941), .A3(
      n_257_76_11943), .ZN(n_257_76_12355));
   INV_X1 i_257_76_12377 (.A(n_257_76_12355), .ZN(n_257_76_12356));
   NAND2_X1 i_257_76_12378 (.A1(n_257_76_18063), .A2(n_257_76_12356), .ZN(
      n_257_76_12357));
   NAND3_X1 i_257_76_12379 (.A1(n_257_76_12333), .A2(n_257_76_12345), .A3(
      n_257_76_12357), .ZN(n_257_76_12358));
   NAND2_X1 i_257_76_12380 (.A1(n_257_76_12021), .A2(n_257_424), .ZN(
      n_257_76_12359));
   INV_X1 i_257_76_12381 (.A(n_257_76_12359), .ZN(n_257_76_12360));
   NAND3_X1 i_257_76_12382 (.A1(n_257_76_12020), .A2(n_257_76_18011), .A3(
      n_257_76_12360), .ZN(n_257_76_12361));
   NOR2_X1 i_257_76_12383 (.A1(n_257_76_12046), .A2(n_257_76_12361), .ZN(
      n_257_76_12362));
   NAND3_X1 i_257_76_12384 (.A1(n_257_522), .A2(n_257_76_12018), .A3(
      n_257_76_11970), .ZN(n_257_76_12363));
   INV_X1 i_257_76_12385 (.A(n_257_76_12363), .ZN(n_257_76_12364));
   NAND4_X1 i_257_76_12386 (.A1(n_257_76_12362), .A2(n_257_76_12364), .A3(
      n_257_76_12026), .A4(n_257_76_11961), .ZN(n_257_76_12365));
   INV_X1 i_257_76_12387 (.A(n_257_76_12004), .ZN(n_257_76_12366));
   NOR2_X1 i_257_76_12388 (.A1(n_257_76_12365), .A2(n_257_76_12366), .ZN(
      n_257_76_12367));
   NAND4_X1 i_257_76_12389 (.A1(n_257_76_12367), .A2(n_257_76_12012), .A3(
      n_257_76_12014), .A4(n_257_76_12097), .ZN(n_257_76_12368));
   INV_X1 i_257_76_12390 (.A(n_257_76_12368), .ZN(n_257_76_12369));
   NAND4_X1 i_257_76_12391 (.A1(n_257_76_12369), .A2(n_257_76_12310), .A3(
      n_257_76_11941), .A4(n_257_76_11943), .ZN(n_257_76_12370));
   INV_X1 i_257_76_12392 (.A(n_257_76_12370), .ZN(n_257_76_12371));
   NAND2_X1 i_257_76_12393 (.A1(n_257_76_18062), .A2(n_257_76_12371), .ZN(
      n_257_76_12372));
   INV_X1 i_257_76_12394 (.A(n_257_76_12266), .ZN(n_257_76_12373));
   NAND3_X1 i_257_76_12395 (.A1(n_257_76_12010), .A2(n_257_76_12008), .A3(
      n_257_76_12300), .ZN(n_257_76_12374));
   NAND2_X1 i_257_76_12396 (.A1(n_257_76_12005), .A2(n_257_76_11978), .ZN(
      n_257_76_12375));
   NOR2_X1 i_257_76_12397 (.A1(n_257_76_12374), .A2(n_257_76_12375), .ZN(
      n_257_76_12376));
   NAND2_X1 i_257_76_12398 (.A1(n_257_76_12029), .A2(n_257_76_11964), .ZN(
      n_257_76_12377));
   INV_X1 i_257_76_12399 (.A(n_257_76_12377), .ZN(n_257_76_12378));
   NAND2_X1 i_257_76_12400 (.A1(n_257_76_11965), .A2(n_257_76_11966), .ZN(
      n_257_76_12379));
   INV_X1 i_257_76_12401 (.A(n_257_76_12379), .ZN(n_257_76_12380));
   NAND4_X1 i_257_76_12402 (.A1(n_257_76_12018), .A2(n_257_76_11970), .A3(
      n_257_76_11971), .A4(n_257_76_11972), .ZN(n_257_76_12381));
   INV_X1 i_257_76_12403 (.A(n_257_76_12381), .ZN(n_257_76_12382));
   NAND3_X1 i_257_76_12404 (.A1(n_257_76_12378), .A2(n_257_76_12380), .A3(
      n_257_76_12382), .ZN(n_257_76_12383));
   NAND2_X1 i_257_76_12405 (.A1(n_257_422), .A2(n_257_76_12021), .ZN(
      n_257_76_12384));
   INV_X1 i_257_76_12406 (.A(n_257_76_12384), .ZN(n_257_76_12385));
   NAND4_X1 i_257_76_12407 (.A1(n_257_76_12020), .A2(n_257_331), .A3(
      n_257_76_18011), .A4(n_257_76_12385), .ZN(n_257_76_12386));
   INV_X1 i_257_76_12408 (.A(n_257_76_12386), .ZN(n_257_76_12387));
   NAND4_X1 i_257_76_12409 (.A1(n_257_76_11944), .A2(n_257_76_12387), .A3(
      n_257_76_12026), .A4(n_257_76_11961), .ZN(n_257_76_12388));
   NOR2_X1 i_257_76_12410 (.A1(n_257_76_12383), .A2(n_257_76_12388), .ZN(
      n_257_76_12389));
   NAND4_X1 i_257_76_12411 (.A1(n_257_76_12373), .A2(n_257_76_12014), .A3(
      n_257_76_12376), .A4(n_257_76_12389), .ZN(n_257_76_12390));
   INV_X1 i_257_76_12412 (.A(n_257_76_12390), .ZN(n_257_76_12391));
   NAND4_X1 i_257_76_12413 (.A1(n_257_76_12391), .A2(n_257_76_11941), .A3(
      n_257_76_12310), .A4(n_257_76_11943), .ZN(n_257_76_12392));
   INV_X1 i_257_76_12414 (.A(n_257_76_12392), .ZN(n_257_76_12393));
   NAND2_X1 i_257_76_12415 (.A1(n_257_342), .A2(n_257_76_12393), .ZN(
      n_257_76_12394));
   NAND2_X1 i_257_76_12416 (.A1(n_257_76_12032), .A2(n_257_76_12365), .ZN(
      n_257_76_12395));
   INV_X1 i_257_76_12417 (.A(n_257_76_12395), .ZN(n_257_76_12396));
   NAND2_X1 i_257_76_12418 (.A1(n_257_754), .A2(n_257_76_17935), .ZN(
      n_257_76_12397));
   NAND2_X1 i_257_76_12419 (.A1(n_257_818), .A2(n_257_76_17952), .ZN(
      n_257_76_12398));
   NAND2_X1 i_257_76_12420 (.A1(n_257_76_12397), .A2(n_257_76_12398), .ZN(
      n_257_76_12399));
   NAND2_X1 i_257_76_12421 (.A1(n_257_134), .A2(n_257_76_17925), .ZN(
      n_257_76_12400));
   NAND2_X1 i_257_76_12422 (.A1(n_257_920), .A2(n_257_76_17940), .ZN(
      n_257_76_12401));
   NAND2_X1 i_257_76_12423 (.A1(n_257_650), .A2(n_257_76_17928), .ZN(
      n_257_76_12402));
   NAND3_X1 i_257_76_12424 (.A1(n_257_76_12400), .A2(n_257_76_12401), .A3(
      n_257_76_12402), .ZN(n_257_76_12403));
   NOR2_X1 i_257_76_12425 (.A1(n_257_76_12399), .A2(n_257_76_12403), .ZN(
      n_257_76_12404));
   NAND3_X1 i_257_76_12426 (.A1(n_257_438), .A2(n_257_1086), .A3(n_257_442), 
      .ZN(n_257_76_12405));
   NAND2_X1 i_257_76_12427 (.A1(n_257_722), .A2(n_257_76_15655), .ZN(
      n_257_76_12406));
   NAND3_X1 i_257_76_12428 (.A1(n_257_76_12405), .A2(n_257_76_12406), .A3(
      n_257_76_11947), .ZN(n_257_76_12407));
   INV_X1 i_257_76_12429 (.A(n_257_76_12196), .ZN(n_257_76_12408));
   NAND2_X1 i_257_76_12430 (.A1(n_257_447), .A2(n_257_76_12408), .ZN(
      n_257_76_12409));
   INV_X1 i_257_76_12431 (.A(n_257_76_12409), .ZN(n_257_76_12410));
   NOR2_X1 i_257_76_12432 (.A1(n_257_76_12407), .A2(n_257_76_12410), .ZN(
      n_257_76_12411));
   NAND2_X1 i_257_76_12433 (.A1(n_257_76_12336), .A2(n_257_76_12386), .ZN(
      n_257_76_12412));
   INV_X1 i_257_76_12434 (.A(n_257_76_12412), .ZN(n_257_76_12413));
   NAND2_X1 i_257_76_12435 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[21]), 
      .ZN(n_257_76_12414));
   NAND2_X1 i_257_76_12436 (.A1(n_257_586), .A2(n_257_428), .ZN(n_257_76_12415));
   INV_X1 i_257_76_12437 (.A(Small_Packet_Data_Size[21]), .ZN(n_257_76_12416));
   NAND3_X1 i_257_76_12438 (.A1(n_257_76_12415), .A2(n_257_76_18015), .A3(
      n_257_76_12021), .ZN(n_257_76_12417));
   OAI21_X1 i_257_76_12439 (.A(n_257_76_12414), .B1(n_257_76_12417), .B2(
      n_257_1080), .ZN(n_257_76_12418));
   INV_X1 i_257_76_12440 (.A(n_257_76_11987), .ZN(n_257_76_12419));
   NAND2_X1 i_257_76_12441 (.A1(n_257_446), .A2(n_257_76_12419), .ZN(
      n_257_76_12420));
   NAND2_X1 i_257_76_12442 (.A1(n_257_449), .A2(n_257_76_12169), .ZN(
      n_257_76_12421));
   NAND3_X1 i_257_76_12443 (.A1(n_257_76_12418), .A2(n_257_76_12420), .A3(
      n_257_76_12421), .ZN(n_257_76_12422));
   INV_X1 i_257_76_12444 (.A(n_257_76_12422), .ZN(n_257_76_12423));
   NAND3_X1 i_257_76_12445 (.A1(n_257_76_12411), .A2(n_257_76_12413), .A3(
      n_257_76_12423), .ZN(n_257_76_12424));
   NAND3_X1 i_257_76_12446 (.A1(n_257_441), .A2(n_257_984), .A3(n_257_442), 
      .ZN(n_257_76_12425));
   NAND2_X1 i_257_76_12447 (.A1(n_257_56), .A2(n_257_76_17918), .ZN(
      n_257_76_12426));
   NAND2_X1 i_257_76_12448 (.A1(n_257_882), .A2(n_257_76_17903), .ZN(
      n_257_76_12427));
   NAND4_X1 i_257_76_12449 (.A1(n_257_76_12425), .A2(n_257_76_12298), .A3(
      n_257_76_12426), .A4(n_257_76_12427), .ZN(n_257_76_12428));
   NOR2_X1 i_257_76_12450 (.A1(n_257_76_12424), .A2(n_257_76_12428), .ZN(
      n_257_76_12429));
   NAND2_X1 i_257_76_12451 (.A1(n_257_173), .A2(n_257_76_17331), .ZN(
      n_257_76_12430));
   NAND4_X1 i_257_76_12452 (.A1(n_257_76_12396), .A2(n_257_76_12404), .A3(
      n_257_76_12429), .A4(n_257_76_12430), .ZN(n_257_76_12431));
   INV_X1 i_257_76_12453 (.A(n_257_754), .ZN(n_257_76_12432));
   NAND2_X1 i_257_76_12454 (.A1(n_257_76_12432), .A2(n_257_442), .ZN(
      n_257_76_12433));
   INV_X1 i_257_76_12455 (.A(n_257_818), .ZN(n_257_76_12434));
   NAND2_X1 i_257_76_12456 (.A1(n_257_76_12434), .A2(n_257_442), .ZN(
      n_257_76_12435));
   INV_X1 i_257_76_12457 (.A(n_257_920), .ZN(n_257_76_12436));
   NAND2_X1 i_257_76_12458 (.A1(n_257_76_12436), .A2(n_257_442), .ZN(
      n_257_76_12437));
   NAND4_X1 i_257_76_12459 (.A1(n_257_76_12433), .A2(n_257_76_12435), .A3(
      n_257_76_12437), .A4(n_257_76_13029), .ZN(n_257_76_12438));
   INV_X1 i_257_76_12460 (.A(n_257_76_12010), .ZN(n_257_76_12439));
   NAND2_X1 i_257_76_12461 (.A1(n_257_76_12438), .A2(n_257_76_12439), .ZN(
      n_257_76_12440));
   NAND2_X1 i_257_76_12462 (.A1(n_257_690), .A2(n_257_76_17958), .ZN(
      n_257_76_12441));
   NAND2_X1 i_257_76_12463 (.A1(n_257_96), .A2(n_257_76_17932), .ZN(
      n_257_76_12442));
   NAND3_X1 i_257_76_12464 (.A1(n_257_76_12440), .A2(n_257_76_12441), .A3(
      n_257_76_12442), .ZN(n_257_76_12443));
   NOR2_X1 i_257_76_12465 (.A1(n_257_76_12431), .A2(n_257_76_12443), .ZN(
      n_257_76_12444));
   NAND2_X1 i_257_76_12466 (.A1(n_257_1048), .A2(n_257_76_17969), .ZN(
      n_257_76_12445));
   INV_X1 i_257_76_12467 (.A(n_257_76_12445), .ZN(n_257_76_12446));
   INV_X1 i_257_76_12468 (.A(n_257_1016), .ZN(n_257_76_12447));
   OAI21_X1 i_257_76_12469 (.A(n_257_76_12100), .B1(n_257_76_12447), .B2(
      n_257_76_17963), .ZN(n_257_76_12448));
   NOR2_X1 i_257_76_12470 (.A1(n_257_76_12446), .A2(n_257_76_12448), .ZN(
      n_257_76_12449));
   NAND4_X1 i_257_76_12471 (.A1(n_257_76_12444), .A2(n_257_76_12449), .A3(
      n_257_76_12331), .A4(n_257_76_12269), .ZN(n_257_76_12450));
   INV_X1 i_257_76_12472 (.A(n_257_76_12450), .ZN(n_257_76_12451));
   NAND3_X1 i_257_76_12473 (.A1(n_257_484), .A2(n_257_409), .A3(n_257_442), 
      .ZN(n_257_76_12452));
   INV_X1 i_257_76_12474 (.A(n_257_76_12452), .ZN(n_257_76_12453));
   NAND3_X1 i_257_76_12475 (.A1(n_257_76_12415), .A2(n_257_76_12021), .A3(
      n_257_76_12453), .ZN(n_257_76_12454));
   INV_X1 i_257_76_12476 (.A(n_257_76_12454), .ZN(n_257_76_12455));
   NAND2_X1 i_257_76_12477 (.A1(n_257_420), .A2(n_257_490), .ZN(n_257_76_12456));
   NAND3_X1 i_257_76_12478 (.A1(n_257_76_12455), .A2(n_257_76_12020), .A3(
      n_257_76_12456), .ZN(n_257_76_12457));
   NOR2_X1 i_257_76_12479 (.A1(n_257_76_12457), .A2(n_257_76_12046), .ZN(
      n_257_76_12458));
   INV_X1 i_257_76_12480 (.A(n_257_76_12319), .ZN(n_257_76_12459));
   NAND3_X1 i_257_76_12481 (.A1(n_257_76_12458), .A2(n_257_76_12380), .A3(
      n_257_76_12459), .ZN(n_257_76_12460));
   NAND4_X1 i_257_76_12482 (.A1(n_257_76_12026), .A2(n_257_76_11961), .A3(
      n_257_76_12029), .A4(n_257_76_11964), .ZN(n_257_76_12461));
   NOR2_X1 i_257_76_12483 (.A1(n_257_76_12460), .A2(n_257_76_12461), .ZN(
      n_257_76_12462));
   NAND3_X1 i_257_76_12484 (.A1(n_257_76_12462), .A2(n_257_76_12013), .A3(
      n_257_76_12014), .ZN(n_257_76_12463));
   NAND4_X1 i_257_76_12485 (.A1(n_257_76_12010), .A2(n_257_76_12008), .A3(
      n_257_76_12300), .A4(n_257_76_11944), .ZN(n_257_76_12464));
   INV_X1 i_257_76_12486 (.A(n_257_76_12464), .ZN(n_257_76_12465));
   NAND4_X1 i_257_76_12487 (.A1(n_257_76_12305), .A2(n_257_76_12465), .A3(
      n_257_76_12306), .A4(n_257_76_12291), .ZN(n_257_76_12466));
   NOR2_X1 i_257_76_12488 (.A1(n_257_76_12463), .A2(n_257_76_12466), .ZN(
      n_257_76_12467));
   NAND4_X1 i_257_76_12489 (.A1(n_257_76_12467), .A2(n_257_76_11941), .A3(
      n_257_76_11943), .A4(n_257_76_12070), .ZN(n_257_76_12468));
   INV_X1 i_257_76_12490 (.A(n_257_76_12468), .ZN(n_257_76_12469));
   AOI21_X1 i_257_76_12491 (.A(n_257_76_12451), .B1(n_257_76_18060), .B2(
      n_257_76_12469), .ZN(n_257_76_12470));
   NAND3_X1 i_257_76_12492 (.A1(n_257_76_12372), .A2(n_257_76_12394), .A3(
      n_257_76_12470), .ZN(n_257_76_12471));
   NOR2_X1 i_257_76_12493 (.A1(n_257_76_12358), .A2(n_257_76_12471), .ZN(
      n_257_76_12472));
   NAND3_X1 i_257_76_12494 (.A1(n_257_76_12218), .A2(n_257_76_12315), .A3(
      n_257_76_12472), .ZN(n_257_76_12473));
   INV_X1 i_257_76_12495 (.A(n_257_76_12473), .ZN(n_257_76_12474));
   NAND2_X1 i_257_76_12496 (.A1(n_257_76_12153), .A2(n_257_76_12474), .ZN(n_21));
   NAND2_X1 i_257_76_12497 (.A1(n_257_1017), .A2(n_257_444), .ZN(n_257_76_12475));
   NAND2_X1 i_257_76_12498 (.A1(n_257_441), .A2(n_257_985), .ZN(n_257_76_12476));
   INV_X1 i_257_76_12499 (.A(n_257_1081), .ZN(n_257_76_12477));
   NAND2_X1 i_257_76_12500 (.A1(n_257_953), .A2(n_257_442), .ZN(n_257_76_12478));
   INV_X1 i_257_76_12501 (.A(n_257_76_12478), .ZN(n_257_76_12479));
   NAND3_X1 i_257_76_12502 (.A1(n_257_440), .A2(n_257_76_12477), .A3(
      n_257_76_12479), .ZN(n_257_76_12480));
   INV_X1 i_257_76_12503 (.A(n_257_76_12480), .ZN(n_257_76_12481));
   NAND2_X1 i_257_76_12504 (.A1(n_257_76_12476), .A2(n_257_76_12481), .ZN(
      n_257_76_12482));
   INV_X1 i_257_76_12505 (.A(n_257_76_12482), .ZN(n_257_76_12483));
   NAND2_X1 i_257_76_12506 (.A1(n_257_76_12475), .A2(n_257_76_12483), .ZN(
      n_257_76_12484));
   INV_X1 i_257_76_12507 (.A(n_257_76_12484), .ZN(n_257_76_12485));
   NAND2_X1 i_257_76_12508 (.A1(n_257_1049), .A2(n_257_443), .ZN(n_257_76_12486));
   NAND2_X1 i_257_76_12509 (.A1(n_257_76_12485), .A2(n_257_76_12486), .ZN(
      n_257_76_12487));
   INV_X1 i_257_76_12510 (.A(n_257_76_12487), .ZN(n_257_76_12488));
   NAND2_X1 i_257_76_12511 (.A1(n_257_17), .A2(n_257_76_12488), .ZN(
      n_257_76_12489));
   NOR2_X1 i_257_76_12512 (.A1(n_257_1081), .A2(n_257_76_17412), .ZN(
      n_257_76_12490));
   INV_X1 i_257_76_12513 (.A(n_257_76_12490), .ZN(n_257_76_12491));
   NOR2_X1 i_257_76_12514 (.A1(n_257_76_12491), .A2(n_257_76_15197), .ZN(
      n_257_76_12492));
   NAND2_X1 i_257_76_12515 (.A1(n_257_1049), .A2(n_257_76_12492), .ZN(
      n_257_76_12493));
   INV_X1 i_257_76_12516 (.A(n_257_76_12493), .ZN(n_257_76_12494));
   NAND2_X1 i_257_76_12517 (.A1(n_257_76_18072), .A2(n_257_76_12494), .ZN(
      n_257_76_12495));
   NAND2_X1 i_257_76_12518 (.A1(n_257_449), .A2(n_257_897), .ZN(n_257_76_12496));
   NAND2_X1 i_257_76_12519 (.A1(n_257_447), .A2(n_257_787), .ZN(n_257_76_12497));
   NAND2_X1 i_257_76_12520 (.A1(n_257_883), .A2(n_257_445), .ZN(n_257_76_12498));
   NAND3_X1 i_257_76_12521 (.A1(n_257_76_12496), .A2(n_257_76_12497), .A3(
      n_257_76_12498), .ZN(n_257_76_12499));
   INV_X1 i_257_76_12522 (.A(n_257_76_12499), .ZN(n_257_76_12500));
   NAND2_X1 i_257_76_12523 (.A1(n_257_446), .A2(n_257_851), .ZN(n_257_76_12501));
   NAND2_X1 i_257_76_12524 (.A1(n_257_651), .A2(n_257_76_12501), .ZN(
      n_257_76_12502));
   INV_X1 i_257_76_12525 (.A(n_257_76_12502), .ZN(n_257_76_12503));
   NAND2_X1 i_257_76_12526 (.A1(n_257_438), .A2(n_257_1087), .ZN(n_257_76_12504));
   NAND2_X1 i_257_76_12527 (.A1(n_257_723), .A2(n_257_435), .ZN(n_257_76_12505));
   NAND3_X1 i_257_76_12528 (.A1(n_257_76_12504), .A2(n_257_76_12505), .A3(
      n_257_450), .ZN(n_257_76_12506));
   NAND2_X1 i_257_76_12529 (.A1(n_257_440), .A2(n_257_953), .ZN(n_257_76_12507));
   NAND2_X1 i_257_76_12530 (.A1(n_257_76_12507), .A2(n_257_76_12490), .ZN(
      n_257_76_12508));
   NOR2_X1 i_257_76_12531 (.A1(n_257_76_12506), .A2(n_257_76_12508), .ZN(
      n_257_76_12509));
   NAND3_X1 i_257_76_12532 (.A1(n_257_76_12500), .A2(n_257_76_12503), .A3(
      n_257_76_12509), .ZN(n_257_76_12510));
   NAND2_X1 i_257_76_12533 (.A1(n_257_755), .A2(n_257_436), .ZN(n_257_76_12511));
   NAND2_X1 i_257_76_12534 (.A1(n_257_921), .A2(n_257_439), .ZN(n_257_76_12512));
   NAND2_X1 i_257_76_12535 (.A1(n_257_819), .A2(n_257_437), .ZN(n_257_76_12513));
   NAND4_X1 i_257_76_12536 (.A1(n_257_76_12511), .A2(n_257_76_12476), .A3(
      n_257_76_12512), .A4(n_257_76_12513), .ZN(n_257_76_12514));
   NOR2_X1 i_257_76_12537 (.A1(n_257_76_12510), .A2(n_257_76_12514), .ZN(
      n_257_76_12515));
   NAND2_X1 i_257_76_12538 (.A1(n_257_691), .A2(n_257_448), .ZN(n_257_76_12516));
   NAND3_X1 i_257_76_12539 (.A1(n_257_76_12515), .A2(n_257_76_12475), .A3(
      n_257_76_12516), .ZN(n_257_76_12517));
   INV_X1 i_257_76_12540 (.A(n_257_76_12486), .ZN(n_257_76_12518));
   NOR2_X1 i_257_76_12541 (.A1(n_257_76_12517), .A2(n_257_76_12518), .ZN(
      n_257_76_12519));
   NAND2_X1 i_257_76_12542 (.A1(n_257_28), .A2(n_257_76_12519), .ZN(
      n_257_76_12520));
   NAND3_X1 i_257_76_12543 (.A1(n_257_76_12489), .A2(n_257_76_12495), .A3(
      n_257_76_12520), .ZN(n_257_76_12521));
   NAND2_X1 i_257_76_12544 (.A1(n_257_76_12476), .A2(n_257_76_12512), .ZN(
      n_257_76_12522));
   NAND2_X1 i_257_76_12545 (.A1(n_257_446), .A2(n_257_76_12507), .ZN(
      n_257_76_12523));
   INV_X1 i_257_76_12546 (.A(n_257_76_12523), .ZN(n_257_76_12524));
   NAND2_X1 i_257_76_12547 (.A1(n_257_851), .A2(n_257_442), .ZN(n_257_76_12525));
   NOR2_X1 i_257_76_12548 (.A1(n_257_1081), .A2(n_257_76_12525), .ZN(
      n_257_76_12526));
   NAND2_X1 i_257_76_12549 (.A1(n_257_76_12504), .A2(n_257_76_12526), .ZN(
      n_257_76_12527));
   INV_X1 i_257_76_12550 (.A(n_257_76_12527), .ZN(n_257_76_12528));
   NAND3_X1 i_257_76_12551 (.A1(n_257_76_12524), .A2(n_257_76_12528), .A3(
      n_257_76_12498), .ZN(n_257_76_12529));
   NOR2_X1 i_257_76_12552 (.A1(n_257_76_12522), .A2(n_257_76_12529), .ZN(
      n_257_76_12530));
   NAND2_X1 i_257_76_12553 (.A1(n_257_76_12475), .A2(n_257_76_12530), .ZN(
      n_257_76_12531));
   INV_X1 i_257_76_12554 (.A(n_257_76_12531), .ZN(n_257_76_12532));
   NAND2_X1 i_257_76_12555 (.A1(n_257_76_12532), .A2(n_257_76_12486), .ZN(
      n_257_76_12533));
   INV_X1 i_257_76_12556 (.A(n_257_76_12533), .ZN(n_257_76_12534));
   NAND2_X1 i_257_76_12557 (.A1(n_257_76_18070), .A2(n_257_76_12534), .ZN(
      n_257_76_12535));
   NAND3_X1 i_257_76_12558 (.A1(n_257_76_12507), .A2(n_257_76_12490), .A3(
      n_257_439), .ZN(n_257_76_12536));
   INV_X1 i_257_76_12559 (.A(n_257_76_12536), .ZN(n_257_76_12537));
   NAND3_X1 i_257_76_12560 (.A1(n_257_76_12476), .A2(n_257_921), .A3(
      n_257_76_12537), .ZN(n_257_76_12538));
   INV_X1 i_257_76_12561 (.A(n_257_76_12538), .ZN(n_257_76_12539));
   NAND2_X1 i_257_76_12562 (.A1(n_257_76_12475), .A2(n_257_76_12539), .ZN(
      n_257_76_12540));
   INV_X1 i_257_76_12563 (.A(n_257_76_12540), .ZN(n_257_76_12541));
   NAND2_X1 i_257_76_12564 (.A1(n_257_76_12541), .A2(n_257_76_12486), .ZN(
      n_257_76_12542));
   INV_X1 i_257_76_12565 (.A(n_257_76_12542), .ZN(n_257_76_12543));
   NAND2_X1 i_257_76_12566 (.A1(n_257_76_18084), .A2(n_257_76_12543), .ZN(
      n_257_76_12544));
   NAND3_X1 i_257_76_12567 (.A1(n_257_76_12512), .A2(n_257_76_12513), .A3(
      n_257_76_12501), .ZN(n_257_76_12545));
   NAND2_X1 i_257_76_12568 (.A1(n_257_76_12507), .A2(n_257_76_12504), .ZN(
      n_257_76_12546));
   INV_X1 i_257_76_12569 (.A(n_257_76_12546), .ZN(n_257_76_12547));
   NAND4_X1 i_257_76_12570 (.A1(n_257_76_12547), .A2(n_257_76_12496), .A3(
      n_257_76_12497), .A4(n_257_76_12498), .ZN(n_257_76_12548));
   NOR2_X1 i_257_76_12571 (.A1(n_257_76_12545), .A2(n_257_76_12548), .ZN(
      n_257_76_12549));
   NAND2_X1 i_257_76_12572 (.A1(n_257_555), .A2(n_257_426), .ZN(n_257_76_12550));
   NAND2_X1 i_257_76_12573 (.A1(n_257_135), .A2(n_257_430), .ZN(n_257_76_12551));
   NAND2_X1 i_257_76_12574 (.A1(n_257_651), .A2(n_257_450), .ZN(n_257_76_12552));
   NAND3_X1 i_257_76_12575 (.A1(n_257_76_12550), .A2(n_257_76_12551), .A3(
      n_257_76_12552), .ZN(n_257_76_12553));
   INV_X1 i_257_76_12576 (.A(n_257_76_12553), .ZN(n_257_76_12554));
   NAND2_X1 i_257_76_12577 (.A1(n_257_97), .A2(n_257_431), .ZN(n_257_76_12555));
   NAND2_X1 i_257_76_12578 (.A1(n_257_474), .A2(n_257_451), .ZN(n_257_76_12556));
   NAND3_X1 i_257_76_12579 (.A1(n_257_76_12511), .A2(n_257_76_12476), .A3(
      n_257_76_12556), .ZN(n_257_76_12557));
   INV_X1 i_257_76_12580 (.A(n_257_76_12557), .ZN(n_257_76_12558));
   NAND4_X1 i_257_76_12581 (.A1(n_257_76_12549), .A2(n_257_76_12554), .A3(
      n_257_76_12555), .A4(n_257_76_12558), .ZN(n_257_76_12559));
   NAND2_X1 i_257_76_12582 (.A1(n_257_174), .A2(n_257_429), .ZN(n_257_76_12560));
   NAND2_X1 i_257_76_12583 (.A1(n_257_214), .A2(n_257_427), .ZN(n_257_76_12561));
   NAND2_X1 i_257_76_12584 (.A1(n_257_76_12505), .A2(n_257_76_12561), .ZN(
      n_257_76_12562));
   NAND2_X1 i_257_76_12585 (.A1(n_257_432), .A2(n_257_619), .ZN(n_257_76_12563));
   NAND2_X1 i_257_76_12586 (.A1(n_257_76_12563), .A2(n_257_423), .ZN(
      n_257_76_12564));
   INV_X1 i_257_76_12587 (.A(n_257_76_12564), .ZN(n_257_76_12565));
   NAND3_X1 i_257_76_12588 (.A1(n_257_76_12565), .A2(n_257_76_12477), .A3(
      n_257_76_18008), .ZN(n_257_76_12566));
   NOR2_X1 i_257_76_12589 (.A1(n_257_76_12562), .A2(n_257_76_12566), .ZN(
      n_257_76_12567));
   NAND2_X1 i_257_76_12590 (.A1(n_257_523), .A2(n_257_424), .ZN(n_257_76_12568));
   NAND2_X1 i_257_76_12591 (.A1(n_257_76_12568), .A2(n_257_294), .ZN(
      n_257_76_12569));
   INV_X1 i_257_76_12592 (.A(n_257_76_12569), .ZN(n_257_76_12570));
   NAND2_X1 i_257_76_12593 (.A1(n_257_57), .A2(n_257_433), .ZN(n_257_76_12571));
   NAND3_X1 i_257_76_12594 (.A1(n_257_76_12567), .A2(n_257_76_12570), .A3(
      n_257_76_12571), .ZN(n_257_76_12572));
   INV_X1 i_257_76_12595 (.A(n_257_76_12572), .ZN(n_257_76_12573));
   NAND3_X1 i_257_76_12596 (.A1(n_257_76_12516), .A2(n_257_76_12560), .A3(
      n_257_76_12573), .ZN(n_257_76_12574));
   NOR2_X1 i_257_76_12597 (.A1(n_257_76_12559), .A2(n_257_76_12574), .ZN(
      n_257_76_12575));
   NAND2_X1 i_257_76_12598 (.A1(n_257_254), .A2(n_257_425), .ZN(n_257_76_12576));
   NAND2_X1 i_257_76_12599 (.A1(n_257_76_12576), .A2(n_257_76_12475), .ZN(
      n_257_76_12577));
   INV_X1 i_257_76_12600 (.A(n_257_76_12577), .ZN(n_257_76_12578));
   NAND3_X1 i_257_76_12601 (.A1(n_257_76_12575), .A2(n_257_76_12578), .A3(
      n_257_76_12486), .ZN(n_257_76_12579));
   INV_X1 i_257_76_12602 (.A(n_257_76_12579), .ZN(n_257_76_12580));
   NAND2_X1 i_257_76_12603 (.A1(n_257_76_18066), .A2(n_257_76_12580), .ZN(
      n_257_76_12581));
   NAND3_X1 i_257_76_12604 (.A1(n_257_76_12535), .A2(n_257_76_12544), .A3(
      n_257_76_12581), .ZN(n_257_76_12582));
   NOR2_X1 i_257_76_12605 (.A1(n_257_76_12521), .A2(n_257_76_12582), .ZN(
      n_257_76_12583));
   NAND2_X1 i_257_76_12606 (.A1(n_257_985), .A2(n_257_76_12490), .ZN(
      n_257_76_12584));
   NOR2_X1 i_257_76_12607 (.A1(n_257_76_13147), .A2(n_257_76_12584), .ZN(
      n_257_76_12585));
   NAND2_X1 i_257_76_12608 (.A1(n_257_76_12475), .A2(n_257_76_12585), .ZN(
      n_257_76_12586));
   INV_X1 i_257_76_12609 (.A(n_257_76_12586), .ZN(n_257_76_12587));
   NAND2_X1 i_257_76_12610 (.A1(n_257_76_12587), .A2(n_257_76_12486), .ZN(
      n_257_76_12588));
   INV_X1 i_257_76_12611 (.A(n_257_76_12588), .ZN(n_257_76_12589));
   NAND2_X1 i_257_76_12612 (.A1(n_257_76_18071), .A2(n_257_76_12589), .ZN(
      n_257_76_12590));
   NAND3_X1 i_257_76_12613 (.A1(n_257_76_12477), .A2(n_257_723), .A3(
      n_257_76_15655), .ZN(n_257_76_12591));
   INV_X1 i_257_76_12614 (.A(n_257_76_12591), .ZN(n_257_76_12592));
   NAND3_X1 i_257_76_12615 (.A1(n_257_76_12592), .A2(n_257_76_12507), .A3(
      n_257_76_12504), .ZN(n_257_76_12593));
   INV_X1 i_257_76_12616 (.A(n_257_76_12593), .ZN(n_257_76_12594));
   NAND4_X1 i_257_76_12617 (.A1(n_257_76_12594), .A2(n_257_76_12501), .A3(
      n_257_76_12497), .A4(n_257_76_12498), .ZN(n_257_76_12595));
   NOR2_X1 i_257_76_12618 (.A1(n_257_76_12514), .A2(n_257_76_12595), .ZN(
      n_257_76_12596));
   NAND2_X1 i_257_76_12619 (.A1(n_257_76_12475), .A2(n_257_76_12596), .ZN(
      n_257_76_12597));
   INV_X1 i_257_76_12620 (.A(n_257_76_12597), .ZN(n_257_76_12598));
   NAND2_X1 i_257_76_12621 (.A1(n_257_76_12598), .A2(n_257_76_12486), .ZN(
      n_257_76_12599));
   INV_X1 i_257_76_12622 (.A(n_257_76_12599), .ZN(n_257_76_12600));
   NAND2_X1 i_257_76_12623 (.A1(n_257_76_18078), .A2(n_257_76_12600), .ZN(
      n_257_76_12601));
   NAND3_X1 i_257_76_12624 (.A1(n_257_76_12551), .A2(n_257_76_12552), .A3(
      n_257_76_12511), .ZN(n_257_76_12602));
   NAND3_X1 i_257_76_12625 (.A1(n_257_76_12476), .A2(n_257_76_12556), .A3(
      n_257_76_12512), .ZN(n_257_76_12603));
   NOR2_X1 i_257_76_12626 (.A1(n_257_76_12602), .A2(n_257_76_12603), .ZN(
      n_257_76_12604));
   NAND3_X1 i_257_76_12627 (.A1(n_257_76_12497), .A2(n_257_76_12571), .A3(
      n_257_76_12498), .ZN(n_257_76_12605));
   INV_X1 i_257_76_12628 (.A(n_257_76_12605), .ZN(n_257_76_12606));
   NAND2_X1 i_257_76_12629 (.A1(n_257_428), .A2(n_257_442), .ZN(n_257_76_12607));
   INV_X1 i_257_76_12630 (.A(n_257_76_12607), .ZN(n_257_76_12608));
   NAND3_X1 i_257_76_12631 (.A1(n_257_76_12563), .A2(n_257_587), .A3(
      n_257_76_12608), .ZN(n_257_76_12609));
   NOR2_X1 i_257_76_12632 (.A1(n_257_76_12609), .A2(n_257_1081), .ZN(
      n_257_76_12610));
   NAND4_X1 i_257_76_12633 (.A1(n_257_76_12610), .A2(n_257_76_12507), .A3(
      n_257_76_12504), .A4(n_257_76_12505), .ZN(n_257_76_12611));
   INV_X1 i_257_76_12634 (.A(n_257_76_12611), .ZN(n_257_76_12612));
   NAND2_X1 i_257_76_12635 (.A1(n_257_76_12501), .A2(n_257_76_12496), .ZN(
      n_257_76_12613));
   INV_X1 i_257_76_12636 (.A(n_257_76_12613), .ZN(n_257_76_12614));
   NAND4_X1 i_257_76_12637 (.A1(n_257_76_12606), .A2(n_257_76_12612), .A3(
      n_257_76_12614), .A4(n_257_76_12513), .ZN(n_257_76_12615));
   INV_X1 i_257_76_12638 (.A(n_257_76_12615), .ZN(n_257_76_12616));
   NAND4_X1 i_257_76_12639 (.A1(n_257_76_12604), .A2(n_257_76_12616), .A3(
      n_257_76_12560), .A4(n_257_76_12555), .ZN(n_257_76_12617));
   INV_X1 i_257_76_12640 (.A(n_257_76_12617), .ZN(n_257_76_12618));
   NAND2_X1 i_257_76_12641 (.A1(n_257_76_12475), .A2(n_257_76_12516), .ZN(
      n_257_76_12619));
   INV_X1 i_257_76_12642 (.A(n_257_76_12619), .ZN(n_257_76_12620));
   NAND3_X1 i_257_76_12643 (.A1(n_257_76_12618), .A2(n_257_76_12620), .A3(
      n_257_76_12486), .ZN(n_257_76_12621));
   INV_X1 i_257_76_12644 (.A(n_257_76_12621), .ZN(n_257_76_12622));
   NAND2_X1 i_257_76_12645 (.A1(n_257_76_18074), .A2(n_257_76_12622), .ZN(
      n_257_76_12623));
   NAND3_X1 i_257_76_12646 (.A1(n_257_76_12590), .A2(n_257_76_12601), .A3(
      n_257_76_12623), .ZN(n_257_76_12624));
   NAND2_X1 i_257_76_12647 (.A1(n_257_1081), .A2(n_257_442), .ZN(n_257_76_12625));
   INV_X1 i_257_76_12648 (.A(n_257_76_12625), .ZN(n_257_76_12626));
   NAND2_X1 i_257_76_12649 (.A1(n_257_13), .A2(n_257_76_12626), .ZN(
      n_257_76_12627));
   NAND3_X1 i_257_76_12650 (.A1(n_257_76_12504), .A2(n_257_883), .A3(n_257_445), 
      .ZN(n_257_76_12628));
   NOR2_X1 i_257_76_12651 (.A1(n_257_76_12628), .A2(n_257_76_12508), .ZN(
      n_257_76_12629));
   NAND3_X1 i_257_76_12652 (.A1(n_257_76_12629), .A2(n_257_76_12476), .A3(
      n_257_76_12512), .ZN(n_257_76_12630));
   INV_X1 i_257_76_12653 (.A(n_257_76_12630), .ZN(n_257_76_12631));
   NAND2_X1 i_257_76_12654 (.A1(n_257_76_12475), .A2(n_257_76_12631), .ZN(
      n_257_76_12632));
   INV_X1 i_257_76_12655 (.A(n_257_76_12632), .ZN(n_257_76_12633));
   NAND2_X1 i_257_76_12656 (.A1(n_257_76_12633), .A2(n_257_76_12486), .ZN(
      n_257_76_12634));
   INV_X1 i_257_76_12657 (.A(n_257_76_12634), .ZN(n_257_76_12635));
   NAND2_X1 i_257_76_12658 (.A1(n_257_76_18077), .A2(n_257_76_12635), .ZN(
      n_257_76_12636));
   NAND2_X1 i_257_76_12659 (.A1(n_257_76_12627), .A2(n_257_76_12636), .ZN(
      n_257_76_12637));
   NOR2_X1 i_257_76_12660 (.A1(n_257_76_12624), .A2(n_257_76_12637), .ZN(
      n_257_76_12638));
   INV_X1 i_257_76_12661 (.A(n_257_76_12475), .ZN(n_257_76_12639));
   NAND4_X1 i_257_76_12662 (.A1(n_257_76_12496), .A2(n_257_76_12497), .A3(
      n_257_76_12571), .A4(n_257_76_12498), .ZN(n_257_76_12640));
   INV_X1 i_257_76_12663 (.A(n_257_76_12562), .ZN(n_257_76_12641));
   NAND2_X1 i_257_76_12664 (.A1(n_257_76_12563), .A2(n_257_426), .ZN(
      n_257_76_12642));
   INV_X1 i_257_76_12665 (.A(n_257_76_12642), .ZN(n_257_76_12643));
   NAND3_X1 i_257_76_12666 (.A1(n_257_76_12643), .A2(n_257_76_12477), .A3(
      n_257_76_18008), .ZN(n_257_76_12644));
   INV_X1 i_257_76_12667 (.A(n_257_76_12644), .ZN(n_257_76_12645));
   NAND4_X1 i_257_76_12668 (.A1(n_257_76_12641), .A2(n_257_76_12645), .A3(
      n_257_76_12507), .A4(n_257_76_12504), .ZN(n_257_76_12646));
   NOR2_X1 i_257_76_12669 (.A1(n_257_76_12640), .A2(n_257_76_12646), .ZN(
      n_257_76_12647));
   INV_X1 i_257_76_12670 (.A(n_257_76_12602), .ZN(n_257_76_12648));
   NAND4_X1 i_257_76_12671 (.A1(n_257_76_12512), .A2(n_257_76_12513), .A3(
      n_257_555), .A4(n_257_76_12501), .ZN(n_257_76_12649));
   INV_X1 i_257_76_12672 (.A(n_257_76_12649), .ZN(n_257_76_12650));
   NAND3_X1 i_257_76_12673 (.A1(n_257_76_12647), .A2(n_257_76_12648), .A3(
      n_257_76_12650), .ZN(n_257_76_12651));
   NOR2_X1 i_257_76_12674 (.A1(n_257_76_12639), .A2(n_257_76_12651), .ZN(
      n_257_76_12652));
   NAND2_X1 i_257_76_12675 (.A1(n_257_76_12476), .A2(n_257_76_12556), .ZN(
      n_257_76_12653));
   INV_X1 i_257_76_12676 (.A(n_257_76_12653), .ZN(n_257_76_12654));
   NAND2_X1 i_257_76_12677 (.A1(n_257_76_12555), .A2(n_257_76_12654), .ZN(
      n_257_76_12655));
   INV_X1 i_257_76_12678 (.A(n_257_76_12655), .ZN(n_257_76_12656));
   NAND3_X1 i_257_76_12679 (.A1(n_257_76_12656), .A2(n_257_76_12516), .A3(
      n_257_76_12560), .ZN(n_257_76_12657));
   INV_X1 i_257_76_12680 (.A(n_257_76_12657), .ZN(n_257_76_12658));
   NAND3_X1 i_257_76_12681 (.A1(n_257_76_12652), .A2(n_257_76_12486), .A3(
      n_257_76_12658), .ZN(n_257_76_12659));
   INV_X1 i_257_76_12682 (.A(n_257_76_12659), .ZN(n_257_76_12660));
   NAND2_X1 i_257_76_12683 (.A1(n_257_76_18076), .A2(n_257_76_12660), .ZN(
      n_257_76_12661));
   NAND2_X1 i_257_76_12684 (.A1(n_257_755), .A2(n_257_76_12501), .ZN(
      n_257_76_12662));
   INV_X1 i_257_76_12685 (.A(n_257_76_12662), .ZN(n_257_76_12663));
   NAND2_X1 i_257_76_12686 (.A1(n_257_76_12497), .A2(n_257_76_12498), .ZN(
      n_257_76_12664));
   INV_X1 i_257_76_12687 (.A(n_257_76_12664), .ZN(n_257_76_12665));
   NOR2_X1 i_257_76_12688 (.A1(n_257_1081), .A2(n_257_76_17934), .ZN(
      n_257_76_12666));
   NAND3_X1 i_257_76_12689 (.A1(n_257_76_12507), .A2(n_257_76_12504), .A3(
      n_257_76_12666), .ZN(n_257_76_12667));
   INV_X1 i_257_76_12690 (.A(n_257_76_12667), .ZN(n_257_76_12668));
   NAND3_X1 i_257_76_12691 (.A1(n_257_76_12663), .A2(n_257_76_12665), .A3(
      n_257_76_12668), .ZN(n_257_76_12669));
   NAND3_X1 i_257_76_12692 (.A1(n_257_76_12476), .A2(n_257_76_12512), .A3(
      n_257_76_12513), .ZN(n_257_76_12670));
   NOR2_X1 i_257_76_12693 (.A1(n_257_76_12669), .A2(n_257_76_12670), .ZN(
      n_257_76_12671));
   NAND2_X1 i_257_76_12694 (.A1(n_257_76_12475), .A2(n_257_76_12671), .ZN(
      n_257_76_12672));
   INV_X1 i_257_76_12695 (.A(n_257_76_12672), .ZN(n_257_76_12673));
   NAND2_X1 i_257_76_12696 (.A1(n_257_76_12673), .A2(n_257_76_12486), .ZN(
      n_257_76_12674));
   INV_X1 i_257_76_12697 (.A(n_257_76_12674), .ZN(n_257_76_12675));
   NAND2_X1 i_257_76_12698 (.A1(n_257_76_18069), .A2(n_257_76_12675), .ZN(
      n_257_76_12676));
   NAND2_X1 i_257_76_12699 (.A1(n_257_619), .A2(n_257_442), .ZN(n_257_76_12677));
   INV_X1 i_257_76_12700 (.A(n_257_76_12677), .ZN(n_257_76_12678));
   NAND2_X1 i_257_76_12701 (.A1(n_257_76_12678), .A2(n_257_432), .ZN(
      n_257_76_12679));
   NOR2_X1 i_257_76_12702 (.A1(n_257_1081), .A2(n_257_76_12679), .ZN(
      n_257_76_12680));
   NAND2_X1 i_257_76_12703 (.A1(n_257_76_12505), .A2(n_257_76_12680), .ZN(
      n_257_76_12681));
   INV_X1 i_257_76_12704 (.A(n_257_76_12681), .ZN(n_257_76_12682));
   NAND4_X1 i_257_76_12705 (.A1(n_257_76_12547), .A2(n_257_76_12682), .A3(
      n_257_76_12571), .A4(n_257_76_12498), .ZN(n_257_76_12683));
   NAND3_X1 i_257_76_12706 (.A1(n_257_76_12501), .A2(n_257_76_12496), .A3(
      n_257_76_12497), .ZN(n_257_76_12684));
   NOR2_X1 i_257_76_12707 (.A1(n_257_76_12683), .A2(n_257_76_12684), .ZN(
      n_257_76_12685));
   NAND3_X1 i_257_76_12708 (.A1(n_257_76_12552), .A2(n_257_76_12511), .A3(
      n_257_76_12476), .ZN(n_257_76_12686));
   INV_X1 i_257_76_12709 (.A(n_257_76_12686), .ZN(n_257_76_12687));
   NAND3_X1 i_257_76_12710 (.A1(n_257_76_12556), .A2(n_257_76_12512), .A3(
      n_257_76_12513), .ZN(n_257_76_12688));
   INV_X1 i_257_76_12711 (.A(n_257_76_12688), .ZN(n_257_76_12689));
   NAND3_X1 i_257_76_12712 (.A1(n_257_76_12685), .A2(n_257_76_12687), .A3(
      n_257_76_12689), .ZN(n_257_76_12690));
   INV_X1 i_257_76_12713 (.A(n_257_76_12690), .ZN(n_257_76_12691));
   NAND3_X1 i_257_76_12714 (.A1(n_257_76_12691), .A2(n_257_76_12475), .A3(
      n_257_76_12516), .ZN(n_257_76_12692));
   NOR2_X1 i_257_76_12715 (.A1(n_257_76_12692), .A2(n_257_76_12518), .ZN(
      n_257_76_12693));
   NAND2_X1 i_257_76_12716 (.A1(n_257_68), .A2(n_257_76_12693), .ZN(
      n_257_76_12694));
   NAND3_X1 i_257_76_12717 (.A1(n_257_76_12661), .A2(n_257_76_12676), .A3(
      n_257_76_12694), .ZN(n_257_76_12695));
   NOR2_X1 i_257_76_12718 (.A1(n_257_1081), .A2(n_257_76_17951), .ZN(
      n_257_76_12696));
   NAND3_X1 i_257_76_12719 (.A1(n_257_76_12507), .A2(n_257_76_12504), .A3(
      n_257_76_12696), .ZN(n_257_76_12697));
   INV_X1 i_257_76_12720 (.A(n_257_76_12697), .ZN(n_257_76_12698));
   NAND4_X1 i_257_76_12721 (.A1(n_257_76_12698), .A2(n_257_76_12501), .A3(
      n_257_819), .A4(n_257_76_12498), .ZN(n_257_76_12699));
   NOR2_X1 i_257_76_12722 (.A1(n_257_76_12699), .A2(n_257_76_12522), .ZN(
      n_257_76_12700));
   NAND2_X1 i_257_76_12723 (.A1(n_257_76_12475), .A2(n_257_76_12700), .ZN(
      n_257_76_12701));
   INV_X1 i_257_76_12724 (.A(n_257_76_12701), .ZN(n_257_76_12702));
   NAND2_X1 i_257_76_12725 (.A1(n_257_76_12702), .A2(n_257_76_12486), .ZN(
      n_257_76_12703));
   INV_X1 i_257_76_12726 (.A(n_257_76_12703), .ZN(n_257_76_12704));
   NAND2_X1 i_257_76_12727 (.A1(n_257_22), .A2(n_257_76_12704), .ZN(
      n_257_76_12705));
   NAND2_X1 i_257_76_12728 (.A1(n_257_444), .A2(n_257_76_12490), .ZN(
      n_257_76_12706));
   INV_X1 i_257_76_12729 (.A(n_257_76_12706), .ZN(n_257_76_12707));
   NAND2_X1 i_257_76_12730 (.A1(n_257_1017), .A2(n_257_76_12707), .ZN(
      n_257_76_12708));
   INV_X1 i_257_76_12731 (.A(n_257_76_12708), .ZN(n_257_76_12709));
   NAND2_X1 i_257_76_12732 (.A1(n_257_76_12486), .A2(n_257_76_12709), .ZN(
      n_257_76_12710));
   INV_X1 i_257_76_12733 (.A(n_257_76_12710), .ZN(n_257_76_12711));
   NAND2_X1 i_257_76_12734 (.A1(n_257_76_18075), .A2(n_257_76_12711), .ZN(
      n_257_76_12712));
   NAND2_X1 i_257_76_12735 (.A1(n_257_76_12705), .A2(n_257_76_12712), .ZN(
      n_257_76_12713));
   NOR2_X1 i_257_76_12736 (.A1(n_257_76_12695), .A2(n_257_76_12713), .ZN(
      n_257_76_12714));
   NAND3_X1 i_257_76_12737 (.A1(n_257_76_12583), .A2(n_257_76_12638), .A3(
      n_257_76_12714), .ZN(n_257_76_12715));
   INV_X1 i_257_76_12738 (.A(n_257_76_12715), .ZN(n_257_76_12716));
   NOR2_X1 i_257_76_12739 (.A1(n_257_1081), .A2(n_257_76_17633), .ZN(
      n_257_76_12717));
   NAND3_X1 i_257_76_12740 (.A1(n_257_76_12717), .A2(n_257_57), .A3(
      n_257_76_12505), .ZN(n_257_76_12718));
   INV_X1 i_257_76_12741 (.A(n_257_76_12718), .ZN(n_257_76_12719));
   NAND3_X1 i_257_76_12742 (.A1(n_257_76_12719), .A2(n_257_76_12547), .A3(
      n_257_76_12498), .ZN(n_257_76_12720));
   NOR2_X1 i_257_76_12743 (.A1(n_257_76_12720), .A2(n_257_76_12684), .ZN(
      n_257_76_12721));
   NAND3_X1 i_257_76_12744 (.A1(n_257_76_12721), .A2(n_257_76_12687), .A3(
      n_257_76_12689), .ZN(n_257_76_12722));
   INV_X1 i_257_76_12745 (.A(n_257_76_12722), .ZN(n_257_76_12723));
   NAND3_X1 i_257_76_12746 (.A1(n_257_76_12723), .A2(n_257_76_12475), .A3(
      n_257_76_12516), .ZN(n_257_76_12724));
   NOR2_X1 i_257_76_12747 (.A1(n_257_76_12724), .A2(n_257_76_12518), .ZN(
      n_257_76_12725));
   NAND2_X1 i_257_76_12748 (.A1(n_257_76_18081), .A2(n_257_76_12725), .ZN(
      n_257_76_12726));
   NAND2_X1 i_257_76_12749 (.A1(n_257_76_12501), .A2(n_257_76_12497), .ZN(
      n_257_76_12727));
   INV_X1 i_257_76_12750 (.A(n_257_76_12727), .ZN(n_257_76_12728));
   NOR2_X1 i_257_76_12751 (.A1(n_257_1081), .A2(n_257_76_17119), .ZN(
      n_257_76_12729));
   NAND4_X1 i_257_76_12752 (.A1(n_257_76_12507), .A2(n_257_76_12504), .A3(
      n_257_76_12729), .A4(n_257_76_12505), .ZN(n_257_76_12730));
   INV_X1 i_257_76_12753 (.A(n_257_76_12730), .ZN(n_257_76_12731));
   NAND2_X1 i_257_76_12754 (.A1(n_257_76_12498), .A2(n_257_449), .ZN(
      n_257_76_12732));
   INV_X1 i_257_76_12755 (.A(n_257_76_12732), .ZN(n_257_76_12733));
   NAND3_X1 i_257_76_12756 (.A1(n_257_76_12728), .A2(n_257_76_12731), .A3(
      n_257_76_12733), .ZN(n_257_76_12734));
   NOR2_X1 i_257_76_12757 (.A1(n_257_76_12514), .A2(n_257_76_12734), .ZN(
      n_257_76_12735));
   NAND3_X1 i_257_76_12758 (.A1(n_257_76_12475), .A2(n_257_76_12735), .A3(
      n_257_76_12516), .ZN(n_257_76_12736));
   NOR2_X1 i_257_76_12759 (.A1(n_257_76_12736), .A2(n_257_76_12518), .ZN(
      n_257_76_12737));
   NAND2_X1 i_257_76_12760 (.A1(n_257_76_18083), .A2(n_257_76_12737), .ZN(
      n_257_76_12738));
   INV_X1 i_257_76_12761 (.A(n_257_619), .ZN(n_257_76_12739));
   NAND2_X1 i_257_76_12762 (.A1(n_257_76_12739), .A2(n_257_442), .ZN(
      n_257_76_12740));
   OAI21_X1 i_257_76_12763 (.A(n_257_76_12740), .B1(n_257_432), .B2(
      n_257_76_17412), .ZN(n_257_76_12741));
   NAND3_X1 i_257_76_12764 (.A1(n_257_76_12477), .A2(n_257_76_12741), .A3(
      n_257_429), .ZN(n_257_76_12742));
   INV_X1 i_257_76_12765 (.A(n_257_76_12742), .ZN(n_257_76_12743));
   NAND4_X1 i_257_76_12766 (.A1(n_257_76_12743), .A2(n_257_76_12507), .A3(
      n_257_76_12504), .A4(n_257_76_12505), .ZN(n_257_76_12744));
   INV_X1 i_257_76_12767 (.A(n_257_76_12744), .ZN(n_257_76_12745));
   NAND4_X1 i_257_76_12768 (.A1(n_257_76_12606), .A2(n_257_76_12614), .A3(
      n_257_76_12745), .A4(n_257_76_12513), .ZN(n_257_76_12746));
   NAND4_X1 i_257_76_12769 (.A1(n_257_76_12511), .A2(n_257_76_12476), .A3(
      n_257_76_12556), .A4(n_257_76_12512), .ZN(n_257_76_12747));
   NOR2_X1 i_257_76_12770 (.A1(n_257_76_12746), .A2(n_257_76_12747), .ZN(
      n_257_76_12748));
   NAND2_X1 i_257_76_12771 (.A1(n_257_76_12551), .A2(n_257_76_12552), .ZN(
      n_257_76_12749));
   INV_X1 i_257_76_12772 (.A(n_257_76_12749), .ZN(n_257_76_12750));
   NAND3_X1 i_257_76_12773 (.A1(n_257_76_12750), .A2(n_257_76_12555), .A3(
      n_257_174), .ZN(n_257_76_12751));
   INV_X1 i_257_76_12774 (.A(n_257_76_12751), .ZN(n_257_76_12752));
   NAND4_X1 i_257_76_12775 (.A1(n_257_76_12748), .A2(n_257_76_12475), .A3(
      n_257_76_12516), .A4(n_257_76_12752), .ZN(n_257_76_12753));
   NOR2_X1 i_257_76_12776 (.A1(n_257_76_12753), .A2(n_257_76_12518), .ZN(
      n_257_76_12754));
   NAND2_X1 i_257_76_12777 (.A1(n_257_76_18061), .A2(n_257_76_12754), .ZN(
      n_257_76_12755));
   NAND3_X1 i_257_76_12778 (.A1(n_257_76_12726), .A2(n_257_76_12738), .A3(
      n_257_76_12755), .ZN(n_257_76_12756));
   INV_X1 i_257_76_12779 (.A(n_257_76_12756), .ZN(n_257_76_12757));
   INV_X1 i_257_76_12780 (.A(n_257_76_12504), .ZN(n_257_76_12758));
   NAND3_X1 i_257_76_12781 (.A1(n_257_76_12758), .A2(n_257_76_12507), .A3(
      n_257_76_12490), .ZN(n_257_76_12759));
   INV_X1 i_257_76_12782 (.A(n_257_76_12759), .ZN(n_257_76_12760));
   NAND3_X1 i_257_76_12783 (.A1(n_257_76_12476), .A2(n_257_76_12512), .A3(
      n_257_76_12760), .ZN(n_257_76_12761));
   INV_X1 i_257_76_12784 (.A(n_257_76_12761), .ZN(n_257_76_12762));
   NAND2_X1 i_257_76_12785 (.A1(n_257_76_12475), .A2(n_257_76_12762), .ZN(
      n_257_76_12763));
   INV_X1 i_257_76_12786 (.A(n_257_76_12763), .ZN(n_257_76_12764));
   NAND2_X1 i_257_76_12787 (.A1(n_257_76_12764), .A2(n_257_76_12486), .ZN(
      n_257_76_12765));
   INV_X1 i_257_76_12788 (.A(n_257_76_12765), .ZN(n_257_76_12766));
   NAND2_X1 i_257_76_12789 (.A1(n_257_76_18067), .A2(n_257_76_12766), .ZN(
      n_257_76_12767));
   NAND2_X1 i_257_76_12790 (.A1(n_257_332), .A2(n_257_422), .ZN(n_257_76_12768));
   NAND4_X1 i_257_76_12791 (.A1(n_257_76_12768), .A2(n_257_76_12504), .A3(
      n_257_76_12505), .A4(n_257_76_12561), .ZN(n_257_76_12769));
   NAND2_X1 i_257_76_12792 (.A1(n_257_76_12568), .A2(n_257_76_12507), .ZN(
      n_257_76_12770));
   NOR2_X1 i_257_76_12793 (.A1(n_257_76_12769), .A2(n_257_76_12770), .ZN(
      n_257_76_12771));
   NAND2_X1 i_257_76_12794 (.A1(n_257_294), .A2(n_257_423), .ZN(n_257_76_12772));
   NAND3_X1 i_257_76_12795 (.A1(n_257_76_12772), .A2(n_257_76_12501), .A3(
      n_257_76_12496), .ZN(n_257_76_12773));
   INV_X1 i_257_76_12796 (.A(n_257_76_12773), .ZN(n_257_76_12774));
   NAND2_X1 i_257_76_12797 (.A1(n_257_76_12563), .A2(n_257_420), .ZN(
      n_257_76_12775));
   INV_X1 i_257_76_12798 (.A(n_257_76_12775), .ZN(n_257_76_12776));
   NAND2_X1 i_257_76_12799 (.A1(n_257_442), .A2(n_257_491), .ZN(n_257_76_12777));
   NAND3_X1 i_257_76_12800 (.A1(n_257_76_12776), .A2(n_257_76_12477), .A3(
      n_257_76_18009), .ZN(n_257_76_12778));
   INV_X1 i_257_76_12801 (.A(n_257_76_12778), .ZN(n_257_76_12779));
   NAND4_X1 i_257_76_12802 (.A1(n_257_76_12497), .A2(n_257_76_12571), .A3(
      n_257_76_12498), .A4(n_257_76_12779), .ZN(n_257_76_12780));
   INV_X1 i_257_76_12803 (.A(n_257_76_12780), .ZN(n_257_76_12781));
   NAND3_X1 i_257_76_12804 (.A1(n_257_76_12771), .A2(n_257_76_12774), .A3(
      n_257_76_12781), .ZN(n_257_76_12782));
   INV_X1 i_257_76_12805 (.A(n_257_76_12782), .ZN(n_257_76_12783));
   NAND2_X1 i_257_76_12806 (.A1(n_257_371), .A2(n_257_421), .ZN(n_257_76_12784));
   NAND4_X1 i_257_76_12807 (.A1(n_257_76_12550), .A2(n_257_76_12551), .A3(
      n_257_76_12784), .A4(n_257_76_12552), .ZN(n_257_76_12785));
   INV_X1 i_257_76_12808 (.A(n_257_76_12785), .ZN(n_257_76_12786));
   NAND2_X1 i_257_76_12809 (.A1(n_257_76_12511), .A2(n_257_76_12476), .ZN(
      n_257_76_12787));
   NOR2_X1 i_257_76_12810 (.A1(n_257_76_12688), .A2(n_257_76_12787), .ZN(
      n_257_76_12788));
   NAND3_X1 i_257_76_12811 (.A1(n_257_76_12783), .A2(n_257_76_12786), .A3(
      n_257_76_12788), .ZN(n_257_76_12789));
   NAND3_X1 i_257_76_12812 (.A1(n_257_76_12516), .A2(n_257_76_12560), .A3(
      n_257_76_12555), .ZN(n_257_76_12790));
   NOR2_X1 i_257_76_12813 (.A1(n_257_76_12789), .A2(n_257_76_12790), .ZN(
      n_257_76_12791));
   NAND3_X1 i_257_76_12814 (.A1(n_257_76_12791), .A2(n_257_76_12578), .A3(
      n_257_76_12486), .ZN(n_257_76_12792));
   INV_X1 i_257_76_12815 (.A(n_257_76_12792), .ZN(n_257_76_12793));
   NAND2_X1 i_257_76_12816 (.A1(n_257_76_18073), .A2(n_257_76_12793), .ZN(
      n_257_76_12794));
   INV_X1 i_257_76_12817 (.A(n_257_76_12603), .ZN(n_257_76_12795));
   NAND2_X1 i_257_76_12818 (.A1(n_257_76_12552), .A2(n_257_76_12511), .ZN(
      n_257_76_12796));
   INV_X1 i_257_76_12819 (.A(n_257_76_12796), .ZN(n_257_76_12797));
   NAND3_X1 i_257_76_12820 (.A1(n_257_76_12795), .A2(n_257_76_12555), .A3(
      n_257_76_12797), .ZN(n_257_76_12798));
   INV_X1 i_257_76_12821 (.A(n_257_76_12798), .ZN(n_257_76_12799));
   NAND3_X1 i_257_76_12822 (.A1(n_257_76_12477), .A2(n_257_76_12741), .A3(
      n_257_430), .ZN(n_257_76_12800));
   INV_X1 i_257_76_12823 (.A(n_257_76_12800), .ZN(n_257_76_12801));
   NAND4_X1 i_257_76_12824 (.A1(n_257_76_12801), .A2(n_257_76_12507), .A3(
      n_257_76_12504), .A4(n_257_76_12505), .ZN(n_257_76_12802));
   INV_X1 i_257_76_12825 (.A(n_257_76_12802), .ZN(n_257_76_12803));
   NAND2_X1 i_257_76_12826 (.A1(n_257_76_12571), .A2(n_257_76_12498), .ZN(
      n_257_76_12804));
   INV_X1 i_257_76_12827 (.A(n_257_76_12804), .ZN(n_257_76_12805));
   NAND3_X1 i_257_76_12828 (.A1(n_257_76_12803), .A2(n_257_76_12805), .A3(
      n_257_76_12497), .ZN(n_257_76_12806));
   NAND4_X1 i_257_76_12829 (.A1(n_257_76_12513), .A2(n_257_135), .A3(
      n_257_76_12501), .A4(n_257_76_12496), .ZN(n_257_76_12807));
   NOR2_X1 i_257_76_12830 (.A1(n_257_76_12806), .A2(n_257_76_12807), .ZN(
      n_257_76_12808));
   NAND4_X1 i_257_76_12831 (.A1(n_257_76_12475), .A2(n_257_76_12799), .A3(
      n_257_76_12808), .A4(n_257_76_12516), .ZN(n_257_76_12809));
   NOR2_X1 i_257_76_12832 (.A1(n_257_76_12809), .A2(n_257_76_12518), .ZN(
      n_257_76_12810));
   NAND2_X1 i_257_76_12833 (.A1(n_257_76_18068), .A2(n_257_76_12810), .ZN(
      n_257_76_12811));
   NAND3_X1 i_257_76_12834 (.A1(n_257_76_12767), .A2(n_257_76_12794), .A3(
      n_257_76_12811), .ZN(n_257_76_12812));
   INV_X1 i_257_76_12835 (.A(n_257_76_12812), .ZN(n_257_76_12813));
   NAND2_X1 i_257_76_12836 (.A1(n_257_447), .A2(n_257_76_12507), .ZN(
      n_257_76_12814));
   INV_X1 i_257_76_12837 (.A(n_257_76_12814), .ZN(n_257_76_12815));
   NAND2_X1 i_257_76_12838 (.A1(n_257_787), .A2(n_257_442), .ZN(n_257_76_12816));
   NOR2_X1 i_257_76_12839 (.A1(n_257_1081), .A2(n_257_76_12816), .ZN(
      n_257_76_12817));
   NAND2_X1 i_257_76_12840 (.A1(n_257_76_12504), .A2(n_257_76_12817), .ZN(
      n_257_76_12818));
   INV_X1 i_257_76_12841 (.A(n_257_76_12818), .ZN(n_257_76_12819));
   NAND4_X1 i_257_76_12842 (.A1(n_257_76_12815), .A2(n_257_76_12819), .A3(
      n_257_76_12501), .A4(n_257_76_12498), .ZN(n_257_76_12820));
   NOR2_X1 i_257_76_12843 (.A1(n_257_76_12670), .A2(n_257_76_12820), .ZN(
      n_257_76_12821));
   NAND2_X1 i_257_76_12844 (.A1(n_257_76_12475), .A2(n_257_76_12821), .ZN(
      n_257_76_12822));
   INV_X1 i_257_76_12845 (.A(n_257_76_12822), .ZN(n_257_76_12823));
   NAND2_X1 i_257_76_12846 (.A1(n_257_76_12823), .A2(n_257_76_12486), .ZN(
      n_257_76_12824));
   INV_X1 i_257_76_12847 (.A(n_257_76_12824), .ZN(n_257_76_12825));
   NAND2_X1 i_257_76_12848 (.A1(n_257_76_12496), .A2(n_257_76_12497), .ZN(
      n_257_76_12826));
   INV_X1 i_257_76_12849 (.A(n_257_76_12826), .ZN(n_257_76_12827));
   NAND3_X1 i_257_76_12850 (.A1(n_257_76_12477), .A2(n_257_76_12741), .A3(
      n_257_431), .ZN(n_257_76_12828));
   INV_X1 i_257_76_12851 (.A(n_257_76_12828), .ZN(n_257_76_12829));
   NAND4_X1 i_257_76_12852 (.A1(n_257_76_12829), .A2(n_257_76_12507), .A3(
      n_257_76_12504), .A4(n_257_76_12505), .ZN(n_257_76_12830));
   INV_X1 i_257_76_12853 (.A(n_257_76_12830), .ZN(n_257_76_12831));
   NAND3_X1 i_257_76_12854 (.A1(n_257_76_12827), .A2(n_257_76_12831), .A3(
      n_257_76_12805), .ZN(n_257_76_12832));
   NOR2_X1 i_257_76_12855 (.A1(n_257_76_12832), .A2(n_257_76_12545), .ZN(
      n_257_76_12833));
   NAND2_X1 i_257_76_12856 (.A1(n_257_97), .A2(n_257_76_12552), .ZN(
      n_257_76_12834));
   NOR2_X1 i_257_76_12857 (.A1(n_257_76_12834), .A2(n_257_76_12557), .ZN(
      n_257_76_12835));
   NAND3_X1 i_257_76_12858 (.A1(n_257_76_12833), .A2(n_257_76_12516), .A3(
      n_257_76_12835), .ZN(n_257_76_12836));
   INV_X1 i_257_76_12859 (.A(n_257_76_12836), .ZN(n_257_76_12837));
   NAND3_X1 i_257_76_12860 (.A1(n_257_76_12837), .A2(n_257_76_12486), .A3(
      n_257_76_12475), .ZN(n_257_76_12838));
   INV_X1 i_257_76_12861 (.A(n_257_76_12838), .ZN(n_257_76_12839));
   AOI22_X1 i_257_76_12862 (.A1(n_257_76_18085), .A2(n_257_76_12825), .B1(
      n_257_76_18080), .B2(n_257_76_12839), .ZN(n_257_76_12840));
   NAND3_X1 i_257_76_12863 (.A1(n_257_76_12757), .A2(n_257_76_12813), .A3(
      n_257_76_12840), .ZN(n_257_76_12841));
   INV_X1 i_257_76_12864 (.A(n_257_723), .ZN(n_257_76_12842));
   NAND2_X1 i_257_76_12865 (.A1(n_257_76_12842), .A2(n_257_442), .ZN(
      n_257_76_12843));
   AOI21_X1 i_257_76_12866 (.A(n_257_1081), .B1(n_257_76_12843), .B2(
      n_257_76_17761), .ZN(n_257_76_12844));
   NAND3_X1 i_257_76_12867 (.A1(n_257_76_12844), .A2(n_257_76_12501), .A3(
      n_257_76_12497), .ZN(n_257_76_12845));
   NAND4_X1 i_257_76_12868 (.A1(n_257_76_12498), .A2(n_257_76_12507), .A3(
      n_257_76_12504), .A4(n_257_448), .ZN(n_257_76_12846));
   NOR2_X1 i_257_76_12869 (.A1(n_257_76_12845), .A2(n_257_76_12846), .ZN(
      n_257_76_12847));
   INV_X1 i_257_76_12870 (.A(n_257_76_12514), .ZN(n_257_76_12848));
   NAND3_X1 i_257_76_12871 (.A1(n_257_76_12847), .A2(n_257_691), .A3(
      n_257_76_12848), .ZN(n_257_76_12849));
   INV_X1 i_257_76_12872 (.A(n_257_76_12849), .ZN(n_257_76_12850));
   NAND2_X1 i_257_76_12873 (.A1(n_257_76_12850), .A2(n_257_76_12475), .ZN(
      n_257_76_12851));
   NOR2_X1 i_257_76_12874 (.A1(n_257_76_12851), .A2(n_257_76_12518), .ZN(
      n_257_76_12852));
   NAND2_X1 i_257_76_12875 (.A1(n_257_76_18079), .A2(n_257_76_12852), .ZN(
      n_257_76_12853));
   NAND2_X1 i_257_76_12876 (.A1(n_257_254), .A2(n_257_76_12516), .ZN(
      n_257_76_12854));
   INV_X1 i_257_76_12877 (.A(n_257_76_12854), .ZN(n_257_76_12855));
   NAND3_X1 i_257_76_12878 (.A1(n_257_76_12507), .A2(n_257_76_12504), .A3(
      n_257_76_12505), .ZN(n_257_76_12856));
   INV_X1 i_257_76_12879 (.A(n_257_76_18008), .ZN(n_257_76_12857));
   NOR2_X1 i_257_76_12880 (.A1(n_257_1081), .A2(n_257_76_12857), .ZN(
      n_257_76_12858));
   NAND2_X1 i_257_76_12881 (.A1(n_257_76_12563), .A2(n_257_425), .ZN(
      n_257_76_12859));
   INV_X1 i_257_76_12882 (.A(n_257_76_12859), .ZN(n_257_76_12860));
   NAND3_X1 i_257_76_12883 (.A1(n_257_76_12858), .A2(n_257_76_12561), .A3(
      n_257_76_12860), .ZN(n_257_76_12861));
   NOR2_X1 i_257_76_12884 (.A1(n_257_76_12856), .A2(n_257_76_12861), .ZN(
      n_257_76_12862));
   NAND4_X1 i_257_76_12885 (.A1(n_257_76_12862), .A2(n_257_76_12606), .A3(
      n_257_76_12614), .A4(n_257_76_12513), .ZN(n_257_76_12863));
   NOR2_X1 i_257_76_12886 (.A1(n_257_76_12863), .A2(n_257_76_12747), .ZN(
      n_257_76_12864));
   NAND3_X1 i_257_76_12887 (.A1(n_257_76_12560), .A2(n_257_76_12555), .A3(
      n_257_76_12554), .ZN(n_257_76_12865));
   INV_X1 i_257_76_12888 (.A(n_257_76_12865), .ZN(n_257_76_12866));
   NAND3_X1 i_257_76_12889 (.A1(n_257_76_12855), .A2(n_257_76_12864), .A3(
      n_257_76_12866), .ZN(n_257_76_12867));
   NAND2_X1 i_257_76_12890 (.A1(n_257_76_12486), .A2(n_257_76_12475), .ZN(
      n_257_76_12868));
   NOR2_X1 i_257_76_12891 (.A1(n_257_76_12867), .A2(n_257_76_12868), .ZN(
      n_257_76_12869));
   NAND2_X1 i_257_76_12892 (.A1(n_257_76_18064), .A2(n_257_76_12869), .ZN(
      n_257_76_12870));
   INV_X1 i_257_76_12893 (.A(n_257_76_12560), .ZN(n_257_76_12871));
   NOR2_X1 i_257_76_12894 (.A1(n_257_76_12871), .A2(n_257_76_12655), .ZN(
      n_257_76_12872));
   NAND4_X1 i_257_76_12895 (.A1(n_257_76_12872), .A2(n_257_76_12576), .A3(
      n_257_76_12475), .A4(n_257_76_12516), .ZN(n_257_76_12873));
   NAND3_X1 i_257_76_12896 (.A1(n_257_371), .A2(n_257_76_12772), .A3(
      n_257_76_12501), .ZN(n_257_76_12874));
   NAND3_X1 i_257_76_12897 (.A1(n_257_76_12496), .A2(n_257_76_12497), .A3(
      n_257_76_12571), .ZN(n_257_76_12875));
   NOR2_X1 i_257_76_12898 (.A1(n_257_76_12874), .A2(n_257_76_12875), .ZN(
      n_257_76_12876));
   NAND4_X1 i_257_76_12899 (.A1(n_257_76_12498), .A2(n_257_76_12568), .A3(
      n_257_76_12507), .A4(n_257_76_12768), .ZN(n_257_76_12877));
   NAND2_X1 i_257_76_12900 (.A1(n_257_76_12563), .A2(n_257_421), .ZN(
      n_257_76_12878));
   INV_X1 i_257_76_12901 (.A(n_257_76_12878), .ZN(n_257_76_12879));
   NAND3_X1 i_257_76_12902 (.A1(n_257_76_12879), .A2(n_257_76_12477), .A3(
      n_257_76_18008), .ZN(n_257_76_12880));
   INV_X1 i_257_76_12903 (.A(n_257_76_12880), .ZN(n_257_76_12881));
   NAND3_X1 i_257_76_12904 (.A1(n_257_76_12641), .A2(n_257_76_12504), .A3(
      n_257_76_12881), .ZN(n_257_76_12882));
   NOR2_X1 i_257_76_12905 (.A1(n_257_76_12877), .A2(n_257_76_12882), .ZN(
      n_257_76_12883));
   NAND3_X1 i_257_76_12906 (.A1(n_257_76_12511), .A2(n_257_76_12512), .A3(
      n_257_76_12513), .ZN(n_257_76_12884));
   INV_X1 i_257_76_12907 (.A(n_257_76_12884), .ZN(n_257_76_12885));
   NAND4_X1 i_257_76_12908 (.A1(n_257_76_12876), .A2(n_257_76_12554), .A3(
      n_257_76_12883), .A4(n_257_76_12885), .ZN(n_257_76_12886));
   INV_X1 i_257_76_12909 (.A(n_257_76_12886), .ZN(n_257_76_12887));
   NAND2_X1 i_257_76_12910 (.A1(n_257_76_12486), .A2(n_257_76_12887), .ZN(
      n_257_76_12888));
   NOR2_X1 i_257_76_12911 (.A1(n_257_76_12873), .A2(n_257_76_12888), .ZN(
      n_257_76_12889));
   NAND2_X1 i_257_76_12912 (.A1(n_257_76_18082), .A2(n_257_76_12889), .ZN(
      n_257_76_12890));
   NAND3_X1 i_257_76_12913 (.A1(n_257_76_12853), .A2(n_257_76_12870), .A3(
      n_257_76_12890), .ZN(n_257_76_12891));
   INV_X1 i_257_76_12914 (.A(n_257_76_12891), .ZN(n_257_76_12892));
   NAND2_X1 i_257_76_12915 (.A1(n_257_76_12477), .A2(n_257_214), .ZN(
      n_257_76_12893));
   NAND3_X1 i_257_76_12916 (.A1(n_257_76_18008), .A2(n_257_427), .A3(
      n_257_76_12563), .ZN(n_257_76_12894));
   NOR2_X1 i_257_76_12917 (.A1(n_257_76_12893), .A2(n_257_76_12894), .ZN(
      n_257_76_12895));
   NAND4_X1 i_257_76_12918 (.A1(n_257_76_12513), .A2(n_257_76_12895), .A3(
      n_257_76_12501), .A4(n_257_76_12496), .ZN(n_257_76_12896));
   INV_X1 i_257_76_12919 (.A(n_257_76_12856), .ZN(n_257_76_12897));
   NAND4_X1 i_257_76_12920 (.A1(n_257_76_12897), .A2(n_257_76_12497), .A3(
      n_257_76_12571), .A4(n_257_76_12498), .ZN(n_257_76_12898));
   NOR2_X1 i_257_76_12921 (.A1(n_257_76_12896), .A2(n_257_76_12898), .ZN(
      n_257_76_12899));
   NAND4_X1 i_257_76_12922 (.A1(n_257_76_12560), .A2(n_257_76_12604), .A3(
      n_257_76_12899), .A4(n_257_76_12555), .ZN(n_257_76_12900));
   INV_X1 i_257_76_12923 (.A(n_257_76_12900), .ZN(n_257_76_12901));
   NAND3_X1 i_257_76_12924 (.A1(n_257_76_12901), .A2(n_257_76_12620), .A3(
      n_257_76_12486), .ZN(n_257_76_12902));
   INV_X1 i_257_76_12925 (.A(n_257_76_12902), .ZN(n_257_76_12903));
   NAND2_X1 i_257_76_12926 (.A1(n_257_76_18065), .A2(n_257_76_12903), .ZN(
      n_257_76_12904));
   NAND4_X1 i_257_76_12927 (.A1(n_257_76_12547), .A2(n_257_474), .A3(n_257_451), 
      .A4(n_257_76_12498), .ZN(n_257_76_12905));
   NOR2_X1 i_257_76_12928 (.A1(n_257_76_12905), .A2(n_257_76_12684), .ZN(
      n_257_76_12906));
   NAND3_X1 i_257_76_12929 (.A1(n_257_76_12512), .A2(n_257_76_12513), .A3(
      n_257_76_12844), .ZN(n_257_76_12907));
   INV_X1 i_257_76_12930 (.A(n_257_76_12907), .ZN(n_257_76_12908));
   NAND3_X1 i_257_76_12931 (.A1(n_257_76_12906), .A2(n_257_76_12687), .A3(
      n_257_76_12908), .ZN(n_257_76_12909));
   INV_X1 i_257_76_12932 (.A(n_257_76_12909), .ZN(n_257_76_12910));
   NAND3_X1 i_257_76_12933 (.A1(n_257_76_12910), .A2(n_257_76_12475), .A3(
      n_257_76_12516), .ZN(n_257_76_12911));
   NOR2_X1 i_257_76_12934 (.A1(n_257_76_12911), .A2(n_257_76_12518), .ZN(
      n_257_76_12912));
   NAND2_X1 i_257_76_12935 (.A1(n_257_76_18063), .A2(n_257_76_12912), .ZN(
      n_257_76_12913));
   INV_X1 i_257_76_12936 (.A(n_257_76_12790), .ZN(n_257_76_12914));
   NAND2_X1 i_257_76_12937 (.A1(n_257_523), .A2(n_257_76_12561), .ZN(
      n_257_76_12915));
   INV_X1 i_257_76_12938 (.A(n_257_76_12915), .ZN(n_257_76_12916));
   NAND2_X1 i_257_76_12939 (.A1(n_257_76_12563), .A2(n_257_424), .ZN(
      n_257_76_12917));
   INV_X1 i_257_76_12940 (.A(n_257_76_12917), .ZN(n_257_76_12918));
   NAND3_X1 i_257_76_12941 (.A1(n_257_76_12918), .A2(n_257_76_12477), .A3(
      n_257_76_18008), .ZN(n_257_76_12919));
   INV_X1 i_257_76_12942 (.A(n_257_76_12919), .ZN(n_257_76_12920));
   NAND4_X1 i_257_76_12943 (.A1(n_257_76_12916), .A2(n_257_76_12571), .A3(
      n_257_76_12920), .A4(n_257_76_12505), .ZN(n_257_76_12921));
   INV_X1 i_257_76_12944 (.A(n_257_76_12921), .ZN(n_257_76_12922));
   NAND3_X1 i_257_76_12945 (.A1(n_257_76_12922), .A2(n_257_76_12550), .A3(
      n_257_76_12551), .ZN(n_257_76_12923));
   INV_X1 i_257_76_12946 (.A(n_257_76_12923), .ZN(n_257_76_12924));
   NAND4_X1 i_257_76_12947 (.A1(n_257_76_12552), .A2(n_257_76_12511), .A3(
      n_257_76_12476), .A4(n_257_76_12556), .ZN(n_257_76_12925));
   INV_X1 i_257_76_12948 (.A(n_257_76_12925), .ZN(n_257_76_12926));
   NAND3_X1 i_257_76_12949 (.A1(n_257_76_12549), .A2(n_257_76_12924), .A3(
      n_257_76_12926), .ZN(n_257_76_12927));
   INV_X1 i_257_76_12950 (.A(n_257_76_12927), .ZN(n_257_76_12928));
   NAND2_X1 i_257_76_12951 (.A1(n_257_76_12914), .A2(n_257_76_12928), .ZN(
      n_257_76_12929));
   NOR3_X1 i_257_76_12952 (.A1(n_257_76_12929), .A2(n_257_76_12518), .A3(
      n_257_76_12577), .ZN(n_257_76_12930));
   NAND2_X1 i_257_76_12953 (.A1(n_257_76_18062), .A2(n_257_76_12930), .ZN(
      n_257_76_12931));
   NAND3_X1 i_257_76_12954 (.A1(n_257_76_12904), .A2(n_257_76_12913), .A3(
      n_257_76_12931), .ZN(n_257_76_12932));
   INV_X1 i_257_76_12955 (.A(n_257_76_12932), .ZN(n_257_76_12933));
   NAND2_X1 i_257_76_12956 (.A1(n_257_76_12563), .A2(n_257_422), .ZN(
      n_257_76_12934));
   INV_X1 i_257_76_12957 (.A(n_257_76_12934), .ZN(n_257_76_12935));
   NAND4_X1 i_257_76_12958 (.A1(n_257_76_12935), .A2(n_257_332), .A3(
      n_257_76_12477), .A4(n_257_76_18008), .ZN(n_257_76_12936));
   NOR2_X1 i_257_76_12959 (.A1(n_257_76_12936), .A2(n_257_76_12562), .ZN(
      n_257_76_12937));
   NAND2_X1 i_257_76_12960 (.A1(n_257_76_12571), .A2(n_257_76_12568), .ZN(
      n_257_76_12938));
   INV_X1 i_257_76_12961 (.A(n_257_76_12938), .ZN(n_257_76_12939));
   NAND3_X1 i_257_76_12962 (.A1(n_257_76_12937), .A2(n_257_76_12939), .A3(
      n_257_76_12772), .ZN(n_257_76_12940));
   INV_X1 i_257_76_12963 (.A(n_257_76_12940), .ZN(n_257_76_12941));
   NAND3_X1 i_257_76_12964 (.A1(n_257_76_12516), .A2(n_257_76_12560), .A3(
      n_257_76_12941), .ZN(n_257_76_12942));
   NOR2_X1 i_257_76_12965 (.A1(n_257_76_12559), .A2(n_257_76_12942), .ZN(
      n_257_76_12943));
   NAND3_X1 i_257_76_12966 (.A1(n_257_76_12943), .A2(n_257_76_12578), .A3(
      n_257_76_12486), .ZN(n_257_76_12944));
   INV_X1 i_257_76_12967 (.A(n_257_76_12944), .ZN(n_257_76_12945));
   NAND2_X1 i_257_76_12968 (.A1(n_257_342), .A2(n_257_76_12945), .ZN(
      n_257_76_12946));
   NAND2_X1 i_257_76_12969 (.A1(n_257_420), .A2(n_257_491), .ZN(n_257_76_12947));
   INV_X1 i_257_76_12970 (.A(n_257_76_12947), .ZN(n_257_76_12948));
   NOR2_X1 i_257_76_12971 (.A1(n_257_76_12948), .A2(n_257_1081), .ZN(
      n_257_76_12949));
   NAND2_X1 i_257_76_12972 (.A1(n_257_587), .A2(n_257_428), .ZN(n_257_76_12950));
   NAND3_X1 i_257_76_12973 (.A1(n_257_484), .A2(n_257_410), .A3(n_257_442), 
      .ZN(n_257_76_12951));
   INV_X1 i_257_76_12974 (.A(n_257_76_12951), .ZN(n_257_76_12952));
   NAND3_X1 i_257_76_12975 (.A1(n_257_76_12563), .A2(n_257_76_12950), .A3(
      n_257_76_12952), .ZN(n_257_76_12953));
   INV_X1 i_257_76_12976 (.A(n_257_76_12953), .ZN(n_257_76_12954));
   NAND4_X1 i_257_76_12977 (.A1(n_257_76_12949), .A2(n_257_76_12505), .A3(
      n_257_76_12561), .A4(n_257_76_12954), .ZN(n_257_76_12955));
   INV_X1 i_257_76_12978 (.A(n_257_76_12955), .ZN(n_257_76_12956));
   NAND2_X1 i_257_76_12979 (.A1(n_257_76_12498), .A2(n_257_76_12568), .ZN(
      n_257_76_12957));
   INV_X1 i_257_76_12980 (.A(n_257_76_12957), .ZN(n_257_76_12958));
   NAND3_X1 i_257_76_12981 (.A1(n_257_76_12507), .A2(n_257_76_12768), .A3(
      n_257_76_12504), .ZN(n_257_76_12959));
   INV_X1 i_257_76_12982 (.A(n_257_76_12959), .ZN(n_257_76_12960));
   NAND3_X1 i_257_76_12983 (.A1(n_257_76_12956), .A2(n_257_76_12958), .A3(
      n_257_76_12960), .ZN(n_257_76_12961));
   NAND4_X1 i_257_76_12984 (.A1(n_257_76_12501), .A2(n_257_76_12496), .A3(
      n_257_76_12497), .A4(n_257_76_12571), .ZN(n_257_76_12962));
   NOR2_X1 i_257_76_12985 (.A1(n_257_76_12961), .A2(n_257_76_12962), .ZN(
      n_257_76_12963));
   NAND3_X1 i_257_76_12986 (.A1(n_257_76_12963), .A2(n_257_76_12516), .A3(
      n_257_76_12560), .ZN(n_257_76_12964));
   NAND4_X1 i_257_76_12987 (.A1(n_257_76_12556), .A2(n_257_76_12512), .A3(
      n_257_76_12513), .A4(n_257_76_12772), .ZN(n_257_76_12965));
   INV_X1 i_257_76_12988 (.A(n_257_76_12965), .ZN(n_257_76_12966));
   NAND3_X1 i_257_76_12989 (.A1(n_257_76_12550), .A2(n_257_76_12551), .A3(
      n_257_76_12784), .ZN(n_257_76_12967));
   INV_X1 i_257_76_12990 (.A(n_257_76_12967), .ZN(n_257_76_12968));
   NAND4_X1 i_257_76_12991 (.A1(n_257_76_12966), .A2(n_257_76_12968), .A3(
      n_257_76_12555), .A4(n_257_76_12687), .ZN(n_257_76_12969));
   NOR2_X1 i_257_76_12992 (.A1(n_257_76_12964), .A2(n_257_76_12969), .ZN(
      n_257_76_12970));
   NAND3_X1 i_257_76_12993 (.A1(n_257_76_12970), .A2(n_257_76_12578), .A3(
      n_257_76_12486), .ZN(n_257_76_12971));
   INV_X1 i_257_76_12994 (.A(n_257_76_12971), .ZN(n_257_76_12972));
   NAND2_X1 i_257_76_12995 (.A1(n_257_76_18060), .A2(n_257_76_12972), .ZN(
      n_257_76_12973));
   NAND2_X1 i_257_76_12996 (.A1(n_257_135), .A2(n_257_76_17925), .ZN(
      n_257_76_12974));
   NAND2_X1 i_257_76_12997 (.A1(n_257_985), .A2(n_257_442), .ZN(n_257_76_12975));
   INV_X1 i_257_76_12998 (.A(n_257_76_12975), .ZN(n_257_76_12976));
   NAND2_X1 i_257_76_12999 (.A1(n_257_76_12976), .A2(n_257_441), .ZN(
      n_257_76_12977));
   NAND2_X1 i_257_76_13000 (.A1(n_257_651), .A2(n_257_76_17928), .ZN(
      n_257_76_12978));
   NAND3_X1 i_257_76_13001 (.A1(n_257_76_12974), .A2(n_257_76_12977), .A3(
      n_257_76_12978), .ZN(n_257_76_12979));
   NAND2_X1 i_257_76_13002 (.A1(n_257_755), .A2(n_257_76_17935), .ZN(
      n_257_76_12980));
   NAND2_X1 i_257_76_13003 (.A1(n_257_921), .A2(n_257_76_17940), .ZN(
      n_257_76_12981));
   NAND2_X1 i_257_76_13004 (.A1(n_257_819), .A2(n_257_76_17952), .ZN(
      n_257_76_12982));
   NAND3_X1 i_257_76_13005 (.A1(n_257_76_12980), .A2(n_257_76_12981), .A3(
      n_257_76_12982), .ZN(n_257_76_12983));
   NOR2_X1 i_257_76_13006 (.A1(n_257_76_12979), .A2(n_257_76_12983), .ZN(
      n_257_76_12984));
   NAND2_X1 i_257_76_13007 (.A1(n_257_76_12572), .A2(n_257_76_12921), .ZN(
      n_257_76_12985));
   INV_X1 i_257_76_13008 (.A(n_257_76_12985), .ZN(n_257_76_12986));
   NAND2_X1 i_257_76_13009 (.A1(n_257_883), .A2(n_257_76_17903), .ZN(
      n_257_76_12987));
   NAND2_X1 i_257_76_13010 (.A1(n_257_76_12987), .A2(n_257_76_12778), .ZN(
      n_257_76_12988));
   NAND3_X1 i_257_76_13011 (.A1(n_257_438), .A2(n_257_1087), .A3(n_257_442), 
      .ZN(n_257_76_12989));
   NAND2_X1 i_257_76_13012 (.A1(n_257_440), .A2(n_257_76_12479), .ZN(
      n_257_76_12990));
   NAND2_X1 i_257_76_13013 (.A1(n_257_723), .A2(n_257_76_15655), .ZN(
      n_257_76_12991));
   NAND3_X1 i_257_76_13014 (.A1(n_257_76_12989), .A2(n_257_76_12990), .A3(
      n_257_76_12991), .ZN(n_257_76_12992));
   NOR2_X1 i_257_76_13015 (.A1(n_257_76_12988), .A2(n_257_76_12992), .ZN(
      n_257_76_12993));
   INV_X1 i_257_76_13016 (.A(n_257_76_12525), .ZN(n_257_76_12994));
   NAND2_X1 i_257_76_13017 (.A1(n_257_446), .A2(n_257_76_12994), .ZN(
      n_257_76_12995));
   NAND2_X1 i_257_76_13018 (.A1(n_257_449), .A2(n_257_76_17387), .ZN(
      n_257_76_12996));
   INV_X1 i_257_76_13019 (.A(Small_Packet_Data_Size[22]), .ZN(n_257_76_12997));
   NAND2_X1 i_257_76_13020 (.A1(n_257_76_12950), .A2(n_257_76_18010), .ZN(
      n_257_76_12998));
   INV_X1 i_257_76_13021 (.A(n_257_76_12998), .ZN(n_257_76_12999));
   NAND3_X1 i_257_76_13022 (.A1(n_257_76_12477), .A2(n_257_76_12999), .A3(
      n_257_76_12563), .ZN(n_257_76_13000));
   NAND2_X1 i_257_76_13023 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[22]), 
      .ZN(n_257_76_13001));
   NAND2_X1 i_257_76_13024 (.A1(n_257_76_13000), .A2(n_257_76_13001), .ZN(
      n_257_76_13002));
   NAND3_X1 i_257_76_13025 (.A1(n_257_76_12995), .A2(n_257_76_12996), .A3(
      n_257_76_13002), .ZN(n_257_76_13003));
   INV_X1 i_257_76_13026 (.A(n_257_76_13003), .ZN(n_257_76_13004));
   INV_X1 i_257_76_13027 (.A(n_257_76_12895), .ZN(n_257_76_13005));
   INV_X1 i_257_76_13028 (.A(n_257_76_12816), .ZN(n_257_76_13006));
   NAND2_X1 i_257_76_13029 (.A1(n_257_447), .A2(n_257_76_13006), .ZN(
      n_257_76_13007));
   NAND2_X1 i_257_76_13030 (.A1(n_257_57), .A2(n_257_76_17918), .ZN(
      n_257_76_13008));
   NAND3_X1 i_257_76_13031 (.A1(n_257_76_13005), .A2(n_257_76_13007), .A3(
      n_257_76_13008), .ZN(n_257_76_13009));
   INV_X1 i_257_76_13032 (.A(n_257_76_13009), .ZN(n_257_76_13010));
   NAND3_X1 i_257_76_13033 (.A1(n_257_76_12993), .A2(n_257_76_13004), .A3(
      n_257_76_13010), .ZN(n_257_76_13011));
   INV_X1 i_257_76_13034 (.A(n_257_76_13011), .ZN(n_257_76_13012));
   NAND3_X1 i_257_76_13035 (.A1(n_257_76_12984), .A2(n_257_76_12986), .A3(
      n_257_76_13012), .ZN(n_257_76_13013));
   NAND2_X1 i_257_76_13036 (.A1(n_257_97), .A2(n_257_76_17932), .ZN(
      n_257_76_13014));
   NAND2_X1 i_257_76_13037 (.A1(n_257_76_12940), .A2(n_257_76_13014), .ZN(
      n_257_76_13015));
   INV_X1 i_257_76_13038 (.A(n_257_76_13015), .ZN(n_257_76_13016));
   NAND2_X1 i_257_76_13039 (.A1(n_257_691), .A2(n_257_76_17958), .ZN(
      n_257_76_13017));
   NAND2_X1 i_257_76_13040 (.A1(n_257_174), .A2(n_257_76_17331), .ZN(
      n_257_76_13018));
   NAND3_X1 i_257_76_13041 (.A1(n_257_76_13016), .A2(n_257_76_13017), .A3(
      n_257_76_13018), .ZN(n_257_76_13019));
   NOR2_X1 i_257_76_13042 (.A1(n_257_76_13013), .A2(n_257_76_13019), .ZN(
      n_257_76_13020));
   NAND2_X1 i_257_76_13043 (.A1(n_257_1017), .A2(n_257_76_17964), .ZN(
      n_257_76_13021));
   INV_X1 i_257_76_13044 (.A(n_257_755), .ZN(n_257_76_13022));
   NAND2_X1 i_257_76_13045 (.A1(n_257_76_13022), .A2(n_257_442), .ZN(
      n_257_76_13023));
   INV_X1 i_257_76_13046 (.A(n_257_921), .ZN(n_257_76_13024));
   NAND2_X1 i_257_76_13047 (.A1(n_257_76_13024), .A2(n_257_442), .ZN(
      n_257_76_13025));
   INV_X1 i_257_76_13048 (.A(n_257_819), .ZN(n_257_76_13026));
   NAND2_X1 i_257_76_13049 (.A1(n_257_76_13026), .A2(n_257_442), .ZN(
      n_257_76_13027));
   INV_X1 i_257_76_13050 (.A(n_257_439), .ZN(n_257_76_13028));
   NAND2_X1 i_257_76_13051 (.A1(n_257_76_13028), .A2(n_257_442), .ZN(
      n_257_76_13029));
   NAND4_X1 i_257_76_13052 (.A1(n_257_76_13023), .A2(n_257_76_13025), .A3(
      n_257_76_13027), .A4(n_257_76_13029), .ZN(n_257_76_13030));
   INV_X1 i_257_76_13053 (.A(n_257_76_12556), .ZN(n_257_76_13031));
   NAND2_X1 i_257_76_13054 (.A1(n_257_76_13030), .A2(n_257_76_13031), .ZN(
      n_257_76_13032));
   NAND4_X1 i_257_76_13055 (.A1(n_257_76_12886), .A2(n_257_76_13021), .A3(
      n_257_76_12651), .A4(n_257_76_13032), .ZN(n_257_76_13033));
   INV_X1 i_257_76_13056 (.A(n_257_76_13033), .ZN(n_257_76_13034));
   NAND2_X1 i_257_76_13057 (.A1(n_257_1049), .A2(n_257_76_17969), .ZN(
      n_257_76_13035));
   NAND4_X1 i_257_76_13058 (.A1(n_257_76_13020), .A2(n_257_76_13034), .A3(
      n_257_76_12867), .A4(n_257_76_13035), .ZN(n_257_76_13036));
   NAND3_X1 i_257_76_13059 (.A1(n_257_76_12946), .A2(n_257_76_12973), .A3(
      n_257_76_13036), .ZN(n_257_76_13037));
   INV_X1 i_257_76_13060 (.A(n_257_76_13037), .ZN(n_257_76_13038));
   NAND3_X1 i_257_76_13061 (.A1(n_257_76_12892), .A2(n_257_76_12933), .A3(
      n_257_76_13038), .ZN(n_257_76_13039));
   NOR2_X1 i_257_76_13062 (.A1(n_257_76_12841), .A2(n_257_76_13039), .ZN(
      n_257_76_13040));
   NAND2_X1 i_257_76_13063 (.A1(n_257_76_12716), .A2(n_257_76_13040), .ZN(n_22));
   NAND2_X1 i_257_76_13064 (.A1(n_257_1018), .A2(n_257_444), .ZN(n_257_76_13041));
   NAND2_X1 i_257_76_13065 (.A1(n_257_441), .A2(n_257_986), .ZN(n_257_76_13042));
   INV_X1 i_257_76_13066 (.A(n_257_1082), .ZN(n_257_76_13043));
   NAND2_X1 i_257_76_13067 (.A1(n_257_954), .A2(n_257_442), .ZN(n_257_76_13044));
   INV_X1 i_257_76_13068 (.A(n_257_76_13044), .ZN(n_257_76_13045));
   NAND3_X1 i_257_76_13069 (.A1(n_257_440), .A2(n_257_76_13043), .A3(
      n_257_76_13045), .ZN(n_257_76_13046));
   INV_X1 i_257_76_13070 (.A(n_257_76_13046), .ZN(n_257_76_13047));
   NAND2_X1 i_257_76_13071 (.A1(n_257_76_13042), .A2(n_257_76_13047), .ZN(
      n_257_76_13048));
   INV_X1 i_257_76_13072 (.A(n_257_76_13048), .ZN(n_257_76_13049));
   NAND2_X1 i_257_76_13073 (.A1(n_257_76_13041), .A2(n_257_76_13049), .ZN(
      n_257_76_13050));
   INV_X1 i_257_76_13074 (.A(n_257_76_13050), .ZN(n_257_76_13051));
   NAND2_X1 i_257_76_13075 (.A1(n_257_1050), .A2(n_257_443), .ZN(n_257_76_13052));
   NAND2_X1 i_257_76_13076 (.A1(n_257_76_13051), .A2(n_257_76_13052), .ZN(
      n_257_76_13053));
   INV_X1 i_257_76_13077 (.A(n_257_76_13053), .ZN(n_257_76_13054));
   NAND2_X1 i_257_76_13078 (.A1(n_257_17), .A2(n_257_76_13054), .ZN(
      n_257_76_13055));
   NOR2_X1 i_257_76_13079 (.A1(n_257_1082), .A2(n_257_76_17412), .ZN(
      n_257_76_13056));
   INV_X1 i_257_76_13080 (.A(n_257_76_13056), .ZN(n_257_76_13057));
   NOR2_X1 i_257_76_13081 (.A1(n_257_76_13057), .A2(n_257_76_15197), .ZN(
      n_257_76_13058));
   NAND2_X1 i_257_76_13082 (.A1(n_257_1050), .A2(n_257_76_13058), .ZN(
      n_257_76_13059));
   INV_X1 i_257_76_13083 (.A(n_257_76_13059), .ZN(n_257_76_13060));
   NAND2_X1 i_257_76_13084 (.A1(n_257_76_18072), .A2(n_257_76_13060), .ZN(
      n_257_76_13061));
   INV_X1 i_257_76_13085 (.A(n_257_76_13052), .ZN(n_257_76_13062));
   NAND2_X1 i_257_76_13086 (.A1(n_257_756), .A2(n_257_436), .ZN(n_257_76_13063));
   NAND2_X1 i_257_76_13087 (.A1(n_257_922), .A2(n_257_439), .ZN(n_257_76_13064));
   NAND2_X1 i_257_76_13088 (.A1(n_257_820), .A2(n_257_437), .ZN(n_257_76_13065));
   NAND4_X1 i_257_76_13089 (.A1(n_257_76_13063), .A2(n_257_76_13064), .A3(
      n_257_76_13042), .A4(n_257_76_13065), .ZN(n_257_76_13066));
   NAND2_X1 i_257_76_13090 (.A1(n_257_447), .A2(n_257_788), .ZN(n_257_76_13067));
   NAND2_X1 i_257_76_13091 (.A1(n_257_884), .A2(n_257_445), .ZN(n_257_76_13068));
   NAND3_X1 i_257_76_13092 (.A1(n_257_76_13067), .A2(n_257_76_13068), .A3(
      n_257_652), .ZN(n_257_76_13069));
   INV_X1 i_257_76_13093 (.A(n_257_76_13069), .ZN(n_257_76_13070));
   NAND2_X1 i_257_76_13094 (.A1(n_257_446), .A2(n_257_852), .ZN(n_257_76_13071));
   NAND2_X1 i_257_76_13095 (.A1(n_257_449), .A2(n_257_898), .ZN(n_257_76_13072));
   NAND2_X1 i_257_76_13096 (.A1(n_257_76_13071), .A2(n_257_76_13072), .ZN(
      n_257_76_13073));
   INV_X1 i_257_76_13097 (.A(n_257_76_13073), .ZN(n_257_76_13074));
   NOR2_X1 i_257_76_13098 (.A1(n_257_1082), .A2(n_257_76_17927), .ZN(
      n_257_76_13075));
   NAND2_X1 i_257_76_13099 (.A1(n_257_440), .A2(n_257_954), .ZN(n_257_76_13076));
   NAND2_X1 i_257_76_13100 (.A1(n_257_438), .A2(n_257_1088), .ZN(n_257_76_13077));
   NAND2_X1 i_257_76_13101 (.A1(n_257_724), .A2(n_257_435), .ZN(n_257_76_13078));
   NAND4_X1 i_257_76_13102 (.A1(n_257_76_13075), .A2(n_257_76_13076), .A3(
      n_257_76_13077), .A4(n_257_76_13078), .ZN(n_257_76_13079));
   INV_X1 i_257_76_13103 (.A(n_257_76_13079), .ZN(n_257_76_13080));
   NAND3_X1 i_257_76_13104 (.A1(n_257_76_13070), .A2(n_257_76_13074), .A3(
      n_257_76_13080), .ZN(n_257_76_13081));
   NOR2_X1 i_257_76_13105 (.A1(n_257_76_13066), .A2(n_257_76_13081), .ZN(
      n_257_76_13082));
   NAND2_X1 i_257_76_13106 (.A1(n_257_692), .A2(n_257_448), .ZN(n_257_76_13083));
   NAND3_X1 i_257_76_13107 (.A1(n_257_76_13082), .A2(n_257_76_13041), .A3(
      n_257_76_13083), .ZN(n_257_76_13084));
   NOR2_X1 i_257_76_13108 (.A1(n_257_76_13062), .A2(n_257_76_13084), .ZN(
      n_257_76_13085));
   NAND2_X1 i_257_76_13109 (.A1(n_257_28), .A2(n_257_76_13085), .ZN(
      n_257_76_13086));
   NAND3_X1 i_257_76_13110 (.A1(n_257_76_13055), .A2(n_257_76_13061), .A3(
      n_257_76_13086), .ZN(n_257_76_13087));
   NAND2_X1 i_257_76_13111 (.A1(n_257_76_13064), .A2(n_257_76_13042), .ZN(
      n_257_76_13088));
   NAND2_X1 i_257_76_13112 (.A1(n_257_446), .A2(n_257_76_13076), .ZN(
      n_257_76_13089));
   INV_X1 i_257_76_13113 (.A(n_257_76_13089), .ZN(n_257_76_13090));
   NAND2_X1 i_257_76_13114 (.A1(n_257_852), .A2(n_257_442), .ZN(n_257_76_13091));
   NOR2_X1 i_257_76_13115 (.A1(n_257_1082), .A2(n_257_76_13091), .ZN(
      n_257_76_13092));
   NAND2_X1 i_257_76_13116 (.A1(n_257_76_13077), .A2(n_257_76_13092), .ZN(
      n_257_76_13093));
   INV_X1 i_257_76_13117 (.A(n_257_76_13093), .ZN(n_257_76_13094));
   NAND3_X1 i_257_76_13118 (.A1(n_257_76_13090), .A2(n_257_76_13094), .A3(
      n_257_76_13068), .ZN(n_257_76_13095));
   NOR2_X1 i_257_76_13119 (.A1(n_257_76_13088), .A2(n_257_76_13095), .ZN(
      n_257_76_13096));
   NAND2_X1 i_257_76_13120 (.A1(n_257_76_13041), .A2(n_257_76_13096), .ZN(
      n_257_76_13097));
   INV_X1 i_257_76_13121 (.A(n_257_76_13097), .ZN(n_257_76_13098));
   NAND2_X1 i_257_76_13122 (.A1(n_257_76_13098), .A2(n_257_76_13052), .ZN(
      n_257_76_13099));
   INV_X1 i_257_76_13123 (.A(n_257_76_13099), .ZN(n_257_76_13100));
   NAND2_X1 i_257_76_13124 (.A1(n_257_76_18070), .A2(n_257_76_13100), .ZN(
      n_257_76_13101));
   NAND3_X1 i_257_76_13125 (.A1(n_257_76_13056), .A2(n_257_76_13076), .A3(
      n_257_439), .ZN(n_257_76_13102));
   INV_X1 i_257_76_13126 (.A(n_257_76_13102), .ZN(n_257_76_13103));
   NAND3_X1 i_257_76_13127 (.A1(n_257_76_13042), .A2(n_257_922), .A3(
      n_257_76_13103), .ZN(n_257_76_13104));
   INV_X1 i_257_76_13128 (.A(n_257_76_13104), .ZN(n_257_76_13105));
   NAND2_X1 i_257_76_13129 (.A1(n_257_76_13041), .A2(n_257_76_13105), .ZN(
      n_257_76_13106));
   INV_X1 i_257_76_13130 (.A(n_257_76_13106), .ZN(n_257_76_13107));
   NAND2_X1 i_257_76_13131 (.A1(n_257_76_13107), .A2(n_257_76_13052), .ZN(
      n_257_76_13108));
   INV_X1 i_257_76_13132 (.A(n_257_76_13108), .ZN(n_257_76_13109));
   NAND2_X1 i_257_76_13133 (.A1(n_257_76_18084), .A2(n_257_76_13109), .ZN(
      n_257_76_13110));
   NAND2_X1 i_257_76_13134 (.A1(n_257_451), .A2(n_257_475), .ZN(n_257_76_13111));
   NAND2_X1 i_257_76_13135 (.A1(n_257_76_13042), .A2(n_257_76_13111), .ZN(
      n_257_76_13112));
   NAND3_X1 i_257_76_13136 (.A1(n_257_76_13071), .A2(n_257_76_13072), .A3(
      n_257_76_13067), .ZN(n_257_76_13113));
   NOR2_X1 i_257_76_13137 (.A1(n_257_76_13112), .A2(n_257_76_13113), .ZN(
      n_257_76_13114));
   NAND2_X1 i_257_76_13138 (.A1(n_257_255), .A2(n_257_425), .ZN(n_257_76_13115));
   NAND2_X1 i_257_76_13139 (.A1(n_257_175), .A2(n_257_429), .ZN(n_257_76_13116));
   NAND2_X1 i_257_76_13140 (.A1(n_257_98), .A2(n_257_431), .ZN(n_257_76_13117));
   NAND4_X1 i_257_76_13141 (.A1(n_257_76_13114), .A2(n_257_76_13115), .A3(
      n_257_76_13116), .A4(n_257_76_13117), .ZN(n_257_76_13118));
   NAND2_X1 i_257_76_13142 (.A1(n_257_556), .A2(n_257_426), .ZN(n_257_76_13119));
   NAND2_X1 i_257_76_13143 (.A1(n_257_76_13083), .A2(n_257_76_13119), .ZN(
      n_257_76_13120));
   NOR2_X1 i_257_76_13144 (.A1(n_257_76_13118), .A2(n_257_76_13120), .ZN(
      n_257_76_13121));
   INV_X1 i_257_76_13145 (.A(n_257_76_13041), .ZN(n_257_76_13122));
   NAND2_X1 i_257_76_13146 (.A1(n_257_432), .A2(n_257_620), .ZN(n_257_76_13123));
   NAND3_X1 i_257_76_13147 (.A1(n_257_76_18002), .A2(n_257_76_13123), .A3(
      n_257_423), .ZN(n_257_76_13124));
   NOR2_X1 i_257_76_13148 (.A1(n_257_76_13124), .A2(n_257_1082), .ZN(
      n_257_76_13125));
   NAND2_X1 i_257_76_13149 (.A1(n_257_215), .A2(n_257_427), .ZN(n_257_76_13126));
   NAND4_X1 i_257_76_13150 (.A1(n_257_76_13125), .A2(n_257_76_13077), .A3(
      n_257_76_13126), .A4(n_257_76_13078), .ZN(n_257_76_13127));
   NAND2_X1 i_257_76_13151 (.A1(n_257_58), .A2(n_257_433), .ZN(n_257_76_13128));
   NAND3_X1 i_257_76_13152 (.A1(n_257_76_13128), .A2(n_257_295), .A3(
      n_257_76_13076), .ZN(n_257_76_13129));
   NOR2_X1 i_257_76_13153 (.A1(n_257_76_13127), .A2(n_257_76_13129), .ZN(
      n_257_76_13130));
   NAND2_X1 i_257_76_13154 (.A1(n_257_136), .A2(n_257_430), .ZN(n_257_76_13131));
   NAND3_X1 i_257_76_13155 (.A1(n_257_76_13063), .A2(n_257_76_13131), .A3(
      n_257_76_13064), .ZN(n_257_76_13132));
   INV_X1 i_257_76_13156 (.A(n_257_76_13132), .ZN(n_257_76_13133));
   NAND2_X1 i_257_76_13157 (.A1(n_257_524), .A2(n_257_424), .ZN(n_257_76_13134));
   NAND2_X1 i_257_76_13158 (.A1(n_257_76_13068), .A2(n_257_76_13134), .ZN(
      n_257_76_13135));
   INV_X1 i_257_76_13159 (.A(n_257_76_13135), .ZN(n_257_76_13136));
   NAND2_X1 i_257_76_13160 (.A1(n_257_652), .A2(n_257_450), .ZN(n_257_76_13137));
   NAND3_X1 i_257_76_13161 (.A1(n_257_76_13136), .A2(n_257_76_13065), .A3(
      n_257_76_13137), .ZN(n_257_76_13138));
   INV_X1 i_257_76_13162 (.A(n_257_76_13138), .ZN(n_257_76_13139));
   NAND3_X1 i_257_76_13163 (.A1(n_257_76_13130), .A2(n_257_76_13133), .A3(
      n_257_76_13139), .ZN(n_257_76_13140));
   NOR2_X1 i_257_76_13164 (.A1(n_257_76_13122), .A2(n_257_76_13140), .ZN(
      n_257_76_13141));
   NAND3_X1 i_257_76_13165 (.A1(n_257_76_13121), .A2(n_257_76_13141), .A3(
      n_257_76_13052), .ZN(n_257_76_13142));
   INV_X1 i_257_76_13166 (.A(n_257_76_13142), .ZN(n_257_76_13143));
   NAND2_X1 i_257_76_13167 (.A1(n_257_76_18066), .A2(n_257_76_13143), .ZN(
      n_257_76_13144));
   NAND3_X1 i_257_76_13168 (.A1(n_257_76_13101), .A2(n_257_76_13110), .A3(
      n_257_76_13144), .ZN(n_257_76_13145));
   NOR2_X1 i_257_76_13169 (.A1(n_257_76_13087), .A2(n_257_76_13145), .ZN(
      n_257_76_13146));
   INV_X1 i_257_76_13170 (.A(n_257_441), .ZN(n_257_76_13147));
   NAND2_X1 i_257_76_13171 (.A1(n_257_986), .A2(n_257_76_13056), .ZN(
      n_257_76_13148));
   NOR2_X1 i_257_76_13172 (.A1(n_257_76_13147), .A2(n_257_76_13148), .ZN(
      n_257_76_13149));
   NAND2_X1 i_257_76_13173 (.A1(n_257_76_13041), .A2(n_257_76_13149), .ZN(
      n_257_76_13150));
   INV_X1 i_257_76_13174 (.A(n_257_76_13150), .ZN(n_257_76_13151));
   NAND2_X1 i_257_76_13175 (.A1(n_257_76_13151), .A2(n_257_76_13052), .ZN(
      n_257_76_13152));
   INV_X1 i_257_76_13176 (.A(n_257_76_13152), .ZN(n_257_76_13153));
   NAND2_X1 i_257_76_13177 (.A1(n_257_76_18071), .A2(n_257_76_13153), .ZN(
      n_257_76_13154));
   NAND2_X1 i_257_76_13178 (.A1(n_257_76_13067), .A2(n_257_76_13068), .ZN(
      n_257_76_13155));
   INV_X1 i_257_76_13179 (.A(n_257_76_13155), .ZN(n_257_76_13156));
   NAND2_X1 i_257_76_13180 (.A1(n_257_724), .A2(n_257_76_15655), .ZN(
      n_257_76_13157));
   INV_X1 i_257_76_13181 (.A(n_257_76_13157), .ZN(n_257_76_13158));
   NAND4_X1 i_257_76_13182 (.A1(n_257_76_13076), .A2(n_257_76_13077), .A3(
      n_257_76_13158), .A4(n_257_76_13043), .ZN(n_257_76_13159));
   INV_X1 i_257_76_13183 (.A(n_257_76_13159), .ZN(n_257_76_13160));
   NAND4_X1 i_257_76_13184 (.A1(n_257_76_13156), .A2(n_257_76_13160), .A3(
      n_257_76_13065), .A4(n_257_76_13071), .ZN(n_257_76_13161));
   NAND3_X1 i_257_76_13185 (.A1(n_257_76_13063), .A2(n_257_76_13064), .A3(
      n_257_76_13042), .ZN(n_257_76_13162));
   NOR2_X1 i_257_76_13186 (.A1(n_257_76_13161), .A2(n_257_76_13162), .ZN(
      n_257_76_13163));
   NAND2_X1 i_257_76_13187 (.A1(n_257_76_13041), .A2(n_257_76_13163), .ZN(
      n_257_76_13164));
   INV_X1 i_257_76_13188 (.A(n_257_76_13164), .ZN(n_257_76_13165));
   NAND2_X1 i_257_76_13189 (.A1(n_257_76_13165), .A2(n_257_76_13052), .ZN(
      n_257_76_13166));
   INV_X1 i_257_76_13190 (.A(n_257_76_13166), .ZN(n_257_76_13167));
   NAND2_X1 i_257_76_13191 (.A1(n_257_76_18078), .A2(n_257_76_13167), .ZN(
      n_257_76_13168));
   NAND2_X1 i_257_76_13192 (.A1(n_257_76_13076), .A2(n_257_76_13077), .ZN(
      n_257_76_13169));
   INV_X1 i_257_76_13193 (.A(n_257_76_13169), .ZN(n_257_76_13170));
   NAND3_X1 i_257_76_13194 (.A1(n_257_588), .A2(n_257_428), .A3(n_257_442), 
      .ZN(n_257_76_13171));
   INV_X1 i_257_76_13195 (.A(n_257_76_13171), .ZN(n_257_76_13172));
   NAND2_X1 i_257_76_13196 (.A1(n_257_76_13172), .A2(n_257_76_13123), .ZN(
      n_257_76_13173));
   INV_X1 i_257_76_13197 (.A(n_257_76_13173), .ZN(n_257_76_13174));
   NAND3_X1 i_257_76_13198 (.A1(n_257_76_13078), .A2(n_257_76_13174), .A3(
      n_257_76_13043), .ZN(n_257_76_13175));
   INV_X1 i_257_76_13199 (.A(n_257_76_13175), .ZN(n_257_76_13176));
   NAND4_X1 i_257_76_13200 (.A1(n_257_76_13170), .A2(n_257_76_13176), .A3(
      n_257_76_13068), .A4(n_257_76_13128), .ZN(n_257_76_13177));
   NOR2_X1 i_257_76_13201 (.A1(n_257_76_13177), .A2(n_257_76_13113), .ZN(
      n_257_76_13178));
   NAND4_X1 i_257_76_13202 (.A1(n_257_76_13042), .A2(n_257_76_13065), .A3(
      n_257_76_13111), .A4(n_257_76_13137), .ZN(n_257_76_13179));
   INV_X1 i_257_76_13203 (.A(n_257_76_13179), .ZN(n_257_76_13180));
   NAND3_X1 i_257_76_13204 (.A1(n_257_76_13178), .A2(n_257_76_13180), .A3(
      n_257_76_13133), .ZN(n_257_76_13181));
   NAND2_X1 i_257_76_13205 (.A1(n_257_76_13116), .A2(n_257_76_13117), .ZN(
      n_257_76_13182));
   NOR2_X1 i_257_76_13206 (.A1(n_257_76_13181), .A2(n_257_76_13182), .ZN(
      n_257_76_13183));
   NAND2_X1 i_257_76_13207 (.A1(n_257_76_13041), .A2(n_257_76_13083), .ZN(
      n_257_76_13184));
   INV_X1 i_257_76_13208 (.A(n_257_76_13184), .ZN(n_257_76_13185));
   NAND3_X1 i_257_76_13209 (.A1(n_257_76_13183), .A2(n_257_76_13185), .A3(
      n_257_76_13052), .ZN(n_257_76_13186));
   INV_X1 i_257_76_13210 (.A(n_257_76_13186), .ZN(n_257_76_13187));
   NAND2_X1 i_257_76_13211 (.A1(n_257_76_18074), .A2(n_257_76_13187), .ZN(
      n_257_76_13188));
   NAND3_X1 i_257_76_13212 (.A1(n_257_76_13154), .A2(n_257_76_13168), .A3(
      n_257_76_13188), .ZN(n_257_76_13189));
   NAND2_X1 i_257_76_13213 (.A1(n_257_1082), .A2(n_257_442), .ZN(n_257_76_13190));
   INV_X1 i_257_76_13214 (.A(n_257_76_13190), .ZN(n_257_76_13191));
   NAND2_X1 i_257_76_13215 (.A1(n_257_13), .A2(n_257_76_13191), .ZN(
      n_257_76_13192));
   NOR2_X1 i_257_76_13216 (.A1(n_257_76_17902), .A2(n_257_1082), .ZN(
      n_257_76_13193));
   NAND4_X1 i_257_76_13217 (.A1(n_257_76_13193), .A2(n_257_76_13076), .A3(
      n_257_884), .A4(n_257_76_13077), .ZN(n_257_76_13194));
   INV_X1 i_257_76_13218 (.A(n_257_76_13194), .ZN(n_257_76_13195));
   NAND3_X1 i_257_76_13219 (.A1(n_257_76_13195), .A2(n_257_76_13064), .A3(
      n_257_76_13042), .ZN(n_257_76_13196));
   INV_X1 i_257_76_13220 (.A(n_257_76_13196), .ZN(n_257_76_13197));
   NAND2_X1 i_257_76_13221 (.A1(n_257_76_13041), .A2(n_257_76_13197), .ZN(
      n_257_76_13198));
   INV_X1 i_257_76_13222 (.A(n_257_76_13198), .ZN(n_257_76_13199));
   NAND2_X1 i_257_76_13223 (.A1(n_257_76_13199), .A2(n_257_76_13052), .ZN(
      n_257_76_13200));
   INV_X1 i_257_76_13224 (.A(n_257_76_13200), .ZN(n_257_76_13201));
   NAND2_X1 i_257_76_13225 (.A1(n_257_76_18077), .A2(n_257_76_13201), .ZN(
      n_257_76_13202));
   NAND2_X1 i_257_76_13226 (.A1(n_257_76_13192), .A2(n_257_76_13202), .ZN(
      n_257_76_13203));
   NOR2_X1 i_257_76_13227 (.A1(n_257_76_13189), .A2(n_257_76_13203), .ZN(
      n_257_76_13204));
   NAND2_X1 i_257_76_13228 (.A1(n_257_76_13052), .A2(n_257_76_13041), .ZN(
      n_257_76_13205));
   NAND3_X1 i_257_76_13229 (.A1(n_257_76_13076), .A2(n_257_76_13077), .A3(
      n_257_76_13126), .ZN(n_257_76_13206));
   NAND2_X1 i_257_76_13230 (.A1(n_257_76_13123), .A2(n_257_426), .ZN(
      n_257_76_13207));
   INV_X1 i_257_76_13231 (.A(n_257_76_13207), .ZN(n_257_76_13208));
   NAND4_X1 i_257_76_13232 (.A1(n_257_76_13078), .A2(n_257_76_13208), .A3(
      n_257_76_13043), .A4(n_257_76_18002), .ZN(n_257_76_13209));
   NOR2_X1 i_257_76_13233 (.A1(n_257_76_13206), .A2(n_257_76_13209), .ZN(
      n_257_76_13210));
   NAND3_X1 i_257_76_13234 (.A1(n_257_76_13067), .A2(n_257_76_13068), .A3(
      n_257_76_13128), .ZN(n_257_76_13211));
   INV_X1 i_257_76_13235 (.A(n_257_76_13211), .ZN(n_257_76_13212));
   NAND3_X1 i_257_76_13236 (.A1(n_257_76_13210), .A2(n_257_76_13212), .A3(
      n_257_76_13074), .ZN(n_257_76_13213));
   NOR2_X1 i_257_76_13237 (.A1(n_257_76_13213), .A2(n_257_76_13179), .ZN(
      n_257_76_13214));
   NAND3_X1 i_257_76_13238 (.A1(n_257_76_13133), .A2(n_257_76_13117), .A3(
      n_257_556), .ZN(n_257_76_13215));
   INV_X1 i_257_76_13239 (.A(n_257_76_13215), .ZN(n_257_76_13216));
   NAND4_X1 i_257_76_13240 (.A1(n_257_76_13214), .A2(n_257_76_13216), .A3(
      n_257_76_13083), .A4(n_257_76_13116), .ZN(n_257_76_13217));
   NOR2_X1 i_257_76_13241 (.A1(n_257_76_13205), .A2(n_257_76_13217), .ZN(
      n_257_76_13218));
   NAND2_X1 i_257_76_13242 (.A1(n_257_76_18076), .A2(n_257_76_13218), .ZN(
      n_257_76_13219));
   NAND2_X1 i_257_76_13243 (.A1(n_257_756), .A2(n_257_76_13071), .ZN(
      n_257_76_13220));
   INV_X1 i_257_76_13244 (.A(n_257_76_13220), .ZN(n_257_76_13221));
   NOR2_X1 i_257_76_13245 (.A1(n_257_1082), .A2(n_257_76_17934), .ZN(
      n_257_76_13222));
   NAND3_X1 i_257_76_13246 (.A1(n_257_76_13222), .A2(n_257_76_13076), .A3(
      n_257_76_13077), .ZN(n_257_76_13223));
   INV_X1 i_257_76_13247 (.A(n_257_76_13223), .ZN(n_257_76_13224));
   NAND3_X1 i_257_76_13248 (.A1(n_257_76_13221), .A2(n_257_76_13156), .A3(
      n_257_76_13224), .ZN(n_257_76_13225));
   NAND3_X1 i_257_76_13249 (.A1(n_257_76_13064), .A2(n_257_76_13042), .A3(
      n_257_76_13065), .ZN(n_257_76_13226));
   NOR2_X1 i_257_76_13250 (.A1(n_257_76_13225), .A2(n_257_76_13226), .ZN(
      n_257_76_13227));
   NAND2_X1 i_257_76_13251 (.A1(n_257_76_13041), .A2(n_257_76_13227), .ZN(
      n_257_76_13228));
   INV_X1 i_257_76_13252 (.A(n_257_76_13228), .ZN(n_257_76_13229));
   NAND2_X1 i_257_76_13253 (.A1(n_257_76_13229), .A2(n_257_76_13052), .ZN(
      n_257_76_13230));
   INV_X1 i_257_76_13254 (.A(n_257_76_13230), .ZN(n_257_76_13231));
   NAND2_X1 i_257_76_13255 (.A1(n_257_76_18069), .A2(n_257_76_13231), .ZN(
      n_257_76_13232));
   NAND2_X1 i_257_76_13256 (.A1(n_257_620), .A2(n_257_442), .ZN(n_257_76_13233));
   INV_X1 i_257_76_13257 (.A(n_257_76_13233), .ZN(n_257_76_13234));
   NAND2_X1 i_257_76_13258 (.A1(n_257_76_13234), .A2(n_257_432), .ZN(
      n_257_76_13235));
   INV_X1 i_257_76_13259 (.A(n_257_76_13235), .ZN(n_257_76_13236));
   NAND3_X1 i_257_76_13260 (.A1(n_257_76_13078), .A2(n_257_76_13043), .A3(
      n_257_76_13236), .ZN(n_257_76_13237));
   INV_X1 i_257_76_13261 (.A(n_257_76_13237), .ZN(n_257_76_13238));
   NAND4_X1 i_257_76_13262 (.A1(n_257_76_13170), .A2(n_257_76_13238), .A3(
      n_257_76_13068), .A4(n_257_76_13128), .ZN(n_257_76_13239));
   NOR2_X1 i_257_76_13263 (.A1(n_257_76_13239), .A2(n_257_76_13113), .ZN(
      n_257_76_13240));
   INV_X1 i_257_76_13264 (.A(n_257_76_13162), .ZN(n_257_76_13241));
   NAND3_X1 i_257_76_13265 (.A1(n_257_76_13065), .A2(n_257_76_13111), .A3(
      n_257_76_13137), .ZN(n_257_76_13242));
   INV_X1 i_257_76_13266 (.A(n_257_76_13242), .ZN(n_257_76_13243));
   NAND3_X1 i_257_76_13267 (.A1(n_257_76_13240), .A2(n_257_76_13241), .A3(
      n_257_76_13243), .ZN(n_257_76_13244));
   INV_X1 i_257_76_13268 (.A(n_257_76_13244), .ZN(n_257_76_13245));
   NAND3_X1 i_257_76_13269 (.A1(n_257_76_13245), .A2(n_257_76_13041), .A3(
      n_257_76_13083), .ZN(n_257_76_13246));
   NOR2_X1 i_257_76_13270 (.A1(n_257_76_13246), .A2(n_257_76_13062), .ZN(
      n_257_76_13247));
   NAND2_X1 i_257_76_13271 (.A1(n_257_68), .A2(n_257_76_13247), .ZN(
      n_257_76_13248));
   NAND3_X1 i_257_76_13272 (.A1(n_257_76_13219), .A2(n_257_76_13232), .A3(
      n_257_76_13248), .ZN(n_257_76_13249));
   NOR2_X1 i_257_76_13273 (.A1(n_257_1082), .A2(n_257_76_17951), .ZN(
      n_257_76_13250));
   NAND3_X1 i_257_76_13274 (.A1(n_257_76_13250), .A2(n_257_76_13076), .A3(
      n_257_76_13077), .ZN(n_257_76_13251));
   INV_X1 i_257_76_13275 (.A(n_257_76_13251), .ZN(n_257_76_13252));
   NAND4_X1 i_257_76_13276 (.A1(n_257_76_13252), .A2(n_257_76_13071), .A3(
      n_257_820), .A4(n_257_76_13068), .ZN(n_257_76_13253));
   NOR2_X1 i_257_76_13277 (.A1(n_257_76_13253), .A2(n_257_76_13088), .ZN(
      n_257_76_13254));
   NAND2_X1 i_257_76_13278 (.A1(n_257_76_13041), .A2(n_257_76_13254), .ZN(
      n_257_76_13255));
   INV_X1 i_257_76_13279 (.A(n_257_76_13255), .ZN(n_257_76_13256));
   NAND2_X1 i_257_76_13280 (.A1(n_257_76_13256), .A2(n_257_76_13052), .ZN(
      n_257_76_13257));
   INV_X1 i_257_76_13281 (.A(n_257_76_13257), .ZN(n_257_76_13258));
   NAND2_X1 i_257_76_13282 (.A1(n_257_22), .A2(n_257_76_13258), .ZN(
      n_257_76_13259));
   NAND2_X1 i_257_76_13283 (.A1(n_257_444), .A2(n_257_76_13056), .ZN(
      n_257_76_13260));
   INV_X1 i_257_76_13284 (.A(n_257_76_13260), .ZN(n_257_76_13261));
   NAND2_X1 i_257_76_13285 (.A1(n_257_1018), .A2(n_257_76_13261), .ZN(
      n_257_76_13262));
   INV_X1 i_257_76_13286 (.A(n_257_76_13262), .ZN(n_257_76_13263));
   NAND2_X1 i_257_76_13287 (.A1(n_257_76_13052), .A2(n_257_76_13263), .ZN(
      n_257_76_13264));
   INV_X1 i_257_76_13288 (.A(n_257_76_13264), .ZN(n_257_76_13265));
   NAND2_X1 i_257_76_13289 (.A1(n_257_76_18075), .A2(n_257_76_13265), .ZN(
      n_257_76_13266));
   NAND2_X1 i_257_76_13290 (.A1(n_257_76_13259), .A2(n_257_76_13266), .ZN(
      n_257_76_13267));
   NOR2_X1 i_257_76_13291 (.A1(n_257_76_13249), .A2(n_257_76_13267), .ZN(
      n_257_76_13268));
   NAND3_X1 i_257_76_13292 (.A1(n_257_76_13146), .A2(n_257_76_13204), .A3(
      n_257_76_13268), .ZN(n_257_76_13269));
   INV_X1 i_257_76_13293 (.A(n_257_76_13269), .ZN(n_257_76_13270));
   NOR2_X1 i_257_76_13294 (.A1(n_257_1082), .A2(n_257_76_17633), .ZN(
      n_257_76_13271));
   NAND3_X1 i_257_76_13295 (.A1(n_257_76_13271), .A2(n_257_58), .A3(
      n_257_76_13078), .ZN(n_257_76_13272));
   INV_X1 i_257_76_13296 (.A(n_257_76_13272), .ZN(n_257_76_13273));
   NAND3_X1 i_257_76_13297 (.A1(n_257_76_13273), .A2(n_257_76_13170), .A3(
      n_257_76_13068), .ZN(n_257_76_13274));
   INV_X1 i_257_76_13298 (.A(n_257_76_13274), .ZN(n_257_76_13275));
   INV_X1 i_257_76_13299 (.A(n_257_76_13113), .ZN(n_257_76_13276));
   NAND2_X1 i_257_76_13300 (.A1(n_257_76_13275), .A2(n_257_76_13276), .ZN(
      n_257_76_13277));
   NOR3_X1 i_257_76_13301 (.A1(n_257_76_13277), .A2(n_257_76_13162), .A3(
      n_257_76_13242), .ZN(n_257_76_13278));
   NAND3_X1 i_257_76_13302 (.A1(n_257_76_13278), .A2(n_257_76_13041), .A3(
      n_257_76_13083), .ZN(n_257_76_13279));
   NOR2_X1 i_257_76_13303 (.A1(n_257_76_13279), .A2(n_257_76_13062), .ZN(
      n_257_76_13280));
   NAND2_X1 i_257_76_13304 (.A1(n_257_76_18081), .A2(n_257_76_13280), .ZN(
      n_257_76_13281));
   NAND2_X1 i_257_76_13305 (.A1(n_257_76_13071), .A2(n_257_76_13067), .ZN(
      n_257_76_13282));
   INV_X1 i_257_76_13306 (.A(n_257_76_13282), .ZN(n_257_76_13283));
   NOR2_X1 i_257_76_13307 (.A1(n_257_1082), .A2(n_257_76_17675), .ZN(
      n_257_76_13284));
   NAND4_X1 i_257_76_13308 (.A1(n_257_76_13284), .A2(n_257_76_13076), .A3(
      n_257_76_13077), .A4(n_257_76_13078), .ZN(n_257_76_13285));
   INV_X1 i_257_76_13309 (.A(n_257_76_13285), .ZN(n_257_76_13286));
   NAND2_X1 i_257_76_13310 (.A1(n_257_76_13068), .A2(n_257_449), .ZN(
      n_257_76_13287));
   INV_X1 i_257_76_13311 (.A(n_257_76_13287), .ZN(n_257_76_13288));
   NAND3_X1 i_257_76_13312 (.A1(n_257_76_13283), .A2(n_257_76_13286), .A3(
      n_257_76_13288), .ZN(n_257_76_13289));
   NOR2_X1 i_257_76_13313 (.A1(n_257_76_13066), .A2(n_257_76_13289), .ZN(
      n_257_76_13290));
   NAND3_X1 i_257_76_13314 (.A1(n_257_76_13041), .A2(n_257_76_13290), .A3(
      n_257_76_13083), .ZN(n_257_76_13291));
   NOR2_X1 i_257_76_13315 (.A1(n_257_76_13062), .A2(n_257_76_13291), .ZN(
      n_257_76_13292));
   NAND2_X1 i_257_76_13316 (.A1(n_257_76_18083), .A2(n_257_76_13292), .ZN(
      n_257_76_13293));
   NAND3_X1 i_257_76_13317 (.A1(n_257_76_18003), .A2(n_257_76_13078), .A3(
      n_257_76_13043), .ZN(n_257_76_13294));
   NOR2_X1 i_257_76_13318 (.A1(n_257_76_13169), .A2(n_257_76_13294), .ZN(
      n_257_76_13295));
   NAND3_X1 i_257_76_13319 (.A1(n_257_76_13212), .A2(n_257_76_13074), .A3(
      n_257_76_13295), .ZN(n_257_76_13296));
   NOR2_X1 i_257_76_13320 (.A1(n_257_76_13296), .A2(n_257_76_13179), .ZN(
      n_257_76_13297));
   NAND3_X1 i_257_76_13321 (.A1(n_257_76_13133), .A2(n_257_76_13117), .A3(
      n_257_175), .ZN(n_257_76_13298));
   INV_X1 i_257_76_13322 (.A(n_257_76_13298), .ZN(n_257_76_13299));
   NAND4_X1 i_257_76_13323 (.A1(n_257_76_13041), .A2(n_257_76_13297), .A3(
      n_257_76_13083), .A4(n_257_76_13299), .ZN(n_257_76_13300));
   NOR2_X1 i_257_76_13324 (.A1(n_257_76_13300), .A2(n_257_76_13062), .ZN(
      n_257_76_13301));
   NAND2_X1 i_257_76_13325 (.A1(n_257_76_18061), .A2(n_257_76_13301), .ZN(
      n_257_76_13302));
   NAND3_X1 i_257_76_13326 (.A1(n_257_76_13281), .A2(n_257_76_13293), .A3(
      n_257_76_13302), .ZN(n_257_76_13303));
   INV_X1 i_257_76_13327 (.A(n_257_76_13303), .ZN(n_257_76_13304));
   NAND3_X1 i_257_76_13328 (.A1(n_257_438), .A2(n_257_76_13043), .A3(
      n_257_76_16422), .ZN(n_257_76_13305));
   INV_X1 i_257_76_13329 (.A(n_257_76_13076), .ZN(n_257_76_13306));
   NOR2_X1 i_257_76_13330 (.A1(n_257_76_13305), .A2(n_257_76_13306), .ZN(
      n_257_76_13307));
   NAND3_X1 i_257_76_13331 (.A1(n_257_76_13307), .A2(n_257_76_13064), .A3(
      n_257_76_13042), .ZN(n_257_76_13308));
   INV_X1 i_257_76_13332 (.A(n_257_76_13308), .ZN(n_257_76_13309));
   NAND2_X1 i_257_76_13333 (.A1(n_257_76_13041), .A2(n_257_76_13309), .ZN(
      n_257_76_13310));
   INV_X1 i_257_76_13334 (.A(n_257_76_13310), .ZN(n_257_76_13311));
   NAND2_X1 i_257_76_13335 (.A1(n_257_76_13311), .A2(n_257_76_13052), .ZN(
      n_257_76_13312));
   INV_X1 i_257_76_13336 (.A(n_257_76_13312), .ZN(n_257_76_13313));
   NAND2_X1 i_257_76_13337 (.A1(n_257_76_18067), .A2(n_257_76_13313), .ZN(
      n_257_76_13314));
   NAND2_X1 i_257_76_13338 (.A1(n_257_76_13119), .A2(n_257_76_13115), .ZN(
      n_257_76_13315));
   NOR2_X1 i_257_76_13339 (.A1(n_257_76_13315), .A2(n_257_76_13182), .ZN(
      n_257_76_13316));
   NAND2_X1 i_257_76_13340 (.A1(n_257_76_13063), .A2(n_257_76_13131), .ZN(
      n_257_76_13317));
   NAND2_X1 i_257_76_13341 (.A1(n_257_372), .A2(n_257_421), .ZN(n_257_76_13318));
   NAND2_X1 i_257_76_13342 (.A1(n_257_76_13318), .A2(n_257_76_13064), .ZN(
      n_257_76_13319));
   NOR2_X1 i_257_76_13343 (.A1(n_257_76_13317), .A2(n_257_76_13319), .ZN(
      n_257_76_13320));
   NAND2_X1 i_257_76_13344 (.A1(n_257_76_13042), .A2(n_257_76_13065), .ZN(
      n_257_76_13321));
   NAND2_X1 i_257_76_13345 (.A1(n_257_76_13111), .A2(n_257_76_13137), .ZN(
      n_257_76_13322));
   NOR2_X1 i_257_76_13346 (.A1(n_257_76_13321), .A2(n_257_76_13322), .ZN(
      n_257_76_13323));
   NAND2_X1 i_257_76_13347 (.A1(n_257_76_13320), .A2(n_257_76_13323), .ZN(
      n_257_76_13324));
   NAND2_X1 i_257_76_13348 (.A1(n_257_333), .A2(n_257_422), .ZN(n_257_76_13325));
   NAND2_X1 i_257_76_13349 (.A1(n_257_76_13325), .A2(n_257_76_13126), .ZN(
      n_257_76_13326));
   INV_X1 i_257_76_13350 (.A(n_257_76_13077), .ZN(n_257_76_13327));
   NOR2_X1 i_257_76_13351 (.A1(n_257_76_13326), .A2(n_257_76_13327), .ZN(
      n_257_76_13328));
   NAND2_X1 i_257_76_13352 (.A1(n_257_76_13078), .A2(n_257_76_13043), .ZN(
      n_257_76_13329));
   NAND2_X1 i_257_76_13353 (.A1(n_257_76_13123), .A2(n_257_420), .ZN(
      n_257_76_13330));
   INV_X1 i_257_76_13354 (.A(n_257_76_13330), .ZN(n_257_76_13331));
   NAND2_X1 i_257_76_13355 (.A1(n_257_442), .A2(n_257_492), .ZN(n_257_76_13332));
   NAND2_X1 i_257_76_13356 (.A1(n_257_76_13331), .A2(n_257_76_18004), .ZN(
      n_257_76_13333));
   NOR2_X1 i_257_76_13357 (.A1(n_257_76_13329), .A2(n_257_76_13333), .ZN(
      n_257_76_13334));
   NAND2_X1 i_257_76_13358 (.A1(n_257_76_13328), .A2(n_257_76_13334), .ZN(
      n_257_76_13335));
   INV_X1 i_257_76_13359 (.A(n_257_76_13335), .ZN(n_257_76_13336));
   NAND2_X1 i_257_76_13360 (.A1(n_257_76_13128), .A2(n_257_76_13076), .ZN(
      n_257_76_13337));
   NOR2_X1 i_257_76_13361 (.A1(n_257_76_13135), .A2(n_257_76_13337), .ZN(
      n_257_76_13338));
   NAND2_X1 i_257_76_13362 (.A1(n_257_76_13336), .A2(n_257_76_13338), .ZN(
      n_257_76_13339));
   INV_X1 i_257_76_13363 (.A(n_257_76_13339), .ZN(n_257_76_13340));
   NAND2_X1 i_257_76_13364 (.A1(n_257_295), .A2(n_257_423), .ZN(n_257_76_13341));
   NAND2_X1 i_257_76_13365 (.A1(n_257_76_13341), .A2(n_257_76_13071), .ZN(
      n_257_76_13342));
   NAND2_X1 i_257_76_13366 (.A1(n_257_76_13072), .A2(n_257_76_13067), .ZN(
      n_257_76_13343));
   NOR2_X1 i_257_76_13367 (.A1(n_257_76_13342), .A2(n_257_76_13343), .ZN(
      n_257_76_13344));
   NAND2_X1 i_257_76_13368 (.A1(n_257_76_13340), .A2(n_257_76_13344), .ZN(
      n_257_76_13345));
   NOR2_X1 i_257_76_13369 (.A1(n_257_76_13324), .A2(n_257_76_13345), .ZN(
      n_257_76_13346));
   NAND2_X1 i_257_76_13370 (.A1(n_257_76_13316), .A2(n_257_76_13346), .ZN(
      n_257_76_13347));
   NAND2_X1 i_257_76_13371 (.A1(n_257_76_13185), .A2(n_257_76_13052), .ZN(
      n_257_76_13348));
   NOR2_X1 i_257_76_13372 (.A1(n_257_76_13347), .A2(n_257_76_13348), .ZN(
      n_257_76_13349));
   NAND2_X1 i_257_76_13373 (.A1(n_257_76_18073), .A2(n_257_76_13349), .ZN(
      n_257_76_13350));
   NAND3_X1 i_257_76_13374 (.A1(n_257_76_13078), .A2(n_257_76_18005), .A3(
      n_257_76_13043), .ZN(n_257_76_13351));
   NOR2_X1 i_257_76_13375 (.A1(n_257_76_13169), .A2(n_257_76_13351), .ZN(
      n_257_76_13352));
   NAND3_X1 i_257_76_13376 (.A1(n_257_76_13212), .A2(n_257_76_13074), .A3(
      n_257_76_13352), .ZN(n_257_76_13353));
   NAND4_X1 i_257_76_13377 (.A1(n_257_76_13065), .A2(n_257_76_13111), .A3(
      n_257_76_13137), .A4(n_257_136), .ZN(n_257_76_13354));
   NOR2_X1 i_257_76_13378 (.A1(n_257_76_13353), .A2(n_257_76_13354), .ZN(
      n_257_76_13355));
   NAND2_X1 i_257_76_13379 (.A1(n_257_76_13241), .A2(n_257_76_13117), .ZN(
      n_257_76_13356));
   INV_X1 i_257_76_13380 (.A(n_257_76_13356), .ZN(n_257_76_13357));
   NAND3_X1 i_257_76_13381 (.A1(n_257_76_13355), .A2(n_257_76_13357), .A3(
      n_257_76_13083), .ZN(n_257_76_13358));
   INV_X1 i_257_76_13382 (.A(n_257_76_13358), .ZN(n_257_76_13359));
   NAND3_X1 i_257_76_13383 (.A1(n_257_76_13359), .A2(n_257_76_13052), .A3(
      n_257_76_13041), .ZN(n_257_76_13360));
   INV_X1 i_257_76_13384 (.A(n_257_76_13360), .ZN(n_257_76_13361));
   NAND2_X1 i_257_76_13385 (.A1(n_257_76_18068), .A2(n_257_76_13361), .ZN(
      n_257_76_13362));
   NAND3_X1 i_257_76_13386 (.A1(n_257_76_13314), .A2(n_257_76_13350), .A3(
      n_257_76_13362), .ZN(n_257_76_13363));
   INV_X1 i_257_76_13387 (.A(n_257_76_13363), .ZN(n_257_76_13364));
   NAND2_X1 i_257_76_13388 (.A1(n_257_788), .A2(n_257_442), .ZN(n_257_76_13365));
   NOR2_X1 i_257_76_13389 (.A1(n_257_1082), .A2(n_257_76_13365), .ZN(
      n_257_76_13366));
   NAND2_X1 i_257_76_13390 (.A1(n_257_76_13077), .A2(n_257_76_13366), .ZN(
      n_257_76_13367));
   INV_X1 i_257_76_13391 (.A(n_257_76_13367), .ZN(n_257_76_13368));
   NAND2_X1 i_257_76_13392 (.A1(n_257_447), .A2(n_257_76_13076), .ZN(
      n_257_76_13369));
   INV_X1 i_257_76_13393 (.A(n_257_76_13369), .ZN(n_257_76_13370));
   NAND4_X1 i_257_76_13394 (.A1(n_257_76_13368), .A2(n_257_76_13370), .A3(
      n_257_76_13071), .A4(n_257_76_13068), .ZN(n_257_76_13371));
   NOR2_X1 i_257_76_13395 (.A1(n_257_76_13226), .A2(n_257_76_13371), .ZN(
      n_257_76_13372));
   NAND2_X1 i_257_76_13396 (.A1(n_257_76_13041), .A2(n_257_76_13372), .ZN(
      n_257_76_13373));
   INV_X1 i_257_76_13397 (.A(n_257_76_13373), .ZN(n_257_76_13374));
   NAND2_X1 i_257_76_13398 (.A1(n_257_76_13374), .A2(n_257_76_13052), .ZN(
      n_257_76_13375));
   INV_X1 i_257_76_13399 (.A(n_257_76_13375), .ZN(n_257_76_13376));
   NAND3_X1 i_257_76_13400 (.A1(n_257_76_13078), .A2(n_257_76_18006), .A3(
      n_257_76_13043), .ZN(n_257_76_13377));
   NOR2_X1 i_257_76_13401 (.A1(n_257_76_13169), .A2(n_257_76_13377), .ZN(
      n_257_76_13378));
   NAND2_X1 i_257_76_13402 (.A1(n_257_76_13068), .A2(n_257_76_13128), .ZN(
      n_257_76_13379));
   INV_X1 i_257_76_13403 (.A(n_257_76_13379), .ZN(n_257_76_13380));
   NAND3_X1 i_257_76_13404 (.A1(n_257_76_13378), .A2(n_257_76_13380), .A3(
      n_257_76_13067), .ZN(n_257_76_13381));
   NAND4_X1 i_257_76_13405 (.A1(n_257_76_13111), .A2(n_257_76_13137), .A3(
      n_257_76_13071), .A4(n_257_76_13072), .ZN(n_257_76_13382));
   NOR2_X1 i_257_76_13406 (.A1(n_257_76_13381), .A2(n_257_76_13382), .ZN(
      n_257_76_13383));
   NAND2_X1 i_257_76_13407 (.A1(n_257_98), .A2(n_257_76_13063), .ZN(
      n_257_76_13384));
   NOR2_X1 i_257_76_13408 (.A1(n_257_76_13384), .A2(n_257_76_13226), .ZN(
      n_257_76_13385));
   NAND3_X1 i_257_76_13409 (.A1(n_257_76_13083), .A2(n_257_76_13383), .A3(
      n_257_76_13385), .ZN(n_257_76_13386));
   INV_X1 i_257_76_13410 (.A(n_257_76_13386), .ZN(n_257_76_13387));
   NAND3_X1 i_257_76_13411 (.A1(n_257_76_13387), .A2(n_257_76_13052), .A3(
      n_257_76_13041), .ZN(n_257_76_13388));
   INV_X1 i_257_76_13412 (.A(n_257_76_13388), .ZN(n_257_76_13389));
   AOI22_X1 i_257_76_13413 (.A1(n_257_76_18085), .A2(n_257_76_13376), .B1(
      n_257_76_18080), .B2(n_257_76_13389), .ZN(n_257_76_13390));
   NAND3_X1 i_257_76_13414 (.A1(n_257_76_13304), .A2(n_257_76_13364), .A3(
      n_257_76_13390), .ZN(n_257_76_13391));
   OAI21_X1 i_257_76_13415 (.A(n_257_76_17761), .B1(n_257_724), .B2(
      n_257_76_17412), .ZN(n_257_76_13392));
   NAND2_X1 i_257_76_13416 (.A1(n_257_76_13068), .A2(n_257_76_13392), .ZN(
      n_257_76_13393));
   INV_X1 i_257_76_13417 (.A(n_257_76_13393), .ZN(n_257_76_13394));
   NAND3_X1 i_257_76_13418 (.A1(n_257_76_13076), .A2(n_257_76_13077), .A3(
      n_257_76_13043), .ZN(n_257_76_13395));
   INV_X1 i_257_76_13419 (.A(n_257_76_13395), .ZN(n_257_76_13396));
   NAND3_X1 i_257_76_13420 (.A1(n_257_76_13394), .A2(n_257_76_13065), .A3(
      n_257_76_13396), .ZN(n_257_76_13397));
   NAND2_X1 i_257_76_13421 (.A1(n_257_76_13063), .A2(n_257_76_13064), .ZN(
      n_257_76_13398));
   NOR2_X1 i_257_76_13422 (.A1(n_257_76_13397), .A2(n_257_76_13398), .ZN(
      n_257_76_13399));
   NAND3_X1 i_257_76_13423 (.A1(n_257_76_13071), .A2(n_257_76_13067), .A3(
      n_257_448), .ZN(n_257_76_13400));
   INV_X1 i_257_76_13424 (.A(n_257_76_13042), .ZN(n_257_76_13401));
   NOR2_X1 i_257_76_13425 (.A1(n_257_76_13400), .A2(n_257_76_13401), .ZN(
      n_257_76_13402));
   NAND2_X1 i_257_76_13426 (.A1(n_257_692), .A2(n_257_76_13402), .ZN(
      n_257_76_13403));
   INV_X1 i_257_76_13427 (.A(n_257_76_13403), .ZN(n_257_76_13404));
   NAND3_X1 i_257_76_13428 (.A1(n_257_76_13041), .A2(n_257_76_13399), .A3(
      n_257_76_13404), .ZN(n_257_76_13405));
   NOR2_X1 i_257_76_13429 (.A1(n_257_76_13062), .A2(n_257_76_13405), .ZN(
      n_257_76_13406));
   NAND2_X1 i_257_76_13430 (.A1(n_257_76_18079), .A2(n_257_76_13406), .ZN(
      n_257_76_13407));
   INV_X1 i_257_76_13431 (.A(n_257_76_18002), .ZN(n_257_76_13408));
   NOR2_X1 i_257_76_13432 (.A1(n_257_76_13408), .A2(n_257_1082), .ZN(
      n_257_76_13409));
   NAND2_X1 i_257_76_13433 (.A1(n_257_76_13123), .A2(n_257_425), .ZN(
      n_257_76_13410));
   INV_X1 i_257_76_13434 (.A(n_257_76_13410), .ZN(n_257_76_13411));
   NAND4_X1 i_257_76_13435 (.A1(n_257_76_13409), .A2(n_257_76_13126), .A3(
      n_257_76_13078), .A4(n_257_76_13411), .ZN(n_257_76_13412));
   NAND3_X1 i_257_76_13436 (.A1(n_257_76_13128), .A2(n_257_76_13076), .A3(
      n_257_76_13077), .ZN(n_257_76_13413));
   NOR2_X1 i_257_76_13437 (.A1(n_257_76_13412), .A2(n_257_76_13413), .ZN(
      n_257_76_13414));
   NAND2_X1 i_257_76_13438 (.A1(n_257_76_13137), .A2(n_257_76_13071), .ZN(
      n_257_76_13415));
   INV_X1 i_257_76_13439 (.A(n_257_76_13415), .ZN(n_257_76_13416));
   NAND3_X1 i_257_76_13440 (.A1(n_257_76_13072), .A2(n_257_76_13067), .A3(
      n_257_76_13068), .ZN(n_257_76_13417));
   INV_X1 i_257_76_13441 (.A(n_257_76_13417), .ZN(n_257_76_13418));
   NAND3_X1 i_257_76_13442 (.A1(n_257_76_13414), .A2(n_257_76_13416), .A3(
      n_257_76_13418), .ZN(n_257_76_13419));
   NAND4_X1 i_257_76_13443 (.A1(n_257_76_13064), .A2(n_257_76_13042), .A3(
      n_257_76_13065), .A4(n_257_76_13111), .ZN(n_257_76_13420));
   NOR2_X1 i_257_76_13444 (.A1(n_257_76_13419), .A2(n_257_76_13420), .ZN(
      n_257_76_13421));
   NAND2_X1 i_257_76_13445 (.A1(n_257_76_13119), .A2(n_257_76_13116), .ZN(
      n_257_76_13422));
   INV_X1 i_257_76_13446 (.A(n_257_76_13422), .ZN(n_257_76_13423));
   INV_X1 i_257_76_13447 (.A(n_257_76_13317), .ZN(n_257_76_13424));
   NAND3_X1 i_257_76_13448 (.A1(n_257_76_13117), .A2(n_257_255), .A3(
      n_257_76_13424), .ZN(n_257_76_13425));
   INV_X1 i_257_76_13449 (.A(n_257_76_13425), .ZN(n_257_76_13426));
   NAND4_X1 i_257_76_13450 (.A1(n_257_76_13421), .A2(n_257_76_13423), .A3(
      n_257_76_13083), .A4(n_257_76_13426), .ZN(n_257_76_13427));
   NOR2_X1 i_257_76_13451 (.A1(n_257_76_13427), .A2(n_257_76_13205), .ZN(
      n_257_76_13428));
   NAND2_X1 i_257_76_13452 (.A1(n_257_76_18064), .A2(n_257_76_13428), .ZN(
      n_257_76_13429));
   NAND3_X1 i_257_76_13453 (.A1(n_257_76_13068), .A2(n_257_76_13134), .A3(
      n_257_76_13128), .ZN(n_257_76_13430));
   INV_X1 i_257_76_13454 (.A(n_257_76_13430), .ZN(n_257_76_13431));
   NAND2_X1 i_257_76_13455 (.A1(n_257_76_13123), .A2(n_257_421), .ZN(
      n_257_76_13432));
   INV_X1 i_257_76_13456 (.A(n_257_76_13432), .ZN(n_257_76_13433));
   NAND4_X1 i_257_76_13457 (.A1(n_257_76_13409), .A2(n_257_76_13126), .A3(
      n_257_76_13078), .A4(n_257_76_13433), .ZN(n_257_76_13434));
   INV_X1 i_257_76_13458 (.A(n_257_76_13434), .ZN(n_257_76_13435));
   NAND3_X1 i_257_76_13459 (.A1(n_257_76_13076), .A2(n_257_76_13077), .A3(
      n_257_76_13325), .ZN(n_257_76_13436));
   INV_X1 i_257_76_13460 (.A(n_257_76_13436), .ZN(n_257_76_13437));
   NAND3_X1 i_257_76_13461 (.A1(n_257_76_13431), .A2(n_257_76_13435), .A3(
      n_257_76_13437), .ZN(n_257_76_13438));
   INV_X1 i_257_76_13462 (.A(n_257_76_13438), .ZN(n_257_76_13439));
   NAND4_X1 i_257_76_13463 (.A1(n_257_76_13065), .A2(n_257_76_13137), .A3(
      n_257_76_13341), .A4(n_257_372), .ZN(n_257_76_13440));
   INV_X1 i_257_76_13464 (.A(n_257_76_13440), .ZN(n_257_76_13441));
   NAND3_X1 i_257_76_13465 (.A1(n_257_76_13439), .A2(n_257_76_13133), .A3(
      n_257_76_13441), .ZN(n_257_76_13442));
   INV_X1 i_257_76_13466 (.A(n_257_76_13442), .ZN(n_257_76_13443));
   NAND2_X1 i_257_76_13467 (.A1(n_257_76_13041), .A2(n_257_76_13443), .ZN(
      n_257_76_13444));
   INV_X1 i_257_76_13468 (.A(n_257_76_13444), .ZN(n_257_76_13445));
   NAND3_X1 i_257_76_13469 (.A1(n_257_76_13121), .A2(n_257_76_13445), .A3(
      n_257_76_13052), .ZN(n_257_76_13446));
   INV_X1 i_257_76_13470 (.A(n_257_76_13446), .ZN(n_257_76_13447));
   NAND2_X1 i_257_76_13471 (.A1(n_257_76_18082), .A2(n_257_76_13447), .ZN(
      n_257_76_13448));
   NAND3_X1 i_257_76_13472 (.A1(n_257_76_13407), .A2(n_257_76_13429), .A3(
      n_257_76_13448), .ZN(n_257_76_13449));
   INV_X1 i_257_76_13473 (.A(n_257_76_13449), .ZN(n_257_76_13450));
   NAND3_X1 i_257_76_13474 (.A1(n_257_76_13042), .A2(n_257_76_13065), .A3(
      n_257_76_13111), .ZN(n_257_76_13451));
   NOR2_X1 i_257_76_13475 (.A1(n_257_76_13132), .A2(n_257_76_13451), .ZN(
      n_257_76_13452));
   NAND2_X1 i_257_76_13476 (.A1(n_257_427), .A2(n_257_76_13123), .ZN(
      n_257_76_13453));
   INV_X1 i_257_76_13477 (.A(n_257_76_13453), .ZN(n_257_76_13454));
   NAND4_X1 i_257_76_13478 (.A1(n_257_76_13454), .A2(n_257_76_13043), .A3(
      n_257_215), .A4(n_257_76_18002), .ZN(n_257_76_13455));
   INV_X1 i_257_76_13479 (.A(n_257_76_13455), .ZN(n_257_76_13456));
   NAND4_X1 i_257_76_13480 (.A1(n_257_76_13137), .A2(n_257_76_13456), .A3(
      n_257_76_13071), .A4(n_257_76_13072), .ZN(n_257_76_13457));
   NAND3_X1 i_257_76_13481 (.A1(n_257_76_13076), .A2(n_257_76_13077), .A3(
      n_257_76_13078), .ZN(n_257_76_13458));
   INV_X1 i_257_76_13482 (.A(n_257_76_13458), .ZN(n_257_76_13459));
   NAND4_X1 i_257_76_13483 (.A1(n_257_76_13459), .A2(n_257_76_13067), .A3(
      n_257_76_13068), .A4(n_257_76_13128), .ZN(n_257_76_13460));
   NOR2_X1 i_257_76_13484 (.A1(n_257_76_13457), .A2(n_257_76_13460), .ZN(
      n_257_76_13461));
   NAND4_X1 i_257_76_13485 (.A1(n_257_76_13116), .A2(n_257_76_13452), .A3(
      n_257_76_13461), .A4(n_257_76_13117), .ZN(n_257_76_13462));
   INV_X1 i_257_76_13486 (.A(n_257_76_13462), .ZN(n_257_76_13463));
   NAND3_X1 i_257_76_13487 (.A1(n_257_76_13463), .A2(n_257_76_13185), .A3(
      n_257_76_13052), .ZN(n_257_76_13464));
   INV_X1 i_257_76_13488 (.A(n_257_76_13464), .ZN(n_257_76_13465));
   NAND2_X1 i_257_76_13489 (.A1(n_257_76_18065), .A2(n_257_76_13465), .ZN(
      n_257_76_13466));
   NAND3_X1 i_257_76_13490 (.A1(n_257_76_13042), .A2(n_257_76_13137), .A3(
      n_257_76_13071), .ZN(n_257_76_13467));
   NAND4_X1 i_257_76_13491 (.A1(n_257_76_13072), .A2(n_257_76_13067), .A3(
      n_257_451), .A4(n_257_475), .ZN(n_257_76_13468));
   NOR2_X1 i_257_76_13492 (.A1(n_257_76_13467), .A2(n_257_76_13468), .ZN(
      n_257_76_13469));
   NAND3_X1 i_257_76_13493 (.A1(n_257_76_13083), .A2(n_257_76_13399), .A3(
      n_257_76_13469), .ZN(n_257_76_13470));
   INV_X1 i_257_76_13494 (.A(n_257_76_13470), .ZN(n_257_76_13471));
   NAND3_X1 i_257_76_13495 (.A1(n_257_76_13052), .A2(n_257_76_13471), .A3(
      n_257_76_13041), .ZN(n_257_76_13472));
   INV_X1 i_257_76_13496 (.A(n_257_76_13472), .ZN(n_257_76_13473));
   NAND2_X1 i_257_76_13497 (.A1(n_257_76_18063), .A2(n_257_76_13473), .ZN(
      n_257_76_13474));
   NAND4_X1 i_257_76_13498 (.A1(n_257_76_13063), .A2(n_257_76_13131), .A3(
      n_257_76_13064), .A4(n_257_76_13042), .ZN(n_257_76_13475));
   INV_X1 i_257_76_13499 (.A(n_257_76_13475), .ZN(n_257_76_13476));
   NAND2_X1 i_257_76_13500 (.A1(n_257_76_13126), .A2(n_257_76_13078), .ZN(
      n_257_76_13477));
   INV_X1 i_257_76_13501 (.A(n_257_76_13477), .ZN(n_257_76_13478));
   NAND4_X1 i_257_76_13502 (.A1(n_257_76_13170), .A2(n_257_76_13478), .A3(
      n_257_76_13068), .A4(n_257_76_13128), .ZN(n_257_76_13479));
   NOR2_X1 i_257_76_13503 (.A1(n_257_76_13479), .A2(n_257_76_13113), .ZN(
      n_257_76_13480));
   NAND3_X1 i_257_76_13504 (.A1(n_257_76_18002), .A2(n_257_76_13123), .A3(
      n_257_424), .ZN(n_257_76_13481));
   INV_X1 i_257_76_13505 (.A(n_257_76_13481), .ZN(n_257_76_13482));
   NAND3_X1 i_257_76_13506 (.A1(n_257_76_13482), .A2(n_257_524), .A3(
      n_257_76_13043), .ZN(n_257_76_13483));
   INV_X1 i_257_76_13507 (.A(n_257_76_13483), .ZN(n_257_76_13484));
   NAND4_X1 i_257_76_13508 (.A1(n_257_76_13065), .A2(n_257_76_13111), .A3(
      n_257_76_13484), .A4(n_257_76_13137), .ZN(n_257_76_13485));
   INV_X1 i_257_76_13509 (.A(n_257_76_13485), .ZN(n_257_76_13486));
   NAND4_X1 i_257_76_13510 (.A1(n_257_76_13476), .A2(n_257_76_13480), .A3(
      n_257_76_13486), .A4(n_257_76_13117), .ZN(n_257_76_13487));
   NAND3_X1 i_257_76_13511 (.A1(n_257_76_13119), .A2(n_257_76_13115), .A3(
      n_257_76_13116), .ZN(n_257_76_13488));
   NOR2_X1 i_257_76_13512 (.A1(n_257_76_13487), .A2(n_257_76_13488), .ZN(
      n_257_76_13489));
   NAND3_X1 i_257_76_13513 (.A1(n_257_76_13489), .A2(n_257_76_13185), .A3(
      n_257_76_13052), .ZN(n_257_76_13490));
   INV_X1 i_257_76_13514 (.A(n_257_76_13490), .ZN(n_257_76_13491));
   NAND2_X1 i_257_76_13515 (.A1(n_257_76_18062), .A2(n_257_76_13491), .ZN(
      n_257_76_13492));
   NAND3_X1 i_257_76_13516 (.A1(n_257_76_13466), .A2(n_257_76_13474), .A3(
      n_257_76_13492), .ZN(n_257_76_13493));
   INV_X1 i_257_76_13517 (.A(n_257_76_13493), .ZN(n_257_76_13494));
   NOR2_X1 i_257_76_13518 (.A1(n_257_76_13242), .A2(n_257_76_13088), .ZN(
      n_257_76_13495));
   NAND4_X1 i_257_76_13519 (.A1(n_257_76_13341), .A2(n_257_76_13071), .A3(
      n_257_76_13072), .A4(n_257_76_13067), .ZN(n_257_76_13496));
   NOR2_X1 i_257_76_13520 (.A1(n_257_76_13496), .A2(n_257_76_13479), .ZN(
      n_257_76_13497));
   INV_X1 i_257_76_13521 (.A(n_257_333), .ZN(n_257_76_13498));
   NOR2_X1 i_257_76_13522 (.A1(n_257_76_13498), .A2(n_257_1082), .ZN(
      n_257_76_13499));
   NAND3_X1 i_257_76_13523 (.A1(n_257_76_18002), .A2(n_257_76_13123), .A3(
      n_257_422), .ZN(n_257_76_13500));
   INV_X1 i_257_76_13524 (.A(n_257_76_13500), .ZN(n_257_76_13501));
   NAND3_X1 i_257_76_13525 (.A1(n_257_76_13134), .A2(n_257_76_13499), .A3(
      n_257_76_13501), .ZN(n_257_76_13502));
   INV_X1 i_257_76_13526 (.A(n_257_76_13502), .ZN(n_257_76_13503));
   NAND3_X1 i_257_76_13527 (.A1(n_257_76_13503), .A2(n_257_76_13063), .A3(
      n_257_76_13131), .ZN(n_257_76_13504));
   INV_X1 i_257_76_13528 (.A(n_257_76_13504), .ZN(n_257_76_13505));
   NAND4_X1 i_257_76_13529 (.A1(n_257_76_13495), .A2(n_257_76_13497), .A3(
      n_257_76_13505), .A4(n_257_76_13117), .ZN(n_257_76_13506));
   NOR2_X1 i_257_76_13530 (.A1(n_257_76_13506), .A2(n_257_76_13488), .ZN(
      n_257_76_13507));
   NAND3_X1 i_257_76_13531 (.A1(n_257_76_13507), .A2(n_257_76_13185), .A3(
      n_257_76_13052), .ZN(n_257_76_13508));
   INV_X1 i_257_76_13532 (.A(n_257_76_13508), .ZN(n_257_76_13509));
   NAND2_X1 i_257_76_13533 (.A1(n_257_342), .A2(n_257_76_13509), .ZN(
      n_257_76_13510));
   NAND3_X1 i_257_76_13534 (.A1(n_257_76_13115), .A2(n_257_76_13116), .A3(
      n_257_76_13117), .ZN(n_257_76_13511));
   NAND3_X1 i_257_76_13535 (.A1(n_257_76_13063), .A2(n_257_76_13131), .A3(
      n_257_76_13318), .ZN(n_257_76_13512));
   INV_X1 i_257_76_13536 (.A(n_257_76_13512), .ZN(n_257_76_13513));
   INV_X1 i_257_76_13537 (.A(n_257_76_13226), .ZN(n_257_76_13514));
   NAND3_X1 i_257_76_13538 (.A1(n_257_76_13111), .A2(n_257_76_13137), .A3(
      n_257_76_13341), .ZN(n_257_76_13515));
   INV_X1 i_257_76_13539 (.A(n_257_76_13515), .ZN(n_257_76_13516));
   NAND3_X1 i_257_76_13540 (.A1(n_257_76_13513), .A2(n_257_76_13514), .A3(
      n_257_76_13516), .ZN(n_257_76_13517));
   NOR2_X1 i_257_76_13541 (.A1(n_257_76_13511), .A2(n_257_76_13517), .ZN(
      n_257_76_13518));
   NAND2_X1 i_257_76_13542 (.A1(n_257_420), .A2(n_257_492), .ZN(n_257_76_13519));
   INV_X1 i_257_76_13543 (.A(n_257_76_13519), .ZN(n_257_76_13520));
   NOR2_X1 i_257_76_13544 (.A1(n_257_76_13520), .A2(n_257_1082), .ZN(
      n_257_76_13521));
   NAND2_X1 i_257_76_13545 (.A1(n_257_588), .A2(n_257_428), .ZN(n_257_76_13522));
   NAND3_X1 i_257_76_13546 (.A1(n_257_411), .A2(n_257_484), .A3(n_257_442), 
      .ZN(n_257_76_13523));
   INV_X1 i_257_76_13547 (.A(n_257_76_13523), .ZN(n_257_76_13524));
   NAND3_X1 i_257_76_13548 (.A1(n_257_76_13123), .A2(n_257_76_13522), .A3(
      n_257_76_13524), .ZN(n_257_76_13525));
   INV_X1 i_257_76_13549 (.A(n_257_76_13525), .ZN(n_257_76_13526));
   NAND4_X1 i_257_76_13550 (.A1(n_257_76_13521), .A2(n_257_76_13126), .A3(
      n_257_76_13078), .A4(n_257_76_13526), .ZN(n_257_76_13527));
   INV_X1 i_257_76_13551 (.A(n_257_76_13527), .ZN(n_257_76_13528));
   NAND2_X1 i_257_76_13552 (.A1(n_257_76_13134), .A2(n_257_76_13128), .ZN(
      n_257_76_13529));
   INV_X1 i_257_76_13553 (.A(n_257_76_13529), .ZN(n_257_76_13530));
   NAND3_X1 i_257_76_13554 (.A1(n_257_76_13528), .A2(n_257_76_13530), .A3(
      n_257_76_13437), .ZN(n_257_76_13531));
   NAND4_X1 i_257_76_13555 (.A1(n_257_76_13071), .A2(n_257_76_13072), .A3(
      n_257_76_13067), .A4(n_257_76_13068), .ZN(n_257_76_13532));
   NOR2_X1 i_257_76_13556 (.A1(n_257_76_13531), .A2(n_257_76_13532), .ZN(
      n_257_76_13533));
   NAND3_X1 i_257_76_13557 (.A1(n_257_76_13533), .A2(n_257_76_13083), .A3(
      n_257_76_13119), .ZN(n_257_76_13534));
   INV_X1 i_257_76_13558 (.A(n_257_76_13534), .ZN(n_257_76_13535));
   NAND4_X1 i_257_76_13559 (.A1(n_257_76_13518), .A2(n_257_76_13535), .A3(
      n_257_76_13052), .A4(n_257_76_13041), .ZN(n_257_76_13536));
   INV_X1 i_257_76_13560 (.A(n_257_76_13536), .ZN(n_257_76_13537));
   NAND2_X1 i_257_76_13561 (.A1(n_257_76_18060), .A2(n_257_76_13537), .ZN(
      n_257_76_13538));
   AOI22_X1 i_257_76_13562 (.A1(n_257_438), .A2(n_257_76_16422), .B1(n_257_724), 
      .B2(n_257_76_15655), .ZN(n_257_76_13539));
   NAND2_X1 i_257_76_13563 (.A1(n_257_884), .A2(n_257_76_17903), .ZN(
      n_257_76_13540));
   NAND2_X1 i_257_76_13564 (.A1(n_257_58), .A2(n_257_76_17918), .ZN(
      n_257_76_13541));
   NAND2_X1 i_257_76_13565 (.A1(n_257_440), .A2(n_257_76_13045), .ZN(
      n_257_76_13542));
   NAND4_X1 i_257_76_13566 (.A1(n_257_76_13539), .A2(n_257_76_13540), .A3(
      n_257_76_13541), .A4(n_257_76_13542), .ZN(n_257_76_13543));
   INV_X1 i_257_76_13567 (.A(n_257_76_13091), .ZN(n_257_76_13544));
   NAND2_X1 i_257_76_13568 (.A1(n_257_446), .A2(n_257_76_13544), .ZN(
      n_257_76_13545));
   NAND2_X1 i_257_76_13569 (.A1(n_257_449), .A2(n_257_76_17923), .ZN(
      n_257_76_13546));
   INV_X1 i_257_76_13570 (.A(n_257_76_13365), .ZN(n_257_76_13547));
   NAND2_X1 i_257_76_13571 (.A1(n_257_447), .A2(n_257_76_13547), .ZN(
      n_257_76_13548));
   NAND3_X1 i_257_76_13572 (.A1(n_257_76_13545), .A2(n_257_76_13546), .A3(
      n_257_76_13548), .ZN(n_257_76_13549));
   NOR2_X1 i_257_76_13573 (.A1(n_257_76_13543), .A2(n_257_76_13549), .ZN(
      n_257_76_13550));
   NAND2_X1 i_257_76_13574 (.A1(n_257_922), .A2(n_257_76_17940), .ZN(
      n_257_76_13551));
   NAND2_X1 i_257_76_13575 (.A1(n_257_820), .A2(n_257_76_17952), .ZN(
      n_257_76_13552));
   NAND3_X1 i_257_76_13576 (.A1(n_257_76_13551), .A2(n_257_76_13502), .A3(
      n_257_76_13552), .ZN(n_257_76_13553));
   INV_X1 i_257_76_13577 (.A(n_257_76_13553), .ZN(n_257_76_13554));
   INV_X1 i_257_76_13578 (.A(Small_Packet_Data_Size[23]), .ZN(n_257_76_13555));
   NAND2_X1 i_257_76_13579 (.A1(n_257_76_13522), .A2(n_257_76_18007), .ZN(
      n_257_76_13556));
   INV_X1 i_257_76_13580 (.A(n_257_76_13556), .ZN(n_257_76_13557));
   NAND4_X1 i_257_76_13581 (.A1(n_257_76_13043), .A2(n_257_76_13557), .A3(
      n_257_76_13519), .A4(n_257_76_13123), .ZN(n_257_76_13558));
   NAND2_X1 i_257_76_13582 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[23]), 
      .ZN(n_257_76_13559));
   NAND2_X1 i_257_76_13583 (.A1(n_257_76_13558), .A2(n_257_76_13559), .ZN(
      n_257_76_13560));
   NAND2_X1 i_257_76_13584 (.A1(n_257_652), .A2(n_257_76_17928), .ZN(
      n_257_76_13561));
   NAND4_X1 i_257_76_13585 (.A1(n_257_76_13560), .A2(n_257_76_13561), .A3(
      n_257_76_13483), .A4(n_257_76_13455), .ZN(n_257_76_13562));
   INV_X1 i_257_76_13586 (.A(n_257_76_13562), .ZN(n_257_76_13563));
   NAND3_X1 i_257_76_13587 (.A1(n_257_76_13550), .A2(n_257_76_13554), .A3(
      n_257_76_13563), .ZN(n_257_76_13564));
   INV_X1 i_257_76_13588 (.A(n_257_76_13564), .ZN(n_257_76_13565));
   NAND3_X1 i_257_76_13589 (.A1(n_257_441), .A2(n_257_986), .A3(n_257_442), 
      .ZN(n_257_76_13566));
   NAND2_X1 i_257_76_13590 (.A1(n_257_756), .A2(n_257_76_17935), .ZN(
      n_257_76_13567));
   NAND2_X1 i_257_76_13591 (.A1(n_257_136), .A2(n_257_76_17925), .ZN(
      n_257_76_13568));
   NAND3_X1 i_257_76_13592 (.A1(n_257_76_13566), .A2(n_257_76_13567), .A3(
      n_257_76_13568), .ZN(n_257_76_13569));
   INV_X1 i_257_76_13593 (.A(n_257_76_13569), .ZN(n_257_76_13570));
   NAND2_X1 i_257_76_13594 (.A1(n_257_98), .A2(n_257_76_17932), .ZN(
      n_257_76_13571));
   NAND2_X1 i_257_76_13595 (.A1(n_257_76_13570), .A2(n_257_76_13571), .ZN(
      n_257_76_13572));
   INV_X1 i_257_76_13596 (.A(n_257_76_13572), .ZN(n_257_76_13573));
   NAND2_X1 i_257_76_13597 (.A1(n_257_692), .A2(n_257_76_17958), .ZN(
      n_257_76_13574));
   NAND2_X1 i_257_76_13598 (.A1(n_257_175), .A2(n_257_76_17331), .ZN(
      n_257_76_13575));
   NAND4_X1 i_257_76_13599 (.A1(n_257_76_13565), .A2(n_257_76_13573), .A3(
      n_257_76_13574), .A4(n_257_76_13575), .ZN(n_257_76_13576));
   NAND2_X1 i_257_76_13600 (.A1(n_257_1018), .A2(n_257_76_17964), .ZN(
      n_257_76_13577));
   INV_X1 i_257_76_13601 (.A(n_257_756), .ZN(n_257_76_13578));
   NAND2_X1 i_257_76_13602 (.A1(n_257_76_13578), .A2(n_257_442), .ZN(
      n_257_76_13579));
   INV_X1 i_257_76_13603 (.A(n_257_922), .ZN(n_257_76_13580));
   NAND2_X1 i_257_76_13604 (.A1(n_257_76_13580), .A2(n_257_442), .ZN(
      n_257_76_13581));
   INV_X1 i_257_76_13605 (.A(n_257_820), .ZN(n_257_76_13582));
   NAND2_X1 i_257_76_13606 (.A1(n_257_76_13582), .A2(n_257_442), .ZN(
      n_257_76_13583));
   NOR2_X1 i_257_76_13607 (.A1(n_257_439), .A2(n_257_76_17412), .ZN(
      n_257_76_13584));
   INV_X1 i_257_76_13608 (.A(n_257_884), .ZN(n_257_76_13585));
   AOI21_X1 i_257_76_13609 (.A(n_257_76_13584), .B1(n_257_76_13585), .B2(
      n_257_442), .ZN(n_257_76_13586));
   NAND4_X1 i_257_76_13610 (.A1(n_257_76_13579), .A2(n_257_76_13581), .A3(
      n_257_76_13583), .A4(n_257_76_13586), .ZN(n_257_76_13587));
   INV_X1 i_257_76_13611 (.A(n_257_76_13111), .ZN(n_257_76_13588));
   NAND2_X1 i_257_76_13612 (.A1(n_257_76_13587), .A2(n_257_76_13588), .ZN(
      n_257_76_13589));
   NAND4_X1 i_257_76_13613 (.A1(n_257_76_13577), .A2(n_257_76_13140), .A3(
      n_257_76_13589), .A4(n_257_76_13442), .ZN(n_257_76_13590));
   NOR2_X1 i_257_76_13614 (.A1(n_257_76_13576), .A2(n_257_76_13590), .ZN(
      n_257_76_13591));
   NAND2_X1 i_257_76_13615 (.A1(n_257_1050), .A2(n_257_76_17969), .ZN(
      n_257_76_13592));
   NAND2_X1 i_257_76_13616 (.A1(n_257_76_13217), .A2(n_257_76_13592), .ZN(
      n_257_76_13593));
   INV_X1 i_257_76_13617 (.A(n_257_76_13593), .ZN(n_257_76_13594));
   NAND3_X1 i_257_76_13618 (.A1(n_257_76_13591), .A2(n_257_76_13594), .A3(
      n_257_76_13427), .ZN(n_257_76_13595));
   NAND3_X1 i_257_76_13619 (.A1(n_257_76_13510), .A2(n_257_76_13538), .A3(
      n_257_76_13595), .ZN(n_257_76_13596));
   INV_X1 i_257_76_13620 (.A(n_257_76_13596), .ZN(n_257_76_13597));
   NAND3_X1 i_257_76_13621 (.A1(n_257_76_13450), .A2(n_257_76_13494), .A3(
      n_257_76_13597), .ZN(n_257_76_13598));
   NOR2_X1 i_257_76_13622 (.A1(n_257_76_13391), .A2(n_257_76_13598), .ZN(
      n_257_76_13599));
   NAND2_X1 i_257_76_13623 (.A1(n_257_76_13270), .A2(n_257_76_13599), .ZN(n_23));
   NAND2_X1 i_257_76_13624 (.A1(n_257_1051), .A2(n_257_443), .ZN(n_257_76_13600));
   INV_X1 i_257_76_13625 (.A(n_257_76_13600), .ZN(n_257_76_13601));
   NAND2_X1 i_257_76_13626 (.A1(n_257_1019), .A2(n_257_444), .ZN(n_257_76_13602));
   NAND2_X1 i_257_76_13627 (.A1(n_257_987), .A2(n_257_441), .ZN(n_257_76_13603));
   INV_X1 i_257_76_13628 (.A(n_257_1083), .ZN(n_257_76_13604));
   NAND2_X1 i_257_76_13629 (.A1(n_257_955), .A2(n_257_442), .ZN(n_257_76_13605));
   INV_X1 i_257_76_13630 (.A(n_257_76_13605), .ZN(n_257_76_13606));
   NAND3_X1 i_257_76_13631 (.A1(n_257_440), .A2(n_257_76_13604), .A3(
      n_257_76_13606), .ZN(n_257_76_13607));
   INV_X1 i_257_76_13632 (.A(n_257_76_13607), .ZN(n_257_76_13608));
   NAND2_X1 i_257_76_13633 (.A1(n_257_76_13603), .A2(n_257_76_13608), .ZN(
      n_257_76_13609));
   INV_X1 i_257_76_13634 (.A(n_257_76_13609), .ZN(n_257_76_13610));
   NAND2_X1 i_257_76_13635 (.A1(n_257_76_13602), .A2(n_257_76_13610), .ZN(
      n_257_76_13611));
   NOR2_X1 i_257_76_13636 (.A1(n_257_76_13601), .A2(n_257_76_13611), .ZN(
      n_257_76_13612));
   NAND2_X1 i_257_76_13637 (.A1(n_257_17), .A2(n_257_76_13612), .ZN(
      n_257_76_13613));
   NOR2_X1 i_257_76_13638 (.A1(n_257_1083), .A2(n_257_76_17412), .ZN(
      n_257_76_13614));
   INV_X1 i_257_76_13639 (.A(n_257_76_13614), .ZN(n_257_76_13615));
   NOR2_X1 i_257_76_13640 (.A1(n_257_76_13615), .A2(n_257_76_15197), .ZN(
      n_257_76_13616));
   NAND2_X1 i_257_76_13641 (.A1(n_257_1051), .A2(n_257_76_13616), .ZN(
      n_257_76_13617));
   INV_X1 i_257_76_13642 (.A(n_257_76_13617), .ZN(n_257_76_13618));
   NAND2_X1 i_257_76_13643 (.A1(n_257_76_18072), .A2(n_257_76_13618), .ZN(
      n_257_76_13619));
   NAND2_X1 i_257_76_13644 (.A1(n_257_725), .A2(n_257_435), .ZN(n_257_76_13620));
   NAND2_X1 i_257_76_13645 (.A1(n_257_440), .A2(n_257_955), .ZN(n_257_76_13621));
   NAND2_X1 i_257_76_13646 (.A1(n_257_76_13620), .A2(n_257_76_13621), .ZN(
      n_257_76_13622));
   INV_X1 i_257_76_13647 (.A(n_257_76_13622), .ZN(n_257_76_13623));
   NAND2_X1 i_257_76_13648 (.A1(n_257_438), .A2(n_257_1089), .ZN(n_257_76_13624));
   NOR2_X1 i_257_76_13649 (.A1(n_257_1083), .A2(n_257_76_17927), .ZN(
      n_257_76_13625));
   NAND2_X1 i_257_76_13650 (.A1(n_257_76_13624), .A2(n_257_76_13625), .ZN(
      n_257_76_13626));
   INV_X1 i_257_76_13651 (.A(n_257_76_13626), .ZN(n_257_76_13627));
   NAND3_X1 i_257_76_13652 (.A1(n_257_76_13623), .A2(n_257_76_13627), .A3(
      n_257_653), .ZN(n_257_76_13628));
   NAND2_X1 i_257_76_13653 (.A1(n_257_446), .A2(n_257_853), .ZN(n_257_76_13629));
   NAND2_X1 i_257_76_13654 (.A1(n_257_449), .A2(n_257_661), .ZN(n_257_76_13630));
   NAND2_X1 i_257_76_13655 (.A1(n_257_447), .A2(n_257_789), .ZN(n_257_76_13631));
   NAND3_X1 i_257_76_13656 (.A1(n_257_76_13629), .A2(n_257_76_13630), .A3(
      n_257_76_13631), .ZN(n_257_76_13632));
   NOR2_X1 i_257_76_13657 (.A1(n_257_76_13628), .A2(n_257_76_13632), .ZN(
      n_257_76_13633));
   NAND2_X1 i_257_76_13658 (.A1(n_257_885), .A2(n_257_445), .ZN(n_257_76_13634));
   NAND2_X1 i_257_76_13659 (.A1(n_257_76_13634), .A2(n_257_76_13603), .ZN(
      n_257_76_13635));
   INV_X1 i_257_76_13660 (.A(n_257_76_13635), .ZN(n_257_76_13636));
   NAND2_X1 i_257_76_13661 (.A1(n_257_923), .A2(n_257_439), .ZN(n_257_76_13637));
   NAND3_X1 i_257_76_13662 (.A1(n_257_76_13633), .A2(n_257_76_13636), .A3(
      n_257_76_13637), .ZN(n_257_76_13638));
   NAND2_X1 i_257_76_13663 (.A1(n_257_757), .A2(n_257_436), .ZN(n_257_76_13639));
   NAND2_X1 i_257_76_13664 (.A1(n_257_821), .A2(n_257_437), .ZN(n_257_76_13640));
   NAND2_X1 i_257_76_13665 (.A1(n_257_76_13639), .A2(n_257_76_13640), .ZN(
      n_257_76_13641));
   NOR2_X1 i_257_76_13666 (.A1(n_257_76_13638), .A2(n_257_76_13641), .ZN(
      n_257_76_13642));
   NAND2_X1 i_257_76_13667 (.A1(n_257_693), .A2(n_257_448), .ZN(n_257_76_13643));
   NAND4_X1 i_257_76_13668 (.A1(n_257_76_13642), .A2(n_257_76_13600), .A3(
      n_257_76_13602), .A4(n_257_76_13643), .ZN(n_257_76_13644));
   INV_X1 i_257_76_13669 (.A(n_257_76_13644), .ZN(n_257_76_13645));
   NAND2_X1 i_257_76_13670 (.A1(n_257_28), .A2(n_257_76_13645), .ZN(
      n_257_76_13646));
   NAND3_X1 i_257_76_13671 (.A1(n_257_76_13613), .A2(n_257_76_13619), .A3(
      n_257_76_13646), .ZN(n_257_76_13647));
   NAND2_X1 i_257_76_13672 (.A1(n_257_853), .A2(n_257_442), .ZN(n_257_76_13648));
   NOR2_X1 i_257_76_13673 (.A1(n_257_76_13648), .A2(n_257_1083), .ZN(
      n_257_76_13649));
   NAND4_X1 i_257_76_13674 (.A1(n_257_446), .A2(n_257_76_13649), .A3(
      n_257_76_13621), .A4(n_257_76_13624), .ZN(n_257_76_13650));
   INV_X1 i_257_76_13675 (.A(n_257_76_13650), .ZN(n_257_76_13651));
   NAND3_X1 i_257_76_13676 (.A1(n_257_76_13634), .A2(n_257_76_13651), .A3(
      n_257_76_13603), .ZN(n_257_76_13652));
   INV_X1 i_257_76_13677 (.A(n_257_76_13637), .ZN(n_257_76_13653));
   NOR2_X1 i_257_76_13678 (.A1(n_257_76_13652), .A2(n_257_76_13653), .ZN(
      n_257_76_13654));
   NAND2_X1 i_257_76_13679 (.A1(n_257_76_13602), .A2(n_257_76_13654), .ZN(
      n_257_76_13655));
   NOR2_X1 i_257_76_13680 (.A1(n_257_76_13601), .A2(n_257_76_13655), .ZN(
      n_257_76_13656));
   NAND2_X1 i_257_76_13681 (.A1(n_257_76_18070), .A2(n_257_76_13656), .ZN(
      n_257_76_13657));
   NAND3_X1 i_257_76_13682 (.A1(n_257_76_13621), .A2(n_257_76_13614), .A3(
      n_257_439), .ZN(n_257_76_13658));
   INV_X1 i_257_76_13683 (.A(n_257_76_13658), .ZN(n_257_76_13659));
   NAND3_X1 i_257_76_13684 (.A1(n_257_76_13603), .A2(n_257_923), .A3(
      n_257_76_13659), .ZN(n_257_76_13660));
   INV_X1 i_257_76_13685 (.A(n_257_76_13660), .ZN(n_257_76_13661));
   NAND2_X1 i_257_76_13686 (.A1(n_257_76_13602), .A2(n_257_76_13661), .ZN(
      n_257_76_13662));
   NOR2_X1 i_257_76_13687 (.A1(n_257_76_13601), .A2(n_257_76_13662), .ZN(
      n_257_76_13663));
   NAND2_X1 i_257_76_13688 (.A1(n_257_76_18084), .A2(n_257_76_13663), .ZN(
      n_257_76_13664));
   INV_X1 i_257_76_13689 (.A(n_257_76_17997), .ZN(n_257_76_13665));
   NOR2_X1 i_257_76_13690 (.A1(n_257_76_13665), .A2(n_257_1083), .ZN(
      n_257_76_13666));
   NAND2_X1 i_257_76_13691 (.A1(n_257_216), .A2(n_257_427), .ZN(n_257_76_13667));
   NAND2_X1 i_257_76_13692 (.A1(n_257_432), .A2(n_257_621), .ZN(n_257_76_13668));
   NAND2_X1 i_257_76_13693 (.A1(n_257_76_13668), .A2(n_257_423), .ZN(
      n_257_76_13669));
   INV_X1 i_257_76_13694 (.A(n_257_76_13669), .ZN(n_257_76_13670));
   NAND3_X1 i_257_76_13695 (.A1(n_257_76_13666), .A2(n_257_76_13667), .A3(
      n_257_76_13670), .ZN(n_257_76_13671));
   NAND3_X1 i_257_76_13696 (.A1(n_257_76_13620), .A2(n_257_76_13621), .A3(
      n_257_76_13624), .ZN(n_257_76_13672));
   NOR2_X1 i_257_76_13697 (.A1(n_257_76_13671), .A2(n_257_76_13672), .ZN(
      n_257_76_13673));
   NAND2_X1 i_257_76_13698 (.A1(n_257_525), .A2(n_257_424), .ZN(n_257_76_13674));
   NAND2_X1 i_257_76_13699 (.A1(n_257_59), .A2(n_257_433), .ZN(n_257_76_13675));
   NAND3_X1 i_257_76_13700 (.A1(n_257_76_13674), .A2(n_257_76_13675), .A3(
      n_257_296), .ZN(n_257_76_13676));
   INV_X1 i_257_76_13701 (.A(n_257_76_13676), .ZN(n_257_76_13677));
   NAND2_X1 i_257_76_13702 (.A1(n_257_653), .A2(n_257_450), .ZN(n_257_76_13678));
   NAND2_X1 i_257_76_13703 (.A1(n_257_137), .A2(n_257_430), .ZN(n_257_76_13679));
   NAND4_X1 i_257_76_13704 (.A1(n_257_76_13673), .A2(n_257_76_13677), .A3(
      n_257_76_13678), .A4(n_257_76_13679), .ZN(n_257_76_13680));
   INV_X1 i_257_76_13705 (.A(n_257_76_13680), .ZN(n_257_76_13681));
   NAND2_X1 i_257_76_13706 (.A1(n_257_176), .A2(n_257_429), .ZN(n_257_76_13682));
   NAND3_X1 i_257_76_13707 (.A1(n_257_76_13681), .A2(n_257_76_13682), .A3(
      n_257_76_13639), .ZN(n_257_76_13683));
   INV_X1 i_257_76_13708 (.A(n_257_76_13683), .ZN(n_257_76_13684));
   NAND2_X1 i_257_76_13709 (.A1(n_257_451), .A2(n_257_476), .ZN(n_257_76_13685));
   NAND2_X1 i_257_76_13710 (.A1(n_257_76_13603), .A2(n_257_76_13685), .ZN(
      n_257_76_13686));
   INV_X1 i_257_76_13711 (.A(n_257_76_13686), .ZN(n_257_76_13687));
   NAND2_X1 i_257_76_13712 (.A1(n_257_557), .A2(n_257_426), .ZN(n_257_76_13688));
   INV_X1 i_257_76_13713 (.A(n_257_76_13632), .ZN(n_257_76_13689));
   NAND4_X1 i_257_76_13714 (.A1(n_257_76_13687), .A2(n_257_76_13688), .A3(
      n_257_76_13634), .A4(n_257_76_13689), .ZN(n_257_76_13690));
   NAND2_X1 i_257_76_13715 (.A1(n_257_99), .A2(n_257_431), .ZN(n_257_76_13691));
   NAND3_X1 i_257_76_13716 (.A1(n_257_76_13691), .A2(n_257_76_13640), .A3(
      n_257_76_13637), .ZN(n_257_76_13692));
   NOR2_X1 i_257_76_13717 (.A1(n_257_76_13690), .A2(n_257_76_13692), .ZN(
      n_257_76_13693));
   NAND4_X1 i_257_76_13718 (.A1(n_257_76_13684), .A2(n_257_76_13693), .A3(
      n_257_76_13602), .A4(n_257_76_13643), .ZN(n_257_76_13694));
   NAND2_X1 i_257_76_13719 (.A1(n_257_256), .A2(n_257_425), .ZN(n_257_76_13695));
   NAND2_X1 i_257_76_13720 (.A1(n_257_76_13600), .A2(n_257_76_13695), .ZN(
      n_257_76_13696));
   NOR2_X1 i_257_76_13721 (.A1(n_257_76_13694), .A2(n_257_76_13696), .ZN(
      n_257_76_13697));
   NAND2_X1 i_257_76_13722 (.A1(n_257_76_18066), .A2(n_257_76_13697), .ZN(
      n_257_76_13698));
   NAND3_X1 i_257_76_13723 (.A1(n_257_76_13657), .A2(n_257_76_13664), .A3(
      n_257_76_13698), .ZN(n_257_76_13699));
   NOR2_X1 i_257_76_13724 (.A1(n_257_76_13647), .A2(n_257_76_13699), .ZN(
      n_257_76_13700));
   NAND3_X1 i_257_76_13725 (.A1(n_257_987), .A2(n_257_441), .A3(n_257_76_13614), 
      .ZN(n_257_76_13701));
   INV_X1 i_257_76_13726 (.A(n_257_76_13701), .ZN(n_257_76_13702));
   NAND2_X1 i_257_76_13727 (.A1(n_257_76_13602), .A2(n_257_76_13702), .ZN(
      n_257_76_13703));
   NOR2_X1 i_257_76_13728 (.A1(n_257_76_13601), .A2(n_257_76_13703), .ZN(
      n_257_76_13704));
   NAND2_X1 i_257_76_13729 (.A1(n_257_76_18071), .A2(n_257_76_13704), .ZN(
      n_257_76_13705));
   NAND2_X1 i_257_76_13730 (.A1(n_257_76_13629), .A2(n_257_76_13631), .ZN(
      n_257_76_13706));
   INV_X1 i_257_76_13731 (.A(n_257_76_13706), .ZN(n_257_76_13707));
   NOR2_X1 i_257_76_13732 (.A1(n_257_1083), .A2(n_257_76_15289), .ZN(
      n_257_76_13708));
   NAND4_X1 i_257_76_13733 (.A1(n_257_76_13621), .A2(n_257_76_13624), .A3(
      n_257_76_13708), .A4(n_257_725), .ZN(n_257_76_13709));
   INV_X1 i_257_76_13734 (.A(n_257_76_13709), .ZN(n_257_76_13710));
   NAND4_X1 i_257_76_13735 (.A1(n_257_76_13634), .A2(n_257_76_13707), .A3(
      n_257_76_13710), .A4(n_257_76_13603), .ZN(n_257_76_13711));
   INV_X1 i_257_76_13736 (.A(n_257_76_13711), .ZN(n_257_76_13712));
   NAND2_X1 i_257_76_13737 (.A1(n_257_76_13640), .A2(n_257_76_13637), .ZN(
      n_257_76_13713));
   INV_X1 i_257_76_13738 (.A(n_257_76_13713), .ZN(n_257_76_13714));
   NAND3_X1 i_257_76_13739 (.A1(n_257_76_13712), .A2(n_257_76_13714), .A3(
      n_257_76_13639), .ZN(n_257_76_13715));
   INV_X1 i_257_76_13740 (.A(n_257_76_13715), .ZN(n_257_76_13716));
   NAND3_X1 i_257_76_13741 (.A1(n_257_76_13600), .A2(n_257_76_13602), .A3(
      n_257_76_13716), .ZN(n_257_76_13717));
   INV_X1 i_257_76_13742 (.A(n_257_76_13717), .ZN(n_257_76_13718));
   NAND2_X1 i_257_76_13743 (.A1(n_257_76_18078), .A2(n_257_76_13718), .ZN(
      n_257_76_13719));
   NAND3_X1 i_257_76_13744 (.A1(n_257_589), .A2(n_257_428), .A3(n_257_442), 
      .ZN(n_257_76_13720));
   INV_X1 i_257_76_13745 (.A(n_257_76_13720), .ZN(n_257_76_13721));
   NAND2_X1 i_257_76_13746 (.A1(n_257_76_13721), .A2(n_257_76_13668), .ZN(
      n_257_76_13722));
   NOR2_X1 i_257_76_13747 (.A1(n_257_76_13722), .A2(n_257_1083), .ZN(
      n_257_76_13723));
   NAND2_X1 i_257_76_13748 (.A1(n_257_76_13624), .A2(n_257_76_13723), .ZN(
      n_257_76_13724));
   INV_X1 i_257_76_13749 (.A(n_257_76_13724), .ZN(n_257_76_13725));
   NAND4_X1 i_257_76_13750 (.A1(n_257_76_13725), .A2(n_257_76_13623), .A3(
      n_257_76_13631), .A4(n_257_76_13675), .ZN(n_257_76_13726));
   NAND3_X1 i_257_76_13751 (.A1(n_257_76_13679), .A2(n_257_76_13629), .A3(
      n_257_76_13630), .ZN(n_257_76_13727));
   NOR2_X1 i_257_76_13752 (.A1(n_257_76_13726), .A2(n_257_76_13727), .ZN(
      n_257_76_13728));
   NAND4_X1 i_257_76_13753 (.A1(n_257_76_13634), .A2(n_257_76_13603), .A3(
      n_257_76_13678), .A4(n_257_76_13685), .ZN(n_257_76_13729));
   INV_X1 i_257_76_13754 (.A(n_257_76_13729), .ZN(n_257_76_13730));
   NAND3_X1 i_257_76_13755 (.A1(n_257_76_13728), .A2(n_257_76_13714), .A3(
      n_257_76_13730), .ZN(n_257_76_13731));
   NAND3_X1 i_257_76_13756 (.A1(n_257_76_13682), .A2(n_257_76_13639), .A3(
      n_257_76_13691), .ZN(n_257_76_13732));
   NOR2_X1 i_257_76_13757 (.A1(n_257_76_13731), .A2(n_257_76_13732), .ZN(
      n_257_76_13733));
   NAND2_X1 i_257_76_13758 (.A1(n_257_76_13602), .A2(n_257_76_13643), .ZN(
      n_257_76_13734));
   INV_X1 i_257_76_13759 (.A(n_257_76_13734), .ZN(n_257_76_13735));
   NAND3_X1 i_257_76_13760 (.A1(n_257_76_13733), .A2(n_257_76_13735), .A3(
      n_257_76_13600), .ZN(n_257_76_13736));
   INV_X1 i_257_76_13761 (.A(n_257_76_13736), .ZN(n_257_76_13737));
   NAND2_X1 i_257_76_13762 (.A1(n_257_76_18074), .A2(n_257_76_13737), .ZN(
      n_257_76_13738));
   NAND3_X1 i_257_76_13763 (.A1(n_257_76_13705), .A2(n_257_76_13719), .A3(
      n_257_76_13738), .ZN(n_257_76_13739));
   NAND2_X1 i_257_76_13764 (.A1(n_257_1083), .A2(n_257_442), .ZN(n_257_76_13740));
   INV_X1 i_257_76_13765 (.A(n_257_76_13740), .ZN(n_257_76_13741));
   NAND2_X1 i_257_76_13766 (.A1(n_257_13), .A2(n_257_76_13741), .ZN(
      n_257_76_13742));
   INV_X1 i_257_76_13767 (.A(n_257_885), .ZN(n_257_76_13743));
   NOR2_X1 i_257_76_13768 (.A1(n_257_76_17902), .A2(n_257_1083), .ZN(
      n_257_76_13744));
   NAND3_X1 i_257_76_13769 (.A1(n_257_76_13744), .A2(n_257_76_13621), .A3(
      n_257_76_13624), .ZN(n_257_76_13745));
   NOR2_X1 i_257_76_13770 (.A1(n_257_76_13743), .A2(n_257_76_13745), .ZN(
      n_257_76_13746));
   NAND3_X1 i_257_76_13771 (.A1(n_257_76_13746), .A2(n_257_76_13637), .A3(
      n_257_76_13603), .ZN(n_257_76_13747));
   INV_X1 i_257_76_13772 (.A(n_257_76_13747), .ZN(n_257_76_13748));
   NAND2_X1 i_257_76_13773 (.A1(n_257_76_13602), .A2(n_257_76_13748), .ZN(
      n_257_76_13749));
   NOR2_X1 i_257_76_13774 (.A1(n_257_76_13601), .A2(n_257_76_13749), .ZN(
      n_257_76_13750));
   NAND2_X1 i_257_76_13775 (.A1(n_257_76_18077), .A2(n_257_76_13750), .ZN(
      n_257_76_13751));
   NAND2_X1 i_257_76_13776 (.A1(n_257_76_13742), .A2(n_257_76_13751), .ZN(
      n_257_76_13752));
   NOR2_X1 i_257_76_13777 (.A1(n_257_76_13739), .A2(n_257_76_13752), .ZN(
      n_257_76_13753));
   NAND2_X1 i_257_76_13778 (.A1(n_257_76_13682), .A2(n_257_76_13639), .ZN(
      n_257_76_13754));
   INV_X1 i_257_76_13779 (.A(n_257_76_13754), .ZN(n_257_76_13755));
   NAND3_X1 i_257_76_13780 (.A1(n_257_76_13602), .A2(n_257_76_13643), .A3(
      n_257_76_13755), .ZN(n_257_76_13756));
   INV_X1 i_257_76_13781 (.A(n_257_76_13756), .ZN(n_257_76_13757));
   NAND4_X1 i_257_76_13782 (.A1(n_257_76_13679), .A2(n_257_557), .A3(
      n_257_76_13629), .A4(n_257_76_13630), .ZN(n_257_76_13758));
   NAND2_X1 i_257_76_13783 (.A1(n_257_76_13668), .A2(n_257_426), .ZN(
      n_257_76_13759));
   INV_X1 i_257_76_13784 (.A(n_257_76_13759), .ZN(n_257_76_13760));
   NAND3_X1 i_257_76_13785 (.A1(n_257_76_13666), .A2(n_257_76_13667), .A3(
      n_257_76_13760), .ZN(n_257_76_13761));
   INV_X1 i_257_76_13786 (.A(n_257_76_13761), .ZN(n_257_76_13762));
   INV_X1 i_257_76_13787 (.A(n_257_76_13672), .ZN(n_257_76_13763));
   NAND4_X1 i_257_76_13788 (.A1(n_257_76_13762), .A2(n_257_76_13763), .A3(
      n_257_76_13631), .A4(n_257_76_13675), .ZN(n_257_76_13764));
   NOR2_X1 i_257_76_13789 (.A1(n_257_76_13758), .A2(n_257_76_13764), .ZN(
      n_257_76_13765));
   NAND4_X1 i_257_76_13790 (.A1(n_257_76_13765), .A2(n_257_76_13714), .A3(
      n_257_76_13691), .A4(n_257_76_13730), .ZN(n_257_76_13766));
   INV_X1 i_257_76_13791 (.A(n_257_76_13766), .ZN(n_257_76_13767));
   NAND3_X1 i_257_76_13792 (.A1(n_257_76_13757), .A2(n_257_76_13767), .A3(
      n_257_76_13600), .ZN(n_257_76_13768));
   INV_X1 i_257_76_13793 (.A(n_257_76_13768), .ZN(n_257_76_13769));
   NAND2_X1 i_257_76_13794 (.A1(n_257_76_18076), .A2(n_257_76_13769), .ZN(
      n_257_76_13770));
   NAND3_X1 i_257_76_13795 (.A1(n_257_76_13640), .A2(n_257_76_13637), .A3(
      n_257_757), .ZN(n_257_76_13771));
   NOR2_X1 i_257_76_13796 (.A1(n_257_1083), .A2(n_257_76_17934), .ZN(
      n_257_76_13772));
   NAND3_X1 i_257_76_13797 (.A1(n_257_76_13621), .A2(n_257_76_13624), .A3(
      n_257_76_13772), .ZN(n_257_76_13773));
   INV_X1 i_257_76_13798 (.A(n_257_76_13773), .ZN(n_257_76_13774));
   NAND4_X1 i_257_76_13799 (.A1(n_257_76_13634), .A2(n_257_76_13707), .A3(
      n_257_76_13603), .A4(n_257_76_13774), .ZN(n_257_76_13775));
   NOR2_X1 i_257_76_13800 (.A1(n_257_76_13771), .A2(n_257_76_13775), .ZN(
      n_257_76_13776));
   NAND2_X1 i_257_76_13801 (.A1(n_257_76_13602), .A2(n_257_76_13776), .ZN(
      n_257_76_13777));
   NOR2_X1 i_257_76_13802 (.A1(n_257_76_13777), .A2(n_257_76_13601), .ZN(
      n_257_76_13778));
   NAND2_X1 i_257_76_13803 (.A1(n_257_76_18069), .A2(n_257_76_13778), .ZN(
      n_257_76_13779));
   NAND2_X1 i_257_76_13804 (.A1(n_257_621), .A2(n_257_442), .ZN(n_257_76_13780));
   INV_X1 i_257_76_13805 (.A(n_257_76_13780), .ZN(n_257_76_13781));
   NAND2_X1 i_257_76_13806 (.A1(n_257_76_13781), .A2(n_257_432), .ZN(
      n_257_76_13782));
   NOR2_X1 i_257_76_13807 (.A1(n_257_1083), .A2(n_257_76_13782), .ZN(
      n_257_76_13783));
   NAND2_X1 i_257_76_13808 (.A1(n_257_76_13624), .A2(n_257_76_13783), .ZN(
      n_257_76_13784));
   INV_X1 i_257_76_13809 (.A(n_257_76_13784), .ZN(n_257_76_13785));
   NAND3_X1 i_257_76_13810 (.A1(n_257_76_13623), .A2(n_257_76_13675), .A3(
      n_257_76_13785), .ZN(n_257_76_13786));
   NOR2_X1 i_257_76_13811 (.A1(n_257_76_13786), .A2(n_257_76_13632), .ZN(
      n_257_76_13787));
   NAND4_X1 i_257_76_13812 (.A1(n_257_76_13714), .A2(n_257_76_13730), .A3(
      n_257_76_13787), .A4(n_257_76_13639), .ZN(n_257_76_13788));
   INV_X1 i_257_76_13813 (.A(n_257_76_13788), .ZN(n_257_76_13789));
   NAND4_X1 i_257_76_13814 (.A1(n_257_76_13600), .A2(n_257_76_13789), .A3(
      n_257_76_13602), .A4(n_257_76_13643), .ZN(n_257_76_13790));
   INV_X1 i_257_76_13815 (.A(n_257_76_13790), .ZN(n_257_76_13791));
   NAND2_X1 i_257_76_13816 (.A1(n_257_68), .A2(n_257_76_13791), .ZN(
      n_257_76_13792));
   NAND3_X1 i_257_76_13817 (.A1(n_257_76_13770), .A2(n_257_76_13779), .A3(
      n_257_76_13792), .ZN(n_257_76_13793));
   INV_X1 i_257_76_13818 (.A(n_257_76_13629), .ZN(n_257_76_13794));
   NOR2_X1 i_257_76_13819 (.A1(n_257_1083), .A2(n_257_76_17951), .ZN(
      n_257_76_13795));
   NAND3_X1 i_257_76_13820 (.A1(n_257_76_13621), .A2(n_257_76_13624), .A3(
      n_257_76_13795), .ZN(n_257_76_13796));
   NOR2_X1 i_257_76_13821 (.A1(n_257_76_13794), .A2(n_257_76_13796), .ZN(
      n_257_76_13797));
   NAND3_X1 i_257_76_13822 (.A1(n_257_76_13797), .A2(n_257_821), .A3(
      n_257_76_13603), .ZN(n_257_76_13798));
   NAND2_X1 i_257_76_13823 (.A1(n_257_76_13637), .A2(n_257_76_13634), .ZN(
      n_257_76_13799));
   NOR2_X1 i_257_76_13824 (.A1(n_257_76_13798), .A2(n_257_76_13799), .ZN(
      n_257_76_13800));
   NAND2_X1 i_257_76_13825 (.A1(n_257_76_13602), .A2(n_257_76_13800), .ZN(
      n_257_76_13801));
   NOR2_X1 i_257_76_13826 (.A1(n_257_76_13601), .A2(n_257_76_13801), .ZN(
      n_257_76_13802));
   NAND2_X1 i_257_76_13827 (.A1(n_257_22), .A2(n_257_76_13802), .ZN(
      n_257_76_13803));
   NAND2_X1 i_257_76_13828 (.A1(n_257_444), .A2(n_257_76_13614), .ZN(
      n_257_76_13804));
   INV_X1 i_257_76_13829 (.A(n_257_76_13804), .ZN(n_257_76_13805));
   NAND2_X1 i_257_76_13830 (.A1(n_257_1019), .A2(n_257_76_13805), .ZN(
      n_257_76_13806));
   INV_X1 i_257_76_13831 (.A(n_257_76_13806), .ZN(n_257_76_13807));
   NAND2_X1 i_257_76_13832 (.A1(n_257_76_13600), .A2(n_257_76_13807), .ZN(
      n_257_76_13808));
   INV_X1 i_257_76_13833 (.A(n_257_76_13808), .ZN(n_257_76_13809));
   NAND2_X1 i_257_76_13834 (.A1(n_257_76_18075), .A2(n_257_76_13809), .ZN(
      n_257_76_13810));
   NAND2_X1 i_257_76_13835 (.A1(n_257_76_13803), .A2(n_257_76_13810), .ZN(
      n_257_76_13811));
   NOR2_X1 i_257_76_13836 (.A1(n_257_76_13793), .A2(n_257_76_13811), .ZN(
      n_257_76_13812));
   NAND3_X1 i_257_76_13837 (.A1(n_257_76_13700), .A2(n_257_76_13753), .A3(
      n_257_76_13812), .ZN(n_257_76_13813));
   INV_X1 i_257_76_13838 (.A(n_257_76_13813), .ZN(n_257_76_13814));
   NOR2_X1 i_257_76_13839 (.A1(n_257_1083), .A2(n_257_76_17633), .ZN(
      n_257_76_13815));
   NAND3_X1 i_257_76_13840 (.A1(n_257_76_13624), .A2(n_257_59), .A3(
      n_257_76_13815), .ZN(n_257_76_13816));
   INV_X1 i_257_76_13841 (.A(n_257_76_13816), .ZN(n_257_76_13817));
   NAND2_X1 i_257_76_13842 (.A1(n_257_76_13817), .A2(n_257_76_13623), .ZN(
      n_257_76_13818));
   NOR2_X1 i_257_76_13843 (.A1(n_257_76_13818), .A2(n_257_76_13632), .ZN(
      n_257_76_13819));
   NAND4_X1 i_257_76_13844 (.A1(n_257_76_13714), .A2(n_257_76_13730), .A3(
      n_257_76_13819), .A4(n_257_76_13639), .ZN(n_257_76_13820));
   INV_X1 i_257_76_13845 (.A(n_257_76_13820), .ZN(n_257_76_13821));
   NAND4_X1 i_257_76_13846 (.A1(n_257_76_13600), .A2(n_257_76_13821), .A3(
      n_257_76_13602), .A4(n_257_76_13643), .ZN(n_257_76_13822));
   INV_X1 i_257_76_13847 (.A(n_257_76_13822), .ZN(n_257_76_13823));
   NAND2_X1 i_257_76_13848 (.A1(n_257_76_18081), .A2(n_257_76_13823), .ZN(
      n_257_76_13824));
   NAND2_X1 i_257_76_13849 (.A1(n_257_442), .A2(n_257_661), .ZN(n_257_76_13825));
   NOR2_X1 i_257_76_13850 (.A1(n_257_1083), .A2(n_257_76_13825), .ZN(
      n_257_76_13826));
   NAND3_X1 i_257_76_13851 (.A1(n_257_76_13621), .A2(n_257_76_13624), .A3(
      n_257_76_13826), .ZN(n_257_76_13827));
   INV_X1 i_257_76_13852 (.A(n_257_76_13827), .ZN(n_257_76_13828));
   NAND2_X1 i_257_76_13853 (.A1(n_257_76_13620), .A2(n_257_449), .ZN(
      n_257_76_13829));
   INV_X1 i_257_76_13854 (.A(n_257_76_13829), .ZN(n_257_76_13830));
   NAND4_X1 i_257_76_13855 (.A1(n_257_76_13828), .A2(n_257_76_13830), .A3(
      n_257_76_13629), .A4(n_257_76_13631), .ZN(n_257_76_13831));
   NOR2_X1 i_257_76_13856 (.A1(n_257_76_13635), .A2(n_257_76_13831), .ZN(
      n_257_76_13832));
   NAND3_X1 i_257_76_13857 (.A1(n_257_76_13832), .A2(n_257_76_13714), .A3(
      n_257_76_13639), .ZN(n_257_76_13833));
   INV_X1 i_257_76_13858 (.A(n_257_76_13833), .ZN(n_257_76_13834));
   NAND4_X1 i_257_76_13859 (.A1(n_257_76_13834), .A2(n_257_76_13600), .A3(
      n_257_76_13602), .A4(n_257_76_13643), .ZN(n_257_76_13835));
   INV_X1 i_257_76_13860 (.A(n_257_76_13835), .ZN(n_257_76_13836));
   NAND2_X1 i_257_76_13861 (.A1(n_257_76_18083), .A2(n_257_76_13836), .ZN(
      n_257_76_13837));
   NAND3_X1 i_257_76_13862 (.A1(n_257_76_13630), .A2(n_257_76_13631), .A3(
      n_257_76_13675), .ZN(n_257_76_13838));
   INV_X1 i_257_76_13863 (.A(n_257_621), .ZN(n_257_76_13839));
   NAND2_X1 i_257_76_13864 (.A1(n_257_76_17331), .A2(n_257_76_13839), .ZN(
      n_257_76_13840));
   AOI21_X1 i_257_76_13865 (.A(n_257_1083), .B1(n_257_76_14366), .B2(
      n_257_76_13840), .ZN(n_257_76_13841));
   NAND4_X1 i_257_76_13866 (.A1(n_257_76_13841), .A2(n_257_76_13620), .A3(
      n_257_76_13621), .A4(n_257_76_13624), .ZN(n_257_76_13842));
   NOR2_X1 i_257_76_13867 (.A1(n_257_76_13838), .A2(n_257_76_13842), .ZN(
      n_257_76_13843));
   NAND3_X1 i_257_76_13868 (.A1(n_257_76_13634), .A2(n_257_76_13603), .A3(
      n_257_76_13678), .ZN(n_257_76_13844));
   INV_X1 i_257_76_13869 (.A(n_257_76_13844), .ZN(n_257_76_13845));
   NAND3_X1 i_257_76_13870 (.A1(n_257_76_13685), .A2(n_257_76_13679), .A3(
      n_257_76_13629), .ZN(n_257_76_13846));
   INV_X1 i_257_76_13871 (.A(n_257_76_13846), .ZN(n_257_76_13847));
   NAND4_X1 i_257_76_13872 (.A1(n_257_76_13843), .A2(n_257_76_13845), .A3(
      n_257_76_13637), .A4(n_257_76_13847), .ZN(n_257_76_13848));
   NAND4_X1 i_257_76_13873 (.A1(n_257_76_13639), .A2(n_257_76_13691), .A3(
      n_257_176), .A4(n_257_76_13640), .ZN(n_257_76_13849));
   NOR2_X1 i_257_76_13874 (.A1(n_257_76_13848), .A2(n_257_76_13849), .ZN(
      n_257_76_13850));
   NAND3_X1 i_257_76_13875 (.A1(n_257_76_13850), .A2(n_257_76_13735), .A3(
      n_257_76_13600), .ZN(n_257_76_13851));
   INV_X1 i_257_76_13876 (.A(n_257_76_13851), .ZN(n_257_76_13852));
   NAND2_X1 i_257_76_13877 (.A1(n_257_76_18061), .A2(n_257_76_13852), .ZN(
      n_257_76_13853));
   NAND3_X1 i_257_76_13878 (.A1(n_257_76_13824), .A2(n_257_76_13837), .A3(
      n_257_76_13853), .ZN(n_257_76_13854));
   INV_X1 i_257_76_13879 (.A(n_257_76_13854), .ZN(n_257_76_13855));
   NAND3_X1 i_257_76_13880 (.A1(n_257_76_16992), .A2(n_257_438), .A3(
      n_257_76_13604), .ZN(n_257_76_13856));
   INV_X1 i_257_76_13881 (.A(n_257_76_13621), .ZN(n_257_76_13857));
   NOR2_X1 i_257_76_13882 (.A1(n_257_76_13856), .A2(n_257_76_13857), .ZN(
      n_257_76_13858));
   NAND2_X1 i_257_76_13883 (.A1(n_257_76_13603), .A2(n_257_76_13858), .ZN(
      n_257_76_13859));
   NOR2_X1 i_257_76_13884 (.A1(n_257_76_13653), .A2(n_257_76_13859), .ZN(
      n_257_76_13860));
   NAND2_X1 i_257_76_13885 (.A1(n_257_76_13602), .A2(n_257_76_13860), .ZN(
      n_257_76_13861));
   NOR2_X1 i_257_76_13886 (.A1(n_257_76_13601), .A2(n_257_76_13861), .ZN(
      n_257_76_13862));
   NAND2_X1 i_257_76_13887 (.A1(n_257_76_18067), .A2(n_257_76_13862), .ZN(
      n_257_76_13863));
   NAND2_X1 i_257_76_13888 (.A1(n_257_76_13643), .A2(n_257_76_13755), .ZN(
      n_257_76_13864));
   INV_X1 i_257_76_13889 (.A(n_257_76_13864), .ZN(n_257_76_13865));
   NAND2_X1 i_257_76_13890 (.A1(n_257_76_13674), .A2(n_257_76_13675), .ZN(
      n_257_76_13866));
   NOR2_X1 i_257_76_13891 (.A1(n_257_76_13866), .A2(n_257_76_13622), .ZN(
      n_257_76_13867));
   NAND2_X1 i_257_76_13892 (.A1(n_257_442), .A2(n_257_493), .ZN(n_257_76_13868));
   NAND2_X1 i_257_76_13893 (.A1(n_257_76_13604), .A2(n_257_76_17998), .ZN(
      n_257_76_13869));
   NAND2_X1 i_257_76_13894 (.A1(n_257_76_13668), .A2(n_257_420), .ZN(
      n_257_76_13870));
   NOR2_X1 i_257_76_13895 (.A1(n_257_76_13869), .A2(n_257_76_13870), .ZN(
      n_257_76_13871));
   NAND2_X1 i_257_76_13896 (.A1(n_257_76_13871), .A2(n_257_76_13667), .ZN(
      n_257_76_13872));
   NAND2_X1 i_257_76_13897 (.A1(n_257_334), .A2(n_257_422), .ZN(n_257_76_13873));
   NAND2_X1 i_257_76_13898 (.A1(n_257_76_13624), .A2(n_257_76_13873), .ZN(
      n_257_76_13874));
   NOR2_X1 i_257_76_13899 (.A1(n_257_76_13872), .A2(n_257_76_13874), .ZN(
      n_257_76_13875));
   NAND2_X1 i_257_76_13900 (.A1(n_257_76_13867), .A2(n_257_76_13875), .ZN(
      n_257_76_13876));
   NAND2_X1 i_257_76_13901 (.A1(n_257_296), .A2(n_257_423), .ZN(n_257_76_13877));
   NAND2_X1 i_257_76_13902 (.A1(n_257_76_13877), .A2(n_257_76_13629), .ZN(
      n_257_76_13878));
   INV_X1 i_257_76_13903 (.A(n_257_76_13878), .ZN(n_257_76_13879));
   NAND2_X1 i_257_76_13904 (.A1(n_257_76_13630), .A2(n_257_76_13631), .ZN(
      n_257_76_13880));
   INV_X1 i_257_76_13905 (.A(n_257_76_13880), .ZN(n_257_76_13881));
   NAND2_X1 i_257_76_13906 (.A1(n_257_76_13879), .A2(n_257_76_13881), .ZN(
      n_257_76_13882));
   NOR2_X1 i_257_76_13907 (.A1(n_257_76_13876), .A2(n_257_76_13882), .ZN(
      n_257_76_13883));
   NAND2_X1 i_257_76_13908 (.A1(n_257_76_13603), .A2(n_257_76_13678), .ZN(
      n_257_76_13884));
   NAND2_X1 i_257_76_13909 (.A1(n_257_76_13685), .A2(n_257_76_13679), .ZN(
      n_257_76_13885));
   NOR2_X1 i_257_76_13910 (.A1(n_257_76_13884), .A2(n_257_76_13885), .ZN(
      n_257_76_13886));
   NAND2_X1 i_257_76_13911 (.A1(n_257_76_13883), .A2(n_257_76_13886), .ZN(
      n_257_76_13887));
   NAND2_X1 i_257_76_13912 (.A1(n_257_76_13637), .A2(n_257_76_13688), .ZN(
      n_257_76_13888));
   NAND2_X1 i_257_76_13913 (.A1(n_257_373), .A2(n_257_421), .ZN(n_257_76_13889));
   NAND2_X1 i_257_76_13914 (.A1(n_257_76_13634), .A2(n_257_76_13889), .ZN(
      n_257_76_13890));
   NOR2_X1 i_257_76_13915 (.A1(n_257_76_13888), .A2(n_257_76_13890), .ZN(
      n_257_76_13891));
   NAND2_X1 i_257_76_13916 (.A1(n_257_76_13691), .A2(n_257_76_13640), .ZN(
      n_257_76_13892));
   INV_X1 i_257_76_13917 (.A(n_257_76_13892), .ZN(n_257_76_13893));
   NAND2_X1 i_257_76_13918 (.A1(n_257_76_13891), .A2(n_257_76_13893), .ZN(
      n_257_76_13894));
   NOR2_X1 i_257_76_13919 (.A1(n_257_76_13887), .A2(n_257_76_13894), .ZN(
      n_257_76_13895));
   NAND2_X1 i_257_76_13920 (.A1(n_257_76_13865), .A2(n_257_76_13895), .ZN(
      n_257_76_13896));
   NAND2_X1 i_257_76_13921 (.A1(n_257_76_13695), .A2(n_257_76_13602), .ZN(
      n_257_76_13897));
   INV_X1 i_257_76_13922 (.A(n_257_76_13897), .ZN(n_257_76_13898));
   NAND2_X1 i_257_76_13923 (.A1(n_257_76_13898), .A2(n_257_76_13600), .ZN(
      n_257_76_13899));
   NOR2_X1 i_257_76_13924 (.A1(n_257_76_13896), .A2(n_257_76_13899), .ZN(
      n_257_76_13900));
   NAND2_X1 i_257_76_13925 (.A1(n_257_76_18073), .A2(n_257_76_13900), .ZN(
      n_257_76_13901));
   INV_X1 i_257_76_13926 (.A(n_257_76_13624), .ZN(n_257_76_13902));
   NAND2_X1 i_257_76_13927 (.A1(n_257_76_17999), .A2(n_257_76_13604), .ZN(
      n_257_76_13903));
   NOR2_X1 i_257_76_13928 (.A1(n_257_76_13902), .A2(n_257_76_13903), .ZN(
      n_257_76_13904));
   NAND3_X1 i_257_76_13929 (.A1(n_257_76_13904), .A2(n_257_76_13623), .A3(
      n_257_76_13675), .ZN(n_257_76_13905));
   NAND3_X1 i_257_76_13930 (.A1(n_257_76_13630), .A2(n_257_76_13631), .A3(
      n_257_137), .ZN(n_257_76_13906));
   NOR2_X1 i_257_76_13931 (.A1(n_257_76_13905), .A2(n_257_76_13906), .ZN(
      n_257_76_13907));
   NAND3_X1 i_257_76_13932 (.A1(n_257_76_13678), .A2(n_257_76_13685), .A3(
      n_257_76_13629), .ZN(n_257_76_13908));
   INV_X1 i_257_76_13933 (.A(n_257_76_13908), .ZN(n_257_76_13909));
   NAND3_X1 i_257_76_13934 (.A1(n_257_76_13907), .A2(n_257_76_13636), .A3(
      n_257_76_13909), .ZN(n_257_76_13910));
   NAND4_X1 i_257_76_13935 (.A1(n_257_76_13639), .A2(n_257_76_13691), .A3(
      n_257_76_13640), .A4(n_257_76_13637), .ZN(n_257_76_13911));
   NOR2_X1 i_257_76_13936 (.A1(n_257_76_13910), .A2(n_257_76_13911), .ZN(
      n_257_76_13912));
   NAND3_X1 i_257_76_13937 (.A1(n_257_76_13912), .A2(n_257_76_13735), .A3(
      n_257_76_13600), .ZN(n_257_76_13913));
   INV_X1 i_257_76_13938 (.A(n_257_76_13913), .ZN(n_257_76_13914));
   NAND2_X1 i_257_76_13939 (.A1(n_257_76_18068), .A2(n_257_76_13914), .ZN(
      n_257_76_13915));
   NAND3_X1 i_257_76_13940 (.A1(n_257_76_13863), .A2(n_257_76_13901), .A3(
      n_257_76_13915), .ZN(n_257_76_13916));
   INV_X1 i_257_76_13941 (.A(n_257_76_13916), .ZN(n_257_76_13917));
   NAND2_X1 i_257_76_13942 (.A1(n_257_789), .A2(n_257_442), .ZN(n_257_76_13918));
   NOR2_X1 i_257_76_13943 (.A1(n_257_1083), .A2(n_257_76_13918), .ZN(
      n_257_76_13919));
   NAND4_X1 i_257_76_13944 (.A1(n_257_447), .A2(n_257_76_13621), .A3(
      n_257_76_13624), .A4(n_257_76_13919), .ZN(n_257_76_13920));
   INV_X1 i_257_76_13945 (.A(n_257_76_13920), .ZN(n_257_76_13921));
   NAND4_X1 i_257_76_13946 (.A1(n_257_76_13634), .A2(n_257_76_13921), .A3(
      n_257_76_13603), .A4(n_257_76_13629), .ZN(n_257_76_13922));
   NOR2_X1 i_257_76_13947 (.A1(n_257_76_13922), .A2(n_257_76_13713), .ZN(
      n_257_76_13923));
   NAND2_X1 i_257_76_13948 (.A1(n_257_76_13602), .A2(n_257_76_13923), .ZN(
      n_257_76_13924));
   NOR2_X1 i_257_76_13949 (.A1(n_257_76_13601), .A2(n_257_76_13924), .ZN(
      n_257_76_13925));
   NAND2_X1 i_257_76_13950 (.A1(n_257_76_13604), .A2(n_257_76_18000), .ZN(
      n_257_76_13926));
   NOR2_X1 i_257_76_13951 (.A1(n_257_76_13902), .A2(n_257_76_13926), .ZN(
      n_257_76_13927));
   NAND3_X1 i_257_76_13952 (.A1(n_257_76_13927), .A2(n_257_76_13623), .A3(
      n_257_76_13675), .ZN(n_257_76_13928));
   NOR2_X1 i_257_76_13953 (.A1(n_257_76_13928), .A2(n_257_76_13632), .ZN(
      n_257_76_13929));
   NAND2_X1 i_257_76_13954 (.A1(n_257_99), .A2(n_257_76_13634), .ZN(
      n_257_76_13930));
   INV_X1 i_257_76_13955 (.A(n_257_76_13930), .ZN(n_257_76_13931));
   NAND3_X1 i_257_76_13956 (.A1(n_257_76_13603), .A2(n_257_76_13678), .A3(
      n_257_76_13685), .ZN(n_257_76_13932));
   INV_X1 i_257_76_13957 (.A(n_257_76_13932), .ZN(n_257_76_13933));
   NAND3_X1 i_257_76_13958 (.A1(n_257_76_13929), .A2(n_257_76_13931), .A3(
      n_257_76_13933), .ZN(n_257_76_13934));
   NAND3_X1 i_257_76_13959 (.A1(n_257_76_13639), .A2(n_257_76_13640), .A3(
      n_257_76_13637), .ZN(n_257_76_13935));
   NOR2_X1 i_257_76_13960 (.A1(n_257_76_13934), .A2(n_257_76_13935), .ZN(
      n_257_76_13936));
   NAND4_X1 i_257_76_13961 (.A1(n_257_76_13936), .A2(n_257_76_13600), .A3(
      n_257_76_13602), .A4(n_257_76_13643), .ZN(n_257_76_13937));
   INV_X1 i_257_76_13962 (.A(n_257_76_13937), .ZN(n_257_76_13938));
   AOI22_X1 i_257_76_13963 (.A1(n_257_76_18085), .A2(n_257_76_13925), .B1(
      n_257_76_18080), .B2(n_257_76_13938), .ZN(n_257_76_13939));
   NAND3_X1 i_257_76_13964 (.A1(n_257_76_13855), .A2(n_257_76_13917), .A3(
      n_257_76_13939), .ZN(n_257_76_13940));
   NAND3_X1 i_257_76_13965 (.A1(n_257_76_13629), .A2(n_257_76_13631), .A3(
      n_257_448), .ZN(n_257_76_13941));
   INV_X1 i_257_76_13966 (.A(n_257_76_13941), .ZN(n_257_76_13942));
   NAND3_X1 i_257_76_13967 (.A1(n_257_76_13621), .A2(n_257_76_13624), .A3(
      n_257_76_13604), .ZN(n_257_76_13943));
   OAI21_X1 i_257_76_13968 (.A(n_257_76_17761), .B1(n_257_725), .B2(
      n_257_76_17412), .ZN(n_257_76_13944));
   INV_X1 i_257_76_13969 (.A(n_257_76_13944), .ZN(n_257_76_13945));
   NOR2_X1 i_257_76_13970 (.A1(n_257_76_13943), .A2(n_257_76_13945), .ZN(
      n_257_76_13946));
   NAND4_X1 i_257_76_13971 (.A1(n_257_76_13942), .A2(n_257_76_13946), .A3(
      n_257_76_13634), .A4(n_257_76_13603), .ZN(n_257_76_13947));
   INV_X1 i_257_76_13972 (.A(n_257_76_13947), .ZN(n_257_76_13948));
   NAND4_X1 i_257_76_13973 (.A1(n_257_76_13948), .A2(n_257_693), .A3(
      n_257_76_13639), .A4(n_257_76_13714), .ZN(n_257_76_13949));
   INV_X1 i_257_76_13974 (.A(n_257_76_13949), .ZN(n_257_76_13950));
   NAND3_X1 i_257_76_13975 (.A1(n_257_76_13950), .A2(n_257_76_13600), .A3(
      n_257_76_13602), .ZN(n_257_76_13951));
   INV_X1 i_257_76_13976 (.A(n_257_76_13951), .ZN(n_257_76_13952));
   NAND2_X1 i_257_76_13977 (.A1(n_257_76_18079), .A2(n_257_76_13952), .ZN(
      n_257_76_13953));
   NAND4_X1 i_257_76_13978 (.A1(n_257_76_13604), .A2(n_257_76_17997), .A3(
      n_257_76_13668), .A4(n_257_425), .ZN(n_257_76_13954));
   INV_X1 i_257_76_13979 (.A(n_257_76_13954), .ZN(n_257_76_13955));
   NAND4_X1 i_257_76_13980 (.A1(n_257_76_13955), .A2(n_257_76_13621), .A3(
      n_257_76_13624), .A4(n_257_76_13667), .ZN(n_257_76_13956));
   NAND3_X1 i_257_76_13981 (.A1(n_257_76_13631), .A2(n_257_76_13675), .A3(
      n_257_76_13620), .ZN(n_257_76_13957));
   NOR2_X1 i_257_76_13982 (.A1(n_257_76_13956), .A2(n_257_76_13957), .ZN(
      n_257_76_13958));
   NAND2_X1 i_257_76_13983 (.A1(n_257_76_13678), .A2(n_257_76_13685), .ZN(
      n_257_76_13959));
   INV_X1 i_257_76_13984 (.A(n_257_76_13959), .ZN(n_257_76_13960));
   INV_X1 i_257_76_13985 (.A(n_257_76_13679), .ZN(n_257_76_13961));
   NAND2_X1 i_257_76_13986 (.A1(n_257_76_13629), .A2(n_257_76_13630), .ZN(
      n_257_76_13962));
   NOR2_X1 i_257_76_13987 (.A1(n_257_76_13961), .A2(n_257_76_13962), .ZN(
      n_257_76_13963));
   NAND3_X1 i_257_76_13988 (.A1(n_257_76_13958), .A2(n_257_76_13960), .A3(
      n_257_76_13963), .ZN(n_257_76_13964));
   NAND4_X1 i_257_76_13989 (.A1(n_257_76_13637), .A2(n_257_76_13688), .A3(
      n_257_76_13634), .A4(n_257_76_13603), .ZN(n_257_76_13965));
   NOR2_X1 i_257_76_13990 (.A1(n_257_76_13964), .A2(n_257_76_13965), .ZN(
      n_257_76_13966));
   NAND4_X1 i_257_76_13991 (.A1(n_257_76_13682), .A2(n_257_76_13639), .A3(
      n_257_76_13691), .A4(n_257_76_13640), .ZN(n_257_76_13967));
   INV_X1 i_257_76_13992 (.A(n_257_76_13967), .ZN(n_257_76_13968));
   NAND4_X1 i_257_76_13993 (.A1(n_257_76_13966), .A2(n_257_76_13968), .A3(
      n_257_76_13643), .A4(n_257_256), .ZN(n_257_76_13969));
   NAND2_X1 i_257_76_13994 (.A1(n_257_76_13600), .A2(n_257_76_13602), .ZN(
      n_257_76_13970));
   NOR2_X1 i_257_76_13995 (.A1(n_257_76_13969), .A2(n_257_76_13970), .ZN(
      n_257_76_13971));
   NAND2_X1 i_257_76_13996 (.A1(n_257_76_18064), .A2(n_257_76_13971), .ZN(
      n_257_76_13972));
   NAND4_X1 i_257_76_13997 (.A1(n_257_76_13604), .A2(n_257_76_17997), .A3(
      n_257_76_13668), .A4(n_257_421), .ZN(n_257_76_13973));
   INV_X1 i_257_76_13998 (.A(n_257_76_13973), .ZN(n_257_76_13974));
   NAND4_X1 i_257_76_13999 (.A1(n_257_76_13974), .A2(n_257_76_13624), .A3(
      n_257_76_13873), .A4(n_257_76_13667), .ZN(n_257_76_13975));
   NAND3_X1 i_257_76_14000 (.A1(n_257_76_13675), .A2(n_257_76_13620), .A3(
      n_257_76_13621), .ZN(n_257_76_13976));
   NOR2_X1 i_257_76_14001 (.A1(n_257_76_13975), .A2(n_257_76_13976), .ZN(
      n_257_76_13977));
   NAND2_X1 i_257_76_14002 (.A1(n_257_76_13678), .A2(n_257_76_13679), .ZN(
      n_257_76_13978));
   INV_X1 i_257_76_14003 (.A(n_257_76_13978), .ZN(n_257_76_13979));
   NAND3_X1 i_257_76_14004 (.A1(n_257_76_13877), .A2(n_257_373), .A3(
      n_257_76_13674), .ZN(n_257_76_13980));
   INV_X1 i_257_76_14005 (.A(n_257_76_13980), .ZN(n_257_76_13981));
   NAND3_X1 i_257_76_14006 (.A1(n_257_76_13977), .A2(n_257_76_13979), .A3(
      n_257_76_13981), .ZN(n_257_76_13982));
   INV_X1 i_257_76_14007 (.A(n_257_76_13982), .ZN(n_257_76_13983));
   NAND3_X1 i_257_76_14008 (.A1(n_257_76_13600), .A2(n_257_76_13983), .A3(
      n_257_76_13695), .ZN(n_257_76_13984));
   NAND3_X1 i_257_76_14009 (.A1(n_257_76_13640), .A2(n_257_76_13637), .A3(
      n_257_76_13688), .ZN(n_257_76_13985));
   NAND4_X1 i_257_76_14010 (.A1(n_257_76_13689), .A2(n_257_76_13634), .A3(
      n_257_76_13603), .A4(n_257_76_13685), .ZN(n_257_76_13986));
   NOR2_X1 i_257_76_14011 (.A1(n_257_76_13985), .A2(n_257_76_13986), .ZN(
      n_257_76_13987));
   INV_X1 i_257_76_14012 (.A(n_257_76_13732), .ZN(n_257_76_13988));
   NAND4_X1 i_257_76_14013 (.A1(n_257_76_13987), .A2(n_257_76_13602), .A3(
      n_257_76_13988), .A4(n_257_76_13643), .ZN(n_257_76_13989));
   NOR2_X1 i_257_76_14014 (.A1(n_257_76_13984), .A2(n_257_76_13989), .ZN(
      n_257_76_13990));
   NAND2_X1 i_257_76_14015 (.A1(n_257_76_18082), .A2(n_257_76_13990), .ZN(
      n_257_76_13991));
   NAND3_X1 i_257_76_14016 (.A1(n_257_76_13953), .A2(n_257_76_13972), .A3(
      n_257_76_13991), .ZN(n_257_76_13992));
   INV_X1 i_257_76_14017 (.A(n_257_76_13992), .ZN(n_257_76_13993));
   NAND4_X1 i_257_76_14018 (.A1(n_257_76_13763), .A2(n_257_76_13630), .A3(
      n_257_76_13631), .A4(n_257_76_13675), .ZN(n_257_76_13994));
   NOR2_X1 i_257_76_14019 (.A1(n_257_76_13846), .A2(n_257_76_13994), .ZN(
      n_257_76_13995));
   NAND2_X1 i_257_76_14020 (.A1(n_257_427), .A2(n_257_76_13668), .ZN(
      n_257_76_13996));
   INV_X1 i_257_76_14021 (.A(n_257_76_13996), .ZN(n_257_76_13997));
   NAND3_X1 i_257_76_14022 (.A1(n_257_76_13666), .A2(n_257_76_13997), .A3(
      n_257_216), .ZN(n_257_76_13998));
   INV_X1 i_257_76_14023 (.A(n_257_76_13998), .ZN(n_257_76_13999));
   NAND4_X1 i_257_76_14024 (.A1(n_257_76_13634), .A2(n_257_76_13999), .A3(
      n_257_76_13603), .A4(n_257_76_13678), .ZN(n_257_76_14000));
   INV_X1 i_257_76_14025 (.A(n_257_76_14000), .ZN(n_257_76_14001));
   NAND3_X1 i_257_76_14026 (.A1(n_257_76_13995), .A2(n_257_76_13714), .A3(
      n_257_76_14001), .ZN(n_257_76_14002));
   NOR2_X1 i_257_76_14027 (.A1(n_257_76_14002), .A2(n_257_76_13732), .ZN(
      n_257_76_14003));
   NAND3_X1 i_257_76_14028 (.A1(n_257_76_14003), .A2(n_257_76_13735), .A3(
      n_257_76_13600), .ZN(n_257_76_14004));
   INV_X1 i_257_76_14029 (.A(n_257_76_14004), .ZN(n_257_76_14005));
   NAND2_X1 i_257_76_14030 (.A1(n_257_76_18065), .A2(n_257_76_14005), .ZN(
      n_257_76_14006));
   NAND4_X1 i_257_76_14031 (.A1(n_257_76_13630), .A2(n_257_451), .A3(
      n_257_76_13631), .A4(n_257_476), .ZN(n_257_76_14007));
   NAND2_X1 i_257_76_14032 (.A1(n_257_76_13678), .A2(n_257_76_13629), .ZN(
      n_257_76_14008));
   NOR2_X1 i_257_76_14033 (.A1(n_257_76_14007), .A2(n_257_76_14008), .ZN(
      n_257_76_14009));
   NAND3_X1 i_257_76_14034 (.A1(n_257_76_13946), .A2(n_257_76_13634), .A3(
      n_257_76_13603), .ZN(n_257_76_14010));
   INV_X1 i_257_76_14035 (.A(n_257_76_14010), .ZN(n_257_76_14011));
   NAND4_X1 i_257_76_14036 (.A1(n_257_76_13714), .A2(n_257_76_14009), .A3(
      n_257_76_13639), .A4(n_257_76_14011), .ZN(n_257_76_14012));
   INV_X1 i_257_76_14037 (.A(n_257_76_14012), .ZN(n_257_76_14013));
   NAND4_X1 i_257_76_14038 (.A1(n_257_76_14013), .A2(n_257_76_13600), .A3(
      n_257_76_13602), .A4(n_257_76_13643), .ZN(n_257_76_14014));
   INV_X1 i_257_76_14039 (.A(n_257_76_14014), .ZN(n_257_76_14015));
   NAND2_X1 i_257_76_14040 (.A1(n_257_76_18063), .A2(n_257_76_14015), .ZN(
      n_257_76_14016));
   NAND2_X1 i_257_76_14041 (.A1(n_257_76_13668), .A2(n_257_424), .ZN(
      n_257_76_14017));
   INV_X1 i_257_76_14042 (.A(n_257_76_14017), .ZN(n_257_76_14018));
   NAND3_X1 i_257_76_14043 (.A1(n_257_76_13666), .A2(n_257_76_13667), .A3(
      n_257_76_14018), .ZN(n_257_76_14019));
   NAND3_X1 i_257_76_14044 (.A1(n_257_76_13621), .A2(n_257_76_13624), .A3(
      n_257_525), .ZN(n_257_76_14020));
   NOR2_X1 i_257_76_14045 (.A1(n_257_76_14019), .A2(n_257_76_14020), .ZN(
      n_257_76_14021));
   NAND2_X1 i_257_76_14046 (.A1(n_257_76_13675), .A2(n_257_76_13620), .ZN(
      n_257_76_14022));
   INV_X1 i_257_76_14047 (.A(n_257_76_14022), .ZN(n_257_76_14023));
   NAND4_X1 i_257_76_14048 (.A1(n_257_76_14021), .A2(n_257_76_13678), .A3(
      n_257_76_13679), .A4(n_257_76_14023), .ZN(n_257_76_14024));
   INV_X1 i_257_76_14049 (.A(n_257_76_14024), .ZN(n_257_76_14025));
   NAND3_X1 i_257_76_14050 (.A1(n_257_76_14025), .A2(n_257_76_13682), .A3(
      n_257_76_13639), .ZN(n_257_76_14026));
   INV_X1 i_257_76_14051 (.A(n_257_76_14026), .ZN(n_257_76_14027));
   NAND4_X1 i_257_76_14052 (.A1(n_257_76_14027), .A2(n_257_76_13693), .A3(
      n_257_76_13602), .A4(n_257_76_13643), .ZN(n_257_76_14028));
   NOR2_X1 i_257_76_14053 (.A1(n_257_76_14028), .A2(n_257_76_13696), .ZN(
      n_257_76_14029));
   NAND2_X1 i_257_76_14054 (.A1(n_257_76_18062), .A2(n_257_76_14029), .ZN(
      n_257_76_14030));
   NAND3_X1 i_257_76_14055 (.A1(n_257_76_14006), .A2(n_257_76_14016), .A3(
      n_257_76_14030), .ZN(n_257_76_14031));
   INV_X1 i_257_76_14056 (.A(n_257_76_14031), .ZN(n_257_76_14032));
   NAND3_X1 i_257_76_14057 (.A1(n_257_76_13678), .A2(n_257_76_13685), .A3(
      n_257_76_13679), .ZN(n_257_76_14033));
   INV_X1 i_257_76_14058 (.A(n_257_76_14033), .ZN(n_257_76_14034));
   NAND3_X1 i_257_76_14059 (.A1(n_257_76_13631), .A2(n_257_76_13674), .A3(
      n_257_76_13675), .ZN(n_257_76_14035));
   NAND4_X1 i_257_76_14060 (.A1(n_257_76_13620), .A2(n_257_76_13621), .A3(
      n_257_76_13624), .A4(n_257_76_13667), .ZN(n_257_76_14036));
   NOR2_X1 i_257_76_14061 (.A1(n_257_76_14035), .A2(n_257_76_14036), .ZN(
      n_257_76_14037));
   NAND2_X1 i_257_76_14062 (.A1(n_257_76_13668), .A2(n_257_422), .ZN(
      n_257_76_14038));
   INV_X1 i_257_76_14063 (.A(n_257_76_14038), .ZN(n_257_76_14039));
   NAND4_X1 i_257_76_14064 (.A1(n_257_76_14039), .A2(n_257_334), .A3(
      n_257_76_13604), .A4(n_257_76_17997), .ZN(n_257_76_14040));
   INV_X1 i_257_76_14065 (.A(n_257_76_14040), .ZN(n_257_76_14041));
   NAND4_X1 i_257_76_14066 (.A1(n_257_76_13877), .A2(n_257_76_14041), .A3(
      n_257_76_13629), .A4(n_257_76_13630), .ZN(n_257_76_14042));
   INV_X1 i_257_76_14067 (.A(n_257_76_14042), .ZN(n_257_76_14043));
   NAND3_X1 i_257_76_14068 (.A1(n_257_76_14034), .A2(n_257_76_14037), .A3(
      n_257_76_14043), .ZN(n_257_76_14044));
   NOR2_X1 i_257_76_14069 (.A1(n_257_76_14044), .A2(n_257_76_13965), .ZN(
      n_257_76_14045));
   NAND4_X1 i_257_76_14070 (.A1(n_257_76_14045), .A2(n_257_76_13968), .A3(
      n_257_76_13602), .A4(n_257_76_13643), .ZN(n_257_76_14046));
   NOR2_X1 i_257_76_14071 (.A1(n_257_76_14046), .A2(n_257_76_13696), .ZN(
      n_257_76_14047));
   NAND2_X1 i_257_76_14072 (.A1(n_257_342), .A2(n_257_76_14047), .ZN(
      n_257_76_14048));
   NAND3_X1 i_257_76_14073 (.A1(n_257_76_13637), .A2(n_257_76_13688), .A3(
      n_257_76_13634), .ZN(n_257_76_14049));
   NAND4_X1 i_257_76_14074 (.A1(n_257_76_13889), .A2(n_257_76_13603), .A3(
      n_257_76_13678), .A4(n_257_76_13685), .ZN(n_257_76_14050));
   NOR2_X1 i_257_76_14075 (.A1(n_257_76_14049), .A2(n_257_76_14050), .ZN(
      n_257_76_14051));
   NAND4_X1 i_257_76_14076 (.A1(n_257_76_13968), .A2(n_257_76_13602), .A3(
      n_257_76_13643), .A4(n_257_76_14051), .ZN(n_257_76_14052));
   NAND3_X1 i_257_76_14077 (.A1(n_257_76_13624), .A2(n_257_76_13873), .A3(
      n_257_76_13667), .ZN(n_257_76_14053));
   INV_X1 i_257_76_14078 (.A(n_257_76_13668), .ZN(n_257_76_14054));
   NAND2_X1 i_257_76_14079 (.A1(n_257_412), .A2(n_257_484), .ZN(n_257_76_14055));
   NOR2_X1 i_257_76_14080 (.A1(n_257_76_14054), .A2(n_257_76_14055), .ZN(
      n_257_76_14056));
   NAND2_X1 i_257_76_14081 (.A1(n_257_420), .A2(n_257_493), .ZN(n_257_76_14057));
   NAND4_X1 i_257_76_14082 (.A1(n_257_76_14056), .A2(n_257_76_13604), .A3(
      n_257_76_14057), .A4(n_257_76_17997), .ZN(n_257_76_14058));
   NOR2_X1 i_257_76_14083 (.A1(n_257_76_14053), .A2(n_257_76_14058), .ZN(
      n_257_76_14059));
   NAND2_X1 i_257_76_14084 (.A1(n_257_76_13631), .A2(n_257_76_13674), .ZN(
      n_257_76_14060));
   INV_X1 i_257_76_14085 (.A(n_257_76_14060), .ZN(n_257_76_14061));
   INV_X1 i_257_76_14086 (.A(n_257_76_13976), .ZN(n_257_76_14062));
   NAND3_X1 i_257_76_14087 (.A1(n_257_76_14059), .A2(n_257_76_14061), .A3(
      n_257_76_14062), .ZN(n_257_76_14063));
   NAND4_X1 i_257_76_14088 (.A1(n_257_76_13679), .A2(n_257_76_13877), .A3(
      n_257_76_13629), .A4(n_257_76_13630), .ZN(n_257_76_14064));
   NOR2_X1 i_257_76_14089 (.A1(n_257_76_14063), .A2(n_257_76_14064), .ZN(
      n_257_76_14065));
   NAND3_X1 i_257_76_14090 (.A1(n_257_76_13600), .A2(n_257_76_13695), .A3(
      n_257_76_14065), .ZN(n_257_76_14066));
   NOR2_X1 i_257_76_14091 (.A1(n_257_76_14052), .A2(n_257_76_14066), .ZN(
      n_257_76_14067));
   NAND2_X1 i_257_76_14092 (.A1(n_257_76_18060), .A2(n_257_76_14067), .ZN(
      n_257_76_14068));
   NAND2_X1 i_257_76_14093 (.A1(n_257_59), .A2(n_257_76_17918), .ZN(
      n_257_76_14069));
   NAND2_X1 i_257_76_14094 (.A1(n_257_76_14040), .A2(n_257_76_14069), .ZN(
      n_257_76_14070));
   NAND2_X1 i_257_76_14095 (.A1(n_257_725), .A2(n_257_76_15655), .ZN(
      n_257_76_14071));
   NAND2_X1 i_257_76_14096 (.A1(n_257_76_16992), .A2(n_257_438), .ZN(
      n_257_76_14072));
   NAND2_X1 i_257_76_14097 (.A1(n_257_440), .A2(n_257_76_13606), .ZN(
      n_257_76_14073));
   NAND3_X1 i_257_76_14098 (.A1(n_257_76_14071), .A2(n_257_76_14072), .A3(
      n_257_76_14073), .ZN(n_257_76_14074));
   NOR2_X1 i_257_76_14099 (.A1(n_257_76_14070), .A2(n_257_76_14074), .ZN(
      n_257_76_14075));
   NAND2_X1 i_257_76_14100 (.A1(n_257_76_13668), .A2(n_257_76_14055), .ZN(
      n_257_76_14076));
   INV_X1 i_257_76_14101 (.A(n_257_76_14076), .ZN(n_257_76_14077));
   INV_X1 i_257_76_14102 (.A(Small_Packet_Data_Size[24]), .ZN(n_257_76_14078));
   NAND4_X1 i_257_76_14103 (.A1(n_257_76_14077), .A2(n_257_76_13604), .A3(
      n_257_76_18001), .A4(n_257_76_14057), .ZN(n_257_76_14079));
   NAND2_X1 i_257_76_14104 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[24]), 
      .ZN(n_257_76_14080));
   NAND2_X1 i_257_76_14105 (.A1(n_257_76_14079), .A2(n_257_76_14080), .ZN(
      n_257_76_14081));
   NAND2_X1 i_257_76_14106 (.A1(n_257_76_13998), .A2(n_257_76_14081), .ZN(
      n_257_76_14082));
   INV_X1 i_257_76_14107 (.A(n_257_76_14082), .ZN(n_257_76_14083));
   INV_X1 i_257_76_14108 (.A(n_257_76_13648), .ZN(n_257_76_14084));
   NAND2_X1 i_257_76_14109 (.A1(n_257_446), .A2(n_257_76_14084), .ZN(
      n_257_76_14085));
   INV_X1 i_257_76_14110 (.A(n_257_76_13825), .ZN(n_257_76_14086));
   NAND2_X1 i_257_76_14111 (.A1(n_257_449), .A2(n_257_76_14086), .ZN(
      n_257_76_14087));
   INV_X1 i_257_76_14112 (.A(n_257_76_13918), .ZN(n_257_76_14088));
   NAND2_X1 i_257_76_14113 (.A1(n_257_447), .A2(n_257_76_14088), .ZN(
      n_257_76_14089));
   NAND3_X1 i_257_76_14114 (.A1(n_257_76_14085), .A2(n_257_76_14087), .A3(
      n_257_76_14089), .ZN(n_257_76_14090));
   INV_X1 i_257_76_14115 (.A(n_257_76_14090), .ZN(n_257_76_14091));
   NAND3_X1 i_257_76_14116 (.A1(n_257_76_14075), .A2(n_257_76_14083), .A3(
      n_257_76_14091), .ZN(n_257_76_14092));
   NAND3_X1 i_257_76_14117 (.A1(n_257_987), .A2(n_257_441), .A3(n_257_442), 
      .ZN(n_257_76_14093));
   NAND2_X1 i_257_76_14118 (.A1(n_257_885), .A2(n_257_76_17903), .ZN(
      n_257_76_14094));
   NAND2_X1 i_257_76_14119 (.A1(n_257_653), .A2(n_257_76_17928), .ZN(
      n_257_76_14095));
   NAND2_X1 i_257_76_14120 (.A1(n_257_137), .A2(n_257_76_17925), .ZN(
      n_257_76_14096));
   NAND4_X1 i_257_76_14121 (.A1(n_257_76_14093), .A2(n_257_76_14094), .A3(
      n_257_76_14095), .A4(n_257_76_14096), .ZN(n_257_76_14097));
   NOR2_X1 i_257_76_14122 (.A1(n_257_76_14092), .A2(n_257_76_14097), .ZN(
      n_257_76_14098));
   NAND2_X1 i_257_76_14123 (.A1(n_257_99), .A2(n_257_76_17932), .ZN(
      n_257_76_14099));
   NAND2_X1 i_257_76_14124 (.A1(n_257_821), .A2(n_257_76_17952), .ZN(
      n_257_76_14100));
   NAND2_X1 i_257_76_14125 (.A1(n_257_923), .A2(n_257_76_17940), .ZN(
      n_257_76_14101));
   NAND3_X1 i_257_76_14126 (.A1(n_257_451), .A2(n_257_476), .A3(n_257_76_13944), 
      .ZN(n_257_76_14102));
   NAND4_X1 i_257_76_14127 (.A1(n_257_76_14099), .A2(n_257_76_14100), .A3(
      n_257_76_14101), .A4(n_257_76_14102), .ZN(n_257_76_14103));
   INV_X1 i_257_76_14128 (.A(n_257_76_14103), .ZN(n_257_76_14104));
   AOI22_X1 i_257_76_14129 (.A1(n_257_176), .A2(n_257_76_17331), .B1(n_257_757), 
      .B2(n_257_76_17935), .ZN(n_257_76_14105));
   NAND3_X1 i_257_76_14130 (.A1(n_257_76_14098), .A2(n_257_76_14104), .A3(
      n_257_76_14105), .ZN(n_257_76_14106));
   NAND2_X1 i_257_76_14131 (.A1(n_257_693), .A2(n_257_76_17958), .ZN(
      n_257_76_14107));
   NAND2_X1 i_257_76_14132 (.A1(n_257_76_13680), .A2(n_257_76_14024), .ZN(
      n_257_76_14108));
   INV_X1 i_257_76_14133 (.A(n_257_76_14108), .ZN(n_257_76_14109));
   NAND3_X1 i_257_76_14134 (.A1(n_257_76_14107), .A2(n_257_76_14109), .A3(
      n_257_76_13982), .ZN(n_257_76_14110));
   NOR2_X1 i_257_76_14135 (.A1(n_257_76_14106), .A2(n_257_76_14110), .ZN(
      n_257_76_14111));
   NAND2_X1 i_257_76_14136 (.A1(n_257_1051), .A2(n_257_76_17969), .ZN(
      n_257_76_14112));
   NAND2_X1 i_257_76_14137 (.A1(n_257_1019), .A2(n_257_76_17964), .ZN(
      n_257_76_14113));
   NAND3_X1 i_257_76_14138 (.A1(n_257_76_14112), .A2(n_257_76_13766), .A3(
      n_257_76_14113), .ZN(n_257_76_14114));
   INV_X1 i_257_76_14139 (.A(n_257_76_14114), .ZN(n_257_76_14115));
   NAND3_X1 i_257_76_14140 (.A1(n_257_76_14111), .A2(n_257_76_14115), .A3(
      n_257_76_13969), .ZN(n_257_76_14116));
   NAND3_X1 i_257_76_14141 (.A1(n_257_76_14048), .A2(n_257_76_14068), .A3(
      n_257_76_14116), .ZN(n_257_76_14117));
   INV_X1 i_257_76_14142 (.A(n_257_76_14117), .ZN(n_257_76_14118));
   NAND3_X1 i_257_76_14143 (.A1(n_257_76_13993), .A2(n_257_76_14032), .A3(
      n_257_76_14118), .ZN(n_257_76_14119));
   NOR2_X1 i_257_76_14144 (.A1(n_257_76_13940), .A2(n_257_76_14119), .ZN(
      n_257_76_14120));
   NAND2_X1 i_257_76_14145 (.A1(n_257_76_13814), .A2(n_257_76_14120), .ZN(n_24));
   NAND2_X1 i_257_76_14146 (.A1(n_257_1020), .A2(n_257_444), .ZN(n_257_76_14121));
   NAND2_X1 i_257_76_14147 (.A1(n_257_988), .A2(n_257_441), .ZN(n_257_76_14122));
   INV_X1 i_257_76_14148 (.A(n_257_1084), .ZN(n_257_76_14123));
   NAND2_X1 i_257_76_14149 (.A1(n_257_956), .A2(n_257_442), .ZN(n_257_76_14124));
   INV_X1 i_257_76_14150 (.A(n_257_76_14124), .ZN(n_257_76_14125));
   NAND3_X1 i_257_76_14151 (.A1(n_257_440), .A2(n_257_76_14123), .A3(
      n_257_76_14125), .ZN(n_257_76_14126));
   INV_X1 i_257_76_14152 (.A(n_257_76_14126), .ZN(n_257_76_14127));
   NAND2_X1 i_257_76_14153 (.A1(n_257_76_14122), .A2(n_257_76_14127), .ZN(
      n_257_76_14128));
   INV_X1 i_257_76_14154 (.A(n_257_76_14128), .ZN(n_257_76_14129));
   NAND2_X1 i_257_76_14155 (.A1(n_257_76_14121), .A2(n_257_76_14129), .ZN(
      n_257_76_14130));
   INV_X1 i_257_76_14156 (.A(n_257_76_14130), .ZN(n_257_76_14131));
   NAND2_X1 i_257_76_14157 (.A1(n_257_1052), .A2(n_257_443), .ZN(n_257_76_14132));
   NAND2_X1 i_257_76_14158 (.A1(n_257_76_14131), .A2(n_257_76_14132), .ZN(
      n_257_76_14133));
   INV_X1 i_257_76_14159 (.A(n_257_76_14133), .ZN(n_257_76_14134));
   NAND2_X1 i_257_76_14160 (.A1(n_257_17), .A2(n_257_76_14134), .ZN(
      n_257_76_14135));
   NOR2_X1 i_257_76_14161 (.A1(n_257_1084), .A2(n_257_76_17412), .ZN(
      n_257_76_14136));
   INV_X1 i_257_76_14162 (.A(n_257_76_14136), .ZN(n_257_76_14137));
   NOR2_X1 i_257_76_14163 (.A1(n_257_76_14137), .A2(n_257_76_15197), .ZN(
      n_257_76_14138));
   NAND2_X1 i_257_76_14164 (.A1(n_257_1052), .A2(n_257_76_14138), .ZN(
      n_257_76_14139));
   INV_X1 i_257_76_14165 (.A(n_257_76_14139), .ZN(n_257_76_14140));
   NAND2_X1 i_257_76_14166 (.A1(n_257_76_18072), .A2(n_257_76_14140), .ZN(
      n_257_76_14141));
   NAND2_X1 i_257_76_14167 (.A1(n_257_447), .A2(n_257_790), .ZN(n_257_76_14142));
   NAND2_X1 i_257_76_14168 (.A1(n_257_76_14142), .A2(n_257_654), .ZN(
      n_257_76_14143));
   NAND2_X1 i_257_76_14169 (.A1(n_257_726), .A2(n_257_435), .ZN(n_257_76_14144));
   NOR2_X1 i_257_76_14170 (.A1(n_257_1084), .A2(n_257_76_17927), .ZN(
      n_257_76_14145));
   NAND2_X1 i_257_76_14171 (.A1(n_257_440), .A2(n_257_956), .ZN(n_257_76_14146));
   NAND2_X1 i_257_76_14172 (.A1(n_257_438), .A2(n_257_1090), .ZN(n_257_76_14147));
   NAND4_X1 i_257_76_14173 (.A1(n_257_76_14144), .A2(n_257_76_14145), .A3(
      n_257_76_14146), .A4(n_257_76_14147), .ZN(n_257_76_14148));
   NOR2_X1 i_257_76_14174 (.A1(n_257_76_14143), .A2(n_257_76_14148), .ZN(
      n_257_76_14149));
   NAND2_X1 i_257_76_14175 (.A1(n_257_886), .A2(n_257_445), .ZN(n_257_76_14150));
   NAND2_X1 i_257_76_14176 (.A1(n_257_446), .A2(n_257_854), .ZN(n_257_76_14151));
   NAND2_X1 i_257_76_14177 (.A1(n_257_449), .A2(n_257_662), .ZN(n_257_76_14152));
   NAND2_X1 i_257_76_14178 (.A1(n_257_76_14151), .A2(n_257_76_14152), .ZN(
      n_257_76_14153));
   INV_X1 i_257_76_14179 (.A(n_257_76_14153), .ZN(n_257_76_14154));
   NAND4_X1 i_257_76_14180 (.A1(n_257_76_14149), .A2(n_257_76_14150), .A3(
      n_257_76_14122), .A4(n_257_76_14154), .ZN(n_257_76_14155));
   NAND2_X1 i_257_76_14181 (.A1(n_257_822), .A2(n_257_437), .ZN(n_257_76_14156));
   NAND2_X1 i_257_76_14182 (.A1(n_257_758), .A2(n_257_436), .ZN(n_257_76_14157));
   NAND2_X1 i_257_76_14183 (.A1(n_257_924), .A2(n_257_439), .ZN(n_257_76_14158));
   NAND3_X1 i_257_76_14184 (.A1(n_257_76_14156), .A2(n_257_76_14157), .A3(
      n_257_76_14158), .ZN(n_257_76_14159));
   NOR2_X1 i_257_76_14185 (.A1(n_257_76_14155), .A2(n_257_76_14159), .ZN(
      n_257_76_14160));
   NAND2_X1 i_257_76_14186 (.A1(n_257_694), .A2(n_257_448), .ZN(n_257_76_14161));
   NAND3_X1 i_257_76_14187 (.A1(n_257_76_14160), .A2(n_257_76_14121), .A3(
      n_257_76_14161), .ZN(n_257_76_14162));
   INV_X1 i_257_76_14188 (.A(n_257_76_14132), .ZN(n_257_76_14163));
   NOR2_X1 i_257_76_14189 (.A1(n_257_76_14162), .A2(n_257_76_14163), .ZN(
      n_257_76_14164));
   NAND2_X1 i_257_76_14190 (.A1(n_257_28), .A2(n_257_76_14164), .ZN(
      n_257_76_14165));
   NAND3_X1 i_257_76_14191 (.A1(n_257_76_14135), .A2(n_257_76_14141), .A3(
      n_257_76_14165), .ZN(n_257_76_14166));
   NAND2_X1 i_257_76_14192 (.A1(n_257_854), .A2(n_257_442), .ZN(n_257_76_14167));
   NOR2_X1 i_257_76_14193 (.A1(n_257_76_14167), .A2(n_257_1084), .ZN(
      n_257_76_14168));
   NAND4_X1 i_257_76_14194 (.A1(n_257_76_14168), .A2(n_257_446), .A3(
      n_257_76_14146), .A4(n_257_76_14147), .ZN(n_257_76_14169));
   INV_X1 i_257_76_14195 (.A(n_257_76_14169), .ZN(n_257_76_14170));
   NAND4_X1 i_257_76_14196 (.A1(n_257_76_14158), .A2(n_257_76_14150), .A3(
      n_257_76_14122), .A4(n_257_76_14170), .ZN(n_257_76_14171));
   INV_X1 i_257_76_14197 (.A(n_257_76_14171), .ZN(n_257_76_14172));
   NAND2_X1 i_257_76_14198 (.A1(n_257_76_14121), .A2(n_257_76_14172), .ZN(
      n_257_76_14173));
   INV_X1 i_257_76_14199 (.A(n_257_76_14173), .ZN(n_257_76_14174));
   NAND2_X1 i_257_76_14200 (.A1(n_257_76_14174), .A2(n_257_76_14132), .ZN(
      n_257_76_14175));
   INV_X1 i_257_76_14201 (.A(n_257_76_14175), .ZN(n_257_76_14176));
   NAND2_X1 i_257_76_14202 (.A1(n_257_76_18070), .A2(n_257_76_14176), .ZN(
      n_257_76_14177));
   NAND3_X1 i_257_76_14203 (.A1(n_257_76_14136), .A2(n_257_76_14146), .A3(
      n_257_439), .ZN(n_257_76_14178));
   INV_X1 i_257_76_14204 (.A(n_257_76_14178), .ZN(n_257_76_14179));
   NAND3_X1 i_257_76_14205 (.A1(n_257_76_14122), .A2(n_257_924), .A3(
      n_257_76_14179), .ZN(n_257_76_14180));
   INV_X1 i_257_76_14206 (.A(n_257_76_14180), .ZN(n_257_76_14181));
   NAND2_X1 i_257_76_14207 (.A1(n_257_76_14121), .A2(n_257_76_14181), .ZN(
      n_257_76_14182));
   INV_X1 i_257_76_14208 (.A(n_257_76_14182), .ZN(n_257_76_14183));
   NAND2_X1 i_257_76_14209 (.A1(n_257_76_14183), .A2(n_257_76_14132), .ZN(
      n_257_76_14184));
   INV_X1 i_257_76_14210 (.A(n_257_76_14184), .ZN(n_257_76_14185));
   NAND2_X1 i_257_76_14211 (.A1(n_257_76_18084), .A2(n_257_76_14185), .ZN(
      n_257_76_14186));
   NAND3_X1 i_257_76_14212 (.A1(n_257_76_14144), .A2(n_257_76_14146), .A3(
      n_257_76_14147), .ZN(n_257_76_14187));
   NAND2_X1 i_257_76_14213 (.A1(n_257_432), .A2(n_257_622), .ZN(n_257_76_14188));
   NAND3_X1 i_257_76_14214 (.A1(n_257_76_17993), .A2(n_257_76_14188), .A3(
      n_257_423), .ZN(n_257_76_14189));
   INV_X1 i_257_76_14215 (.A(n_257_76_14189), .ZN(n_257_76_14190));
   NAND2_X1 i_257_76_14216 (.A1(n_257_217), .A2(n_257_427), .ZN(n_257_76_14191));
   NAND3_X1 i_257_76_14217 (.A1(n_257_76_14190), .A2(n_257_76_14191), .A3(
      n_257_76_14123), .ZN(n_257_76_14192));
   NOR2_X1 i_257_76_14218 (.A1(n_257_76_14187), .A2(n_257_76_14192), .ZN(
      n_257_76_14193));
   NAND2_X1 i_257_76_14219 (.A1(n_257_526), .A2(n_257_424), .ZN(n_257_76_14194));
   NAND2_X1 i_257_76_14220 (.A1(n_257_60), .A2(n_257_433), .ZN(n_257_76_14195));
   NAND3_X1 i_257_76_14221 (.A1(n_257_76_14194), .A2(n_257_76_14195), .A3(
      n_257_297), .ZN(n_257_76_14196));
   INV_X1 i_257_76_14222 (.A(n_257_76_14196), .ZN(n_257_76_14197));
   NAND2_X1 i_257_76_14223 (.A1(n_257_654), .A2(n_257_450), .ZN(n_257_76_14198));
   NAND3_X1 i_257_76_14224 (.A1(n_257_76_14193), .A2(n_257_76_14197), .A3(
      n_257_76_14198), .ZN(n_257_76_14199));
   INV_X1 i_257_76_14225 (.A(n_257_76_14199), .ZN(n_257_76_14200));
   NAND2_X1 i_257_76_14226 (.A1(n_257_177), .A2(n_257_429), .ZN(n_257_76_14201));
   NAND2_X1 i_257_76_14227 (.A1(n_257_100), .A2(n_257_431), .ZN(n_257_76_14202));
   NAND3_X1 i_257_76_14228 (.A1(n_257_76_14200), .A2(n_257_76_14201), .A3(
      n_257_76_14202), .ZN(n_257_76_14203));
   NAND2_X1 i_257_76_14229 (.A1(n_257_76_14156), .A2(n_257_76_14157), .ZN(
      n_257_76_14204));
   INV_X1 i_257_76_14230 (.A(n_257_76_14204), .ZN(n_257_76_14205));
   NAND2_X1 i_257_76_14231 (.A1(n_257_558), .A2(n_257_426), .ZN(n_257_76_14206));
   NAND3_X1 i_257_76_14232 (.A1(n_257_76_14158), .A2(n_257_76_14150), .A3(
      n_257_76_14206), .ZN(n_257_76_14207));
   INV_X1 i_257_76_14233 (.A(n_257_76_14207), .ZN(n_257_76_14208));
   NAND3_X1 i_257_76_14234 (.A1(n_257_76_14151), .A2(n_257_76_14152), .A3(
      n_257_76_14142), .ZN(n_257_76_14209));
   INV_X1 i_257_76_14235 (.A(n_257_76_14209), .ZN(n_257_76_14210));
   NAND2_X1 i_257_76_14236 (.A1(n_257_138), .A2(n_257_430), .ZN(n_257_76_14211));
   NAND2_X1 i_257_76_14237 (.A1(n_257_451), .A2(n_257_477), .ZN(n_257_76_14212));
   NAND4_X1 i_257_76_14238 (.A1(n_257_76_14210), .A2(n_257_76_14211), .A3(
      n_257_76_14122), .A4(n_257_76_14212), .ZN(n_257_76_14213));
   INV_X1 i_257_76_14239 (.A(n_257_76_14213), .ZN(n_257_76_14214));
   NAND3_X1 i_257_76_14240 (.A1(n_257_76_14205), .A2(n_257_76_14208), .A3(
      n_257_76_14214), .ZN(n_257_76_14215));
   NOR2_X1 i_257_76_14241 (.A1(n_257_76_14203), .A2(n_257_76_14215), .ZN(
      n_257_76_14216));
   NAND2_X1 i_257_76_14242 (.A1(n_257_257), .A2(n_257_425), .ZN(n_257_76_14217));
   NAND3_X1 i_257_76_14243 (.A1(n_257_76_14217), .A2(n_257_76_14121), .A3(
      n_257_76_14161), .ZN(n_257_76_14218));
   INV_X1 i_257_76_14244 (.A(n_257_76_14218), .ZN(n_257_76_14219));
   NAND3_X1 i_257_76_14245 (.A1(n_257_76_14216), .A2(n_257_76_14219), .A3(
      n_257_76_14132), .ZN(n_257_76_14220));
   INV_X1 i_257_76_14246 (.A(n_257_76_14220), .ZN(n_257_76_14221));
   NAND2_X1 i_257_76_14247 (.A1(n_257_76_18066), .A2(n_257_76_14221), .ZN(
      n_257_76_14222));
   NAND3_X1 i_257_76_14248 (.A1(n_257_76_14177), .A2(n_257_76_14186), .A3(
      n_257_76_14222), .ZN(n_257_76_14223));
   NOR2_X1 i_257_76_14249 (.A1(n_257_76_14166), .A2(n_257_76_14223), .ZN(
      n_257_76_14224));
   NAND3_X1 i_257_76_14250 (.A1(n_257_988), .A2(n_257_441), .A3(n_257_76_14136), 
      .ZN(n_257_76_14225));
   INV_X1 i_257_76_14251 (.A(n_257_76_14225), .ZN(n_257_76_14226));
   NAND2_X1 i_257_76_14252 (.A1(n_257_76_14121), .A2(n_257_76_14226), .ZN(
      n_257_76_14227));
   INV_X1 i_257_76_14253 (.A(n_257_76_14227), .ZN(n_257_76_14228));
   NAND2_X1 i_257_76_14254 (.A1(n_257_76_14228), .A2(n_257_76_14132), .ZN(
      n_257_76_14229));
   INV_X1 i_257_76_14255 (.A(n_257_76_14229), .ZN(n_257_76_14230));
   NAND2_X1 i_257_76_14256 (.A1(n_257_76_18071), .A2(n_257_76_14230), .ZN(
      n_257_76_14231));
   NAND2_X1 i_257_76_14257 (.A1(n_257_76_14151), .A2(n_257_76_14142), .ZN(
      n_257_76_14232));
   INV_X1 i_257_76_14258 (.A(n_257_76_14232), .ZN(n_257_76_14233));
   NOR2_X1 i_257_76_14259 (.A1(n_257_1084), .A2(n_257_76_15289), .ZN(
      n_257_76_14234));
   NAND4_X1 i_257_76_14260 (.A1(n_257_76_14234), .A2(n_257_76_14146), .A3(
      n_257_76_14147), .A4(n_257_726), .ZN(n_257_76_14235));
   INV_X1 i_257_76_14261 (.A(n_257_76_14235), .ZN(n_257_76_14236));
   NAND4_X1 i_257_76_14262 (.A1(n_257_76_14150), .A2(n_257_76_14122), .A3(
      n_257_76_14233), .A4(n_257_76_14236), .ZN(n_257_76_14237));
   NOR2_X1 i_257_76_14263 (.A1(n_257_76_14159), .A2(n_257_76_14237), .ZN(
      n_257_76_14238));
   NAND2_X1 i_257_76_14264 (.A1(n_257_76_14121), .A2(n_257_76_14238), .ZN(
      n_257_76_14239));
   NOR2_X1 i_257_76_14265 (.A1(n_257_76_14163), .A2(n_257_76_14239), .ZN(
      n_257_76_14240));
   NAND2_X1 i_257_76_14266 (.A1(n_257_76_18078), .A2(n_257_76_14240), .ZN(
      n_257_76_14241));
   NAND3_X1 i_257_76_14267 (.A1(n_257_76_14205), .A2(n_257_76_14201), .A3(
      n_257_76_14202), .ZN(n_257_76_14242));
   NAND3_X1 i_257_76_14268 (.A1(n_257_590), .A2(n_257_428), .A3(n_257_442), 
      .ZN(n_257_76_14243));
   INV_X1 i_257_76_14269 (.A(n_257_76_14243), .ZN(n_257_76_14244));
   NAND2_X1 i_257_76_14270 (.A1(n_257_76_14244), .A2(n_257_76_14188), .ZN(
      n_257_76_14245));
   NOR2_X1 i_257_76_14271 (.A1(n_257_76_14245), .A2(n_257_1084), .ZN(
      n_257_76_14246));
   NAND2_X1 i_257_76_14272 (.A1(n_257_76_14147), .A2(n_257_76_14246), .ZN(
      n_257_76_14247));
   INV_X1 i_257_76_14273 (.A(n_257_76_14247), .ZN(n_257_76_14248));
   NAND2_X1 i_257_76_14274 (.A1(n_257_76_14144), .A2(n_257_76_14146), .ZN(
      n_257_76_14249));
   INV_X1 i_257_76_14275 (.A(n_257_76_14249), .ZN(n_257_76_14250));
   NAND3_X1 i_257_76_14276 (.A1(n_257_76_14248), .A2(n_257_76_14250), .A3(
      n_257_76_14195), .ZN(n_257_76_14251));
   NOR2_X1 i_257_76_14277 (.A1(n_257_76_14251), .A2(n_257_76_14209), .ZN(
      n_257_76_14252));
   NAND2_X1 i_257_76_14278 (.A1(n_257_76_14150), .A2(n_257_76_14211), .ZN(
      n_257_76_14253));
   INV_X1 i_257_76_14279 (.A(n_257_76_14253), .ZN(n_257_76_14254));
   NAND3_X1 i_257_76_14280 (.A1(n_257_76_14122), .A2(n_257_76_14212), .A3(
      n_257_76_14198), .ZN(n_257_76_14255));
   INV_X1 i_257_76_14281 (.A(n_257_76_14255), .ZN(n_257_76_14256));
   NAND4_X1 i_257_76_14282 (.A1(n_257_76_14252), .A2(n_257_76_14254), .A3(
      n_257_76_14158), .A4(n_257_76_14256), .ZN(n_257_76_14257));
   NOR2_X1 i_257_76_14283 (.A1(n_257_76_14242), .A2(n_257_76_14257), .ZN(
      n_257_76_14258));
   NAND2_X1 i_257_76_14284 (.A1(n_257_76_14121), .A2(n_257_76_14161), .ZN(
      n_257_76_14259));
   INV_X1 i_257_76_14285 (.A(n_257_76_14259), .ZN(n_257_76_14260));
   NAND3_X1 i_257_76_14286 (.A1(n_257_76_14258), .A2(n_257_76_14260), .A3(
      n_257_76_14132), .ZN(n_257_76_14261));
   INV_X1 i_257_76_14287 (.A(n_257_76_14261), .ZN(n_257_76_14262));
   NAND2_X1 i_257_76_14288 (.A1(n_257_76_18074), .A2(n_257_76_14262), .ZN(
      n_257_76_14263));
   NAND3_X1 i_257_76_14289 (.A1(n_257_76_14231), .A2(n_257_76_14241), .A3(
      n_257_76_14263), .ZN(n_257_76_14264));
   NAND2_X1 i_257_76_14290 (.A1(n_257_1084), .A2(n_257_442), .ZN(n_257_76_14265));
   INV_X1 i_257_76_14291 (.A(n_257_76_14265), .ZN(n_257_76_14266));
   NAND2_X1 i_257_76_14292 (.A1(n_257_13), .A2(n_257_76_14266), .ZN(
      n_257_76_14267));
   INV_X1 i_257_76_14293 (.A(n_257_76_14158), .ZN(n_257_76_14268));
   NOR2_X1 i_257_76_14294 (.A1(n_257_76_17902), .A2(n_257_1084), .ZN(
      n_257_76_14269));
   NAND3_X1 i_257_76_14295 (.A1(n_257_76_14269), .A2(n_257_76_14146), .A3(
      n_257_76_14147), .ZN(n_257_76_14270));
   INV_X1 i_257_76_14296 (.A(n_257_76_14270), .ZN(n_257_76_14271));
   NAND3_X1 i_257_76_14297 (.A1(n_257_76_14122), .A2(n_257_886), .A3(
      n_257_76_14271), .ZN(n_257_76_14272));
   NOR2_X1 i_257_76_14298 (.A1(n_257_76_14268), .A2(n_257_76_14272), .ZN(
      n_257_76_14273));
   NAND2_X1 i_257_76_14299 (.A1(n_257_76_14121), .A2(n_257_76_14273), .ZN(
      n_257_76_14274));
   INV_X1 i_257_76_14300 (.A(n_257_76_14274), .ZN(n_257_76_14275));
   NAND2_X1 i_257_76_14301 (.A1(n_257_76_14275), .A2(n_257_76_14132), .ZN(
      n_257_76_14276));
   INV_X1 i_257_76_14302 (.A(n_257_76_14276), .ZN(n_257_76_14277));
   NAND2_X1 i_257_76_14303 (.A1(n_257_76_18077), .A2(n_257_76_14277), .ZN(
      n_257_76_14278));
   NAND2_X1 i_257_76_14304 (.A1(n_257_76_14267), .A2(n_257_76_14278), .ZN(
      n_257_76_14279));
   NOR2_X1 i_257_76_14305 (.A1(n_257_76_14264), .A2(n_257_76_14279), .ZN(
      n_257_76_14280));
   NAND4_X1 i_257_76_14306 (.A1(n_257_76_14198), .A2(n_257_76_14151), .A3(
      n_257_76_14152), .A4(n_257_76_14142), .ZN(n_257_76_14281));
   NAND3_X1 i_257_76_14307 (.A1(n_257_76_17993), .A2(n_257_76_14188), .A3(
      n_257_426), .ZN(n_257_76_14282));
   NOR2_X1 i_257_76_14308 (.A1(n_257_76_14282), .A2(n_257_1084), .ZN(
      n_257_76_14283));
   NAND2_X1 i_257_76_14309 (.A1(n_257_76_14147), .A2(n_257_76_14191), .ZN(
      n_257_76_14284));
   INV_X1 i_257_76_14310 (.A(n_257_76_14284), .ZN(n_257_76_14285));
   NAND4_X1 i_257_76_14311 (.A1(n_257_76_14250), .A2(n_257_76_14283), .A3(
      n_257_76_14285), .A4(n_257_76_14195), .ZN(n_257_76_14286));
   NOR2_X1 i_257_76_14312 (.A1(n_257_76_14281), .A2(n_257_76_14286), .ZN(
      n_257_76_14287));
   NAND2_X1 i_257_76_14313 (.A1(n_257_76_14158), .A2(n_257_76_14150), .ZN(
      n_257_76_14288));
   INV_X1 i_257_76_14314 (.A(n_257_76_14288), .ZN(n_257_76_14289));
   NAND4_X1 i_257_76_14315 (.A1(n_257_76_14211), .A2(n_257_76_14122), .A3(
      n_257_76_14212), .A4(n_257_558), .ZN(n_257_76_14290));
   INV_X1 i_257_76_14316 (.A(n_257_76_14290), .ZN(n_257_76_14291));
   NAND4_X1 i_257_76_14317 (.A1(n_257_76_14287), .A2(n_257_76_14205), .A3(
      n_257_76_14289), .A4(n_257_76_14291), .ZN(n_257_76_14292));
   INV_X1 i_257_76_14318 (.A(n_257_76_14292), .ZN(n_257_76_14293));
   NAND2_X1 i_257_76_14319 (.A1(n_257_76_14201), .A2(n_257_76_14202), .ZN(
      n_257_76_14294));
   INV_X1 i_257_76_14320 (.A(n_257_76_14294), .ZN(n_257_76_14295));
   NAND4_X1 i_257_76_14321 (.A1(n_257_76_14260), .A2(n_257_76_14293), .A3(
      n_257_76_14132), .A4(n_257_76_14295), .ZN(n_257_76_14296));
   INV_X1 i_257_76_14322 (.A(n_257_76_14296), .ZN(n_257_76_14297));
   NAND2_X1 i_257_76_14323 (.A1(n_257_76_18076), .A2(n_257_76_14297), .ZN(
      n_257_76_14298));
   NAND3_X1 i_257_76_14324 (.A1(n_257_76_14156), .A2(n_257_76_14158), .A3(
      n_257_76_14150), .ZN(n_257_76_14299));
   NOR2_X1 i_257_76_14325 (.A1(n_257_1084), .A2(n_257_76_17934), .ZN(
      n_257_76_14300));
   NAND3_X1 i_257_76_14326 (.A1(n_257_76_14300), .A2(n_257_76_14146), .A3(
      n_257_76_14147), .ZN(n_257_76_14301));
   INV_X1 i_257_76_14327 (.A(n_257_76_14301), .ZN(n_257_76_14302));
   NAND4_X1 i_257_76_14328 (.A1(n_257_758), .A2(n_257_76_14233), .A3(
      n_257_76_14122), .A4(n_257_76_14302), .ZN(n_257_76_14303));
   NOR2_X1 i_257_76_14329 (.A1(n_257_76_14299), .A2(n_257_76_14303), .ZN(
      n_257_76_14304));
   NAND2_X1 i_257_76_14330 (.A1(n_257_76_14121), .A2(n_257_76_14304), .ZN(
      n_257_76_14305));
   NOR2_X1 i_257_76_14331 (.A1(n_257_76_14163), .A2(n_257_76_14305), .ZN(
      n_257_76_14306));
   NAND2_X1 i_257_76_14332 (.A1(n_257_76_18069), .A2(n_257_76_14306), .ZN(
      n_257_76_14307));
   NAND2_X1 i_257_76_14333 (.A1(n_257_76_14142), .A2(n_257_76_14195), .ZN(
      n_257_76_14308));
   NAND2_X1 i_257_76_14334 (.A1(n_257_622), .A2(n_257_442), .ZN(n_257_76_14309));
   INV_X1 i_257_76_14335 (.A(n_257_76_14309), .ZN(n_257_76_14310));
   NAND2_X1 i_257_76_14336 (.A1(n_257_76_14310), .A2(n_257_432), .ZN(
      n_257_76_14311));
   NOR2_X1 i_257_76_14337 (.A1(n_257_1084), .A2(n_257_76_14311), .ZN(
      n_257_76_14312));
   NAND4_X1 i_257_76_14338 (.A1(n_257_76_14144), .A2(n_257_76_14312), .A3(
      n_257_76_14146), .A4(n_257_76_14147), .ZN(n_257_76_14313));
   NOR2_X1 i_257_76_14339 (.A1(n_257_76_14308), .A2(n_257_76_14313), .ZN(
      n_257_76_14314));
   NAND2_X1 i_257_76_14340 (.A1(n_257_76_14122), .A2(n_257_76_14212), .ZN(
      n_257_76_14315));
   INV_X1 i_257_76_14341 (.A(n_257_76_14315), .ZN(n_257_76_14316));
   NAND3_X1 i_257_76_14342 (.A1(n_257_76_14198), .A2(n_257_76_14151), .A3(
      n_257_76_14152), .ZN(n_257_76_14317));
   INV_X1 i_257_76_14343 (.A(n_257_76_14317), .ZN(n_257_76_14318));
   NAND4_X1 i_257_76_14344 (.A1(n_257_76_14314), .A2(n_257_76_14316), .A3(
      n_257_76_14318), .A4(n_257_76_14150), .ZN(n_257_76_14319));
   NOR2_X1 i_257_76_14345 (.A1(n_257_76_14319), .A2(n_257_76_14159), .ZN(
      n_257_76_14320));
   NAND3_X1 i_257_76_14346 (.A1(n_257_76_14320), .A2(n_257_76_14121), .A3(
      n_257_76_14161), .ZN(n_257_76_14321));
   NOR2_X1 i_257_76_14347 (.A1(n_257_76_14321), .A2(n_257_76_14163), .ZN(
      n_257_76_14322));
   NAND2_X1 i_257_76_14348 (.A1(n_257_68), .A2(n_257_76_14322), .ZN(
      n_257_76_14323));
   NAND3_X1 i_257_76_14349 (.A1(n_257_76_14298), .A2(n_257_76_14307), .A3(
      n_257_76_14323), .ZN(n_257_76_14324));
   INV_X1 i_257_76_14350 (.A(n_257_76_14151), .ZN(n_257_76_14325));
   NOR2_X1 i_257_76_14351 (.A1(n_257_1084), .A2(n_257_76_17951), .ZN(
      n_257_76_14326));
   NAND3_X1 i_257_76_14352 (.A1(n_257_76_14326), .A2(n_257_76_14146), .A3(
      n_257_76_14147), .ZN(n_257_76_14327));
   NOR2_X1 i_257_76_14353 (.A1(n_257_76_14325), .A2(n_257_76_14327), .ZN(
      n_257_76_14328));
   NAND3_X1 i_257_76_14354 (.A1(n_257_76_14328), .A2(n_257_822), .A3(
      n_257_76_14122), .ZN(n_257_76_14329));
   NOR2_X1 i_257_76_14355 (.A1(n_257_76_14329), .A2(n_257_76_14288), .ZN(
      n_257_76_14330));
   NAND2_X1 i_257_76_14356 (.A1(n_257_76_14121), .A2(n_257_76_14330), .ZN(
      n_257_76_14331));
   NOR2_X1 i_257_76_14357 (.A1(n_257_76_14163), .A2(n_257_76_14331), .ZN(
      n_257_76_14332));
   NAND2_X1 i_257_76_14358 (.A1(n_257_22), .A2(n_257_76_14332), .ZN(
      n_257_76_14333));
   NAND2_X1 i_257_76_14359 (.A1(n_257_444), .A2(n_257_76_14136), .ZN(
      n_257_76_14334));
   INV_X1 i_257_76_14360 (.A(n_257_76_14334), .ZN(n_257_76_14335));
   NAND2_X1 i_257_76_14361 (.A1(n_257_1020), .A2(n_257_76_14335), .ZN(
      n_257_76_14336));
   INV_X1 i_257_76_14362 (.A(n_257_76_14336), .ZN(n_257_76_14337));
   NAND2_X1 i_257_76_14363 (.A1(n_257_76_14132), .A2(n_257_76_14337), .ZN(
      n_257_76_14338));
   INV_X1 i_257_76_14364 (.A(n_257_76_14338), .ZN(n_257_76_14339));
   NAND2_X1 i_257_76_14365 (.A1(n_257_76_18075), .A2(n_257_76_14339), .ZN(
      n_257_76_14340));
   NAND2_X1 i_257_76_14366 (.A1(n_257_76_14333), .A2(n_257_76_14340), .ZN(
      n_257_76_14341));
   NOR2_X1 i_257_76_14367 (.A1(n_257_76_14324), .A2(n_257_76_14341), .ZN(
      n_257_76_14342));
   NAND3_X1 i_257_76_14368 (.A1(n_257_76_14224), .A2(n_257_76_14280), .A3(
      n_257_76_14342), .ZN(n_257_76_14343));
   INV_X1 i_257_76_14369 (.A(n_257_76_14343), .ZN(n_257_76_14344));
   NAND2_X1 i_257_76_14370 (.A1(n_257_76_14142), .A2(n_257_76_14144), .ZN(
      n_257_76_14345));
   NOR2_X1 i_257_76_14371 (.A1(n_257_1084), .A2(n_257_76_17633), .ZN(
      n_257_76_14346));
   NAND4_X1 i_257_76_14372 (.A1(n_257_76_14346), .A2(n_257_76_14146), .A3(
      n_257_76_14147), .A4(n_257_60), .ZN(n_257_76_14347));
   NOR2_X1 i_257_76_14373 (.A1(n_257_76_14345), .A2(n_257_76_14347), .ZN(
      n_257_76_14348));
   NAND4_X1 i_257_76_14374 (.A1(n_257_76_14348), .A2(n_257_76_14316), .A3(
      n_257_76_14318), .A4(n_257_76_14150), .ZN(n_257_76_14349));
   NOR2_X1 i_257_76_14375 (.A1(n_257_76_14349), .A2(n_257_76_14159), .ZN(
      n_257_76_14350));
   NAND3_X1 i_257_76_14376 (.A1(n_257_76_14350), .A2(n_257_76_14121), .A3(
      n_257_76_14161), .ZN(n_257_76_14351));
   NOR2_X1 i_257_76_14377 (.A1(n_257_76_14351), .A2(n_257_76_14163), .ZN(
      n_257_76_14352));
   NAND2_X1 i_257_76_14378 (.A1(n_257_76_18081), .A2(n_257_76_14352), .ZN(
      n_257_76_14353));
   NAND2_X1 i_257_76_14379 (.A1(n_257_442), .A2(n_257_662), .ZN(n_257_76_14354));
   NOR2_X1 i_257_76_14380 (.A1(n_257_1084), .A2(n_257_76_14354), .ZN(
      n_257_76_14355));
   NAND3_X1 i_257_76_14381 (.A1(n_257_76_14355), .A2(n_257_76_14146), .A3(
      n_257_76_14147), .ZN(n_257_76_14356));
   NAND2_X1 i_257_76_14382 (.A1(n_257_76_14144), .A2(n_257_449), .ZN(
      n_257_76_14357));
   NOR2_X1 i_257_76_14383 (.A1(n_257_76_14356), .A2(n_257_76_14357), .ZN(
      n_257_76_14358));
   NAND4_X1 i_257_76_14384 (.A1(n_257_76_14150), .A2(n_257_76_14358), .A3(
      n_257_76_14122), .A4(n_257_76_14233), .ZN(n_257_76_14359));
   NOR2_X1 i_257_76_14385 (.A1(n_257_76_14159), .A2(n_257_76_14359), .ZN(
      n_257_76_14360));
   NAND3_X1 i_257_76_14386 (.A1(n_257_76_14360), .A2(n_257_76_14121), .A3(
      n_257_76_14161), .ZN(n_257_76_14361));
   NOR2_X1 i_257_76_14387 (.A1(n_257_76_14361), .A2(n_257_76_14163), .ZN(
      n_257_76_14362));
   NAND2_X1 i_257_76_14388 (.A1(n_257_76_18083), .A2(n_257_76_14362), .ZN(
      n_257_76_14363));
   NAND2_X1 i_257_76_14389 (.A1(n_257_76_14146), .A2(n_257_76_14147), .ZN(
      n_257_76_14364));
   INV_X1 i_257_76_14390 (.A(n_257_76_14364), .ZN(n_257_76_14365));
   NAND2_X1 i_257_76_14391 (.A1(n_257_76_17331), .A2(n_257_76_15481), .ZN(
      n_257_76_14366));
   INV_X1 i_257_76_14392 (.A(n_257_622), .ZN(n_257_76_14367));
   NAND2_X1 i_257_76_14393 (.A1(n_257_76_17331), .A2(n_257_76_14367), .ZN(
      n_257_76_14368));
   AOI21_X1 i_257_76_14394 (.A(n_257_1084), .B1(n_257_76_14366), .B2(
      n_257_76_14368), .ZN(n_257_76_14369));
   NAND4_X1 i_257_76_14395 (.A1(n_257_76_14365), .A2(n_257_76_14369), .A3(
      n_257_76_14195), .A4(n_257_76_14144), .ZN(n_257_76_14370));
   NOR2_X1 i_257_76_14396 (.A1(n_257_76_14370), .A2(n_257_76_14209), .ZN(
      n_257_76_14371));
   NAND4_X1 i_257_76_14397 (.A1(n_257_76_14371), .A2(n_257_76_14254), .A3(
      n_257_76_14158), .A4(n_257_76_14256), .ZN(n_257_76_14372));
   NAND3_X1 i_257_76_14398 (.A1(n_257_76_14205), .A2(n_257_76_14202), .A3(
      n_257_177), .ZN(n_257_76_14373));
   NOR2_X1 i_257_76_14399 (.A1(n_257_76_14372), .A2(n_257_76_14373), .ZN(
      n_257_76_14374));
   NAND3_X1 i_257_76_14400 (.A1(n_257_76_14374), .A2(n_257_76_14260), .A3(
      n_257_76_14132), .ZN(n_257_76_14375));
   INV_X1 i_257_76_14401 (.A(n_257_76_14375), .ZN(n_257_76_14376));
   NAND2_X1 i_257_76_14402 (.A1(n_257_76_18061), .A2(n_257_76_14376), .ZN(
      n_257_76_14377));
   NAND3_X1 i_257_76_14403 (.A1(n_257_76_14353), .A2(n_257_76_14363), .A3(
      n_257_76_14377), .ZN(n_257_76_14378));
   INV_X1 i_257_76_14404 (.A(n_257_76_14378), .ZN(n_257_76_14379));
   INV_X1 i_257_76_14405 (.A(n_257_76_14147), .ZN(n_257_76_14380));
   NAND3_X1 i_257_76_14406 (.A1(n_257_76_14380), .A2(n_257_76_14136), .A3(
      n_257_76_14146), .ZN(n_257_76_14381));
   INV_X1 i_257_76_14407 (.A(n_257_76_14381), .ZN(n_257_76_14382));
   NAND2_X1 i_257_76_14408 (.A1(n_257_76_14122), .A2(n_257_76_14382), .ZN(
      n_257_76_14383));
   NOR2_X1 i_257_76_14409 (.A1(n_257_76_14268), .A2(n_257_76_14383), .ZN(
      n_257_76_14384));
   NAND2_X1 i_257_76_14410 (.A1(n_257_76_14121), .A2(n_257_76_14384), .ZN(
      n_257_76_14385));
   INV_X1 i_257_76_14411 (.A(n_257_76_14385), .ZN(n_257_76_14386));
   NAND2_X1 i_257_76_14412 (.A1(n_257_76_14386), .A2(n_257_76_14132), .ZN(
      n_257_76_14387));
   INV_X1 i_257_76_14413 (.A(n_257_76_14387), .ZN(n_257_76_14388));
   NAND2_X1 i_257_76_14414 (.A1(n_257_76_18067), .A2(n_257_76_14388), .ZN(
      n_257_76_14389));
   NAND2_X1 i_257_76_14415 (.A1(n_257_76_14295), .A2(n_257_76_14161), .ZN(
      n_257_76_14390));
   INV_X1 i_257_76_14416 (.A(n_257_76_14390), .ZN(n_257_76_14391));
   NAND2_X1 i_257_76_14417 (.A1(n_257_76_14206), .A2(n_257_76_14211), .ZN(
      n_257_76_14392));
   NOR2_X1 i_257_76_14418 (.A1(n_257_76_14288), .A2(n_257_76_14392), .ZN(
      n_257_76_14393));
   NAND2_X1 i_257_76_14419 (.A1(n_257_76_14393), .A2(n_257_76_14205), .ZN(
      n_257_76_14394));
   NAND2_X1 i_257_76_14420 (.A1(n_257_297), .A2(n_257_423), .ZN(n_257_76_14395));
   NAND2_X1 i_257_76_14421 (.A1(n_257_76_14198), .A2(n_257_76_14395), .ZN(
      n_257_76_14396));
   INV_X1 i_257_76_14422 (.A(n_257_76_14396), .ZN(n_257_76_14397));
   NAND2_X1 i_257_76_14423 (.A1(n_257_76_14397), .A2(n_257_76_14212), .ZN(
      n_257_76_14398));
   NAND2_X1 i_257_76_14424 (.A1(n_257_374), .A2(n_257_421), .ZN(n_257_76_14399));
   NAND2_X1 i_257_76_14425 (.A1(n_257_76_14399), .A2(n_257_76_14122), .ZN(
      n_257_76_14400));
   NOR2_X1 i_257_76_14426 (.A1(n_257_76_14398), .A2(n_257_76_14400), .ZN(
      n_257_76_14401));
   NAND2_X1 i_257_76_14427 (.A1(n_257_76_14195), .A2(n_257_76_14144), .ZN(
      n_257_76_14402));
   NAND2_X1 i_257_76_14428 (.A1(n_257_335), .A2(n_257_422), .ZN(n_257_76_14403));
   NAND2_X1 i_257_76_14429 (.A1(n_257_76_14403), .A2(n_257_76_14146), .ZN(
      n_257_76_14404));
   NOR2_X1 i_257_76_14430 (.A1(n_257_76_14402), .A2(n_257_76_14404), .ZN(
      n_257_76_14405));
   NAND2_X1 i_257_76_14431 (.A1(n_257_442), .A2(n_257_494), .ZN(n_257_76_14406));
   INV_X1 i_257_76_14432 (.A(n_257_76_17994), .ZN(n_257_76_14407));
   NOR2_X1 i_257_76_14433 (.A1(n_257_76_14407), .A2(n_257_1084), .ZN(
      n_257_76_14408));
   NAND2_X1 i_257_76_14434 (.A1(n_257_76_14188), .A2(n_257_420), .ZN(
      n_257_76_14409));
   INV_X1 i_257_76_14435 (.A(n_257_76_14409), .ZN(n_257_76_14410));
   NAND2_X1 i_257_76_14436 (.A1(n_257_76_14408), .A2(n_257_76_14410), .ZN(
      n_257_76_14411));
   NOR2_X1 i_257_76_14437 (.A1(n_257_76_14411), .A2(n_257_76_14284), .ZN(
      n_257_76_14412));
   NAND2_X1 i_257_76_14438 (.A1(n_257_76_14405), .A2(n_257_76_14412), .ZN(
      n_257_76_14413));
   NAND2_X1 i_257_76_14439 (.A1(n_257_76_14142), .A2(n_257_76_14194), .ZN(
      n_257_76_14414));
   INV_X1 i_257_76_14440 (.A(n_257_76_14414), .ZN(n_257_76_14415));
   NAND2_X1 i_257_76_14441 (.A1(n_257_76_14154), .A2(n_257_76_14415), .ZN(
      n_257_76_14416));
   NOR2_X1 i_257_76_14442 (.A1(n_257_76_14413), .A2(n_257_76_14416), .ZN(
      n_257_76_14417));
   NAND2_X1 i_257_76_14443 (.A1(n_257_76_14401), .A2(n_257_76_14417), .ZN(
      n_257_76_14418));
   NOR2_X1 i_257_76_14444 (.A1(n_257_76_14394), .A2(n_257_76_14418), .ZN(
      n_257_76_14419));
   NAND2_X1 i_257_76_14445 (.A1(n_257_76_14391), .A2(n_257_76_14419), .ZN(
      n_257_76_14420));
   NAND2_X1 i_257_76_14446 (.A1(n_257_76_14217), .A2(n_257_76_14121), .ZN(
      n_257_76_14421));
   INV_X1 i_257_76_14447 (.A(n_257_76_14421), .ZN(n_257_76_14422));
   NAND2_X1 i_257_76_14448 (.A1(n_257_76_14422), .A2(n_257_76_14132), .ZN(
      n_257_76_14423));
   NOR2_X1 i_257_76_14449 (.A1(n_257_76_14420), .A2(n_257_76_14423), .ZN(
      n_257_76_14424));
   NAND2_X1 i_257_76_14450 (.A1(n_257_76_18073), .A2(n_257_76_14424), .ZN(
      n_257_76_14425));
   NAND2_X1 i_257_76_14451 (.A1(n_257_76_14123), .A2(n_257_76_17995), .ZN(
      n_257_76_14426));
   NOR2_X1 i_257_76_14452 (.A1(n_257_76_14426), .A2(n_257_76_14380), .ZN(
      n_257_76_14427));
   NAND4_X1 i_257_76_14453 (.A1(n_257_76_14427), .A2(n_257_76_14250), .A3(
      n_257_76_14142), .A4(n_257_76_14195), .ZN(n_257_76_14428));
   NAND4_X1 i_257_76_14454 (.A1(n_257_76_14198), .A2(n_257_138), .A3(
      n_257_76_14151), .A4(n_257_76_14152), .ZN(n_257_76_14429));
   NOR2_X1 i_257_76_14455 (.A1(n_257_76_14428), .A2(n_257_76_14429), .ZN(
      n_257_76_14430));
   NAND4_X1 i_257_76_14456 (.A1(n_257_76_14158), .A2(n_257_76_14150), .A3(
      n_257_76_14122), .A4(n_257_76_14212), .ZN(n_257_76_14431));
   INV_X1 i_257_76_14457 (.A(n_257_76_14431), .ZN(n_257_76_14432));
   NAND4_X1 i_257_76_14458 (.A1(n_257_76_14430), .A2(n_257_76_14432), .A3(
      n_257_76_14205), .A4(n_257_76_14202), .ZN(n_257_76_14433));
   INV_X1 i_257_76_14459 (.A(n_257_76_14433), .ZN(n_257_76_14434));
   NAND3_X1 i_257_76_14460 (.A1(n_257_76_14434), .A2(n_257_76_14260), .A3(
      n_257_76_14132), .ZN(n_257_76_14435));
   INV_X1 i_257_76_14461 (.A(n_257_76_14435), .ZN(n_257_76_14436));
   NAND2_X1 i_257_76_14462 (.A1(n_257_76_18068), .A2(n_257_76_14436), .ZN(
      n_257_76_14437));
   NAND3_X1 i_257_76_14463 (.A1(n_257_76_14389), .A2(n_257_76_14425), .A3(
      n_257_76_14437), .ZN(n_257_76_14438));
   INV_X1 i_257_76_14464 (.A(n_257_76_14438), .ZN(n_257_76_14439));
   NAND2_X1 i_257_76_14465 (.A1(n_257_790), .A2(n_257_442), .ZN(n_257_76_14440));
   NOR2_X1 i_257_76_14466 (.A1(n_257_1084), .A2(n_257_76_14440), .ZN(
      n_257_76_14441));
   NAND4_X1 i_257_76_14467 (.A1(n_257_447), .A2(n_257_76_14441), .A3(
      n_257_76_14146), .A4(n_257_76_14147), .ZN(n_257_76_14442));
   NOR2_X1 i_257_76_14468 (.A1(n_257_76_14442), .A2(n_257_76_14325), .ZN(
      n_257_76_14443));
   NAND3_X1 i_257_76_14469 (.A1(n_257_76_14443), .A2(n_257_76_14150), .A3(
      n_257_76_14122), .ZN(n_257_76_14444));
   NAND2_X1 i_257_76_14470 (.A1(n_257_76_14156), .A2(n_257_76_14158), .ZN(
      n_257_76_14445));
   NOR2_X1 i_257_76_14471 (.A1(n_257_76_14444), .A2(n_257_76_14445), .ZN(
      n_257_76_14446));
   NAND2_X1 i_257_76_14472 (.A1(n_257_76_14121), .A2(n_257_76_14446), .ZN(
      n_257_76_14447));
   NOR2_X1 i_257_76_14473 (.A1(n_257_76_14163), .A2(n_257_76_14447), .ZN(
      n_257_76_14448));
   NAND2_X1 i_257_76_14474 (.A1(n_257_76_17932), .A2(n_257_76_14367), .ZN(
      n_257_76_14449));
   AOI21_X1 i_257_76_14475 (.A(n_257_1084), .B1(n_257_76_15507), .B2(
      n_257_76_14449), .ZN(n_257_76_14450));
   NAND4_X1 i_257_76_14476 (.A1(n_257_76_14450), .A2(n_257_76_14144), .A3(
      n_257_76_14146), .A4(n_257_76_14147), .ZN(n_257_76_14451));
   INV_X1 i_257_76_14477 (.A(n_257_76_14451), .ZN(n_257_76_14452));
   INV_X1 i_257_76_14478 (.A(n_257_76_14308), .ZN(n_257_76_14453));
   NAND4_X1 i_257_76_14479 (.A1(n_257_76_14452), .A2(n_257_76_14154), .A3(
      n_257_76_14453), .A4(n_257_76_14198), .ZN(n_257_76_14454));
   NAND3_X1 i_257_76_14480 (.A1(n_257_76_14150), .A2(n_257_76_14122), .A3(
      n_257_76_14212), .ZN(n_257_76_14455));
   NOR2_X1 i_257_76_14481 (.A1(n_257_76_14454), .A2(n_257_76_14455), .ZN(
      n_257_76_14456));
   NAND4_X1 i_257_76_14482 (.A1(n_257_100), .A2(n_257_76_14156), .A3(
      n_257_76_14157), .A4(n_257_76_14158), .ZN(n_257_76_14457));
   INV_X1 i_257_76_14483 (.A(n_257_76_14457), .ZN(n_257_76_14458));
   NAND4_X1 i_257_76_14484 (.A1(n_257_76_14456), .A2(n_257_76_14121), .A3(
      n_257_76_14161), .A4(n_257_76_14458), .ZN(n_257_76_14459));
   NOR2_X1 i_257_76_14485 (.A1(n_257_76_14459), .A2(n_257_76_14163), .ZN(
      n_257_76_14460));
   AOI22_X1 i_257_76_14486 (.A1(n_257_76_18085), .A2(n_257_76_14448), .B1(
      n_257_76_18080), .B2(n_257_76_14460), .ZN(n_257_76_14461));
   NAND3_X1 i_257_76_14487 (.A1(n_257_76_14379), .A2(n_257_76_14439), .A3(
      n_257_76_14461), .ZN(n_257_76_14462));
   NAND3_X1 i_257_76_14488 (.A1(n_257_76_14151), .A2(n_257_76_14142), .A3(
      n_257_448), .ZN(n_257_76_14463));
   INV_X1 i_257_76_14489 (.A(n_257_76_14463), .ZN(n_257_76_14464));
   NAND3_X1 i_257_76_14490 (.A1(n_257_76_14146), .A2(n_257_76_14147), .A3(
      n_257_76_14123), .ZN(n_257_76_14465));
   OAI21_X1 i_257_76_14491 (.A(n_257_76_17761), .B1(n_257_726), .B2(
      n_257_76_17412), .ZN(n_257_76_14466));
   INV_X1 i_257_76_14492 (.A(n_257_76_14466), .ZN(n_257_76_14467));
   NOR2_X1 i_257_76_14493 (.A1(n_257_76_14465), .A2(n_257_76_14467), .ZN(
      n_257_76_14468));
   NAND4_X1 i_257_76_14494 (.A1(n_257_76_14150), .A2(n_257_76_14464), .A3(
      n_257_76_14468), .A4(n_257_76_14122), .ZN(n_257_76_14469));
   NOR2_X1 i_257_76_14495 (.A1(n_257_76_14469), .A2(n_257_76_14159), .ZN(
      n_257_76_14470));
   NAND3_X1 i_257_76_14496 (.A1(n_257_76_14470), .A2(n_257_76_14121), .A3(
      n_257_694), .ZN(n_257_76_14471));
   NOR2_X1 i_257_76_14497 (.A1(n_257_76_14471), .A2(n_257_76_14163), .ZN(
      n_257_76_14472));
   NAND2_X1 i_257_76_14498 (.A1(n_257_76_18079), .A2(n_257_76_14472), .ZN(
      n_257_76_14473));
   NAND3_X1 i_257_76_14499 (.A1(n_257_76_17993), .A2(n_257_76_14188), .A3(
      n_257_425), .ZN(n_257_76_14474));
   NOR2_X1 i_257_76_14500 (.A1(n_257_76_14474), .A2(n_257_1084), .ZN(
      n_257_76_14475));
   NAND4_X1 i_257_76_14501 (.A1(n_257_76_14475), .A2(n_257_76_14285), .A3(
      n_257_76_14144), .A4(n_257_76_14146), .ZN(n_257_76_14476));
   NAND3_X1 i_257_76_14502 (.A1(n_257_76_14152), .A2(n_257_76_14142), .A3(
      n_257_76_14195), .ZN(n_257_76_14477));
   NOR2_X1 i_257_76_14503 (.A1(n_257_76_14476), .A2(n_257_76_14477), .ZN(
      n_257_76_14478));
   INV_X1 i_257_76_14504 (.A(n_257_76_14392), .ZN(n_257_76_14479));
   NAND4_X1 i_257_76_14505 (.A1(n_257_76_14122), .A2(n_257_76_14212), .A3(
      n_257_76_14198), .A4(n_257_76_14151), .ZN(n_257_76_14480));
   INV_X1 i_257_76_14506 (.A(n_257_76_14480), .ZN(n_257_76_14481));
   NAND3_X1 i_257_76_14507 (.A1(n_257_76_14478), .A2(n_257_76_14479), .A3(
      n_257_76_14481), .ZN(n_257_76_14482));
   NAND4_X1 i_257_76_14508 (.A1(n_257_76_14156), .A2(n_257_76_14157), .A3(
      n_257_76_14158), .A4(n_257_76_14150), .ZN(n_257_76_14483));
   NOR2_X1 i_257_76_14509 (.A1(n_257_76_14482), .A2(n_257_76_14483), .ZN(
      n_257_76_14484));
   NAND3_X1 i_257_76_14510 (.A1(n_257_257), .A2(n_257_76_14201), .A3(
      n_257_76_14202), .ZN(n_257_76_14485));
   INV_X1 i_257_76_14511 (.A(n_257_76_14485), .ZN(n_257_76_14486));
   NAND4_X1 i_257_76_14512 (.A1(n_257_76_14484), .A2(n_257_76_14486), .A3(
      n_257_76_14121), .A4(n_257_76_14161), .ZN(n_257_76_14487));
   NOR2_X1 i_257_76_14513 (.A1(n_257_76_14487), .A2(n_257_76_14163), .ZN(
      n_257_76_14488));
   NAND2_X1 i_257_76_14514 (.A1(n_257_76_18064), .A2(n_257_76_14488), .ZN(
      n_257_76_14489));
   NAND3_X1 i_257_76_14515 (.A1(n_257_76_14403), .A2(n_257_76_14146), .A3(
      n_257_76_14147), .ZN(n_257_76_14490));
   NAND3_X1 i_257_76_14516 (.A1(n_257_76_17993), .A2(n_257_76_14188), .A3(
      n_257_421), .ZN(n_257_76_14491));
   INV_X1 i_257_76_14517 (.A(n_257_76_14491), .ZN(n_257_76_14492));
   NAND3_X1 i_257_76_14518 (.A1(n_257_76_14492), .A2(n_257_76_14191), .A3(
      n_257_76_14123), .ZN(n_257_76_14493));
   NOR2_X1 i_257_76_14519 (.A1(n_257_76_14490), .A2(n_257_76_14493), .ZN(
      n_257_76_14494));
   NAND2_X1 i_257_76_14520 (.A1(n_257_76_14152), .A2(n_257_76_14142), .ZN(
      n_257_76_14495));
   INV_X1 i_257_76_14521 (.A(n_257_76_14495), .ZN(n_257_76_14496));
   NAND3_X1 i_257_76_14522 (.A1(n_257_76_14194), .A2(n_257_76_14195), .A3(
      n_257_76_14144), .ZN(n_257_76_14497));
   INV_X1 i_257_76_14523 (.A(n_257_76_14497), .ZN(n_257_76_14498));
   NAND3_X1 i_257_76_14524 (.A1(n_257_76_14494), .A2(n_257_76_14496), .A3(
      n_257_76_14498), .ZN(n_257_76_14499));
   NAND4_X1 i_257_76_14525 (.A1(n_257_76_14198), .A2(n_257_76_14395), .A3(
      n_257_374), .A4(n_257_76_14151), .ZN(n_257_76_14500));
   NOR2_X1 i_257_76_14526 (.A1(n_257_76_14499), .A2(n_257_76_14500), .ZN(
      n_257_76_14501));
   INV_X1 i_257_76_14527 (.A(n_257_76_14159), .ZN(n_257_76_14502));
   NAND2_X1 i_257_76_14528 (.A1(n_257_76_14150), .A2(n_257_76_14206), .ZN(
      n_257_76_14503));
   NAND3_X1 i_257_76_14529 (.A1(n_257_76_14211), .A2(n_257_76_14122), .A3(
      n_257_76_14212), .ZN(n_257_76_14504));
   NOR2_X1 i_257_76_14530 (.A1(n_257_76_14503), .A2(n_257_76_14504), .ZN(
      n_257_76_14505));
   NAND3_X1 i_257_76_14531 (.A1(n_257_76_14501), .A2(n_257_76_14502), .A3(
      n_257_76_14505), .ZN(n_257_76_14506));
   INV_X1 i_257_76_14532 (.A(n_257_76_14506), .ZN(n_257_76_14507));
   NAND2_X1 i_257_76_14533 (.A1(n_257_76_14132), .A2(n_257_76_14507), .ZN(
      n_257_76_14508));
   NAND4_X1 i_257_76_14534 (.A1(n_257_76_14217), .A2(n_257_76_14295), .A3(
      n_257_76_14121), .A4(n_257_76_14161), .ZN(n_257_76_14509));
   NOR2_X1 i_257_76_14535 (.A1(n_257_76_14508), .A2(n_257_76_14509), .ZN(
      n_257_76_14510));
   NAND2_X1 i_257_76_14536 (.A1(n_257_76_18082), .A2(n_257_76_14510), .ZN(
      n_257_76_14511));
   NAND3_X1 i_257_76_14537 (.A1(n_257_76_14473), .A2(n_257_76_14489), .A3(
      n_257_76_14511), .ZN(n_257_76_14512));
   INV_X1 i_257_76_14538 (.A(n_257_76_14512), .ZN(n_257_76_14513));
   NAND4_X1 i_257_76_14539 (.A1(n_257_76_14365), .A2(n_257_76_14142), .A3(
      n_257_76_14195), .A4(n_257_76_14144), .ZN(n_257_76_14514));
   NAND2_X1 i_257_76_14540 (.A1(n_257_427), .A2(n_257_76_14188), .ZN(
      n_257_76_14515));
   INV_X1 i_257_76_14541 (.A(n_257_76_14515), .ZN(n_257_76_14516));
   NAND4_X1 i_257_76_14542 (.A1(n_257_76_14516), .A2(n_257_76_14123), .A3(
      n_257_217), .A4(n_257_76_17993), .ZN(n_257_76_14517));
   INV_X1 i_257_76_14543 (.A(n_257_76_14517), .ZN(n_257_76_14518));
   NAND3_X1 i_257_76_14544 (.A1(n_257_76_14518), .A2(n_257_76_14151), .A3(
      n_257_76_14152), .ZN(n_257_76_14519));
   NOR2_X1 i_257_76_14545 (.A1(n_257_76_14514), .A2(n_257_76_14519), .ZN(
      n_257_76_14520));
   NAND4_X1 i_257_76_14546 (.A1(n_257_76_14211), .A2(n_257_76_14122), .A3(
      n_257_76_14212), .A4(n_257_76_14198), .ZN(n_257_76_14521));
   INV_X1 i_257_76_14547 (.A(n_257_76_14521), .ZN(n_257_76_14522));
   NAND3_X1 i_257_76_14548 (.A1(n_257_76_14289), .A2(n_257_76_14520), .A3(
      n_257_76_14522), .ZN(n_257_76_14523));
   NOR2_X1 i_257_76_14549 (.A1(n_257_76_14242), .A2(n_257_76_14523), .ZN(
      n_257_76_14524));
   NAND3_X1 i_257_76_14550 (.A1(n_257_76_14524), .A2(n_257_76_14260), .A3(
      n_257_76_14132), .ZN(n_257_76_14525));
   INV_X1 i_257_76_14551 (.A(n_257_76_14525), .ZN(n_257_76_14526));
   NAND2_X1 i_257_76_14552 (.A1(n_257_76_18065), .A2(n_257_76_14526), .ZN(
      n_257_76_14527));
   NAND4_X1 i_257_76_14553 (.A1(n_257_76_14156), .A2(n_257_76_14157), .A3(
      n_257_76_14158), .A4(n_257_76_14468), .ZN(n_257_76_14528));
   NAND4_X1 i_257_76_14554 (.A1(n_257_451), .A2(n_257_76_14152), .A3(
      n_257_76_14142), .A4(n_257_477), .ZN(n_257_76_14529));
   INV_X1 i_257_76_14555 (.A(n_257_76_14529), .ZN(n_257_76_14530));
   NAND2_X1 i_257_76_14556 (.A1(n_257_76_14198), .A2(n_257_76_14151), .ZN(
      n_257_76_14531));
   INV_X1 i_257_76_14557 (.A(n_257_76_14531), .ZN(n_257_76_14532));
   NAND4_X1 i_257_76_14558 (.A1(n_257_76_14530), .A2(n_257_76_14532), .A3(
      n_257_76_14150), .A4(n_257_76_14122), .ZN(n_257_76_14533));
   NOR2_X1 i_257_76_14559 (.A1(n_257_76_14528), .A2(n_257_76_14533), .ZN(
      n_257_76_14534));
   NAND3_X1 i_257_76_14560 (.A1(n_257_76_14534), .A2(n_257_76_14121), .A3(
      n_257_76_14161), .ZN(n_257_76_14535));
   NOR2_X1 i_257_76_14561 (.A1(n_257_76_14535), .A2(n_257_76_14163), .ZN(
      n_257_76_14536));
   NAND2_X1 i_257_76_14562 (.A1(n_257_76_18063), .A2(n_257_76_14536), .ZN(
      n_257_76_14537));
   INV_X1 i_257_76_14563 (.A(n_257_76_14402), .ZN(n_257_76_14538));
   NAND3_X1 i_257_76_14564 (.A1(n_257_76_17993), .A2(n_257_76_14188), .A3(
      n_257_424), .ZN(n_257_76_14539));
   INV_X1 i_257_76_14565 (.A(n_257_76_14539), .ZN(n_257_76_14540));
   NAND3_X1 i_257_76_14566 (.A1(n_257_76_14540), .A2(n_257_76_14191), .A3(
      n_257_76_14123), .ZN(n_257_76_14541));
   INV_X1 i_257_76_14567 (.A(n_257_76_14541), .ZN(n_257_76_14542));
   NAND3_X1 i_257_76_14568 (.A1(n_257_76_14146), .A2(n_257_526), .A3(
      n_257_76_14147), .ZN(n_257_76_14543));
   INV_X1 i_257_76_14569 (.A(n_257_76_14543), .ZN(n_257_76_14544));
   NAND4_X1 i_257_76_14570 (.A1(n_257_76_14538), .A2(n_257_76_14542), .A3(
      n_257_76_14198), .A4(n_257_76_14544), .ZN(n_257_76_14545));
   INV_X1 i_257_76_14571 (.A(n_257_76_14545), .ZN(n_257_76_14546));
   NAND3_X1 i_257_76_14572 (.A1(n_257_76_14201), .A2(n_257_76_14202), .A3(
      n_257_76_14546), .ZN(n_257_76_14547));
   NOR2_X1 i_257_76_14573 (.A1(n_257_76_14215), .A2(n_257_76_14547), .ZN(
      n_257_76_14548));
   NAND3_X1 i_257_76_14574 (.A1(n_257_76_14548), .A2(n_257_76_14219), .A3(
      n_257_76_14132), .ZN(n_257_76_14549));
   INV_X1 i_257_76_14575 (.A(n_257_76_14549), .ZN(n_257_76_14550));
   NAND2_X1 i_257_76_14576 (.A1(n_257_76_18062), .A2(n_257_76_14550), .ZN(
      n_257_76_14551));
   NAND3_X1 i_257_76_14577 (.A1(n_257_76_14527), .A2(n_257_76_14537), .A3(
      n_257_76_14551), .ZN(n_257_76_14552));
   INV_X1 i_257_76_14578 (.A(n_257_76_14552), .ZN(n_257_76_14553));
   NAND2_X1 i_257_76_14579 (.A1(n_257_76_14188), .A2(n_257_422), .ZN(
      n_257_76_14554));
   INV_X1 i_257_76_14580 (.A(n_257_76_14554), .ZN(n_257_76_14555));
   NAND4_X1 i_257_76_14581 (.A1(n_257_335), .A2(n_257_76_14555), .A3(
      n_257_76_14123), .A4(n_257_76_17993), .ZN(n_257_76_14556));
   INV_X1 i_257_76_14582 (.A(n_257_76_14556), .ZN(n_257_76_14557));
   NAND3_X1 i_257_76_14583 (.A1(n_257_76_14395), .A2(n_257_76_14557), .A3(
      n_257_76_14151), .ZN(n_257_76_14558));
   INV_X1 i_257_76_14584 (.A(n_257_76_14558), .ZN(n_257_76_14559));
   NAND3_X1 i_257_76_14585 (.A1(n_257_76_14146), .A2(n_257_76_14147), .A3(
      n_257_76_14191), .ZN(n_257_76_14560));
   NOR2_X1 i_257_76_14586 (.A1(n_257_76_14402), .A2(n_257_76_14560), .ZN(
      n_257_76_14561));
   NAND3_X1 i_257_76_14587 (.A1(n_257_76_14152), .A2(n_257_76_14142), .A3(
      n_257_76_14194), .ZN(n_257_76_14562));
   INV_X1 i_257_76_14588 (.A(n_257_76_14562), .ZN(n_257_76_14563));
   NAND3_X1 i_257_76_14589 (.A1(n_257_76_14559), .A2(n_257_76_14561), .A3(
      n_257_76_14563), .ZN(n_257_76_14564));
   INV_X1 i_257_76_14590 (.A(n_257_76_14564), .ZN(n_257_76_14565));
   NAND3_X1 i_257_76_14591 (.A1(n_257_76_14565), .A2(n_257_76_14208), .A3(
      n_257_76_14522), .ZN(n_257_76_14566));
   NOR2_X1 i_257_76_14592 (.A1(n_257_76_14566), .A2(n_257_76_14242), .ZN(
      n_257_76_14567));
   NAND3_X1 i_257_76_14593 (.A1(n_257_76_14567), .A2(n_257_76_14219), .A3(
      n_257_76_14132), .ZN(n_257_76_14568));
   INV_X1 i_257_76_14594 (.A(n_257_76_14568), .ZN(n_257_76_14569));
   NAND2_X1 i_257_76_14595 (.A1(n_257_342), .A2(n_257_76_14569), .ZN(
      n_257_76_14570));
   NAND2_X1 i_257_76_14596 (.A1(n_257_420), .A2(n_257_494), .ZN(n_257_76_14571));
   NAND2_X1 i_257_76_14597 (.A1(n_257_590), .A2(n_257_428), .ZN(n_257_76_14572));
   NAND3_X1 i_257_76_14598 (.A1(n_257_413), .A2(n_257_484), .A3(n_257_442), 
      .ZN(n_257_76_14573));
   INV_X1 i_257_76_14599 (.A(n_257_76_14573), .ZN(n_257_76_14574));
   NAND2_X1 i_257_76_14600 (.A1(n_257_76_14572), .A2(n_257_76_14574), .ZN(
      n_257_76_14575));
   INV_X1 i_257_76_14601 (.A(n_257_76_14575), .ZN(n_257_76_14576));
   NAND4_X1 i_257_76_14602 (.A1(n_257_76_14123), .A2(n_257_76_14571), .A3(
      n_257_76_14576), .A4(n_257_76_14188), .ZN(n_257_76_14577));
   NOR2_X1 i_257_76_14603 (.A1(n_257_76_14284), .A2(n_257_76_14577), .ZN(
      n_257_76_14578));
   NAND2_X1 i_257_76_14604 (.A1(n_257_76_14194), .A2(n_257_76_14195), .ZN(
      n_257_76_14579));
   INV_X1 i_257_76_14605 (.A(n_257_76_14579), .ZN(n_257_76_14580));
   NAND3_X1 i_257_76_14606 (.A1(n_257_76_14144), .A2(n_257_76_14403), .A3(
      n_257_76_14146), .ZN(n_257_76_14581));
   INV_X1 i_257_76_14607 (.A(n_257_76_14581), .ZN(n_257_76_14582));
   NAND3_X1 i_257_76_14608 (.A1(n_257_76_14578), .A2(n_257_76_14580), .A3(
      n_257_76_14582), .ZN(n_257_76_14583));
   NAND4_X1 i_257_76_14609 (.A1(n_257_76_14395), .A2(n_257_76_14151), .A3(
      n_257_76_14152), .A4(n_257_76_14142), .ZN(n_257_76_14584));
   NOR2_X1 i_257_76_14610 (.A1(n_257_76_14583), .A2(n_257_76_14584), .ZN(
      n_257_76_14585));
   NAND3_X1 i_257_76_14611 (.A1(n_257_76_14585), .A2(n_257_76_14201), .A3(
      n_257_76_14202), .ZN(n_257_76_14586));
   NAND2_X1 i_257_76_14612 (.A1(n_257_76_14211), .A2(n_257_76_14399), .ZN(
      n_257_76_14587));
   NOR2_X1 i_257_76_14613 (.A1(n_257_76_14255), .A2(n_257_76_14587), .ZN(
      n_257_76_14588));
   NAND3_X1 i_257_76_14614 (.A1(n_257_76_14588), .A2(n_257_76_14205), .A3(
      n_257_76_14208), .ZN(n_257_76_14589));
   NOR2_X1 i_257_76_14615 (.A1(n_257_76_14586), .A2(n_257_76_14589), .ZN(
      n_257_76_14590));
   NAND3_X1 i_257_76_14616 (.A1(n_257_76_14590), .A2(n_257_76_14219), .A3(
      n_257_76_14132), .ZN(n_257_76_14591));
   INV_X1 i_257_76_14617 (.A(n_257_76_14591), .ZN(n_257_76_14592));
   NAND2_X1 i_257_76_14618 (.A1(n_257_76_18060), .A2(n_257_76_14592), .ZN(
      n_257_76_14593));
   INV_X1 i_257_76_14619 (.A(Small_Packet_Data_Size[25]), .ZN(n_257_76_14594));
   NAND2_X1 i_257_76_14620 (.A1(n_257_76_14572), .A2(n_257_76_17996), .ZN(
      n_257_76_14595));
   INV_X1 i_257_76_14621 (.A(n_257_76_14595), .ZN(n_257_76_14596));
   NAND4_X1 i_257_76_14622 (.A1(n_257_76_14123), .A2(n_257_76_14596), .A3(
      n_257_76_14571), .A4(n_257_76_14188), .ZN(n_257_76_14597));
   NAND2_X1 i_257_76_14623 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[25]), 
      .ZN(n_257_76_14598));
   AOI22_X1 i_257_76_14624 (.A1(n_257_654), .A2(n_257_76_17928), .B1(
      n_257_76_14597), .B2(n_257_76_14598), .ZN(n_257_76_14599));
   INV_X1 i_257_76_14625 (.A(n_257_76_14354), .ZN(n_257_76_14600));
   NAND2_X1 i_257_76_14626 (.A1(n_257_449), .A2(n_257_76_14600), .ZN(
      n_257_76_14601));
   INV_X1 i_257_76_14627 (.A(n_257_76_14440), .ZN(n_257_76_14602));
   NAND2_X1 i_257_76_14628 (.A1(n_257_447), .A2(n_257_76_14602), .ZN(
      n_257_76_14603));
   NAND3_X1 i_257_76_14629 (.A1(n_257_76_14601), .A2(n_257_76_14603), .A3(
      n_257_76_14556), .ZN(n_257_76_14604));
   INV_X1 i_257_76_14630 (.A(n_257_76_14604), .ZN(n_257_76_14605));
   INV_X1 i_257_76_14631 (.A(n_257_76_14167), .ZN(n_257_76_14606));
   NAND2_X1 i_257_76_14632 (.A1(n_257_446), .A2(n_257_76_14606), .ZN(
      n_257_76_14607));
   NAND2_X1 i_257_76_14633 (.A1(n_257_76_14517), .A2(n_257_76_14607), .ZN(
      n_257_76_14608));
   INV_X1 i_257_76_14634 (.A(n_257_76_14608), .ZN(n_257_76_14609));
   NAND2_X1 i_257_76_14635 (.A1(n_257_60), .A2(n_257_76_17918), .ZN(
      n_257_76_14610));
   NAND2_X1 i_257_76_14636 (.A1(n_257_726), .A2(n_257_76_15655), .ZN(
      n_257_76_14611));
   NAND3_X1 i_257_76_14637 (.A1(n_257_438), .A2(n_257_1090), .A3(n_257_442), 
      .ZN(n_257_76_14612));
   NAND2_X1 i_257_76_14638 (.A1(n_257_440), .A2(n_257_76_14125), .ZN(
      n_257_76_14613));
   NAND4_X1 i_257_76_14639 (.A1(n_257_76_14610), .A2(n_257_76_14611), .A3(
      n_257_76_14612), .A4(n_257_76_14613), .ZN(n_257_76_14614));
   INV_X1 i_257_76_14640 (.A(n_257_76_14614), .ZN(n_257_76_14615));
   NAND4_X1 i_257_76_14641 (.A1(n_257_76_14599), .A2(n_257_76_14605), .A3(
      n_257_76_14609), .A4(n_257_76_14615), .ZN(n_257_76_14616));
   NAND2_X1 i_257_76_14642 (.A1(n_257_886), .A2(n_257_76_17903), .ZN(
      n_257_76_14617));
   NAND3_X1 i_257_76_14643 (.A1(n_257_988), .A2(n_257_441), .A3(n_257_442), 
      .ZN(n_257_76_14618));
   NAND3_X1 i_257_76_14644 (.A1(n_257_451), .A2(n_257_477), .A3(n_257_76_14466), 
      .ZN(n_257_76_14619));
   NAND2_X1 i_257_76_14645 (.A1(n_257_138), .A2(n_257_76_17925), .ZN(
      n_257_76_14620));
   NAND4_X1 i_257_76_14646 (.A1(n_257_76_14617), .A2(n_257_76_14618), .A3(
      n_257_76_14619), .A4(n_257_76_14620), .ZN(n_257_76_14621));
   NOR2_X1 i_257_76_14647 (.A1(n_257_76_14616), .A2(n_257_76_14621), .ZN(
      n_257_76_14622));
   NAND2_X1 i_257_76_14648 (.A1(n_257_100), .A2(n_257_76_17932), .ZN(
      n_257_76_14623));
   NAND2_X1 i_257_76_14649 (.A1(n_257_76_14199), .A2(n_257_76_14623), .ZN(
      n_257_76_14624));
   INV_X1 i_257_76_14650 (.A(n_257_76_14624), .ZN(n_257_76_14625));
   NAND2_X1 i_257_76_14651 (.A1(n_257_822), .A2(n_257_76_17952), .ZN(
      n_257_76_14626));
   NAND2_X1 i_257_76_14652 (.A1(n_257_758), .A2(n_257_76_17935), .ZN(
      n_257_76_14627));
   NAND2_X1 i_257_76_14653 (.A1(n_257_924), .A2(n_257_76_17940), .ZN(
      n_257_76_14628));
   NAND4_X1 i_257_76_14654 (.A1(n_257_76_14545), .A2(n_257_76_14626), .A3(
      n_257_76_14627), .A4(n_257_76_14628), .ZN(n_257_76_14629));
   INV_X1 i_257_76_14655 (.A(n_257_76_14629), .ZN(n_257_76_14630));
   NAND3_X1 i_257_76_14656 (.A1(n_257_76_14622), .A2(n_257_76_14625), .A3(
      n_257_76_14630), .ZN(n_257_76_14631));
   NAND2_X1 i_257_76_14657 (.A1(n_257_1020), .A2(n_257_76_17964), .ZN(
      n_257_76_14632));
   NAND2_X1 i_257_76_14658 (.A1(n_257_694), .A2(n_257_76_17958), .ZN(
      n_257_76_14633));
   NAND2_X1 i_257_76_14659 (.A1(n_257_177), .A2(n_257_76_17331), .ZN(
      n_257_76_14634));
   NAND3_X1 i_257_76_14660 (.A1(n_257_76_14632), .A2(n_257_76_14633), .A3(
      n_257_76_14634), .ZN(n_257_76_14635));
   NOR2_X1 i_257_76_14661 (.A1(n_257_76_14631), .A2(n_257_76_14635), .ZN(
      n_257_76_14636));
   NAND2_X1 i_257_76_14662 (.A1(n_257_1052), .A2(n_257_76_17969), .ZN(
      n_257_76_14637));
   NAND3_X1 i_257_76_14663 (.A1(n_257_76_14637), .A2(n_257_76_14506), .A3(
      n_257_76_14292), .ZN(n_257_76_14638));
   INV_X1 i_257_76_14664 (.A(n_257_76_14638), .ZN(n_257_76_14639));
   NAND3_X1 i_257_76_14665 (.A1(n_257_76_14636), .A2(n_257_76_14487), .A3(
      n_257_76_14639), .ZN(n_257_76_14640));
   NAND3_X1 i_257_76_14666 (.A1(n_257_76_14570), .A2(n_257_76_14593), .A3(
      n_257_76_14640), .ZN(n_257_76_14641));
   INV_X1 i_257_76_14667 (.A(n_257_76_14641), .ZN(n_257_76_14642));
   NAND3_X1 i_257_76_14668 (.A1(n_257_76_14513), .A2(n_257_76_14553), .A3(
      n_257_76_14642), .ZN(n_257_76_14643));
   NOR2_X1 i_257_76_14669 (.A1(n_257_76_14462), .A2(n_257_76_14643), .ZN(
      n_257_76_14644));
   NAND2_X1 i_257_76_14670 (.A1(n_257_76_14344), .A2(n_257_76_14644), .ZN(n_25));
   NAND2_X1 i_257_76_14671 (.A1(n_257_1021), .A2(n_257_444), .ZN(n_257_76_14645));
   NAND2_X1 i_257_76_14672 (.A1(n_257_989), .A2(n_257_441), .ZN(n_257_76_14646));
   NOR2_X1 i_257_76_14673 (.A1(n_257_1085), .A2(n_257_76_17412), .ZN(
      n_257_76_14647));
   NAND3_X1 i_257_76_14674 (.A1(n_257_76_14647), .A2(n_257_440), .A3(n_257_957), 
      .ZN(n_257_76_14648));
   INV_X1 i_257_76_14675 (.A(n_257_76_14648), .ZN(n_257_76_14649));
   NAND2_X1 i_257_76_14676 (.A1(n_257_76_14646), .A2(n_257_76_14649), .ZN(
      n_257_76_14650));
   INV_X1 i_257_76_14677 (.A(n_257_76_14650), .ZN(n_257_76_14651));
   NAND2_X1 i_257_76_14678 (.A1(n_257_76_14645), .A2(n_257_76_14651), .ZN(
      n_257_76_14652));
   INV_X1 i_257_76_14679 (.A(n_257_76_14652), .ZN(n_257_76_14653));
   NAND2_X1 i_257_76_14680 (.A1(n_257_1053), .A2(n_257_443), .ZN(n_257_76_14654));
   NAND2_X1 i_257_76_14681 (.A1(n_257_76_14653), .A2(n_257_76_14654), .ZN(
      n_257_76_14655));
   INV_X1 i_257_76_14682 (.A(n_257_76_14655), .ZN(n_257_76_14656));
   NAND2_X1 i_257_76_14683 (.A1(n_257_17), .A2(n_257_76_14656), .ZN(
      n_257_76_14657));
   NAND2_X1 i_257_76_14684 (.A1(n_257_695), .A2(n_257_448), .ZN(n_257_76_14658));
   NAND2_X1 i_257_76_14685 (.A1(n_257_823), .A2(n_257_437), .ZN(n_257_76_14659));
   NAND2_X1 i_257_76_14686 (.A1(n_257_759), .A2(n_257_436), .ZN(n_257_76_14660));
   NAND2_X1 i_257_76_14687 (.A1(n_257_887), .A2(n_257_445), .ZN(n_257_76_14661));
   NAND2_X1 i_257_76_14688 (.A1(n_257_925), .A2(n_257_439), .ZN(n_257_76_14662));
   NAND4_X1 i_257_76_14689 (.A1(n_257_76_14659), .A2(n_257_76_14660), .A3(
      n_257_76_14661), .A4(n_257_76_14662), .ZN(n_257_76_14663));
   INV_X1 i_257_76_14690 (.A(n_257_76_14663), .ZN(n_257_76_14664));
   NAND2_X1 i_257_76_14691 (.A1(n_257_446), .A2(n_257_855), .ZN(n_257_76_14665));
   NAND2_X1 i_257_76_14692 (.A1(n_257_449), .A2(n_257_663), .ZN(n_257_76_14666));
   NAND2_X1 i_257_76_14693 (.A1(n_257_76_14665), .A2(n_257_76_14666), .ZN(
      n_257_76_14667));
   INV_X1 i_257_76_14694 (.A(n_257_76_14667), .ZN(n_257_76_14668));
   NAND2_X1 i_257_76_14695 (.A1(n_257_447), .A2(n_257_791), .ZN(n_257_76_14669));
   NAND2_X1 i_257_76_14696 (.A1(n_257_61), .A2(n_257_433), .ZN(n_257_76_14670));
   NAND2_X1 i_257_76_14697 (.A1(n_257_76_14669), .A2(n_257_76_14670), .ZN(
      n_257_76_14671));
   INV_X1 i_257_76_14698 (.A(n_257_76_14671), .ZN(n_257_76_14672));
   NAND2_X1 i_257_76_14699 (.A1(n_257_727), .A2(n_257_435), .ZN(n_257_76_14673));
   NAND2_X1 i_257_76_14700 (.A1(n_257_440), .A2(n_257_957), .ZN(n_257_76_14674));
   NAND2_X1 i_257_76_14701 (.A1(n_257_623), .A2(n_257_442), .ZN(n_257_76_14675));
   INV_X1 i_257_76_14702 (.A(n_257_76_14675), .ZN(n_257_76_14676));
   NAND2_X1 i_257_76_14703 (.A1(n_257_76_14676), .A2(n_257_432), .ZN(
      n_257_76_14677));
   NOR2_X1 i_257_76_14704 (.A1(n_257_76_14677), .A2(n_257_1085), .ZN(
      n_257_76_14678));
   NAND2_X1 i_257_76_14705 (.A1(n_257_438), .A2(n_257_893), .ZN(n_257_76_14679));
   NAND4_X1 i_257_76_14706 (.A1(n_257_76_14673), .A2(n_257_76_14674), .A3(
      n_257_76_14678), .A4(n_257_76_14679), .ZN(n_257_76_14680));
   INV_X1 i_257_76_14707 (.A(n_257_76_14680), .ZN(n_257_76_14681));
   NAND3_X1 i_257_76_14708 (.A1(n_257_76_14668), .A2(n_257_76_14672), .A3(
      n_257_76_14681), .ZN(n_257_76_14682));
   NAND2_X1 i_257_76_14709 (.A1(n_257_451), .A2(n_257_478), .ZN(n_257_76_14683));
   NAND2_X1 i_257_76_14710 (.A1(n_257_655), .A2(n_257_450), .ZN(n_257_76_14684));
   NAND3_X1 i_257_76_14711 (.A1(n_257_76_14646), .A2(n_257_76_14683), .A3(
      n_257_76_14684), .ZN(n_257_76_14685));
   NOR2_X1 i_257_76_14712 (.A1(n_257_76_14682), .A2(n_257_76_14685), .ZN(
      n_257_76_14686));
   NAND4_X1 i_257_76_14713 (.A1(n_257_76_14658), .A2(n_257_76_14645), .A3(
      n_257_76_14664), .A4(n_257_76_14686), .ZN(n_257_76_14687));
   INV_X1 i_257_76_14714 (.A(n_257_76_14654), .ZN(n_257_76_14688));
   NOR2_X1 i_257_76_14715 (.A1(n_257_76_14687), .A2(n_257_76_14688), .ZN(
      n_257_76_14689));
   NAND2_X1 i_257_76_14716 (.A1(n_257_68), .A2(n_257_76_14689), .ZN(
      n_257_76_14690));
   NAND2_X1 i_257_76_14717 (.A1(n_257_76_14674), .A2(n_257_76_14679), .ZN(
      n_257_76_14691));
   INV_X1 i_257_76_14718 (.A(n_257_76_14691), .ZN(n_257_76_14692));
   INV_X1 i_257_76_14719 (.A(n_257_76_14647), .ZN(n_257_76_14693));
   INV_X1 i_257_76_14720 (.A(n_257_450), .ZN(n_257_76_14694));
   NOR2_X1 i_257_76_14721 (.A1(n_257_76_14693), .A2(n_257_76_14694), .ZN(
      n_257_76_14695));
   NAND4_X1 i_257_76_14722 (.A1(n_257_76_14692), .A2(n_257_655), .A3(
      n_257_76_14695), .A4(n_257_76_14673), .ZN(n_257_76_14696));
   INV_X1 i_257_76_14723 (.A(n_257_76_14696), .ZN(n_257_76_14697));
   NAND3_X1 i_257_76_14724 (.A1(n_257_76_14665), .A2(n_257_76_14666), .A3(
      n_257_76_14669), .ZN(n_257_76_14698));
   INV_X1 i_257_76_14725 (.A(n_257_76_14698), .ZN(n_257_76_14699));
   NAND4_X1 i_257_76_14726 (.A1(n_257_76_14662), .A2(n_257_76_14697), .A3(
      n_257_76_14646), .A4(n_257_76_14699), .ZN(n_257_76_14700));
   NAND3_X1 i_257_76_14727 (.A1(n_257_76_14659), .A2(n_257_76_14660), .A3(
      n_257_76_14661), .ZN(n_257_76_14701));
   NOR2_X1 i_257_76_14728 (.A1(n_257_76_14700), .A2(n_257_76_14701), .ZN(
      n_257_76_14702));
   NAND3_X1 i_257_76_14729 (.A1(n_257_76_14702), .A2(n_257_76_14658), .A3(
      n_257_76_14645), .ZN(n_257_76_14703));
   NOR2_X1 i_257_76_14730 (.A1(n_257_76_14703), .A2(n_257_76_14688), .ZN(
      n_257_76_14704));
   NAND2_X1 i_257_76_14731 (.A1(n_257_28), .A2(n_257_76_14704), .ZN(
      n_257_76_14705));
   NAND3_X1 i_257_76_14732 (.A1(n_257_76_14657), .A2(n_257_76_14690), .A3(
      n_257_76_14705), .ZN(n_257_76_14706));
   NAND3_X1 i_257_76_14733 (.A1(n_257_76_14674), .A2(n_257_76_14647), .A3(
      n_257_439), .ZN(n_257_76_14707));
   INV_X1 i_257_76_14734 (.A(n_257_76_14707), .ZN(n_257_76_14708));
   NAND3_X1 i_257_76_14735 (.A1(n_257_76_14646), .A2(n_257_925), .A3(
      n_257_76_14708), .ZN(n_257_76_14709));
   INV_X1 i_257_76_14736 (.A(n_257_76_14709), .ZN(n_257_76_14710));
   NAND2_X1 i_257_76_14737 (.A1(n_257_76_14645), .A2(n_257_76_14710), .ZN(
      n_257_76_14711));
   INV_X1 i_257_76_14738 (.A(n_257_76_14711), .ZN(n_257_76_14712));
   NAND2_X1 i_257_76_14739 (.A1(n_257_76_14712), .A2(n_257_76_14654), .ZN(
      n_257_76_14713));
   INV_X1 i_257_76_14740 (.A(n_257_76_14713), .ZN(n_257_76_14714));
   NAND2_X1 i_257_76_14741 (.A1(n_257_76_18084), .A2(n_257_76_14714), .ZN(
      n_257_76_14715));
   NAND3_X1 i_257_76_14742 (.A1(n_257_76_14679), .A2(n_257_76_14647), .A3(
      n_257_855), .ZN(n_257_76_14716));
   NAND2_X1 i_257_76_14743 (.A1(n_257_446), .A2(n_257_76_14674), .ZN(
      n_257_76_14717));
   NOR2_X1 i_257_76_14744 (.A1(n_257_76_14716), .A2(n_257_76_14717), .ZN(
      n_257_76_14718));
   NAND2_X1 i_257_76_14745 (.A1(n_257_76_14646), .A2(n_257_76_14718), .ZN(
      n_257_76_14719));
   INV_X1 i_257_76_14746 (.A(n_257_76_14719), .ZN(n_257_76_14720));
   NAND3_X1 i_257_76_14747 (.A1(n_257_76_14720), .A2(n_257_76_14661), .A3(
      n_257_76_14662), .ZN(n_257_76_14721));
   INV_X1 i_257_76_14748 (.A(n_257_76_14721), .ZN(n_257_76_14722));
   NAND2_X1 i_257_76_14749 (.A1(n_257_76_14645), .A2(n_257_76_14722), .ZN(
      n_257_76_14723));
   INV_X1 i_257_76_14750 (.A(n_257_76_14723), .ZN(n_257_76_14724));
   NAND2_X1 i_257_76_14751 (.A1(n_257_76_14724), .A2(n_257_76_14654), .ZN(
      n_257_76_14725));
   INV_X1 i_257_76_14752 (.A(n_257_76_14725), .ZN(n_257_76_14726));
   NAND2_X1 i_257_76_14753 (.A1(n_257_76_18070), .A2(n_257_76_14726), .ZN(
      n_257_76_14727));
   NAND2_X1 i_257_76_14754 (.A1(n_257_527), .A2(n_257_424), .ZN(n_257_76_14728));
   NAND3_X1 i_257_76_14755 (.A1(n_257_76_14728), .A2(n_257_76_14665), .A3(
      n_257_76_14666), .ZN(n_257_76_14729));
   INV_X1 i_257_76_14756 (.A(n_257_76_14729), .ZN(n_257_76_14730));
   NAND3_X1 i_257_76_14757 (.A1(n_257_76_14669), .A2(n_257_76_14670), .A3(
      n_257_76_14673), .ZN(n_257_76_14731));
   INV_X1 i_257_76_14758 (.A(n_257_76_14731), .ZN(n_257_76_14732));
   INV_X1 i_257_76_14759 (.A(n_257_1085), .ZN(n_257_76_14733));
   NAND2_X1 i_257_76_14760 (.A1(n_257_432), .A2(n_257_623), .ZN(n_257_76_14734));
   NAND4_X1 i_257_76_14761 (.A1(n_257_76_17990), .A2(n_257_76_14733), .A3(
      n_257_76_14734), .A4(n_257_423), .ZN(n_257_76_14735));
   INV_X1 i_257_76_14762 (.A(n_257_76_14735), .ZN(n_257_76_14736));
   NAND2_X1 i_257_76_14763 (.A1(n_257_218), .A2(n_257_427), .ZN(n_257_76_14737));
   NAND4_X1 i_257_76_14764 (.A1(n_257_76_14736), .A2(n_257_76_14737), .A3(
      n_257_76_14674), .A4(n_257_76_14679), .ZN(n_257_76_14738));
   INV_X1 i_257_76_14765 (.A(n_257_76_14738), .ZN(n_257_76_14739));
   NAND3_X1 i_257_76_14766 (.A1(n_257_76_14730), .A2(n_257_76_14732), .A3(
      n_257_76_14739), .ZN(n_257_76_14740));
   NAND2_X1 i_257_76_14767 (.A1(n_257_139), .A2(n_257_430), .ZN(n_257_76_14741));
   NAND3_X1 i_257_76_14768 (.A1(n_257_298), .A2(n_257_76_14741), .A3(
      n_257_76_14684), .ZN(n_257_76_14742));
   NOR2_X1 i_257_76_14769 (.A1(n_257_76_14740), .A2(n_257_76_14742), .ZN(
      n_257_76_14743));
   INV_X1 i_257_76_14770 (.A(n_257_76_14701), .ZN(n_257_76_14744));
   NAND2_X1 i_257_76_14771 (.A1(n_257_559), .A2(n_257_426), .ZN(n_257_76_14745));
   NAND3_X1 i_257_76_14772 (.A1(n_257_76_14662), .A2(n_257_76_14745), .A3(
      n_257_76_14646), .ZN(n_257_76_14746));
   INV_X1 i_257_76_14773 (.A(n_257_76_14746), .ZN(n_257_76_14747));
   NAND3_X1 i_257_76_14774 (.A1(n_257_76_14743), .A2(n_257_76_14744), .A3(
      n_257_76_14747), .ZN(n_257_76_14748));
   INV_X1 i_257_76_14775 (.A(n_257_76_14748), .ZN(n_257_76_14749));
   NAND2_X1 i_257_76_14776 (.A1(n_257_76_14658), .A2(n_257_76_14645), .ZN(
      n_257_76_14750));
   INV_X1 i_257_76_14777 (.A(n_257_76_14750), .ZN(n_257_76_14751));
   NAND2_X1 i_257_76_14778 (.A1(n_257_178), .A2(n_257_429), .ZN(n_257_76_14752));
   NAND2_X1 i_257_76_14779 (.A1(n_257_258), .A2(n_257_425), .ZN(n_257_76_14753));
   NAND2_X1 i_257_76_14780 (.A1(n_257_101), .A2(n_257_431), .ZN(n_257_76_14754));
   NAND4_X1 i_257_76_14781 (.A1(n_257_76_14752), .A2(n_257_76_14753), .A3(
      n_257_76_14754), .A4(n_257_76_14683), .ZN(n_257_76_14755));
   INV_X1 i_257_76_14782 (.A(n_257_76_14755), .ZN(n_257_76_14756));
   NAND4_X1 i_257_76_14783 (.A1(n_257_76_14749), .A2(n_257_76_14751), .A3(
      n_257_76_14654), .A4(n_257_76_14756), .ZN(n_257_76_14757));
   INV_X1 i_257_76_14784 (.A(n_257_76_14757), .ZN(n_257_76_14758));
   NAND2_X1 i_257_76_14785 (.A1(n_257_76_18066), .A2(n_257_76_14758), .ZN(
      n_257_76_14759));
   NAND3_X1 i_257_76_14786 (.A1(n_257_76_14715), .A2(n_257_76_14727), .A3(
      n_257_76_14759), .ZN(n_257_76_14760));
   NOR2_X1 i_257_76_14787 (.A1(n_257_76_14706), .A2(n_257_76_14760), .ZN(
      n_257_76_14761));
   NAND3_X1 i_257_76_14788 (.A1(n_257_989), .A2(n_257_441), .A3(n_257_76_14647), 
      .ZN(n_257_76_14762));
   INV_X1 i_257_76_14789 (.A(n_257_76_14762), .ZN(n_257_76_14763));
   NAND2_X1 i_257_76_14790 (.A1(n_257_76_14645), .A2(n_257_76_14763), .ZN(
      n_257_76_14764));
   INV_X1 i_257_76_14791 (.A(n_257_76_14764), .ZN(n_257_76_14765));
   NAND2_X1 i_257_76_14792 (.A1(n_257_76_14765), .A2(n_257_76_14654), .ZN(
      n_257_76_14766));
   INV_X1 i_257_76_14793 (.A(n_257_76_14766), .ZN(n_257_76_14767));
   NAND2_X1 i_257_76_14794 (.A1(n_257_76_18071), .A2(n_257_76_14767), .ZN(
      n_257_76_14768));
   NAND3_X1 i_257_76_14795 (.A1(n_257_76_14647), .A2(n_257_727), .A3(n_257_435), 
      .ZN(n_257_76_14769));
   INV_X1 i_257_76_14796 (.A(n_257_76_14769), .ZN(n_257_76_14770));
   NAND4_X1 i_257_76_14797 (.A1(n_257_76_14770), .A2(n_257_76_14692), .A3(
      n_257_76_14665), .A4(n_257_76_14669), .ZN(n_257_76_14771));
   INV_X1 i_257_76_14798 (.A(n_257_76_14771), .ZN(n_257_76_14772));
   NAND3_X1 i_257_76_14799 (.A1(n_257_76_14662), .A2(n_257_76_14772), .A3(
      n_257_76_14646), .ZN(n_257_76_14773));
   NOR2_X1 i_257_76_14800 (.A1(n_257_76_14701), .A2(n_257_76_14773), .ZN(
      n_257_76_14774));
   NAND2_X1 i_257_76_14801 (.A1(n_257_76_14645), .A2(n_257_76_14774), .ZN(
      n_257_76_14775));
   NOR2_X1 i_257_76_14802 (.A1(n_257_76_14775), .A2(n_257_76_14688), .ZN(
      n_257_76_14776));
   NAND2_X1 i_257_76_14803 (.A1(n_257_76_18078), .A2(n_257_76_14776), .ZN(
      n_257_76_14777));
   NAND4_X1 i_257_76_14804 (.A1(n_257_76_14646), .A2(n_257_76_14683), .A3(
      n_257_76_14741), .A4(n_257_76_14684), .ZN(n_257_76_14778));
   NAND3_X1 i_257_76_14805 (.A1(n_257_591), .A2(n_257_428), .A3(n_257_442), 
      .ZN(n_257_76_14779));
   INV_X1 i_257_76_14806 (.A(n_257_76_14779), .ZN(n_257_76_14780));
   NAND3_X1 i_257_76_14807 (.A1(n_257_76_14733), .A2(n_257_76_14734), .A3(
      n_257_76_14780), .ZN(n_257_76_14781));
   INV_X1 i_257_76_14808 (.A(n_257_76_14781), .ZN(n_257_76_14782));
   NAND4_X1 i_257_76_14809 (.A1(n_257_76_14673), .A2(n_257_76_14782), .A3(
      n_257_76_14674), .A4(n_257_76_14679), .ZN(n_257_76_14783));
   INV_X1 i_257_76_14810 (.A(n_257_76_14783), .ZN(n_257_76_14784));
   NAND3_X1 i_257_76_14811 (.A1(n_257_76_14784), .A2(n_257_76_14668), .A3(
      n_257_76_14672), .ZN(n_257_76_14785));
   NOR2_X1 i_257_76_14812 (.A1(n_257_76_14778), .A2(n_257_76_14785), .ZN(
      n_257_76_14786));
   NAND2_X1 i_257_76_14813 (.A1(n_257_76_14754), .A2(n_257_76_14659), .ZN(
      n_257_76_14787));
   INV_X1 i_257_76_14814 (.A(n_257_76_14787), .ZN(n_257_76_14788));
   NAND3_X1 i_257_76_14815 (.A1(n_257_76_14660), .A2(n_257_76_14661), .A3(
      n_257_76_14662), .ZN(n_257_76_14789));
   INV_X1 i_257_76_14816 (.A(n_257_76_14789), .ZN(n_257_76_14790));
   NAND4_X1 i_257_76_14817 (.A1(n_257_76_14786), .A2(n_257_76_14788), .A3(
      n_257_76_14752), .A4(n_257_76_14790), .ZN(n_257_76_14791));
   INV_X1 i_257_76_14818 (.A(n_257_76_14791), .ZN(n_257_76_14792));
   NAND3_X1 i_257_76_14819 (.A1(n_257_76_14792), .A2(n_257_76_14751), .A3(
      n_257_76_14654), .ZN(n_257_76_14793));
   INV_X1 i_257_76_14820 (.A(n_257_76_14793), .ZN(n_257_76_14794));
   NAND2_X1 i_257_76_14821 (.A1(n_257_76_18074), .A2(n_257_76_14794), .ZN(
      n_257_76_14795));
   NAND3_X1 i_257_76_14822 (.A1(n_257_76_14768), .A2(n_257_76_14777), .A3(
      n_257_76_14795), .ZN(n_257_76_14796));
   NAND2_X1 i_257_76_14823 (.A1(n_257_1085), .A2(n_257_442), .ZN(n_257_76_14797));
   INV_X1 i_257_76_14824 (.A(n_257_76_14797), .ZN(n_257_76_14798));
   NAND2_X1 i_257_76_14825 (.A1(n_257_13), .A2(n_257_76_14798), .ZN(
      n_257_76_14799));
   NAND4_X1 i_257_76_14826 (.A1(n_257_76_14674), .A2(n_257_76_14679), .A3(
      n_257_76_14647), .A4(n_257_445), .ZN(n_257_76_14800));
   INV_X1 i_257_76_14827 (.A(n_257_76_14800), .ZN(n_257_76_14801));
   NAND3_X1 i_257_76_14828 (.A1(n_257_887), .A2(n_257_76_14646), .A3(
      n_257_76_14801), .ZN(n_257_76_14802));
   INV_X1 i_257_76_14829 (.A(n_257_76_14662), .ZN(n_257_76_14803));
   NOR2_X1 i_257_76_14830 (.A1(n_257_76_14802), .A2(n_257_76_14803), .ZN(
      n_257_76_14804));
   NAND2_X1 i_257_76_14831 (.A1(n_257_76_14645), .A2(n_257_76_14804), .ZN(
      n_257_76_14805));
   INV_X1 i_257_76_14832 (.A(n_257_76_14805), .ZN(n_257_76_14806));
   NAND2_X1 i_257_76_14833 (.A1(n_257_76_14806), .A2(n_257_76_14654), .ZN(
      n_257_76_14807));
   INV_X1 i_257_76_14834 (.A(n_257_76_14807), .ZN(n_257_76_14808));
   NAND2_X1 i_257_76_14835 (.A1(n_257_76_18077), .A2(n_257_76_14808), .ZN(
      n_257_76_14809));
   NAND2_X1 i_257_76_14836 (.A1(n_257_76_14799), .A2(n_257_76_14809), .ZN(
      n_257_76_14810));
   NOR2_X1 i_257_76_14837 (.A1(n_257_76_14796), .A2(n_257_76_14810), .ZN(
      n_257_76_14811));
   NAND3_X1 i_257_76_14838 (.A1(n_257_76_14659), .A2(n_257_76_14661), .A3(
      n_257_76_14662), .ZN(n_257_76_14812));
   NAND2_X1 i_257_76_14839 (.A1(n_257_76_14665), .A2(n_257_76_14669), .ZN(
      n_257_76_14813));
   INV_X1 i_257_76_14840 (.A(n_257_76_14813), .ZN(n_257_76_14814));
   NAND4_X1 i_257_76_14841 (.A1(n_257_76_14674), .A2(n_257_76_14679), .A3(
      n_257_76_14647), .A4(n_257_436), .ZN(n_257_76_14815));
   INV_X1 i_257_76_14842 (.A(n_257_76_14815), .ZN(n_257_76_14816));
   NAND4_X1 i_257_76_14843 (.A1(n_257_759), .A2(n_257_76_14646), .A3(
      n_257_76_14814), .A4(n_257_76_14816), .ZN(n_257_76_14817));
   NOR2_X1 i_257_76_14844 (.A1(n_257_76_14812), .A2(n_257_76_14817), .ZN(
      n_257_76_14818));
   NAND2_X1 i_257_76_14845 (.A1(n_257_76_14645), .A2(n_257_76_14818), .ZN(
      n_257_76_14819));
   NOR2_X1 i_257_76_14846 (.A1(n_257_76_14819), .A2(n_257_76_14688), .ZN(
      n_257_76_14820));
   NAND2_X1 i_257_76_14847 (.A1(n_257_76_18069), .A2(n_257_76_14820), .ZN(
      n_257_76_14821));
   NAND4_X1 i_257_76_14848 (.A1(n_257_76_17990), .A2(n_257_76_14733), .A3(
      n_257_76_14734), .A4(n_257_426), .ZN(n_257_76_14822));
   INV_X1 i_257_76_14849 (.A(n_257_76_14822), .ZN(n_257_76_14823));
   NAND4_X1 i_257_76_14850 (.A1(n_257_76_14823), .A2(n_257_76_14737), .A3(
      n_257_76_14674), .A4(n_257_76_14679), .ZN(n_257_76_14824));
   INV_X1 i_257_76_14851 (.A(n_257_76_14824), .ZN(n_257_76_14825));
   NAND3_X1 i_257_76_14852 (.A1(n_257_76_14825), .A2(n_257_76_14732), .A3(
      n_257_76_14668), .ZN(n_257_76_14826));
   NAND3_X1 i_257_76_14853 (.A1(n_257_76_14741), .A2(n_257_559), .A3(
      n_257_76_14684), .ZN(n_257_76_14827));
   NOR2_X1 i_257_76_14854 (.A1(n_257_76_14826), .A2(n_257_76_14827), .ZN(
      n_257_76_14828));
   NAND3_X1 i_257_76_14855 (.A1(n_257_76_14661), .A2(n_257_76_14662), .A3(
      n_257_76_14646), .ZN(n_257_76_14829));
   INV_X1 i_257_76_14856 (.A(n_257_76_14829), .ZN(n_257_76_14830));
   NAND2_X1 i_257_76_14857 (.A1(n_257_76_14659), .A2(n_257_76_14660), .ZN(
      n_257_76_14831));
   INV_X1 i_257_76_14858 (.A(n_257_76_14831), .ZN(n_257_76_14832));
   NAND3_X1 i_257_76_14859 (.A1(n_257_76_14828), .A2(n_257_76_14830), .A3(
      n_257_76_14832), .ZN(n_257_76_14833));
   INV_X1 i_257_76_14860 (.A(n_257_76_14833), .ZN(n_257_76_14834));
   NAND2_X1 i_257_76_14861 (.A1(n_257_76_14654), .A2(n_257_76_14834), .ZN(
      n_257_76_14835));
   NAND2_X1 i_257_76_14862 (.A1(n_257_76_14754), .A2(n_257_76_14683), .ZN(
      n_257_76_14836));
   INV_X1 i_257_76_14863 (.A(n_257_76_14836), .ZN(n_257_76_14837));
   NAND4_X1 i_257_76_14864 (.A1(n_257_76_14658), .A2(n_257_76_14645), .A3(
      n_257_76_14752), .A4(n_257_76_14837), .ZN(n_257_76_14838));
   NOR2_X1 i_257_76_14865 (.A1(n_257_76_14835), .A2(n_257_76_14838), .ZN(
      n_257_76_14839));
   NAND2_X1 i_257_76_14866 (.A1(n_257_76_18076), .A2(n_257_76_14839), .ZN(
      n_257_76_14840));
   NOR2_X1 i_257_76_14867 (.A1(n_257_76_14693), .A2(n_257_76_15197), .ZN(
      n_257_76_14841));
   NAND2_X1 i_257_76_14868 (.A1(n_257_1053), .A2(n_257_76_14841), .ZN(
      n_257_76_14842));
   INV_X1 i_257_76_14869 (.A(n_257_76_14842), .ZN(n_257_76_14843));
   NAND2_X1 i_257_76_14870 (.A1(n_257_76_18072), .A2(n_257_76_14843), .ZN(
      n_257_76_14844));
   NAND3_X1 i_257_76_14871 (.A1(n_257_76_14821), .A2(n_257_76_14840), .A3(
      n_257_76_14844), .ZN(n_257_76_14845));
   NAND4_X1 i_257_76_14872 (.A1(n_257_76_14674), .A2(n_257_76_14679), .A3(
      n_257_76_14647), .A4(n_257_437), .ZN(n_257_76_14846));
   INV_X1 i_257_76_14873 (.A(n_257_76_14665), .ZN(n_257_76_14847));
   NOR2_X1 i_257_76_14874 (.A1(n_257_76_14846), .A2(n_257_76_14847), .ZN(
      n_257_76_14848));
   NAND3_X1 i_257_76_14875 (.A1(n_257_76_14848), .A2(n_257_823), .A3(
      n_257_76_14646), .ZN(n_257_76_14849));
   NAND2_X1 i_257_76_14876 (.A1(n_257_76_14661), .A2(n_257_76_14662), .ZN(
      n_257_76_14850));
   NOR2_X1 i_257_76_14877 (.A1(n_257_76_14849), .A2(n_257_76_14850), .ZN(
      n_257_76_14851));
   NAND2_X1 i_257_76_14878 (.A1(n_257_76_14645), .A2(n_257_76_14851), .ZN(
      n_257_76_14852));
   NOR2_X1 i_257_76_14879 (.A1(n_257_76_14688), .A2(n_257_76_14852), .ZN(
      n_257_76_14853));
   NAND2_X1 i_257_76_14880 (.A1(n_257_22), .A2(n_257_76_14853), .ZN(
      n_257_76_14854));
   NAND2_X1 i_257_76_14881 (.A1(n_257_444), .A2(n_257_76_14647), .ZN(
      n_257_76_14855));
   INV_X1 i_257_76_14882 (.A(n_257_76_14855), .ZN(n_257_76_14856));
   NAND2_X1 i_257_76_14883 (.A1(n_257_1021), .A2(n_257_76_14856), .ZN(
      n_257_76_14857));
   INV_X1 i_257_76_14884 (.A(n_257_76_14857), .ZN(n_257_76_14858));
   NAND2_X1 i_257_76_14885 (.A1(n_257_76_14654), .A2(n_257_76_14858), .ZN(
      n_257_76_14859));
   INV_X1 i_257_76_14886 (.A(n_257_76_14859), .ZN(n_257_76_14860));
   NAND2_X1 i_257_76_14887 (.A1(n_257_76_18075), .A2(n_257_76_14860), .ZN(
      n_257_76_14861));
   NAND2_X1 i_257_76_14888 (.A1(n_257_76_14854), .A2(n_257_76_14861), .ZN(
      n_257_76_14862));
   NOR2_X1 i_257_76_14889 (.A1(n_257_76_14845), .A2(n_257_76_14862), .ZN(
      n_257_76_14863));
   NAND3_X1 i_257_76_14890 (.A1(n_257_76_14761), .A2(n_257_76_14811), .A3(
      n_257_76_14863), .ZN(n_257_76_14864));
   INV_X1 i_257_76_14891 (.A(n_257_76_14864), .ZN(n_257_76_14865));
   NAND2_X1 i_257_76_14892 (.A1(n_257_76_14669), .A2(n_257_76_14673), .ZN(
      n_257_76_14866));
   INV_X1 i_257_76_14893 (.A(n_257_76_14866), .ZN(n_257_76_14867));
   NOR2_X1 i_257_76_14894 (.A1(n_257_1085), .A2(n_257_76_17633), .ZN(
      n_257_76_14868));
   NAND4_X1 i_257_76_14895 (.A1(n_257_61), .A2(n_257_76_14674), .A3(
      n_257_76_14679), .A4(n_257_76_14868), .ZN(n_257_76_14869));
   INV_X1 i_257_76_14896 (.A(n_257_76_14869), .ZN(n_257_76_14870));
   NAND3_X1 i_257_76_14897 (.A1(n_257_76_14668), .A2(n_257_76_14867), .A3(
      n_257_76_14870), .ZN(n_257_76_14871));
   NOR2_X1 i_257_76_14898 (.A1(n_257_76_14685), .A2(n_257_76_14871), .ZN(
      n_257_76_14872));
   NAND4_X1 i_257_76_14899 (.A1(n_257_76_14658), .A2(n_257_76_14645), .A3(
      n_257_76_14664), .A4(n_257_76_14872), .ZN(n_257_76_14873));
   NOR2_X1 i_257_76_14900 (.A1(n_257_76_14873), .A2(n_257_76_14688), .ZN(
      n_257_76_14874));
   NAND2_X1 i_257_76_14901 (.A1(n_257_76_18081), .A2(n_257_76_14874), .ZN(
      n_257_76_14875));
   NAND3_X1 i_257_76_14902 (.A1(n_257_101), .A2(n_257_76_14646), .A3(
      n_257_76_14683), .ZN(n_257_76_14876));
   NAND2_X1 i_257_76_14903 (.A1(n_257_76_14734), .A2(n_257_76_17932), .ZN(
      n_257_76_14877));
   NOR2_X1 i_257_76_14904 (.A1(n_257_76_14877), .A2(n_257_1085), .ZN(
      n_257_76_14878));
   NAND4_X1 i_257_76_14905 (.A1(n_257_76_14673), .A2(n_257_76_14878), .A3(
      n_257_76_14674), .A4(n_257_76_14679), .ZN(n_257_76_14879));
   INV_X1 i_257_76_14906 (.A(n_257_76_14879), .ZN(n_257_76_14880));
   NAND4_X1 i_257_76_14907 (.A1(n_257_76_14880), .A2(n_257_76_14668), .A3(
      n_257_76_14672), .A4(n_257_76_14684), .ZN(n_257_76_14881));
   NOR2_X1 i_257_76_14908 (.A1(n_257_76_14876), .A2(n_257_76_14881), .ZN(
      n_257_76_14882));
   NAND4_X1 i_257_76_14909 (.A1(n_257_76_14882), .A2(n_257_76_14658), .A3(
      n_257_76_14664), .A4(n_257_76_14645), .ZN(n_257_76_14883));
   NOR2_X1 i_257_76_14910 (.A1(n_257_76_14883), .A2(n_257_76_14688), .ZN(
      n_257_76_14884));
   NAND2_X1 i_257_76_14911 (.A1(n_257_76_18080), .A2(n_257_76_14884), .ZN(
      n_257_76_14885));
   INV_X1 i_257_76_14912 (.A(n_257_76_14778), .ZN(n_257_76_14886));
   NAND2_X1 i_257_76_14913 (.A1(n_257_76_17331), .A2(n_257_76_14734), .ZN(
      n_257_76_14887));
   NOR2_X1 i_257_76_14914 (.A1(n_257_76_14887), .A2(n_257_1085), .ZN(
      n_257_76_14888));
   NAND4_X1 i_257_76_14915 (.A1(n_257_76_14692), .A2(n_257_76_14670), .A3(
      n_257_76_14673), .A4(n_257_76_14888), .ZN(n_257_76_14889));
   NOR2_X1 i_257_76_14916 (.A1(n_257_76_14889), .A2(n_257_76_14698), .ZN(
      n_257_76_14890));
   NAND4_X1 i_257_76_14917 (.A1(n_257_76_14886), .A2(n_257_76_14890), .A3(
      n_257_76_14661), .A4(n_257_76_14662), .ZN(n_257_76_14891));
   NAND4_X1 i_257_76_14918 (.A1(n_257_76_14754), .A2(n_257_178), .A3(
      n_257_76_14659), .A4(n_257_76_14660), .ZN(n_257_76_14892));
   NOR2_X1 i_257_76_14919 (.A1(n_257_76_14891), .A2(n_257_76_14892), .ZN(
      n_257_76_14893));
   NAND3_X1 i_257_76_14920 (.A1(n_257_76_14893), .A2(n_257_76_14751), .A3(
      n_257_76_14654), .ZN(n_257_76_14894));
   INV_X1 i_257_76_14921 (.A(n_257_76_14894), .ZN(n_257_76_14895));
   NAND2_X1 i_257_76_14922 (.A1(n_257_76_18061), .A2(n_257_76_14895), .ZN(
      n_257_76_14896));
   NAND3_X1 i_257_76_14923 (.A1(n_257_76_14875), .A2(n_257_76_14885), .A3(
      n_257_76_14896), .ZN(n_257_76_14897));
   INV_X1 i_257_76_14924 (.A(n_257_76_14897), .ZN(n_257_76_14898));
   NAND2_X1 i_257_76_14925 (.A1(n_257_442), .A2(n_257_893), .ZN(n_257_76_14899));
   NOR2_X1 i_257_76_14926 (.A1(n_257_1085), .A2(n_257_76_14899), .ZN(
      n_257_76_14900));
   NAND3_X1 i_257_76_14927 (.A1(n_257_76_14674), .A2(n_257_438), .A3(
      n_257_76_14900), .ZN(n_257_76_14901));
   INV_X1 i_257_76_14928 (.A(n_257_76_14901), .ZN(n_257_76_14902));
   NAND2_X1 i_257_76_14929 (.A1(n_257_76_14646), .A2(n_257_76_14902), .ZN(
      n_257_76_14903));
   NOR2_X1 i_257_76_14930 (.A1(n_257_76_14803), .A2(n_257_76_14903), .ZN(
      n_257_76_14904));
   NAND2_X1 i_257_76_14931 (.A1(n_257_76_14645), .A2(n_257_76_14904), .ZN(
      n_257_76_14905));
   INV_X1 i_257_76_14932 (.A(n_257_76_14905), .ZN(n_257_76_14906));
   NAND2_X1 i_257_76_14933 (.A1(n_257_76_14906), .A2(n_257_76_14654), .ZN(
      n_257_76_14907));
   INV_X1 i_257_76_14934 (.A(n_257_76_14907), .ZN(n_257_76_14908));
   NAND2_X1 i_257_76_14935 (.A1(n_257_76_18067), .A2(n_257_76_14908), .ZN(
      n_257_76_14909));
   NAND2_X1 i_257_76_14936 (.A1(n_257_76_14673), .A2(n_257_76_14737), .ZN(
      n_257_76_14910));
   INV_X1 i_257_76_14937 (.A(n_257_76_14670), .ZN(n_257_76_14911));
   NOR2_X1 i_257_76_14938 (.A1(n_257_76_14910), .A2(n_257_76_14911), .ZN(
      n_257_76_14912));
   NAND2_X1 i_257_76_14939 (.A1(n_257_442), .A2(n_257_495), .ZN(n_257_76_14913));
   NAND2_X1 i_257_76_14940 (.A1(n_257_76_14733), .A2(n_257_76_17991), .ZN(
      n_257_76_14914));
   NAND2_X1 i_257_76_14941 (.A1(n_257_420), .A2(n_257_76_14734), .ZN(
      n_257_76_14915));
   NOR2_X1 i_257_76_14942 (.A1(n_257_76_14914), .A2(n_257_76_14915), .ZN(
      n_257_76_14916));
   NAND2_X1 i_257_76_14943 (.A1(n_257_76_14916), .A2(n_257_76_14679), .ZN(
      n_257_76_14917));
   NAND2_X1 i_257_76_14944 (.A1(n_257_336), .A2(n_257_422), .ZN(n_257_76_14918));
   NAND2_X1 i_257_76_14945 (.A1(n_257_76_14918), .A2(n_257_76_14674), .ZN(
      n_257_76_14919));
   NOR2_X1 i_257_76_14946 (.A1(n_257_76_14917), .A2(n_257_76_14919), .ZN(
      n_257_76_14920));
   NAND2_X1 i_257_76_14947 (.A1(n_257_76_14912), .A2(n_257_76_14920), .ZN(
      n_257_76_14921));
   NAND2_X1 i_257_76_14948 (.A1(n_257_76_14728), .A2(n_257_76_14665), .ZN(
      n_257_76_14922));
   INV_X1 i_257_76_14949 (.A(n_257_76_14922), .ZN(n_257_76_14923));
   NAND2_X1 i_257_76_14950 (.A1(n_257_76_14666), .A2(n_257_76_14669), .ZN(
      n_257_76_14924));
   INV_X1 i_257_76_14951 (.A(n_257_76_14924), .ZN(n_257_76_14925));
   NAND2_X1 i_257_76_14952 (.A1(n_257_76_14923), .A2(n_257_76_14925), .ZN(
      n_257_76_14926));
   NOR2_X1 i_257_76_14953 (.A1(n_257_76_14921), .A2(n_257_76_14926), .ZN(
      n_257_76_14927));
   NAND2_X1 i_257_76_14954 (.A1(n_257_76_14646), .A2(n_257_76_14683), .ZN(
      n_257_76_14928));
   NAND2_X1 i_257_76_14955 (.A1(n_257_76_14741), .A2(n_257_76_14684), .ZN(
      n_257_76_14929));
   NOR2_X1 i_257_76_14956 (.A1(n_257_76_14928), .A2(n_257_76_14929), .ZN(
      n_257_76_14930));
   NAND2_X1 i_257_76_14957 (.A1(n_257_76_14927), .A2(n_257_76_14930), .ZN(
      n_257_76_14931));
   NAND2_X1 i_257_76_14958 (.A1(n_257_375), .A2(n_257_421), .ZN(n_257_76_14932));
   NAND2_X1 i_257_76_14959 (.A1(n_257_76_14745), .A2(n_257_76_14932), .ZN(
      n_257_76_14933));
   NOR2_X1 i_257_76_14960 (.A1(n_257_76_14933), .A2(n_257_76_14803), .ZN(
      n_257_76_14934));
   NAND2_X1 i_257_76_14961 (.A1(n_257_298), .A2(n_257_423), .ZN(n_257_76_14935));
   NAND2_X1 i_257_76_14962 (.A1(n_257_76_14935), .A2(n_257_76_14661), .ZN(
      n_257_76_14936));
   INV_X1 i_257_76_14963 (.A(n_257_76_14936), .ZN(n_257_76_14937));
   NAND2_X1 i_257_76_14964 (.A1(n_257_76_14934), .A2(n_257_76_14937), .ZN(
      n_257_76_14938));
   NOR2_X1 i_257_76_14965 (.A1(n_257_76_14931), .A2(n_257_76_14938), .ZN(
      n_257_76_14939));
   NAND2_X1 i_257_76_14966 (.A1(n_257_76_14832), .A2(n_257_76_14754), .ZN(
      n_257_76_14940));
   NAND2_X1 i_257_76_14967 (.A1(n_257_76_14752), .A2(n_257_76_14753), .ZN(
      n_257_76_14941));
   NOR2_X1 i_257_76_14968 (.A1(n_257_76_14940), .A2(n_257_76_14941), .ZN(
      n_257_76_14942));
   NAND2_X1 i_257_76_14969 (.A1(n_257_76_14939), .A2(n_257_76_14942), .ZN(
      n_257_76_14943));
   NAND2_X1 i_257_76_14970 (.A1(n_257_76_14751), .A2(n_257_76_14654), .ZN(
      n_257_76_14944));
   NOR2_X1 i_257_76_14971 (.A1(n_257_76_14943), .A2(n_257_76_14944), .ZN(
      n_257_76_14945));
   NAND2_X1 i_257_76_14972 (.A1(n_257_76_18073), .A2(n_257_76_14945), .ZN(
      n_257_76_14946));
   NAND4_X1 i_257_76_14973 (.A1(n_257_139), .A2(n_257_76_14665), .A3(
      n_257_76_14666), .A4(n_257_76_14669), .ZN(n_257_76_14947));
   NAND2_X1 i_257_76_14974 (.A1(n_257_76_14734), .A2(n_257_76_17925), .ZN(
      n_257_76_14948));
   NOR2_X1 i_257_76_14975 (.A1(n_257_76_14948), .A2(n_257_1085), .ZN(
      n_257_76_14949));
   NAND2_X1 i_257_76_14976 (.A1(n_257_76_14679), .A2(n_257_76_14949), .ZN(
      n_257_76_14950));
   INV_X1 i_257_76_14977 (.A(n_257_76_14950), .ZN(n_257_76_14951));
   NAND4_X1 i_257_76_14978 (.A1(n_257_76_14951), .A2(n_257_76_14670), .A3(
      n_257_76_14673), .A4(n_257_76_14674), .ZN(n_257_76_14952));
   NOR2_X1 i_257_76_14979 (.A1(n_257_76_14947), .A2(n_257_76_14952), .ZN(
      n_257_76_14953));
   INV_X1 i_257_76_14980 (.A(n_257_76_14685), .ZN(n_257_76_14954));
   NAND3_X1 i_257_76_14981 (.A1(n_257_76_14953), .A2(n_257_76_14954), .A3(
      n_257_76_14662), .ZN(n_257_76_14955));
   NAND4_X1 i_257_76_14982 (.A1(n_257_76_14754), .A2(n_257_76_14659), .A3(
      n_257_76_14660), .A4(n_257_76_14661), .ZN(n_257_76_14956));
   NOR2_X1 i_257_76_14983 (.A1(n_257_76_14955), .A2(n_257_76_14956), .ZN(
      n_257_76_14957));
   NAND4_X1 i_257_76_14984 (.A1(n_257_76_14957), .A2(n_257_76_14654), .A3(
      n_257_76_14658), .A4(n_257_76_14645), .ZN(n_257_76_14958));
   INV_X1 i_257_76_14985 (.A(n_257_76_14958), .ZN(n_257_76_14959));
   NAND2_X1 i_257_76_14986 (.A1(n_257_76_18068), .A2(n_257_76_14959), .ZN(
      n_257_76_14960));
   NAND3_X1 i_257_76_14987 (.A1(n_257_76_14909), .A2(n_257_76_14946), .A3(
      n_257_76_14960), .ZN(n_257_76_14961));
   INV_X1 i_257_76_14988 (.A(n_257_76_14961), .ZN(n_257_76_14962));
   INV_X1 i_257_76_14989 (.A(n_257_76_14646), .ZN(n_257_76_14963));
   NAND2_X1 i_257_76_14990 (.A1(n_257_447), .A2(n_257_76_14674), .ZN(
      n_257_76_14964));
   INV_X1 i_257_76_14991 (.A(n_257_76_14964), .ZN(n_257_76_14965));
   NAND2_X1 i_257_76_14992 (.A1(n_257_791), .A2(n_257_442), .ZN(n_257_76_14966));
   NOR2_X1 i_257_76_14993 (.A1(n_257_1085), .A2(n_257_76_14966), .ZN(
      n_257_76_14967));
   NAND2_X1 i_257_76_14994 (.A1(n_257_76_14679), .A2(n_257_76_14967), .ZN(
      n_257_76_14968));
   INV_X1 i_257_76_14995 (.A(n_257_76_14968), .ZN(n_257_76_14969));
   NAND3_X1 i_257_76_14996 (.A1(n_257_76_14965), .A2(n_257_76_14969), .A3(
      n_257_76_14665), .ZN(n_257_76_14970));
   NOR2_X1 i_257_76_14997 (.A1(n_257_76_14963), .A2(n_257_76_14970), .ZN(
      n_257_76_14971));
   NAND4_X1 i_257_76_14998 (.A1(n_257_76_14971), .A2(n_257_76_14659), .A3(
      n_257_76_14661), .A4(n_257_76_14662), .ZN(n_257_76_14972));
   INV_X1 i_257_76_14999 (.A(n_257_76_14972), .ZN(n_257_76_14973));
   NAND2_X1 i_257_76_15000 (.A1(n_257_76_14645), .A2(n_257_76_14973), .ZN(
      n_257_76_14974));
   NOR2_X1 i_257_76_15001 (.A1(n_257_76_14974), .A2(n_257_76_14688), .ZN(
      n_257_76_14975));
   NAND3_X1 i_257_76_15002 (.A1(n_257_76_14665), .A2(n_257_76_14669), .A3(
      n_257_76_14673), .ZN(n_257_76_14976));
   NAND2_X1 i_257_76_15003 (.A1(n_257_442), .A2(n_257_663), .ZN(n_257_76_14977));
   NOR2_X1 i_257_76_15004 (.A1(n_257_1085), .A2(n_257_76_14977), .ZN(
      n_257_76_14978));
   NAND4_X1 i_257_76_15005 (.A1(n_257_449), .A2(n_257_76_14674), .A3(
      n_257_76_14679), .A4(n_257_76_14978), .ZN(n_257_76_14979));
   NOR2_X1 i_257_76_15006 (.A1(n_257_76_14976), .A2(n_257_76_14979), .ZN(
      n_257_76_14980));
   NAND3_X1 i_257_76_15007 (.A1(n_257_76_14980), .A2(n_257_76_14662), .A3(
      n_257_76_14646), .ZN(n_257_76_14981));
   NOR2_X1 i_257_76_15008 (.A1(n_257_76_14981), .A2(n_257_76_14701), .ZN(
      n_257_76_14982));
   NAND3_X1 i_257_76_15009 (.A1(n_257_76_14982), .A2(n_257_76_14658), .A3(
      n_257_76_14645), .ZN(n_257_76_14983));
   NOR2_X1 i_257_76_15010 (.A1(n_257_76_14983), .A2(n_257_76_14688), .ZN(
      n_257_76_14984));
   AOI22_X1 i_257_76_15011 (.A1(n_257_76_18085), .A2(n_257_76_14975), .B1(
      n_257_76_18083), .B2(n_257_76_14984), .ZN(n_257_76_14985));
   NAND3_X1 i_257_76_15012 (.A1(n_257_76_14898), .A2(n_257_76_14962), .A3(
      n_257_76_14985), .ZN(n_257_76_14986));
   INV_X1 i_257_76_15013 (.A(n_257_727), .ZN(n_257_76_14987));
   NAND2_X1 i_257_76_15014 (.A1(n_257_76_14987), .A2(n_257_76_14647), .ZN(
      n_257_76_14988));
   NAND2_X1 i_257_76_15015 (.A1(n_257_76_14647), .A2(n_257_76_17760), .ZN(
      n_257_76_14989));
   AOI21_X1 i_257_76_15016 (.A(n_257_76_14691), .B1(n_257_76_14988), .B2(
      n_257_76_14989), .ZN(n_257_76_14990));
   NAND3_X1 i_257_76_15017 (.A1(n_257_76_14665), .A2(n_257_76_14669), .A3(
      n_257_448), .ZN(n_257_76_14991));
   INV_X1 i_257_76_15018 (.A(n_257_76_14991), .ZN(n_257_76_14992));
   NAND3_X1 i_257_76_15019 (.A1(n_257_76_14990), .A2(n_257_76_14992), .A3(
      n_257_76_14646), .ZN(n_257_76_14993));
   NOR2_X1 i_257_76_15020 (.A1(n_257_76_14993), .A2(n_257_76_14803), .ZN(
      n_257_76_14994));
   NAND3_X1 i_257_76_15021 (.A1(n_257_76_14994), .A2(n_257_76_14744), .A3(
      n_257_695), .ZN(n_257_76_14995));
   INV_X1 i_257_76_15022 (.A(n_257_76_14995), .ZN(n_257_76_14996));
   NAND3_X1 i_257_76_15023 (.A1(n_257_76_14996), .A2(n_257_76_14654), .A3(
      n_257_76_14645), .ZN(n_257_76_14997));
   INV_X1 i_257_76_15024 (.A(n_257_76_14997), .ZN(n_257_76_14998));
   NAND2_X1 i_257_76_15025 (.A1(n_257_76_18079), .A2(n_257_76_14998), .ZN(
      n_257_76_14999));
   NAND3_X1 i_257_76_15026 (.A1(n_257_76_14654), .A2(n_257_76_14658), .A3(
      n_257_76_14645), .ZN(n_257_76_15000));
   NAND3_X1 i_257_76_15027 (.A1(n_257_76_14754), .A2(n_257_76_14659), .A3(
      n_257_258), .ZN(n_257_76_15001));
   INV_X1 i_257_76_15028 (.A(n_257_76_15001), .ZN(n_257_76_15002));
   NAND4_X1 i_257_76_15029 (.A1(n_257_76_17990), .A2(n_257_76_14733), .A3(
      n_257_76_14734), .A4(n_257_425), .ZN(n_257_76_15003));
   INV_X1 i_257_76_15030 (.A(n_257_76_15003), .ZN(n_257_76_15004));
   NAND4_X1 i_257_76_15031 (.A1(n_257_76_15004), .A2(n_257_76_14737), .A3(
      n_257_76_14674), .A4(n_257_76_14679), .ZN(n_257_76_15005));
   INV_X1 i_257_76_15032 (.A(n_257_76_15005), .ZN(n_257_76_15006));
   NAND3_X1 i_257_76_15033 (.A1(n_257_76_15006), .A2(n_257_76_14732), .A3(
      n_257_76_14668), .ZN(n_257_76_15007));
   NOR2_X1 i_257_76_15034 (.A1(n_257_76_14778), .A2(n_257_76_15007), .ZN(
      n_257_76_15008));
   NAND4_X1 i_257_76_15035 (.A1(n_257_76_14660), .A2(n_257_76_14661), .A3(
      n_257_76_14662), .A4(n_257_76_14745), .ZN(n_257_76_15009));
   INV_X1 i_257_76_15036 (.A(n_257_76_15009), .ZN(n_257_76_15010));
   NAND4_X1 i_257_76_15037 (.A1(n_257_76_15002), .A2(n_257_76_15008), .A3(
      n_257_76_15010), .A4(n_257_76_14752), .ZN(n_257_76_15011));
   NOR2_X1 i_257_76_15038 (.A1(n_257_76_15000), .A2(n_257_76_15011), .ZN(
      n_257_76_15012));
   NAND2_X1 i_257_76_15039 (.A1(n_257_76_18064), .A2(n_257_76_15012), .ZN(
      n_257_76_15013));
   NAND3_X1 i_257_76_15040 (.A1(n_257_76_14737), .A2(n_257_76_14918), .A3(
      n_257_76_14674), .ZN(n_257_76_15014));
   NAND2_X1 i_257_76_15041 (.A1(n_257_76_14734), .A2(n_257_421), .ZN(
      n_257_76_15015));
   NOR2_X1 i_257_76_15042 (.A1(n_257_76_15015), .A2(n_257_1085), .ZN(
      n_257_76_15016));
   NAND3_X1 i_257_76_15043 (.A1(n_257_76_15016), .A2(n_257_76_14679), .A3(
      n_257_76_17990), .ZN(n_257_76_15017));
   NOR2_X1 i_257_76_15044 (.A1(n_257_76_15014), .A2(n_257_76_15017), .ZN(
      n_257_76_15018));
   NAND3_X1 i_257_76_15045 (.A1(n_257_76_15018), .A2(n_257_76_14730), .A3(
      n_257_76_14732), .ZN(n_257_76_15019));
   NAND4_X1 i_257_76_15046 (.A1(n_257_76_14646), .A2(n_257_76_14741), .A3(
      n_257_76_14684), .A4(n_257_375), .ZN(n_257_76_15020));
   NOR2_X1 i_257_76_15047 (.A1(n_257_76_15019), .A2(n_257_76_15020), .ZN(
      n_257_76_15021));
   NAND3_X1 i_257_76_15048 (.A1(n_257_76_14659), .A2(n_257_76_14660), .A3(
      n_257_76_14935), .ZN(n_257_76_15022));
   INV_X1 i_257_76_15049 (.A(n_257_76_15022), .ZN(n_257_76_15023));
   NAND3_X1 i_257_76_15050 (.A1(n_257_76_14661), .A2(n_257_76_14662), .A3(
      n_257_76_14745), .ZN(n_257_76_15024));
   INV_X1 i_257_76_15051 (.A(n_257_76_15024), .ZN(n_257_76_15025));
   NAND3_X1 i_257_76_15052 (.A1(n_257_76_15021), .A2(n_257_76_15023), .A3(
      n_257_76_15025), .ZN(n_257_76_15026));
   INV_X1 i_257_76_15053 (.A(n_257_76_15026), .ZN(n_257_76_15027));
   NAND4_X1 i_257_76_15054 (.A1(n_257_76_15027), .A2(n_257_76_14751), .A3(
      n_257_76_14654), .A4(n_257_76_14756), .ZN(n_257_76_15028));
   INV_X1 i_257_76_15055 (.A(n_257_76_15028), .ZN(n_257_76_15029));
   NAND2_X1 i_257_76_15056 (.A1(n_257_76_18082), .A2(n_257_76_15029), .ZN(
      n_257_76_15030));
   NAND3_X1 i_257_76_15057 (.A1(n_257_76_14999), .A2(n_257_76_15013), .A3(
      n_257_76_15030), .ZN(n_257_76_15031));
   INV_X1 i_257_76_15058 (.A(n_257_76_15031), .ZN(n_257_76_15032));
   NAND3_X1 i_257_76_15059 (.A1(n_257_76_14832), .A2(n_257_76_14752), .A3(
      n_257_76_14754), .ZN(n_257_76_15033));
   INV_X1 i_257_76_15060 (.A(n_257_76_14850), .ZN(n_257_76_15034));
   NAND3_X1 i_257_76_15061 (.A1(n_257_76_14684), .A2(n_257_76_14665), .A3(
      n_257_76_14666), .ZN(n_257_76_15035));
   NAND4_X1 i_257_76_15062 (.A1(n_257_76_14692), .A2(n_257_76_14669), .A3(
      n_257_76_14670), .A4(n_257_76_14673), .ZN(n_257_76_15036));
   NOR2_X1 i_257_76_15063 (.A1(n_257_76_15035), .A2(n_257_76_15036), .ZN(
      n_257_76_15037));
   INV_X1 i_257_76_15064 (.A(n_257_76_17990), .ZN(n_257_76_15038));
   NOR2_X1 i_257_76_15065 (.A1(n_257_76_15038), .A2(n_257_1085), .ZN(
      n_257_76_15039));
   NAND2_X1 i_257_76_15066 (.A1(n_257_427), .A2(n_257_76_14734), .ZN(
      n_257_76_15040));
   INV_X1 i_257_76_15067 (.A(n_257_76_15040), .ZN(n_257_76_15041));
   NAND3_X1 i_257_76_15068 (.A1(n_257_76_15039), .A2(n_257_76_15041), .A3(
      n_257_218), .ZN(n_257_76_15042));
   INV_X1 i_257_76_15069 (.A(n_257_76_15042), .ZN(n_257_76_15043));
   NAND4_X1 i_257_76_15070 (.A1(n_257_76_14646), .A2(n_257_76_15043), .A3(
      n_257_76_14683), .A4(n_257_76_14741), .ZN(n_257_76_15044));
   INV_X1 i_257_76_15071 (.A(n_257_76_15044), .ZN(n_257_76_15045));
   NAND3_X1 i_257_76_15072 (.A1(n_257_76_15034), .A2(n_257_76_15037), .A3(
      n_257_76_15045), .ZN(n_257_76_15046));
   NOR2_X1 i_257_76_15073 (.A1(n_257_76_15033), .A2(n_257_76_15046), .ZN(
      n_257_76_15047));
   NAND3_X1 i_257_76_15074 (.A1(n_257_76_15047), .A2(n_257_76_14751), .A3(
      n_257_76_14654), .ZN(n_257_76_15048));
   INV_X1 i_257_76_15075 (.A(n_257_76_15048), .ZN(n_257_76_15049));
   NAND2_X1 i_257_76_15076 (.A1(n_257_76_18065), .A2(n_257_76_15049), .ZN(
      n_257_76_15050));
   NAND3_X1 i_257_76_15077 (.A1(n_257_76_14990), .A2(n_257_76_14646), .A3(
      n_257_76_14684), .ZN(n_257_76_15051));
   INV_X1 i_257_76_15078 (.A(n_257_76_14683), .ZN(n_257_76_15052));
   NAND2_X1 i_257_76_15079 (.A1(n_257_76_14699), .A2(n_257_76_15052), .ZN(
      n_257_76_15053));
   NOR2_X1 i_257_76_15080 (.A1(n_257_76_15051), .A2(n_257_76_15053), .ZN(
      n_257_76_15054));
   NAND4_X1 i_257_76_15081 (.A1(n_257_76_15054), .A2(n_257_76_14658), .A3(
      n_257_76_14664), .A4(n_257_76_14645), .ZN(n_257_76_15055));
   NOR2_X1 i_257_76_15082 (.A1(n_257_76_15055), .A2(n_257_76_14688), .ZN(
      n_257_76_15056));
   NAND2_X1 i_257_76_15083 (.A1(n_257_76_18063), .A2(n_257_76_15056), .ZN(
      n_257_76_15057));
   NAND4_X1 i_257_76_15084 (.A1(n_257_76_17990), .A2(n_257_76_14733), .A3(
      n_257_76_14734), .A4(n_257_424), .ZN(n_257_76_15058));
   INV_X1 i_257_76_15085 (.A(n_257_76_15058), .ZN(n_257_76_15059));
   NAND4_X1 i_257_76_15086 (.A1(n_257_76_15059), .A2(n_257_527), .A3(
      n_257_76_14674), .A4(n_257_76_14679), .ZN(n_257_76_15060));
   INV_X1 i_257_76_15087 (.A(n_257_76_15060), .ZN(n_257_76_15061));
   NAND3_X1 i_257_76_15088 (.A1(n_257_76_14670), .A2(n_257_76_14673), .A3(
      n_257_76_14737), .ZN(n_257_76_15062));
   INV_X1 i_257_76_15089 (.A(n_257_76_15062), .ZN(n_257_76_15063));
   NAND3_X1 i_257_76_15090 (.A1(n_257_76_15061), .A2(n_257_76_15063), .A3(
      n_257_76_14684), .ZN(n_257_76_15064));
   INV_X1 i_257_76_15091 (.A(n_257_76_15064), .ZN(n_257_76_15065));
   NAND3_X1 i_257_76_15092 (.A1(n_257_76_15065), .A2(n_257_76_14754), .A3(
      n_257_76_14659), .ZN(n_257_76_15066));
   NOR2_X1 i_257_76_15093 (.A1(n_257_76_14941), .A2(n_257_76_15066), .ZN(
      n_257_76_15067));
   INV_X1 i_257_76_15094 (.A(n_257_76_14741), .ZN(n_257_76_15068));
   NOR2_X1 i_257_76_15095 (.A1(n_257_76_15068), .A2(n_257_76_14698), .ZN(
      n_257_76_15069));
   INV_X1 i_257_76_15096 (.A(n_257_76_14928), .ZN(n_257_76_15070));
   NAND3_X1 i_257_76_15097 (.A1(n_257_76_15069), .A2(n_257_76_15070), .A3(
      n_257_76_14745), .ZN(n_257_76_15071));
   NOR2_X1 i_257_76_15098 (.A1(n_257_76_15071), .A2(n_257_76_14789), .ZN(
      n_257_76_15072));
   NAND4_X1 i_257_76_15099 (.A1(n_257_76_15067), .A2(n_257_76_14751), .A3(
      n_257_76_14654), .A4(n_257_76_15072), .ZN(n_257_76_15073));
   INV_X1 i_257_76_15100 (.A(n_257_76_15073), .ZN(n_257_76_15074));
   NAND2_X1 i_257_76_15101 (.A1(n_257_76_18062), .A2(n_257_76_15074), .ZN(
      n_257_76_15075));
   NAND3_X1 i_257_76_15102 (.A1(n_257_76_15050), .A2(n_257_76_15057), .A3(
      n_257_76_15075), .ZN(n_257_76_15076));
   INV_X1 i_257_76_15103 (.A(n_257_76_15076), .ZN(n_257_76_15077));
   NAND4_X1 i_257_76_15104 (.A1(n_257_76_14754), .A2(n_257_76_14659), .A3(
      n_257_76_14660), .A4(n_257_76_14935), .ZN(n_257_76_15078));
   NOR2_X1 i_257_76_15105 (.A1(n_257_76_14941), .A2(n_257_76_15078), .ZN(
      n_257_76_15079));
   NAND2_X1 i_257_76_15106 (.A1(n_257_76_14683), .A2(n_257_76_14741), .ZN(
      n_257_76_15080));
   INV_X1 i_257_76_15107 (.A(n_257_76_15080), .ZN(n_257_76_15081));
   NAND3_X1 i_257_76_15108 (.A1(n_257_76_14666), .A2(n_257_76_14669), .A3(
      n_257_76_14670), .ZN(n_257_76_15082));
   NAND4_X1 i_257_76_15109 (.A1(n_257_76_14673), .A2(n_257_76_14737), .A3(
      n_257_76_14674), .A4(n_257_76_14679), .ZN(n_257_76_15083));
   NOR2_X1 i_257_76_15110 (.A1(n_257_76_15082), .A2(n_257_76_15083), .ZN(
      n_257_76_15084));
   NAND2_X1 i_257_76_15111 (.A1(n_257_76_14734), .A2(n_257_422), .ZN(
      n_257_76_15085));
   INV_X1 i_257_76_15112 (.A(n_257_76_15085), .ZN(n_257_76_15086));
   NAND4_X1 i_257_76_15113 (.A1(n_257_336), .A2(n_257_76_15086), .A3(
      n_257_76_17990), .A4(n_257_76_14733), .ZN(n_257_76_15087));
   INV_X1 i_257_76_15114 (.A(n_257_76_15087), .ZN(n_257_76_15088));
   NAND3_X1 i_257_76_15115 (.A1(n_257_76_15088), .A2(n_257_76_14728), .A3(
      n_257_76_14665), .ZN(n_257_76_15089));
   INV_X1 i_257_76_15116 (.A(n_257_76_14684), .ZN(n_257_76_15090));
   NOR2_X1 i_257_76_15117 (.A1(n_257_76_15089), .A2(n_257_76_15090), .ZN(
      n_257_76_15091));
   NAND3_X1 i_257_76_15118 (.A1(n_257_76_15081), .A2(n_257_76_15084), .A3(
      n_257_76_15091), .ZN(n_257_76_15092));
   NAND4_X1 i_257_76_15119 (.A1(n_257_76_14661), .A2(n_257_76_14662), .A3(
      n_257_76_14745), .A4(n_257_76_14646), .ZN(n_257_76_15093));
   NOR2_X1 i_257_76_15120 (.A1(n_257_76_15092), .A2(n_257_76_15093), .ZN(
      n_257_76_15094));
   NAND4_X1 i_257_76_15121 (.A1(n_257_76_15079), .A2(n_257_76_14751), .A3(
      n_257_76_15094), .A4(n_257_76_14654), .ZN(n_257_76_15095));
   INV_X1 i_257_76_15122 (.A(n_257_76_15095), .ZN(n_257_76_15096));
   NAND2_X1 i_257_76_15123 (.A1(n_257_342), .A2(n_257_76_15096), .ZN(
      n_257_76_15097));
   NAND2_X1 i_257_76_15124 (.A1(n_257_695), .A2(n_257_76_17958), .ZN(
      n_257_76_15098));
   NAND2_X1 i_257_76_15125 (.A1(n_257_1021), .A2(n_257_76_17964), .ZN(
      n_257_76_15099));
   NAND2_X1 i_257_76_15126 (.A1(n_257_178), .A2(n_257_76_17331), .ZN(
      n_257_76_15100));
   NAND3_X1 i_257_76_15127 (.A1(n_257_76_15098), .A2(n_257_76_15099), .A3(
      n_257_76_15100), .ZN(n_257_76_15101));
   INV_X1 i_257_76_15128 (.A(n_257_76_15101), .ZN(n_257_76_15102));
   NAND2_X1 i_257_76_15129 (.A1(n_257_727), .A2(n_257_76_15655), .ZN(
      n_257_76_15103));
   NAND2_X1 i_257_76_15130 (.A1(n_257_76_15087), .A2(n_257_76_15103), .ZN(
      n_257_76_15104));
   NAND2_X1 i_257_76_15131 (.A1(n_257_957), .A2(n_257_442), .ZN(n_257_76_15105));
   INV_X1 i_257_76_15132 (.A(n_257_76_15105), .ZN(n_257_76_15106));
   NAND2_X1 i_257_76_15133 (.A1(n_257_440), .A2(n_257_76_15106), .ZN(
      n_257_76_15107));
   INV_X1 i_257_76_15134 (.A(n_257_76_14899), .ZN(n_257_76_15108));
   NAND2_X1 i_257_76_15135 (.A1(n_257_438), .A2(n_257_76_15108), .ZN(
      n_257_76_15109));
   NAND3_X1 i_257_76_15136 (.A1(n_257_76_15107), .A2(n_257_76_15109), .A3(
      n_257_76_14677), .ZN(n_257_76_15110));
   NOR2_X1 i_257_76_15137 (.A1(n_257_76_15104), .A2(n_257_76_15110), .ZN(
      n_257_76_15111));
   NAND2_X1 i_257_76_15138 (.A1(n_257_591), .A2(n_257_428), .ZN(n_257_76_15112));
   INV_X1 i_257_76_15139 (.A(Small_Packet_Data_Size[26]), .ZN(n_257_76_15113));
   NAND2_X1 i_257_76_15140 (.A1(n_257_76_15112), .A2(n_257_76_17992), .ZN(
      n_257_76_15114));
   INV_X1 i_257_76_15141 (.A(n_257_76_15114), .ZN(n_257_76_15115));
   NAND2_X1 i_257_76_15142 (.A1(n_257_420), .A2(n_257_495), .ZN(n_257_76_15116));
   NAND3_X1 i_257_76_15143 (.A1(n_257_76_15115), .A2(n_257_76_15116), .A3(
      n_257_76_14733), .ZN(n_257_76_15117));
   NAND2_X1 i_257_76_15144 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[26]), 
      .ZN(n_257_76_15118));
   NAND2_X1 i_257_76_15145 (.A1(n_257_76_15117), .A2(n_257_76_15118), .ZN(
      n_257_76_15119));
   NAND2_X1 i_257_76_15146 (.A1(n_257_855), .A2(n_257_442), .ZN(n_257_76_15120));
   INV_X1 i_257_76_15147 (.A(n_257_76_15120), .ZN(n_257_76_15121));
   NAND2_X1 i_257_76_15148 (.A1(n_257_446), .A2(n_257_76_15121), .ZN(
      n_257_76_15122));
   NAND3_X1 i_257_76_15149 (.A1(n_257_76_15119), .A2(n_257_76_15042), .A3(
      n_257_76_15122), .ZN(n_257_76_15123));
   INV_X1 i_257_76_15150 (.A(n_257_76_15123), .ZN(n_257_76_15124));
   INV_X1 i_257_76_15151 (.A(n_257_76_14977), .ZN(n_257_76_15125));
   NAND2_X1 i_257_76_15152 (.A1(n_257_449), .A2(n_257_76_15125), .ZN(
      n_257_76_15126));
   INV_X1 i_257_76_15153 (.A(n_257_76_14966), .ZN(n_257_76_15127));
   NAND2_X1 i_257_76_15154 (.A1(n_257_447), .A2(n_257_76_15127), .ZN(
      n_257_76_15128));
   NAND2_X1 i_257_76_15155 (.A1(n_257_61), .A2(n_257_76_17918), .ZN(
      n_257_76_15129));
   NAND3_X1 i_257_76_15156 (.A1(n_257_76_15126), .A2(n_257_76_15128), .A3(
      n_257_76_15129), .ZN(n_257_76_15130));
   INV_X1 i_257_76_15157 (.A(n_257_76_15130), .ZN(n_257_76_15131));
   NAND3_X1 i_257_76_15158 (.A1(n_257_76_15111), .A2(n_257_76_15124), .A3(
      n_257_76_15131), .ZN(n_257_76_15132));
   NAND3_X1 i_257_76_15159 (.A1(n_257_989), .A2(n_257_441), .A3(n_257_442), 
      .ZN(n_257_76_15133));
   NAND3_X1 i_257_76_15160 (.A1(n_257_451), .A2(n_257_478), .A3(n_257_442), 
      .ZN(n_257_76_15134));
   NAND2_X1 i_257_76_15161 (.A1(n_257_139), .A2(n_257_76_17925), .ZN(
      n_257_76_15135));
   NAND2_X1 i_257_76_15162 (.A1(n_257_655), .A2(n_257_76_17928), .ZN(
      n_257_76_15136));
   NAND4_X1 i_257_76_15163 (.A1(n_257_76_15133), .A2(n_257_76_15134), .A3(
      n_257_76_15135), .A4(n_257_76_15136), .ZN(n_257_76_15137));
   NOR2_X1 i_257_76_15164 (.A1(n_257_76_15132), .A2(n_257_76_15137), .ZN(
      n_257_76_15138));
   NAND2_X1 i_257_76_15165 (.A1(n_257_101), .A2(n_257_76_17932), .ZN(
      n_257_76_15139));
   NAND2_X1 i_257_76_15166 (.A1(n_257_823), .A2(n_257_76_17952), .ZN(
      n_257_76_15140));
   NAND3_X1 i_257_76_15167 (.A1(n_257_76_15139), .A2(n_257_76_15064), .A3(
      n_257_76_15140), .ZN(n_257_76_15141));
   INV_X1 i_257_76_15168 (.A(n_257_76_15141), .ZN(n_257_76_15142));
   NAND2_X1 i_257_76_15169 (.A1(n_257_759), .A2(n_257_76_17935), .ZN(
      n_257_76_15143));
   NAND2_X1 i_257_76_15170 (.A1(n_257_887), .A2(n_257_76_17903), .ZN(
      n_257_76_15144));
   NAND2_X1 i_257_76_15171 (.A1(n_257_925), .A2(n_257_76_17940), .ZN(
      n_257_76_15145));
   NAND3_X1 i_257_76_15172 (.A1(n_257_76_15143), .A2(n_257_76_15144), .A3(
      n_257_76_15145), .ZN(n_257_76_15146));
   INV_X1 i_257_76_15173 (.A(n_257_76_15146), .ZN(n_257_76_15147));
   NAND3_X1 i_257_76_15174 (.A1(n_257_76_15138), .A2(n_257_76_15142), .A3(
      n_257_76_15147), .ZN(n_257_76_15148));
   INV_X1 i_257_76_15175 (.A(n_257_76_15148), .ZN(n_257_76_15149));
   NAND2_X1 i_257_76_15176 (.A1(n_257_76_15102), .A2(n_257_76_15149), .ZN(
      n_257_76_15150));
   NAND2_X1 i_257_76_15177 (.A1(n_257_1053), .A2(n_257_76_17969), .ZN(
      n_257_76_15151));
   NAND3_X1 i_257_76_15178 (.A1(n_257_76_15151), .A2(n_257_76_14748), .A3(
      n_257_76_14833), .ZN(n_257_76_15152));
   NAND2_X1 i_257_76_15179 (.A1(n_257_76_15011), .A2(n_257_76_15026), .ZN(
      n_257_76_15153));
   NOR3_X1 i_257_76_15180 (.A1(n_257_76_15150), .A2(n_257_76_15152), .A3(
      n_257_76_15153), .ZN(n_257_76_15154));
   NAND3_X1 i_257_76_15181 (.A1(n_257_414), .A2(n_257_484), .A3(n_257_442), 
      .ZN(n_257_76_15155));
   INV_X1 i_257_76_15182 (.A(n_257_76_15155), .ZN(n_257_76_15156));
   NAND2_X1 i_257_76_15183 (.A1(n_257_76_15112), .A2(n_257_76_15156), .ZN(
      n_257_76_15157));
   INV_X1 i_257_76_15184 (.A(n_257_76_15157), .ZN(n_257_76_15158));
   NAND4_X1 i_257_76_15185 (.A1(n_257_76_15116), .A2(n_257_76_15158), .A3(
      n_257_76_14733), .A4(n_257_76_14734), .ZN(n_257_76_15159));
   NOR2_X1 i_257_76_15186 (.A1(n_257_76_14691), .A2(n_257_76_15159), .ZN(
      n_257_76_15160));
   NAND3_X1 i_257_76_15187 (.A1(n_257_76_14673), .A2(n_257_76_14737), .A3(
      n_257_76_14918), .ZN(n_257_76_15161));
   INV_X1 i_257_76_15188 (.A(n_257_76_15161), .ZN(n_257_76_15162));
   NAND3_X1 i_257_76_15189 (.A1(n_257_76_15160), .A2(n_257_76_14672), .A3(
      n_257_76_15162), .ZN(n_257_76_15163));
   NAND4_X1 i_257_76_15190 (.A1(n_257_76_14684), .A2(n_257_76_14728), .A3(
      n_257_76_14665), .A4(n_257_76_14666), .ZN(n_257_76_15164));
   NOR2_X1 i_257_76_15191 (.A1(n_257_76_15163), .A2(n_257_76_15164), .ZN(
      n_257_76_15165));
   NAND4_X1 i_257_76_15192 (.A1(n_257_76_15165), .A2(n_257_76_14752), .A3(
      n_257_76_14753), .A4(n_257_76_14754), .ZN(n_257_76_15166));
   INV_X1 i_257_76_15193 (.A(n_257_76_15166), .ZN(n_257_76_15167));
   NAND2_X1 i_257_76_15194 (.A1(n_257_76_14932), .A2(n_257_76_14646), .ZN(
      n_257_76_15168));
   INV_X1 i_257_76_15195 (.A(n_257_76_15168), .ZN(n_257_76_15169));
   NAND4_X1 i_257_76_15196 (.A1(n_257_76_15169), .A2(n_257_76_15081), .A3(
      n_257_76_14662), .A4(n_257_76_14745), .ZN(n_257_76_15170));
   NAND4_X1 i_257_76_15197 (.A1(n_257_76_14659), .A2(n_257_76_14660), .A3(
      n_257_76_14935), .A4(n_257_76_14661), .ZN(n_257_76_15171));
   NOR2_X1 i_257_76_15198 (.A1(n_257_76_15170), .A2(n_257_76_15171), .ZN(
      n_257_76_15172));
   NAND4_X1 i_257_76_15199 (.A1(n_257_76_14751), .A2(n_257_76_15167), .A3(
      n_257_76_15172), .A4(n_257_76_14654), .ZN(n_257_76_15173));
   INV_X1 i_257_76_15200 (.A(n_257_76_15173), .ZN(n_257_76_15174));
   AOI21_X1 i_257_76_15201 (.A(n_257_76_15154), .B1(n_257_76_18060), .B2(
      n_257_76_15174), .ZN(n_257_76_15175));
   NAND2_X1 i_257_76_15202 (.A1(n_257_76_15097), .A2(n_257_76_15175), .ZN(
      n_257_76_15176));
   INV_X1 i_257_76_15203 (.A(n_257_76_15176), .ZN(n_257_76_15177));
   NAND3_X1 i_257_76_15204 (.A1(n_257_76_15032), .A2(n_257_76_15077), .A3(
      n_257_76_15177), .ZN(n_257_76_15178));
   NOR2_X1 i_257_76_15205 (.A1(n_257_76_14986), .A2(n_257_76_15178), .ZN(
      n_257_76_15179));
   NAND2_X1 i_257_76_15206 (.A1(n_257_76_14865), .A2(n_257_76_15179), .ZN(n_26));
   NAND2_X1 i_257_76_15207 (.A1(n_257_1022), .A2(n_257_444), .ZN(n_257_76_15180));
   NAND2_X1 i_257_76_15208 (.A1(n_257_990), .A2(n_257_441), .ZN(n_257_76_15181));
   INV_X1 i_257_76_15209 (.A(n_257_1086), .ZN(n_257_76_15182));
   NAND2_X1 i_257_76_15210 (.A1(n_257_958), .A2(n_257_442), .ZN(n_257_76_15183));
   INV_X1 i_257_76_15211 (.A(n_257_76_15183), .ZN(n_257_76_15184));
   NAND3_X1 i_257_76_15212 (.A1(n_257_440), .A2(n_257_76_15182), .A3(
      n_257_76_15184), .ZN(n_257_76_15185));
   INV_X1 i_257_76_15213 (.A(n_257_76_15185), .ZN(n_257_76_15186));
   NAND2_X1 i_257_76_15214 (.A1(n_257_76_15181), .A2(n_257_76_15186), .ZN(
      n_257_76_15187));
   INV_X1 i_257_76_15215 (.A(n_257_76_15187), .ZN(n_257_76_15188));
   NAND2_X1 i_257_76_15216 (.A1(n_257_76_15180), .A2(n_257_76_15188), .ZN(
      n_257_76_15189));
   INV_X1 i_257_76_15217 (.A(n_257_76_15189), .ZN(n_257_76_15190));
   NAND2_X1 i_257_76_15218 (.A1(n_257_1054), .A2(n_257_443), .ZN(n_257_76_15191));
   NAND2_X1 i_257_76_15219 (.A1(n_257_76_15190), .A2(n_257_76_15191), .ZN(
      n_257_76_15192));
   INV_X1 i_257_76_15220 (.A(n_257_76_15192), .ZN(n_257_76_15193));
   NAND2_X1 i_257_76_15221 (.A1(n_257_17), .A2(n_257_76_15193), .ZN(
      n_257_76_15194));
   NOR2_X1 i_257_76_15222 (.A1(n_257_1086), .A2(n_257_76_17412), .ZN(
      n_257_76_15195));
   INV_X1 i_257_76_15223 (.A(n_257_76_15195), .ZN(n_257_76_15196));
   INV_X1 i_257_76_15224 (.A(n_257_443), .ZN(n_257_76_15197));
   NOR2_X1 i_257_76_15225 (.A1(n_257_76_15196), .A2(n_257_76_15197), .ZN(
      n_257_76_15198));
   NAND2_X1 i_257_76_15226 (.A1(n_257_1054), .A2(n_257_76_15198), .ZN(
      n_257_76_15199));
   INV_X1 i_257_76_15227 (.A(n_257_76_15199), .ZN(n_257_76_15200));
   NAND2_X1 i_257_76_15228 (.A1(n_257_76_18072), .A2(n_257_76_15200), .ZN(
      n_257_76_15201));
   NAND2_X1 i_257_76_15229 (.A1(n_257_728), .A2(n_257_435), .ZN(n_257_76_15202));
   NAND2_X1 i_257_76_15230 (.A1(n_257_656), .A2(n_257_76_15202), .ZN(
      n_257_76_15203));
   NAND2_X1 i_257_76_15231 (.A1(n_257_440), .A2(n_257_958), .ZN(n_257_76_15204));
   NAND2_X1 i_257_76_15232 (.A1(n_257_438), .A2(n_257_894), .ZN(n_257_76_15205));
   NOR2_X1 i_257_76_15233 (.A1(n_257_1086), .A2(n_257_76_17927), .ZN(
      n_257_76_15206));
   NAND3_X1 i_257_76_15234 (.A1(n_257_76_15204), .A2(n_257_76_15205), .A3(
      n_257_76_15206), .ZN(n_257_76_15207));
   NOR2_X1 i_257_76_15235 (.A1(n_257_76_15203), .A2(n_257_76_15207), .ZN(
      n_257_76_15208));
   NAND2_X1 i_257_76_15236 (.A1(n_257_888), .A2(n_257_445), .ZN(n_257_76_15209));
   NAND2_X1 i_257_76_15237 (.A1(n_257_446), .A2(n_257_856), .ZN(n_257_76_15210));
   NAND2_X1 i_257_76_15238 (.A1(n_257_449), .A2(n_257_664), .ZN(n_257_76_15211));
   NAND2_X1 i_257_76_15239 (.A1(n_257_447), .A2(n_257_792), .ZN(n_257_76_15212));
   NAND3_X1 i_257_76_15240 (.A1(n_257_76_15210), .A2(n_257_76_15211), .A3(
      n_257_76_15212), .ZN(n_257_76_15213));
   INV_X1 i_257_76_15241 (.A(n_257_76_15213), .ZN(n_257_76_15214));
   NAND4_X1 i_257_76_15242 (.A1(n_257_76_15208), .A2(n_257_76_15209), .A3(
      n_257_76_15214), .A4(n_257_76_15181), .ZN(n_257_76_15215));
   NAND2_X1 i_257_76_15243 (.A1(n_257_760), .A2(n_257_436), .ZN(n_257_76_15216));
   NAND2_X1 i_257_76_15244 (.A1(n_257_926), .A2(n_257_439), .ZN(n_257_76_15217));
   NAND2_X1 i_257_76_15245 (.A1(n_257_824), .A2(n_257_437), .ZN(n_257_76_15218));
   NAND3_X1 i_257_76_15246 (.A1(n_257_76_15216), .A2(n_257_76_15217), .A3(
      n_257_76_15218), .ZN(n_257_76_15219));
   NOR2_X1 i_257_76_15247 (.A1(n_257_76_15215), .A2(n_257_76_15219), .ZN(
      n_257_76_15220));
   NAND2_X1 i_257_76_15248 (.A1(n_257_696), .A2(n_257_448), .ZN(n_257_76_15221));
   NAND3_X1 i_257_76_15249 (.A1(n_257_76_15220), .A2(n_257_76_15221), .A3(
      n_257_76_15180), .ZN(n_257_76_15222));
   INV_X1 i_257_76_15250 (.A(n_257_76_15191), .ZN(n_257_76_15223));
   NOR2_X1 i_257_76_15251 (.A1(n_257_76_15222), .A2(n_257_76_15223), .ZN(
      n_257_76_15224));
   NAND2_X1 i_257_76_15252 (.A1(n_257_28), .A2(n_257_76_15224), .ZN(
      n_257_76_15225));
   NAND3_X1 i_257_76_15253 (.A1(n_257_76_15194), .A2(n_257_76_15201), .A3(
      n_257_76_15225), .ZN(n_257_76_15226));
   NAND3_X1 i_257_76_15254 (.A1(n_257_76_15205), .A2(n_257_76_15195), .A3(
      n_257_856), .ZN(n_257_76_15227));
   NAND2_X1 i_257_76_15255 (.A1(n_257_446), .A2(n_257_76_15204), .ZN(
      n_257_76_15228));
   NOR2_X1 i_257_76_15256 (.A1(n_257_76_15227), .A2(n_257_76_15228), .ZN(
      n_257_76_15229));
   NAND4_X1 i_257_76_15257 (.A1(n_257_76_15217), .A2(n_257_76_15209), .A3(
      n_257_76_15229), .A4(n_257_76_15181), .ZN(n_257_76_15230));
   INV_X1 i_257_76_15258 (.A(n_257_76_15230), .ZN(n_257_76_15231));
   NAND2_X1 i_257_76_15259 (.A1(n_257_76_15180), .A2(n_257_76_15231), .ZN(
      n_257_76_15232));
   INV_X1 i_257_76_15260 (.A(n_257_76_15232), .ZN(n_257_76_15233));
   NAND2_X1 i_257_76_15261 (.A1(n_257_76_15233), .A2(n_257_76_15191), .ZN(
      n_257_76_15234));
   INV_X1 i_257_76_15262 (.A(n_257_76_15234), .ZN(n_257_76_15235));
   NAND2_X1 i_257_76_15263 (.A1(n_257_76_18070), .A2(n_257_76_15235), .ZN(
      n_257_76_15236));
   NAND3_X1 i_257_76_15264 (.A1(n_257_76_15204), .A2(n_257_76_15195), .A3(
      n_257_439), .ZN(n_257_76_15237));
   INV_X1 i_257_76_15265 (.A(n_257_76_15237), .ZN(n_257_76_15238));
   NAND3_X1 i_257_76_15266 (.A1(n_257_76_15181), .A2(n_257_926), .A3(
      n_257_76_15238), .ZN(n_257_76_15239));
   INV_X1 i_257_76_15267 (.A(n_257_76_15239), .ZN(n_257_76_15240));
   NAND2_X1 i_257_76_15268 (.A1(n_257_76_15180), .A2(n_257_76_15240), .ZN(
      n_257_76_15241));
   INV_X1 i_257_76_15269 (.A(n_257_76_15241), .ZN(n_257_76_15242));
   NAND2_X1 i_257_76_15270 (.A1(n_257_76_15242), .A2(n_257_76_15191), .ZN(
      n_257_76_15243));
   INV_X1 i_257_76_15271 (.A(n_257_76_15243), .ZN(n_257_76_15244));
   NAND2_X1 i_257_76_15272 (.A1(n_257_76_18084), .A2(n_257_76_15244), .ZN(
      n_257_76_15245));
   NAND2_X1 i_257_76_15273 (.A1(n_257_179), .A2(n_257_429), .ZN(n_257_76_15246));
   NAND2_X1 i_257_76_15274 (.A1(n_257_140), .A2(n_257_430), .ZN(n_257_76_15247));
   NAND2_X1 i_257_76_15275 (.A1(n_257_102), .A2(n_257_431), .ZN(n_257_76_15248));
   NAND3_X1 i_257_76_15276 (.A1(n_257_76_15246), .A2(n_257_76_15247), .A3(
      n_257_76_15248), .ZN(n_257_76_15249));
   NAND2_X1 i_257_76_15277 (.A1(n_257_259), .A2(n_257_425), .ZN(n_257_76_15250));
   NAND2_X1 i_257_76_15278 (.A1(n_257_219), .A2(n_257_427), .ZN(n_257_76_15251));
   NAND3_X1 i_257_76_15279 (.A1(n_257_76_15202), .A2(n_257_76_15204), .A3(
      n_257_76_15251), .ZN(n_257_76_15252));
   NAND2_X1 i_257_76_15280 (.A1(n_257_432), .A2(n_257_624), .ZN(n_257_76_15253));
   INV_X1 i_257_76_15281 (.A(n_257_76_15253), .ZN(n_257_76_15254));
   NOR2_X1 i_257_76_15282 (.A1(n_257_1086), .A2(n_257_76_15254), .ZN(
      n_257_76_15255));
   NAND2_X1 i_257_76_15283 (.A1(n_257_423), .A2(n_257_442), .ZN(n_257_76_15256));
   NAND3_X1 i_257_76_15284 (.A1(n_257_76_15205), .A2(n_257_76_15255), .A3(
      n_257_76_17981), .ZN(n_257_76_15257));
   NOR2_X1 i_257_76_15285 (.A1(n_257_76_15252), .A2(n_257_76_15257), .ZN(
      n_257_76_15258));
   NAND2_X1 i_257_76_15286 (.A1(n_257_528), .A2(n_257_424), .ZN(n_257_76_15259));
   NAND2_X1 i_257_76_15287 (.A1(n_257_62), .A2(n_257_433), .ZN(n_257_76_15260));
   NAND3_X1 i_257_76_15288 (.A1(n_257_299), .A2(n_257_76_15259), .A3(
      n_257_76_15260), .ZN(n_257_76_15261));
   INV_X1 i_257_76_15289 (.A(n_257_76_15261), .ZN(n_257_76_15262));
   NAND2_X1 i_257_76_15290 (.A1(n_257_656), .A2(n_257_450), .ZN(n_257_76_15263));
   NAND3_X1 i_257_76_15291 (.A1(n_257_76_15258), .A2(n_257_76_15262), .A3(
      n_257_76_15263), .ZN(n_257_76_15264));
   INV_X1 i_257_76_15292 (.A(n_257_76_15264), .ZN(n_257_76_15265));
   NAND2_X1 i_257_76_15293 (.A1(n_257_76_15250), .A2(n_257_76_15265), .ZN(
      n_257_76_15266));
   NOR2_X1 i_257_76_15294 (.A1(n_257_76_15249), .A2(n_257_76_15266), .ZN(
      n_257_76_15267));
   NAND2_X1 i_257_76_15295 (.A1(n_257_76_15221), .A2(n_257_76_15180), .ZN(
      n_257_76_15268));
   INV_X1 i_257_76_15296 (.A(n_257_76_15268), .ZN(n_257_76_15269));
   NAND4_X1 i_257_76_15297 (.A1(n_257_76_15216), .A2(n_257_76_15217), .A3(
      n_257_76_15218), .A4(n_257_76_15209), .ZN(n_257_76_15270));
   NAND2_X1 i_257_76_15298 (.A1(n_257_560), .A2(n_257_426), .ZN(n_257_76_15271));
   NAND2_X1 i_257_76_15299 (.A1(n_257_451), .A2(n_257_479), .ZN(n_257_76_15272));
   NAND4_X1 i_257_76_15300 (.A1(n_257_76_15271), .A2(n_257_76_15214), .A3(
      n_257_76_15181), .A4(n_257_76_15272), .ZN(n_257_76_15273));
   NOR2_X1 i_257_76_15301 (.A1(n_257_76_15270), .A2(n_257_76_15273), .ZN(
      n_257_76_15274));
   NAND4_X1 i_257_76_15302 (.A1(n_257_76_15267), .A2(n_257_76_15269), .A3(
      n_257_76_15191), .A4(n_257_76_15274), .ZN(n_257_76_15275));
   INV_X1 i_257_76_15303 (.A(n_257_76_15275), .ZN(n_257_76_15276));
   NAND2_X1 i_257_76_15304 (.A1(n_257_76_18066), .A2(n_257_76_15276), .ZN(
      n_257_76_15277));
   NAND3_X1 i_257_76_15305 (.A1(n_257_76_15236), .A2(n_257_76_15245), .A3(
      n_257_76_15277), .ZN(n_257_76_15278));
   NOR2_X1 i_257_76_15306 (.A1(n_257_76_15226), .A2(n_257_76_15278), .ZN(
      n_257_76_15279));
   NAND3_X1 i_257_76_15307 (.A1(n_257_990), .A2(n_257_441), .A3(n_257_76_15195), 
      .ZN(n_257_76_15280));
   INV_X1 i_257_76_15308 (.A(n_257_76_15280), .ZN(n_257_76_15281));
   NAND2_X1 i_257_76_15309 (.A1(n_257_76_15180), .A2(n_257_76_15281), .ZN(
      n_257_76_15282));
   INV_X1 i_257_76_15310 (.A(n_257_76_15282), .ZN(n_257_76_15283));
   NAND2_X1 i_257_76_15311 (.A1(n_257_76_15283), .A2(n_257_76_15191), .ZN(
      n_257_76_15284));
   INV_X1 i_257_76_15312 (.A(n_257_76_15284), .ZN(n_257_76_15285));
   NAND2_X1 i_257_76_15313 (.A1(n_257_76_18071), .A2(n_257_76_15285), .ZN(
      n_257_76_15286));
   NAND2_X1 i_257_76_15314 (.A1(n_257_76_15210), .A2(n_257_76_15212), .ZN(
      n_257_76_15287));
   INV_X1 i_257_76_15315 (.A(n_257_76_15287), .ZN(n_257_76_15288));
   NAND2_X1 i_257_76_15316 (.A1(n_257_435), .A2(n_257_442), .ZN(n_257_76_15289));
   NOR2_X1 i_257_76_15317 (.A1(n_257_1086), .A2(n_257_76_15289), .ZN(
      n_257_76_15290));
   NAND4_X1 i_257_76_15318 (.A1(n_257_76_15204), .A2(n_257_76_15205), .A3(
      n_257_76_15290), .A4(n_257_728), .ZN(n_257_76_15291));
   INV_X1 i_257_76_15319 (.A(n_257_76_15291), .ZN(n_257_76_15292));
   NAND4_X1 i_257_76_15320 (.A1(n_257_76_15209), .A2(n_257_76_15181), .A3(
      n_257_76_15288), .A4(n_257_76_15292), .ZN(n_257_76_15293));
   NOR2_X1 i_257_76_15321 (.A1(n_257_76_15219), .A2(n_257_76_15293), .ZN(
      n_257_76_15294));
   NAND2_X1 i_257_76_15322 (.A1(n_257_76_15180), .A2(n_257_76_15294), .ZN(
      n_257_76_15295));
   NOR2_X1 i_257_76_15323 (.A1(n_257_76_15295), .A2(n_257_76_15223), .ZN(
      n_257_76_15296));
   NAND2_X1 i_257_76_15324 (.A1(n_257_76_18078), .A2(n_257_76_15296), .ZN(
      n_257_76_15297));
   INV_X1 i_257_76_15325 (.A(n_257_76_15205), .ZN(n_257_76_15298));
   NAND3_X1 i_257_76_15326 (.A1(n_257_592), .A2(n_257_428), .A3(n_257_442), 
      .ZN(n_257_76_15299));
   INV_X1 i_257_76_15327 (.A(n_257_76_15299), .ZN(n_257_76_15300));
   NAND3_X1 i_257_76_15328 (.A1(n_257_76_15182), .A2(n_257_76_15253), .A3(
      n_257_76_15300), .ZN(n_257_76_15301));
   NOR2_X1 i_257_76_15329 (.A1(n_257_76_15298), .A2(n_257_76_15301), .ZN(
      n_257_76_15302));
   NAND2_X1 i_257_76_15330 (.A1(n_257_76_15202), .A2(n_257_76_15204), .ZN(
      n_257_76_15303));
   INV_X1 i_257_76_15331 (.A(n_257_76_15303), .ZN(n_257_76_15304));
   NAND4_X1 i_257_76_15332 (.A1(n_257_76_15302), .A2(n_257_76_15304), .A3(
      n_257_76_15212), .A4(n_257_76_15260), .ZN(n_257_76_15305));
   NAND3_X1 i_257_76_15333 (.A1(n_257_76_15263), .A2(n_257_76_15210), .A3(
      n_257_76_15211), .ZN(n_257_76_15306));
   NOR2_X1 i_257_76_15334 (.A1(n_257_76_15305), .A2(n_257_76_15306), .ZN(
      n_257_76_15307));
   NAND2_X1 i_257_76_15335 (.A1(n_257_76_15217), .A2(n_257_76_15218), .ZN(
      n_257_76_15308));
   INV_X1 i_257_76_15336 (.A(n_257_76_15308), .ZN(n_257_76_15309));
   NAND3_X1 i_257_76_15337 (.A1(n_257_76_15209), .A2(n_257_76_15181), .A3(
      n_257_76_15272), .ZN(n_257_76_15310));
   INV_X1 i_257_76_15338 (.A(n_257_76_15310), .ZN(n_257_76_15311));
   NAND3_X1 i_257_76_15339 (.A1(n_257_76_15307), .A2(n_257_76_15309), .A3(
      n_257_76_15311), .ZN(n_257_76_15312));
   NAND4_X1 i_257_76_15340 (.A1(n_257_76_15246), .A2(n_257_76_15247), .A3(
      n_257_76_15248), .A4(n_257_76_15216), .ZN(n_257_76_15313));
   NOR2_X1 i_257_76_15341 (.A1(n_257_76_15312), .A2(n_257_76_15313), .ZN(
      n_257_76_15314));
   NAND3_X1 i_257_76_15342 (.A1(n_257_76_15314), .A2(n_257_76_15269), .A3(
      n_257_76_15191), .ZN(n_257_76_15315));
   INV_X1 i_257_76_15343 (.A(n_257_76_15315), .ZN(n_257_76_15316));
   NAND2_X1 i_257_76_15344 (.A1(n_257_76_18074), .A2(n_257_76_15316), .ZN(
      n_257_76_15317));
   NAND3_X1 i_257_76_15345 (.A1(n_257_76_15286), .A2(n_257_76_15297), .A3(
      n_257_76_15317), .ZN(n_257_76_15318));
   NAND2_X1 i_257_76_15346 (.A1(n_257_1086), .A2(n_257_442), .ZN(n_257_76_15319));
   INV_X1 i_257_76_15347 (.A(n_257_76_15319), .ZN(n_257_76_15320));
   NAND2_X1 i_257_76_15348 (.A1(n_257_13), .A2(n_257_76_15320), .ZN(
      n_257_76_15321));
   INV_X1 i_257_76_15349 (.A(n_257_76_15217), .ZN(n_257_76_15322));
   NOR2_X1 i_257_76_15350 (.A1(n_257_76_17902), .A2(n_257_1086), .ZN(
      n_257_76_15323));
   NAND3_X1 i_257_76_15351 (.A1(n_257_76_15323), .A2(n_257_76_15204), .A3(
      n_257_76_15205), .ZN(n_257_76_15324));
   INV_X1 i_257_76_15352 (.A(n_257_76_15324), .ZN(n_257_76_15325));
   NAND3_X1 i_257_76_15353 (.A1(n_257_76_15181), .A2(n_257_888), .A3(
      n_257_76_15325), .ZN(n_257_76_15326));
   NOR2_X1 i_257_76_15354 (.A1(n_257_76_15322), .A2(n_257_76_15326), .ZN(
      n_257_76_15327));
   NAND2_X1 i_257_76_15355 (.A1(n_257_76_15180), .A2(n_257_76_15327), .ZN(
      n_257_76_15328));
   INV_X1 i_257_76_15356 (.A(n_257_76_15328), .ZN(n_257_76_15329));
   NAND2_X1 i_257_76_15357 (.A1(n_257_76_15329), .A2(n_257_76_15191), .ZN(
      n_257_76_15330));
   INV_X1 i_257_76_15358 (.A(n_257_76_15330), .ZN(n_257_76_15331));
   NAND2_X1 i_257_76_15359 (.A1(n_257_76_18077), .A2(n_257_76_15331), .ZN(
      n_257_76_15332));
   NAND2_X1 i_257_76_15360 (.A1(n_257_76_15321), .A2(n_257_76_15332), .ZN(
      n_257_76_15333));
   NOR2_X1 i_257_76_15361 (.A1(n_257_76_15318), .A2(n_257_76_15333), .ZN(
      n_257_76_15334));
   NAND2_X1 i_257_76_15362 (.A1(n_257_426), .A2(n_257_442), .ZN(n_257_76_15335));
   NAND3_X1 i_257_76_15363 (.A1(n_257_76_15205), .A2(n_257_76_15255), .A3(
      n_257_76_17982), .ZN(n_257_76_15336));
   NAND2_X1 i_257_76_15364 (.A1(n_257_76_15204), .A2(n_257_76_15251), .ZN(
      n_257_76_15337));
   NOR2_X1 i_257_76_15365 (.A1(n_257_76_15336), .A2(n_257_76_15337), .ZN(
      n_257_76_15338));
   NAND3_X1 i_257_76_15366 (.A1(n_257_76_15212), .A2(n_257_76_15260), .A3(
      n_257_76_15202), .ZN(n_257_76_15339));
   INV_X1 i_257_76_15367 (.A(n_257_76_15339), .ZN(n_257_76_15340));
   NAND2_X1 i_257_76_15368 (.A1(n_257_76_15210), .A2(n_257_76_15211), .ZN(
      n_257_76_15341));
   INV_X1 i_257_76_15369 (.A(n_257_76_15341), .ZN(n_257_76_15342));
   NAND3_X1 i_257_76_15370 (.A1(n_257_76_15338), .A2(n_257_76_15340), .A3(
      n_257_76_15342), .ZN(n_257_76_15343));
   NAND4_X1 i_257_76_15371 (.A1(n_257_76_15181), .A2(n_257_76_15272), .A3(
      n_257_560), .A4(n_257_76_15263), .ZN(n_257_76_15344));
   NOR2_X1 i_257_76_15372 (.A1(n_257_76_15343), .A2(n_257_76_15344), .ZN(
      n_257_76_15345));
   NAND2_X1 i_257_76_15373 (.A1(n_257_76_15248), .A2(n_257_76_15216), .ZN(
      n_257_76_15346));
   INV_X1 i_257_76_15374 (.A(n_257_76_15346), .ZN(n_257_76_15347));
   NAND3_X1 i_257_76_15375 (.A1(n_257_76_15217), .A2(n_257_76_15218), .A3(
      n_257_76_15209), .ZN(n_257_76_15348));
   INV_X1 i_257_76_15376 (.A(n_257_76_15348), .ZN(n_257_76_15349));
   NAND3_X1 i_257_76_15377 (.A1(n_257_76_15345), .A2(n_257_76_15347), .A3(
      n_257_76_15349), .ZN(n_257_76_15350));
   INV_X1 i_257_76_15378 (.A(n_257_76_15350), .ZN(n_257_76_15351));
   NAND2_X1 i_257_76_15379 (.A1(n_257_76_15246), .A2(n_257_76_15247), .ZN(
      n_257_76_15352));
   INV_X1 i_257_76_15380 (.A(n_257_76_15352), .ZN(n_257_76_15353));
   NAND3_X1 i_257_76_15381 (.A1(n_257_76_15221), .A2(n_257_76_15353), .A3(
      n_257_76_15180), .ZN(n_257_76_15354));
   INV_X1 i_257_76_15382 (.A(n_257_76_15354), .ZN(n_257_76_15355));
   NAND3_X1 i_257_76_15383 (.A1(n_257_76_15351), .A2(n_257_76_15355), .A3(
      n_257_76_15191), .ZN(n_257_76_15356));
   INV_X1 i_257_76_15384 (.A(n_257_76_15356), .ZN(n_257_76_15357));
   NAND2_X1 i_257_76_15385 (.A1(n_257_76_18076), .A2(n_257_76_15357), .ZN(
      n_257_76_15358));
   NOR2_X1 i_257_76_15386 (.A1(n_257_1086), .A2(n_257_76_17934), .ZN(
      n_257_76_15359));
   NAND3_X1 i_257_76_15387 (.A1(n_257_76_15204), .A2(n_257_76_15205), .A3(
      n_257_76_15359), .ZN(n_257_76_15360));
   INV_X1 i_257_76_15388 (.A(n_257_76_15360), .ZN(n_257_76_15361));
   NAND4_X1 i_257_76_15389 (.A1(n_257_760), .A2(n_257_76_15288), .A3(
      n_257_76_15181), .A4(n_257_76_15361), .ZN(n_257_76_15362));
   NOR2_X1 i_257_76_15390 (.A1(n_257_76_15348), .A2(n_257_76_15362), .ZN(
      n_257_76_15363));
   NAND2_X1 i_257_76_15391 (.A1(n_257_76_15180), .A2(n_257_76_15363), .ZN(
      n_257_76_15364));
   NOR2_X1 i_257_76_15392 (.A1(n_257_76_15223), .A2(n_257_76_15364), .ZN(
      n_257_76_15365));
   NAND2_X1 i_257_76_15393 (.A1(n_257_76_18069), .A2(n_257_76_15365), .ZN(
      n_257_76_15366));
   INV_X1 i_257_76_15394 (.A(n_257_76_15270), .ZN(n_257_76_15367));
   NAND2_X1 i_257_76_15395 (.A1(n_257_76_15212), .A2(n_257_76_15260), .ZN(
      n_257_76_15368));
   INV_X1 i_257_76_15396 (.A(n_257_76_15368), .ZN(n_257_76_15369));
   NAND3_X1 i_257_76_15397 (.A1(n_257_432), .A2(n_257_624), .A3(n_257_442), 
      .ZN(n_257_76_15370));
   NOR2_X1 i_257_76_15398 (.A1(n_257_1086), .A2(n_257_76_15370), .ZN(
      n_257_76_15371));
   NAND4_X1 i_257_76_15399 (.A1(n_257_76_15202), .A2(n_257_76_15204), .A3(
      n_257_76_15205), .A4(n_257_76_15371), .ZN(n_257_76_15372));
   INV_X1 i_257_76_15400 (.A(n_257_76_15372), .ZN(n_257_76_15373));
   NAND3_X1 i_257_76_15401 (.A1(n_257_76_15342), .A2(n_257_76_15369), .A3(
      n_257_76_15373), .ZN(n_257_76_15374));
   NAND3_X1 i_257_76_15402 (.A1(n_257_76_15181), .A2(n_257_76_15272), .A3(
      n_257_76_15263), .ZN(n_257_76_15375));
   NOR2_X1 i_257_76_15403 (.A1(n_257_76_15374), .A2(n_257_76_15375), .ZN(
      n_257_76_15376));
   NAND4_X1 i_257_76_15404 (.A1(n_257_76_15221), .A2(n_257_76_15180), .A3(
      n_257_76_15367), .A4(n_257_76_15376), .ZN(n_257_76_15377));
   NOR2_X1 i_257_76_15405 (.A1(n_257_76_15377), .A2(n_257_76_15223), .ZN(
      n_257_76_15378));
   NAND2_X1 i_257_76_15406 (.A1(n_257_68), .A2(n_257_76_15378), .ZN(
      n_257_76_15379));
   NAND3_X1 i_257_76_15407 (.A1(n_257_76_15358), .A2(n_257_76_15366), .A3(
      n_257_76_15379), .ZN(n_257_76_15380));
   INV_X1 i_257_76_15408 (.A(n_257_76_15210), .ZN(n_257_76_15381));
   NOR2_X1 i_257_76_15409 (.A1(n_257_1086), .A2(n_257_76_17951), .ZN(
      n_257_76_15382));
   NAND3_X1 i_257_76_15410 (.A1(n_257_76_15204), .A2(n_257_76_15205), .A3(
      n_257_76_15382), .ZN(n_257_76_15383));
   NOR2_X1 i_257_76_15411 (.A1(n_257_76_15381), .A2(n_257_76_15383), .ZN(
      n_257_76_15384));
   NAND3_X1 i_257_76_15412 (.A1(n_257_76_15384), .A2(n_257_824), .A3(
      n_257_76_15181), .ZN(n_257_76_15385));
   NAND2_X1 i_257_76_15413 (.A1(n_257_76_15217), .A2(n_257_76_15209), .ZN(
      n_257_76_15386));
   NOR2_X1 i_257_76_15414 (.A1(n_257_76_15385), .A2(n_257_76_15386), .ZN(
      n_257_76_15387));
   NAND2_X1 i_257_76_15415 (.A1(n_257_76_15180), .A2(n_257_76_15387), .ZN(
      n_257_76_15388));
   NOR2_X1 i_257_76_15416 (.A1(n_257_76_15223), .A2(n_257_76_15388), .ZN(
      n_257_76_15389));
   NAND2_X1 i_257_76_15417 (.A1(n_257_22), .A2(n_257_76_15389), .ZN(
      n_257_76_15390));
   NAND2_X1 i_257_76_15418 (.A1(n_257_444), .A2(n_257_76_15195), .ZN(
      n_257_76_15391));
   INV_X1 i_257_76_15419 (.A(n_257_76_15391), .ZN(n_257_76_15392));
   NAND2_X1 i_257_76_15420 (.A1(n_257_1022), .A2(n_257_76_15392), .ZN(
      n_257_76_15393));
   INV_X1 i_257_76_15421 (.A(n_257_76_15393), .ZN(n_257_76_15394));
   NAND2_X1 i_257_76_15422 (.A1(n_257_76_15191), .A2(n_257_76_15394), .ZN(
      n_257_76_15395));
   INV_X1 i_257_76_15423 (.A(n_257_76_15395), .ZN(n_257_76_15396));
   NAND2_X1 i_257_76_15424 (.A1(n_257_76_18075), .A2(n_257_76_15396), .ZN(
      n_257_76_15397));
   NAND2_X1 i_257_76_15425 (.A1(n_257_76_15390), .A2(n_257_76_15397), .ZN(
      n_257_76_15398));
   NOR2_X1 i_257_76_15426 (.A1(n_257_76_15380), .A2(n_257_76_15398), .ZN(
      n_257_76_15399));
   NAND3_X1 i_257_76_15427 (.A1(n_257_76_15279), .A2(n_257_76_15334), .A3(
      n_257_76_15399), .ZN(n_257_76_15400));
   INV_X1 i_257_76_15428 (.A(n_257_76_15400), .ZN(n_257_76_15401));
   NAND2_X1 i_257_76_15429 (.A1(n_257_76_15212), .A2(n_257_76_15202), .ZN(
      n_257_76_15402));
   INV_X1 i_257_76_15430 (.A(n_257_76_15402), .ZN(n_257_76_15403));
   NOR2_X1 i_257_76_15431 (.A1(n_257_1086), .A2(n_257_76_17633), .ZN(
      n_257_76_15404));
   NAND4_X1 i_257_76_15432 (.A1(n_257_76_15204), .A2(n_257_62), .A3(
      n_257_76_15205), .A4(n_257_76_15404), .ZN(n_257_76_15405));
   INV_X1 i_257_76_15433 (.A(n_257_76_15405), .ZN(n_257_76_15406));
   NAND3_X1 i_257_76_15434 (.A1(n_257_76_15342), .A2(n_257_76_15403), .A3(
      n_257_76_15406), .ZN(n_257_76_15407));
   NOR2_X1 i_257_76_15435 (.A1(n_257_76_15407), .A2(n_257_76_15375), .ZN(
      n_257_76_15408));
   NAND4_X1 i_257_76_15436 (.A1(n_257_76_15221), .A2(n_257_76_15180), .A3(
      n_257_76_15367), .A4(n_257_76_15408), .ZN(n_257_76_15409));
   NOR2_X1 i_257_76_15437 (.A1(n_257_76_15409), .A2(n_257_76_15223), .ZN(
      n_257_76_15410));
   NAND2_X1 i_257_76_15438 (.A1(n_257_76_18081), .A2(n_257_76_15410), .ZN(
      n_257_76_15411));
   NAND2_X1 i_257_76_15439 (.A1(n_257_442), .A2(n_257_664), .ZN(n_257_76_15412));
   NOR2_X1 i_257_76_15440 (.A1(n_257_1086), .A2(n_257_76_15412), .ZN(
      n_257_76_15413));
   NAND3_X1 i_257_76_15441 (.A1(n_257_76_15204), .A2(n_257_76_15205), .A3(
      n_257_76_15413), .ZN(n_257_76_15414));
   NAND2_X1 i_257_76_15442 (.A1(n_257_76_15202), .A2(n_257_449), .ZN(
      n_257_76_15415));
   NOR2_X1 i_257_76_15443 (.A1(n_257_76_15414), .A2(n_257_76_15415), .ZN(
      n_257_76_15416));
   NAND4_X1 i_257_76_15444 (.A1(n_257_76_15209), .A2(n_257_76_15416), .A3(
      n_257_76_15181), .A4(n_257_76_15288), .ZN(n_257_76_15417));
   NOR2_X1 i_257_76_15445 (.A1(n_257_76_15417), .A2(n_257_76_15219), .ZN(
      n_257_76_15418));
   NAND3_X1 i_257_76_15446 (.A1(n_257_76_15418), .A2(n_257_76_15221), .A3(
      n_257_76_15180), .ZN(n_257_76_15419));
   NOR2_X1 i_257_76_15447 (.A1(n_257_76_15419), .A2(n_257_76_15223), .ZN(
      n_257_76_15420));
   NAND2_X1 i_257_76_15448 (.A1(n_257_76_18083), .A2(n_257_76_15420), .ZN(
      n_257_76_15421));
   NAND3_X1 i_257_76_15449 (.A1(n_257_76_15205), .A2(n_257_76_17983), .A3(
      n_257_76_15182), .ZN(n_257_76_15422));
   INV_X1 i_257_76_15450 (.A(n_257_76_15422), .ZN(n_257_76_15423));
   NAND4_X1 i_257_76_15451 (.A1(n_257_76_15304), .A2(n_257_76_15423), .A3(
      n_257_76_15212), .A4(n_257_76_15260), .ZN(n_257_76_15424));
   NOR2_X1 i_257_76_15452 (.A1(n_257_76_15424), .A2(n_257_76_15306), .ZN(
      n_257_76_15425));
   NAND3_X1 i_257_76_15453 (.A1(n_257_76_15425), .A2(n_257_76_15309), .A3(
      n_257_76_15311), .ZN(n_257_76_15426));
   NAND4_X1 i_257_76_15454 (.A1(n_257_76_15247), .A2(n_257_76_15248), .A3(
      n_257_179), .A4(n_257_76_15216), .ZN(n_257_76_15427));
   NOR2_X1 i_257_76_15455 (.A1(n_257_76_15426), .A2(n_257_76_15427), .ZN(
      n_257_76_15428));
   NAND3_X1 i_257_76_15456 (.A1(n_257_76_15428), .A2(n_257_76_15269), .A3(
      n_257_76_15191), .ZN(n_257_76_15429));
   INV_X1 i_257_76_15457 (.A(n_257_76_15429), .ZN(n_257_76_15430));
   NAND2_X1 i_257_76_15458 (.A1(n_257_76_18061), .A2(n_257_76_15430), .ZN(
      n_257_76_15431));
   NAND3_X1 i_257_76_15459 (.A1(n_257_76_15411), .A2(n_257_76_15421), .A3(
      n_257_76_15431), .ZN(n_257_76_15432));
   INV_X1 i_257_76_15460 (.A(n_257_76_15432), .ZN(n_257_76_15433));
   NAND2_X1 i_257_76_15461 (.A1(n_257_442), .A2(n_257_894), .ZN(n_257_76_15434));
   NOR2_X1 i_257_76_15462 (.A1(n_257_1086), .A2(n_257_76_15434), .ZN(
      n_257_76_15435));
   NAND3_X1 i_257_76_15463 (.A1(n_257_76_15204), .A2(n_257_76_15435), .A3(
      n_257_438), .ZN(n_257_76_15436));
   INV_X1 i_257_76_15464 (.A(n_257_76_15436), .ZN(n_257_76_15437));
   NAND2_X1 i_257_76_15465 (.A1(n_257_76_15181), .A2(n_257_76_15437), .ZN(
      n_257_76_15438));
   NOR2_X1 i_257_76_15466 (.A1(n_257_76_15322), .A2(n_257_76_15438), .ZN(
      n_257_76_15439));
   NAND2_X1 i_257_76_15467 (.A1(n_257_76_15180), .A2(n_257_76_15439), .ZN(
      n_257_76_15440));
   INV_X1 i_257_76_15468 (.A(n_257_76_15440), .ZN(n_257_76_15441));
   NAND2_X1 i_257_76_15469 (.A1(n_257_76_15441), .A2(n_257_76_15191), .ZN(
      n_257_76_15442));
   INV_X1 i_257_76_15470 (.A(n_257_76_15442), .ZN(n_257_76_15443));
   NAND2_X1 i_257_76_15471 (.A1(n_257_76_18067), .A2(n_257_76_15443), .ZN(
      n_257_76_15444));
   NAND2_X1 i_257_76_15472 (.A1(n_257_76_15347), .A2(n_257_76_15247), .ZN(
      n_257_76_15445));
   NAND2_X1 i_257_76_15473 (.A1(n_257_76_15250), .A2(n_257_76_15246), .ZN(
      n_257_76_15446));
   NOR2_X1 i_257_76_15474 (.A1(n_257_76_15445), .A2(n_257_76_15446), .ZN(
      n_257_76_15447));
   NAND2_X1 i_257_76_15475 (.A1(n_257_76_15209), .A2(n_257_76_15271), .ZN(
      n_257_76_15448));
   NAND2_X1 i_257_76_15476 (.A1(n_257_376), .A2(n_257_421), .ZN(n_257_76_15449));
   NAND2_X1 i_257_76_15477 (.A1(n_257_76_15449), .A2(n_257_76_15181), .ZN(
      n_257_76_15450));
   NOR2_X1 i_257_76_15478 (.A1(n_257_76_15448), .A2(n_257_76_15450), .ZN(
      n_257_76_15451));
   NAND2_X1 i_257_76_15479 (.A1(n_257_76_15451), .A2(n_257_76_15309), .ZN(
      n_257_76_15452));
   NAND2_X1 i_257_76_15480 (.A1(n_257_337), .A2(n_257_422), .ZN(n_257_76_15453));
   INV_X1 i_257_76_15481 (.A(n_257_76_15453), .ZN(n_257_76_15454));
   NOR2_X1 i_257_76_15482 (.A1(n_257_76_15337), .A2(n_257_76_15454), .ZN(
      n_257_76_15455));
   NAND2_X1 i_257_76_15483 (.A1(n_257_442), .A2(n_257_496), .ZN(n_257_76_15456));
   NAND2_X1 i_257_76_15484 (.A1(n_257_76_15205), .A2(n_257_76_17984), .ZN(
      n_257_76_15457));
   NAND2_X1 i_257_76_15485 (.A1(n_257_420), .A2(n_257_76_15253), .ZN(
      n_257_76_15458));
   INV_X1 i_257_76_15486 (.A(n_257_76_15458), .ZN(n_257_76_15459));
   NAND2_X1 i_257_76_15487 (.A1(n_257_76_15459), .A2(n_257_76_15182), .ZN(
      n_257_76_15460));
   NOR2_X1 i_257_76_15488 (.A1(n_257_76_15457), .A2(n_257_76_15460), .ZN(
      n_257_76_15461));
   NAND2_X1 i_257_76_15489 (.A1(n_257_76_15455), .A2(n_257_76_15461), .ZN(
      n_257_76_15462));
   NAND2_X1 i_257_76_15490 (.A1(n_257_76_15212), .A2(n_257_76_15259), .ZN(
      n_257_76_15463));
   INV_X1 i_257_76_15491 (.A(n_257_76_15463), .ZN(n_257_76_15464));
   NAND2_X1 i_257_76_15492 (.A1(n_257_76_15260), .A2(n_257_76_15202), .ZN(
      n_257_76_15465));
   INV_X1 i_257_76_15493 (.A(n_257_76_15465), .ZN(n_257_76_15466));
   NAND2_X1 i_257_76_15494 (.A1(n_257_76_15464), .A2(n_257_76_15466), .ZN(
      n_257_76_15467));
   NOR2_X1 i_257_76_15495 (.A1(n_257_76_15462), .A2(n_257_76_15467), .ZN(
      n_257_76_15468));
   NAND2_X1 i_257_76_15496 (.A1(n_257_76_15342), .A2(n_257_76_15263), .ZN(
      n_257_76_15469));
   NAND2_X1 i_257_76_15497 (.A1(n_257_299), .A2(n_257_423), .ZN(n_257_76_15470));
   NAND2_X1 i_257_76_15498 (.A1(n_257_76_15272), .A2(n_257_76_15470), .ZN(
      n_257_76_15471));
   NOR2_X1 i_257_76_15499 (.A1(n_257_76_15469), .A2(n_257_76_15471), .ZN(
      n_257_76_15472));
   NAND2_X1 i_257_76_15500 (.A1(n_257_76_15468), .A2(n_257_76_15472), .ZN(
      n_257_76_15473));
   NOR2_X1 i_257_76_15501 (.A1(n_257_76_15452), .A2(n_257_76_15473), .ZN(
      n_257_76_15474));
   NAND2_X1 i_257_76_15502 (.A1(n_257_76_15447), .A2(n_257_76_15474), .ZN(
      n_257_76_15475));
   NAND2_X1 i_257_76_15503 (.A1(n_257_76_15269), .A2(n_257_76_15191), .ZN(
      n_257_76_15476));
   NOR2_X1 i_257_76_15504 (.A1(n_257_76_15475), .A2(n_257_76_15476), .ZN(
      n_257_76_15477));
   NAND2_X1 i_257_76_15505 (.A1(n_257_76_18073), .A2(n_257_76_15477), .ZN(
      n_257_76_15478));
   NAND2_X1 i_257_76_15506 (.A1(n_257_76_15204), .A2(n_257_76_15205), .ZN(
      n_257_76_15479));
   INV_X1 i_257_76_15507 (.A(n_257_76_15479), .ZN(n_257_76_15480));
   INV_X1 i_257_76_15508 (.A(n_257_432), .ZN(n_257_76_15481));
   NAND2_X1 i_257_76_15509 (.A1(n_257_76_17925), .A2(n_257_76_15481), .ZN(
      n_257_76_15482));
   INV_X1 i_257_76_15510 (.A(n_257_624), .ZN(n_257_76_15483));
   NAND2_X1 i_257_76_15511 (.A1(n_257_76_17925), .A2(n_257_76_15483), .ZN(
      n_257_76_15484));
   AOI21_X1 i_257_76_15512 (.A(n_257_1086), .B1(n_257_76_15482), .B2(
      n_257_76_15484), .ZN(n_257_76_15485));
   NAND4_X1 i_257_76_15513 (.A1(n_257_76_15480), .A2(n_257_76_15260), .A3(
      n_257_76_15485), .A4(n_257_76_15202), .ZN(n_257_76_15486));
   NOR2_X1 i_257_76_15514 (.A1(n_257_76_15486), .A2(n_257_76_15213), .ZN(
      n_257_76_15487));
   NAND2_X1 i_257_76_15515 (.A1(n_257_76_15209), .A2(n_257_140), .ZN(
      n_257_76_15488));
   INV_X1 i_257_76_15516 (.A(n_257_76_15488), .ZN(n_257_76_15489));
   INV_X1 i_257_76_15517 (.A(n_257_76_15375), .ZN(n_257_76_15490));
   NAND3_X1 i_257_76_15518 (.A1(n_257_76_15487), .A2(n_257_76_15489), .A3(
      n_257_76_15490), .ZN(n_257_76_15491));
   NAND4_X1 i_257_76_15519 (.A1(n_257_76_15248), .A2(n_257_76_15216), .A3(
      n_257_76_15217), .A4(n_257_76_15218), .ZN(n_257_76_15492));
   NOR2_X1 i_257_76_15520 (.A1(n_257_76_15491), .A2(n_257_76_15492), .ZN(
      n_257_76_15493));
   NAND4_X1 i_257_76_15521 (.A1(n_257_76_15493), .A2(n_257_76_15191), .A3(
      n_257_76_15221), .A4(n_257_76_15180), .ZN(n_257_76_15494));
   INV_X1 i_257_76_15522 (.A(n_257_76_15494), .ZN(n_257_76_15495));
   NAND2_X1 i_257_76_15523 (.A1(n_257_76_18068), .A2(n_257_76_15495), .ZN(
      n_257_76_15496));
   NAND3_X1 i_257_76_15524 (.A1(n_257_76_15444), .A2(n_257_76_15478), .A3(
      n_257_76_15496), .ZN(n_257_76_15497));
   INV_X1 i_257_76_15525 (.A(n_257_76_15497), .ZN(n_257_76_15498));
   NAND2_X1 i_257_76_15526 (.A1(n_257_792), .A2(n_257_442), .ZN(n_257_76_15499));
   NOR2_X1 i_257_76_15527 (.A1(n_257_1086), .A2(n_257_76_15499), .ZN(
      n_257_76_15500));
   NAND4_X1 i_257_76_15528 (.A1(n_257_447), .A2(n_257_76_15204), .A3(
      n_257_76_15205), .A4(n_257_76_15500), .ZN(n_257_76_15501));
   NOR2_X1 i_257_76_15529 (.A1(n_257_76_15501), .A2(n_257_76_15381), .ZN(
      n_257_76_15502));
   NAND3_X1 i_257_76_15530 (.A1(n_257_76_15502), .A2(n_257_76_15209), .A3(
      n_257_76_15181), .ZN(n_257_76_15503));
   NOR2_X1 i_257_76_15531 (.A1(n_257_76_15503), .A2(n_257_76_15308), .ZN(
      n_257_76_15504));
   NAND2_X1 i_257_76_15532 (.A1(n_257_76_15180), .A2(n_257_76_15504), .ZN(
      n_257_76_15505));
   NOR2_X1 i_257_76_15533 (.A1(n_257_76_15505), .A2(n_257_76_15223), .ZN(
      n_257_76_15506));
   NAND2_X1 i_257_76_15534 (.A1(n_257_76_17932), .A2(n_257_76_15481), .ZN(
      n_257_76_15507));
   NAND2_X1 i_257_76_15535 (.A1(n_257_76_17932), .A2(n_257_76_15483), .ZN(
      n_257_76_15508));
   AOI21_X1 i_257_76_15536 (.A(n_257_1086), .B1(n_257_76_15507), .B2(
      n_257_76_15508), .ZN(n_257_76_15509));
   NAND3_X1 i_257_76_15537 (.A1(n_257_76_15509), .A2(n_257_76_15204), .A3(
      n_257_76_15205), .ZN(n_257_76_15510));
   NOR2_X1 i_257_76_15538 (.A1(n_257_76_15510), .A2(n_257_76_15465), .ZN(
      n_257_76_15511));
   NAND3_X1 i_257_76_15539 (.A1(n_257_76_15511), .A2(n_257_76_15214), .A3(
      n_257_76_15263), .ZN(n_257_76_15512));
   NAND3_X1 i_257_76_15540 (.A1(n_257_102), .A2(n_257_76_15181), .A3(
      n_257_76_15272), .ZN(n_257_76_15513));
   NOR2_X1 i_257_76_15541 (.A1(n_257_76_15512), .A2(n_257_76_15513), .ZN(
      n_257_76_15514));
   NAND4_X1 i_257_76_15542 (.A1(n_257_76_15514), .A2(n_257_76_15221), .A3(
      n_257_76_15180), .A4(n_257_76_15367), .ZN(n_257_76_15515));
   NOR2_X1 i_257_76_15543 (.A1(n_257_76_15515), .A2(n_257_76_15223), .ZN(
      n_257_76_15516));
   AOI22_X1 i_257_76_15544 (.A1(n_257_76_18085), .A2(n_257_76_15506), .B1(
      n_257_76_18080), .B2(n_257_76_15516), .ZN(n_257_76_15517));
   NAND3_X1 i_257_76_15545 (.A1(n_257_76_15433), .A2(n_257_76_15498), .A3(
      n_257_76_15517), .ZN(n_257_76_15518));
   NAND3_X1 i_257_76_15546 (.A1(n_257_76_15204), .A2(n_257_76_15205), .A3(
      n_257_76_15182), .ZN(n_257_76_15519));
   OAI21_X1 i_257_76_15547 (.A(n_257_76_17761), .B1(n_257_728), .B2(
      n_257_76_17412), .ZN(n_257_76_15520));
   INV_X1 i_257_76_15548 (.A(n_257_76_15520), .ZN(n_257_76_15521));
   NOR2_X1 i_257_76_15549 (.A1(n_257_76_15519), .A2(n_257_76_15521), .ZN(
      n_257_76_15522));
   NAND3_X1 i_257_76_15550 (.A1(n_257_76_15210), .A2(n_257_76_15212), .A3(
      n_257_448), .ZN(n_257_76_15523));
   INV_X1 i_257_76_15551 (.A(n_257_76_15523), .ZN(n_257_76_15524));
   NAND4_X1 i_257_76_15552 (.A1(n_257_76_15209), .A2(n_257_76_15522), .A3(
      n_257_76_15524), .A4(n_257_76_15181), .ZN(n_257_76_15525));
   INV_X1 i_257_76_15553 (.A(n_257_76_15525), .ZN(n_257_76_15526));
   INV_X1 i_257_76_15554 (.A(n_257_76_15219), .ZN(n_257_76_15527));
   NAND3_X1 i_257_76_15555 (.A1(n_257_76_15526), .A2(n_257_696), .A3(
      n_257_76_15527), .ZN(n_257_76_15528));
   INV_X1 i_257_76_15556 (.A(n_257_76_15528), .ZN(n_257_76_15529));
   NAND3_X1 i_257_76_15557 (.A1(n_257_76_15191), .A2(n_257_76_15529), .A3(
      n_257_76_15180), .ZN(n_257_76_15530));
   INV_X1 i_257_76_15558 (.A(n_257_76_15530), .ZN(n_257_76_15531));
   NAND2_X1 i_257_76_15559 (.A1(n_257_76_18079), .A2(n_257_76_15531), .ZN(
      n_257_76_15532));
   NAND3_X1 i_257_76_15560 (.A1(n_257_76_15191), .A2(n_257_76_15221), .A3(
      n_257_76_15180), .ZN(n_257_76_15533));
   NAND4_X1 i_257_76_15561 (.A1(n_257_76_15209), .A2(n_257_76_15271), .A3(
      n_257_76_15181), .A4(n_257_76_15272), .ZN(n_257_76_15534));
   NAND2_X1 i_257_76_15562 (.A1(n_257_425), .A2(n_257_442), .ZN(n_257_76_15535));
   NAND3_X1 i_257_76_15563 (.A1(n_257_76_15205), .A2(n_257_76_15255), .A3(
      n_257_76_17985), .ZN(n_257_76_15536));
   NOR2_X1 i_257_76_15564 (.A1(n_257_76_15536), .A2(n_257_76_15337), .ZN(
      n_257_76_15537));
   NAND4_X1 i_257_76_15565 (.A1(n_257_76_15537), .A2(n_257_76_15340), .A3(
      n_257_76_15342), .A4(n_257_76_15263), .ZN(n_257_76_15538));
   NOR2_X1 i_257_76_15566 (.A1(n_257_76_15534), .A2(n_257_76_15538), .ZN(
      n_257_76_15539));
   NAND2_X1 i_257_76_15567 (.A1(n_257_76_15248), .A2(n_257_259), .ZN(
      n_257_76_15540));
   NOR2_X1 i_257_76_15568 (.A1(n_257_76_15219), .A2(n_257_76_15540), .ZN(
      n_257_76_15541));
   NAND3_X1 i_257_76_15569 (.A1(n_257_76_15353), .A2(n_257_76_15539), .A3(
      n_257_76_15541), .ZN(n_257_76_15542));
   NOR2_X1 i_257_76_15570 (.A1(n_257_76_15533), .A2(n_257_76_15542), .ZN(
      n_257_76_15543));
   NAND2_X1 i_257_76_15571 (.A1(n_257_76_18064), .A2(n_257_76_15543), .ZN(
      n_257_76_15544));
   NAND3_X1 i_257_76_15572 (.A1(n_257_76_15453), .A2(n_257_76_15204), .A3(
      n_257_76_15251), .ZN(n_257_76_15545));
   NAND2_X1 i_257_76_15573 (.A1(n_257_421), .A2(n_257_442), .ZN(n_257_76_15546));
   NAND3_X1 i_257_76_15574 (.A1(n_257_76_15205), .A2(n_257_76_15255), .A3(
      n_257_76_17986), .ZN(n_257_76_15547));
   NOR2_X1 i_257_76_15575 (.A1(n_257_76_15545), .A2(n_257_76_15547), .ZN(
      n_257_76_15548));
   NAND3_X1 i_257_76_15576 (.A1(n_257_76_15259), .A2(n_257_76_15260), .A3(
      n_257_76_15202), .ZN(n_257_76_15549));
   INV_X1 i_257_76_15577 (.A(n_257_76_15549), .ZN(n_257_76_15550));
   NAND3_X1 i_257_76_15578 (.A1(n_257_76_15548), .A2(n_257_76_15214), .A3(
      n_257_76_15550), .ZN(n_257_76_15551));
   NAND4_X1 i_257_76_15579 (.A1(n_257_76_15272), .A2(n_257_76_15470), .A3(
      n_257_76_15263), .A4(n_257_376), .ZN(n_257_76_15552));
   NOR2_X1 i_257_76_15580 (.A1(n_257_76_15551), .A2(n_257_76_15552), .ZN(
      n_257_76_15553));
   NAND3_X1 i_257_76_15581 (.A1(n_257_76_15248), .A2(n_257_76_15216), .A3(
      n_257_76_15217), .ZN(n_257_76_15554));
   INV_X1 i_257_76_15582 (.A(n_257_76_15554), .ZN(n_257_76_15555));
   NAND4_X1 i_257_76_15583 (.A1(n_257_76_15218), .A2(n_257_76_15209), .A3(
      n_257_76_15271), .A4(n_257_76_15181), .ZN(n_257_76_15556));
   INV_X1 i_257_76_15584 (.A(n_257_76_15556), .ZN(n_257_76_15557));
   NAND3_X1 i_257_76_15585 (.A1(n_257_76_15553), .A2(n_257_76_15555), .A3(
      n_257_76_15557), .ZN(n_257_76_15558));
   INV_X1 i_257_76_15586 (.A(n_257_76_15558), .ZN(n_257_76_15559));
   NAND3_X1 i_257_76_15587 (.A1(n_257_76_15250), .A2(n_257_76_15246), .A3(
      n_257_76_15247), .ZN(n_257_76_15560));
   INV_X1 i_257_76_15588 (.A(n_257_76_15560), .ZN(n_257_76_15561));
   NAND4_X1 i_257_76_15589 (.A1(n_257_76_15559), .A2(n_257_76_15269), .A3(
      n_257_76_15191), .A4(n_257_76_15561), .ZN(n_257_76_15562));
   INV_X1 i_257_76_15590 (.A(n_257_76_15562), .ZN(n_257_76_15563));
   NAND2_X1 i_257_76_15591 (.A1(n_257_76_18082), .A2(n_257_76_15563), .ZN(
      n_257_76_15564));
   NAND3_X1 i_257_76_15592 (.A1(n_257_76_15532), .A2(n_257_76_15544), .A3(
      n_257_76_15564), .ZN(n_257_76_15565));
   INV_X1 i_257_76_15593 (.A(n_257_76_15565), .ZN(n_257_76_15566));
   NAND2_X1 i_257_76_15594 (.A1(n_257_427), .A2(n_257_76_15253), .ZN(
      n_257_76_15567));
   INV_X1 i_257_76_15595 (.A(n_257_76_15567), .ZN(n_257_76_15568));
   NAND4_X1 i_257_76_15596 (.A1(n_257_76_15568), .A2(n_257_219), .A3(
      n_257_76_17987), .A4(n_257_76_15182), .ZN(n_257_76_15569));
   INV_X1 i_257_76_15597 (.A(n_257_76_15569), .ZN(n_257_76_15570));
   NAND4_X1 i_257_76_15598 (.A1(n_257_76_15181), .A2(n_257_76_15272), .A3(
      n_257_76_15263), .A4(n_257_76_15570), .ZN(n_257_76_15571));
   NAND3_X1 i_257_76_15599 (.A1(n_257_76_15202), .A2(n_257_76_15204), .A3(
      n_257_76_15205), .ZN(n_257_76_15572));
   INV_X1 i_257_76_15600 (.A(n_257_76_15572), .ZN(n_257_76_15573));
   NAND3_X1 i_257_76_15601 (.A1(n_257_76_15342), .A2(n_257_76_15369), .A3(
      n_257_76_15573), .ZN(n_257_76_15574));
   NOR2_X1 i_257_76_15602 (.A1(n_257_76_15571), .A2(n_257_76_15574), .ZN(
      n_257_76_15575));
   NAND3_X1 i_257_76_15603 (.A1(n_257_76_15247), .A2(n_257_76_15248), .A3(
      n_257_76_15216), .ZN(n_257_76_15576));
   INV_X1 i_257_76_15604 (.A(n_257_76_15576), .ZN(n_257_76_15577));
   NAND4_X1 i_257_76_15605 (.A1(n_257_76_15575), .A2(n_257_76_15577), .A3(
      n_257_76_15246), .A4(n_257_76_15349), .ZN(n_257_76_15578));
   INV_X1 i_257_76_15606 (.A(n_257_76_15578), .ZN(n_257_76_15579));
   NAND3_X1 i_257_76_15607 (.A1(n_257_76_15579), .A2(n_257_76_15269), .A3(
      n_257_76_15191), .ZN(n_257_76_15580));
   INV_X1 i_257_76_15608 (.A(n_257_76_15580), .ZN(n_257_76_15581));
   NAND2_X1 i_257_76_15609 (.A1(n_257_76_18065), .A2(n_257_76_15581), .ZN(
      n_257_76_15582));
   NAND3_X1 i_257_76_15610 (.A1(n_257_76_15522), .A2(n_257_76_15181), .A3(
      n_257_76_15263), .ZN(n_257_76_15583));
   NAND3_X1 i_257_76_15611 (.A1(n_257_76_15211), .A2(n_257_479), .A3(
      n_257_76_15212), .ZN(n_257_76_15584));
   INV_X1 i_257_76_15612 (.A(n_257_76_15584), .ZN(n_257_76_15585));
   NAND2_X1 i_257_76_15613 (.A1(n_257_451), .A2(n_257_76_15210), .ZN(
      n_257_76_15586));
   INV_X1 i_257_76_15614 (.A(n_257_76_15586), .ZN(n_257_76_15587));
   NAND2_X1 i_257_76_15615 (.A1(n_257_76_15585), .A2(n_257_76_15587), .ZN(
      n_257_76_15588));
   NOR2_X1 i_257_76_15616 (.A1(n_257_76_15583), .A2(n_257_76_15588), .ZN(
      n_257_76_15589));
   NAND4_X1 i_257_76_15617 (.A1(n_257_76_15221), .A2(n_257_76_15180), .A3(
      n_257_76_15589), .A4(n_257_76_15367), .ZN(n_257_76_15590));
   NOR2_X1 i_257_76_15618 (.A1(n_257_76_15590), .A2(n_257_76_15223), .ZN(
      n_257_76_15591));
   NAND2_X1 i_257_76_15619 (.A1(n_257_76_18063), .A2(n_257_76_15591), .ZN(
      n_257_76_15592));
   NAND2_X1 i_257_76_15620 (.A1(n_257_76_15253), .A2(n_257_424), .ZN(
      n_257_76_15593));
   NOR2_X1 i_257_76_15621 (.A1(n_257_76_15593), .A2(n_257_1086), .ZN(
      n_257_76_15594));
   NAND3_X1 i_257_76_15622 (.A1(n_257_76_15594), .A2(n_257_76_15205), .A3(
      n_257_76_17987), .ZN(n_257_76_15595));
   INV_X1 i_257_76_15623 (.A(n_257_76_15595), .ZN(n_257_76_15596));
   NAND3_X1 i_257_76_15624 (.A1(n_257_528), .A2(n_257_76_15204), .A3(
      n_257_76_15251), .ZN(n_257_76_15597));
   INV_X1 i_257_76_15625 (.A(n_257_76_15597), .ZN(n_257_76_15598));
   NAND4_X1 i_257_76_15626 (.A1(n_257_76_15466), .A2(n_257_76_15596), .A3(
      n_257_76_15263), .A4(n_257_76_15598), .ZN(n_257_76_15599));
   INV_X1 i_257_76_15627 (.A(n_257_76_15599), .ZN(n_257_76_15600));
   NAND4_X1 i_257_76_15628 (.A1(n_257_76_15600), .A2(n_257_76_15247), .A3(
      n_257_76_15248), .A4(n_257_76_15216), .ZN(n_257_76_15601));
   NOR2_X1 i_257_76_15629 (.A1(n_257_76_15601), .A2(n_257_76_15446), .ZN(
      n_257_76_15602));
   NOR2_X1 i_257_76_15630 (.A1(n_257_76_15273), .A2(n_257_76_15348), .ZN(
      n_257_76_15603));
   NAND4_X1 i_257_76_15631 (.A1(n_257_76_15602), .A2(n_257_76_15269), .A3(
      n_257_76_15191), .A4(n_257_76_15603), .ZN(n_257_76_15604));
   INV_X1 i_257_76_15632 (.A(n_257_76_15604), .ZN(n_257_76_15605));
   NAND2_X1 i_257_76_15633 (.A1(n_257_76_18062), .A2(n_257_76_15605), .ZN(
      n_257_76_15606));
   NAND3_X1 i_257_76_15634 (.A1(n_257_76_15582), .A2(n_257_76_15592), .A3(
      n_257_76_15606), .ZN(n_257_76_15607));
   INV_X1 i_257_76_15635 (.A(n_257_76_15607), .ZN(n_257_76_15608));
   NAND2_X1 i_257_76_15636 (.A1(n_257_76_15253), .A2(n_257_422), .ZN(
      n_257_76_15609));
   INV_X1 i_257_76_15637 (.A(n_257_76_15609), .ZN(n_257_76_15610));
   NAND4_X1 i_257_76_15638 (.A1(n_257_337), .A2(n_257_76_15610), .A3(
      n_257_76_17987), .A4(n_257_76_15182), .ZN(n_257_76_15611));
   INV_X1 i_257_76_15639 (.A(n_257_76_15611), .ZN(n_257_76_15612));
   NAND3_X1 i_257_76_15640 (.A1(n_257_76_15612), .A2(n_257_76_15210), .A3(
      n_257_76_15211), .ZN(n_257_76_15613));
   INV_X1 i_257_76_15641 (.A(n_257_76_15263), .ZN(n_257_76_15614));
   NOR2_X1 i_257_76_15642 (.A1(n_257_76_15613), .A2(n_257_76_15614), .ZN(
      n_257_76_15615));
   INV_X1 i_257_76_15643 (.A(n_257_76_15471), .ZN(n_257_76_15616));
   NAND3_X1 i_257_76_15644 (.A1(n_257_76_15212), .A2(n_257_76_15259), .A3(
      n_257_76_15260), .ZN(n_257_76_15617));
   NAND4_X1 i_257_76_15645 (.A1(n_257_76_15202), .A2(n_257_76_15204), .A3(
      n_257_76_15251), .A4(n_257_76_15205), .ZN(n_257_76_15618));
   NOR2_X1 i_257_76_15646 (.A1(n_257_76_15617), .A2(n_257_76_15618), .ZN(
      n_257_76_15619));
   NAND3_X1 i_257_76_15647 (.A1(n_257_76_15615), .A2(n_257_76_15616), .A3(
      n_257_76_15619), .ZN(n_257_76_15620));
   NOR2_X1 i_257_76_15648 (.A1(n_257_76_15620), .A2(n_257_76_15556), .ZN(
      n_257_76_15621));
   INV_X1 i_257_76_15649 (.A(n_257_76_15446), .ZN(n_257_76_15622));
   NAND4_X1 i_257_76_15650 (.A1(n_257_76_15247), .A2(n_257_76_15248), .A3(
      n_257_76_15216), .A4(n_257_76_15217), .ZN(n_257_76_15623));
   INV_X1 i_257_76_15651 (.A(n_257_76_15623), .ZN(n_257_76_15624));
   NAND4_X1 i_257_76_15652 (.A1(n_257_76_15621), .A2(n_257_76_15622), .A3(
      n_257_76_15180), .A4(n_257_76_15624), .ZN(n_257_76_15625));
   NAND2_X1 i_257_76_15653 (.A1(n_257_76_15191), .A2(n_257_76_15221), .ZN(
      n_257_76_15626));
   NOR2_X1 i_257_76_15654 (.A1(n_257_76_15625), .A2(n_257_76_15626), .ZN(
      n_257_76_15627));
   NAND2_X1 i_257_76_15655 (.A1(n_257_342), .A2(n_257_76_15627), .ZN(
      n_257_76_15628));
   NAND4_X1 i_257_76_15656 (.A1(n_257_76_15250), .A2(n_257_76_15246), .A3(
      n_257_76_15247), .A4(n_257_76_15248), .ZN(n_257_76_15629));
   INV_X1 i_257_76_15657 (.A(n_257_76_15629), .ZN(n_257_76_15630));
   INV_X1 i_257_76_15658 (.A(n_257_76_15448), .ZN(n_257_76_15631));
   NAND3_X1 i_257_76_15659 (.A1(n_257_76_15449), .A2(n_257_76_15181), .A3(
      n_257_76_15272), .ZN(n_257_76_15632));
   INV_X1 i_257_76_15660 (.A(n_257_76_15632), .ZN(n_257_76_15633));
   NAND2_X1 i_257_76_15661 (.A1(n_257_76_15631), .A2(n_257_76_15633), .ZN(
      n_257_76_15634));
   NOR2_X1 i_257_76_15662 (.A1(n_257_76_15634), .A2(n_257_76_15219), .ZN(
      n_257_76_15635));
   NAND2_X1 i_257_76_15663 (.A1(n_257_76_15630), .A2(n_257_76_15635), .ZN(
      n_257_76_15636));
   NAND2_X1 i_257_76_15664 (.A1(n_257_76_15253), .A2(n_257_415), .ZN(
      n_257_76_15637));
   NOR2_X1 i_257_76_15665 (.A1(n_257_76_15637), .A2(n_257_1086), .ZN(
      n_257_76_15638));
   NAND2_X1 i_257_76_15666 (.A1(n_257_420), .A2(n_257_496), .ZN(n_257_76_15639));
   NAND2_X1 i_257_76_15667 (.A1(n_257_484), .A2(n_257_442), .ZN(n_257_76_15640));
   NAND2_X1 i_257_76_15668 (.A1(n_257_76_15639), .A2(n_257_76_17988), .ZN(
      n_257_76_15641));
   INV_X1 i_257_76_15669 (.A(n_257_76_15641), .ZN(n_257_76_15642));
   NAND3_X1 i_257_76_15670 (.A1(n_257_76_15638), .A2(n_257_76_15642), .A3(
      n_257_76_15205), .ZN(n_257_76_15643));
   NOR2_X1 i_257_76_15671 (.A1(n_257_76_15643), .A2(n_257_76_15337), .ZN(
      n_257_76_15644));
   NAND3_X1 i_257_76_15672 (.A1(n_257_76_15260), .A2(n_257_76_15202), .A3(
      n_257_76_15453), .ZN(n_257_76_15645));
   INV_X1 i_257_76_15673 (.A(n_257_76_15645), .ZN(n_257_76_15646));
   NAND3_X1 i_257_76_15674 (.A1(n_257_76_15644), .A2(n_257_76_15464), .A3(
      n_257_76_15646), .ZN(n_257_76_15647));
   NAND4_X1 i_257_76_15675 (.A1(n_257_76_15470), .A2(n_257_76_15263), .A3(
      n_257_76_15210), .A4(n_257_76_15211), .ZN(n_257_76_15648));
   NOR2_X1 i_257_76_15676 (.A1(n_257_76_15647), .A2(n_257_76_15648), .ZN(
      n_257_76_15649));
   NAND3_X1 i_257_76_15677 (.A1(n_257_76_15221), .A2(n_257_76_15649), .A3(
      n_257_76_15180), .ZN(n_257_76_15650));
   NOR3_X1 i_257_76_15678 (.A1(n_257_76_15636), .A2(n_257_76_15650), .A3(
      n_257_76_15223), .ZN(n_257_76_15651));
   NAND2_X1 i_257_76_15679 (.A1(n_257_76_18060), .A2(n_257_76_15651), .ZN(
      n_257_76_15652));
   NAND2_X1 i_257_76_15680 (.A1(n_257_62), .A2(n_257_76_17918), .ZN(
      n_257_76_15653));
   NAND2_X1 i_257_76_15681 (.A1(n_257_76_15611), .A2(n_257_76_15653), .ZN(
      n_257_76_15654));
   INV_X1 i_257_76_15682 (.A(n_257_76_15289), .ZN(n_257_76_15655));
   NAND2_X1 i_257_76_15683 (.A1(n_257_728), .A2(n_257_76_15655), .ZN(
      n_257_76_15656));
   NAND2_X1 i_257_76_15684 (.A1(n_257_440), .A2(n_257_76_15184), .ZN(
      n_257_76_15657));
   INV_X1 i_257_76_15685 (.A(n_257_76_15434), .ZN(n_257_76_15658));
   NAND2_X1 i_257_76_15686 (.A1(n_257_438), .A2(n_257_76_15658), .ZN(
      n_257_76_15659));
   NAND3_X1 i_257_76_15687 (.A1(n_257_76_15656), .A2(n_257_76_15657), .A3(
      n_257_76_15659), .ZN(n_257_76_15660));
   NOR2_X1 i_257_76_15688 (.A1(n_257_76_15654), .A2(n_257_76_15660), .ZN(
      n_257_76_15661));
   NAND2_X1 i_257_76_15689 (.A1(n_257_415), .A2(n_257_484), .ZN(n_257_76_15662));
   NAND2_X1 i_257_76_15690 (.A1(n_257_76_15662), .A2(n_257_76_15253), .ZN(
      n_257_76_15663));
   INV_X1 i_257_76_15691 (.A(n_257_76_15663), .ZN(n_257_76_15664));
   INV_X1 i_257_76_15692 (.A(Small_Packet_Data_Size[27]), .ZN(n_257_76_15665));
   NAND4_X1 i_257_76_15693 (.A1(n_257_76_15664), .A2(n_257_76_17989), .A3(
      n_257_76_15639), .A4(n_257_76_15182), .ZN(n_257_76_15666));
   INV_X1 i_257_76_15694 (.A(n_257_76_15666), .ZN(n_257_76_15667));
   NOR2_X1 i_257_76_15695 (.A1(n_257_442), .A2(n_257_76_15665), .ZN(
      n_257_76_15668));
   OAI21_X1 i_257_76_15696 (.A(n_257_76_15569), .B1(n_257_76_15667), .B2(
      n_257_76_15668), .ZN(n_257_76_15669));
   INV_X1 i_257_76_15697 (.A(n_257_76_15669), .ZN(n_257_76_15670));
   NAND2_X1 i_257_76_15698 (.A1(n_257_856), .A2(n_257_442), .ZN(n_257_76_15671));
   INV_X1 i_257_76_15699 (.A(n_257_76_15671), .ZN(n_257_76_15672));
   NAND2_X1 i_257_76_15700 (.A1(n_257_446), .A2(n_257_76_15672), .ZN(
      n_257_76_15673));
   INV_X1 i_257_76_15701 (.A(n_257_76_15412), .ZN(n_257_76_15674));
   NAND2_X1 i_257_76_15702 (.A1(n_257_449), .A2(n_257_76_15674), .ZN(
      n_257_76_15675));
   INV_X1 i_257_76_15703 (.A(n_257_76_15499), .ZN(n_257_76_15676));
   NAND2_X1 i_257_76_15704 (.A1(n_257_447), .A2(n_257_76_15676), .ZN(
      n_257_76_15677));
   NAND3_X1 i_257_76_15705 (.A1(n_257_76_15673), .A2(n_257_76_15675), .A3(
      n_257_76_15677), .ZN(n_257_76_15678));
   INV_X1 i_257_76_15706 (.A(n_257_76_15678), .ZN(n_257_76_15679));
   NAND3_X1 i_257_76_15707 (.A1(n_257_76_15661), .A2(n_257_76_15670), .A3(
      n_257_76_15679), .ZN(n_257_76_15680));
   NAND2_X1 i_257_76_15708 (.A1(n_257_888), .A2(n_257_76_17903), .ZN(
      n_257_76_15681));
   NAND3_X1 i_257_76_15709 (.A1(n_257_990), .A2(n_257_441), .A3(n_257_442), 
      .ZN(n_257_76_15682));
   NAND3_X1 i_257_76_15710 (.A1(n_257_451), .A2(n_257_479), .A3(n_257_76_15520), 
      .ZN(n_257_76_15683));
   NAND2_X1 i_257_76_15711 (.A1(n_257_656), .A2(n_257_76_17928), .ZN(
      n_257_76_15684));
   NAND4_X1 i_257_76_15712 (.A1(n_257_76_15681), .A2(n_257_76_15682), .A3(
      n_257_76_15683), .A4(n_257_76_15684), .ZN(n_257_76_15685));
   NOR2_X1 i_257_76_15713 (.A1(n_257_76_15680), .A2(n_257_76_15685), .ZN(
      n_257_76_15686));
   NAND2_X1 i_257_76_15714 (.A1(n_257_140), .A2(n_257_76_17925), .ZN(
      n_257_76_15687));
   NAND2_X1 i_257_76_15715 (.A1(n_257_102), .A2(n_257_76_17932), .ZN(
      n_257_76_15688));
   NAND3_X1 i_257_76_15716 (.A1(n_257_76_15599), .A2(n_257_76_15687), .A3(
      n_257_76_15688), .ZN(n_257_76_15689));
   INV_X1 i_257_76_15717 (.A(n_257_76_15689), .ZN(n_257_76_15690));
   NAND2_X1 i_257_76_15718 (.A1(n_257_760), .A2(n_257_76_17935), .ZN(
      n_257_76_15691));
   NAND2_X1 i_257_76_15719 (.A1(n_257_926), .A2(n_257_76_17940), .ZN(
      n_257_76_15692));
   NAND2_X1 i_257_76_15720 (.A1(n_257_824), .A2(n_257_76_17952), .ZN(
      n_257_76_15693));
   NAND3_X1 i_257_76_15721 (.A1(n_257_76_15691), .A2(n_257_76_15692), .A3(
      n_257_76_15693), .ZN(n_257_76_15694));
   INV_X1 i_257_76_15722 (.A(n_257_76_15694), .ZN(n_257_76_15695));
   NAND3_X1 i_257_76_15723 (.A1(n_257_76_15686), .A2(n_257_76_15690), .A3(
      n_257_76_15695), .ZN(n_257_76_15696));
   NAND2_X1 i_257_76_15724 (.A1(n_257_696), .A2(n_257_76_17958), .ZN(
      n_257_76_15697));
   INV_X1 i_257_76_15725 (.A(n_257_179), .ZN(n_257_76_15698));
   OAI21_X1 i_257_76_15726 (.A(n_257_76_15264), .B1(n_257_76_15698), .B2(
      n_257_76_17660), .ZN(n_257_76_15699));
   INV_X1 i_257_76_15727 (.A(n_257_76_15699), .ZN(n_257_76_15700));
   NAND2_X1 i_257_76_15728 (.A1(n_257_1022), .A2(n_257_76_17964), .ZN(
      n_257_76_15701));
   NAND3_X1 i_257_76_15729 (.A1(n_257_76_15697), .A2(n_257_76_15700), .A3(
      n_257_76_15701), .ZN(n_257_76_15702));
   NOR2_X1 i_257_76_15730 (.A1(n_257_76_15696), .A2(n_257_76_15702), .ZN(
      n_257_76_15703));
   NAND2_X1 i_257_76_15731 (.A1(n_257_1054), .A2(n_257_76_17969), .ZN(
      n_257_76_15704));
   NAND3_X1 i_257_76_15732 (.A1(n_257_76_15704), .A2(n_257_76_15558), .A3(
      n_257_76_15350), .ZN(n_257_76_15705));
   INV_X1 i_257_76_15733 (.A(n_257_76_15705), .ZN(n_257_76_15706));
   NAND3_X1 i_257_76_15734 (.A1(n_257_76_15703), .A2(n_257_76_15706), .A3(
      n_257_76_15542), .ZN(n_257_76_15707));
   NAND3_X1 i_257_76_15735 (.A1(n_257_76_15628), .A2(n_257_76_15652), .A3(
      n_257_76_15707), .ZN(n_257_76_15708));
   INV_X1 i_257_76_15736 (.A(n_257_76_15708), .ZN(n_257_76_15709));
   NAND3_X1 i_257_76_15737 (.A1(n_257_76_15566), .A2(n_257_76_15608), .A3(
      n_257_76_15709), .ZN(n_257_76_15710));
   NOR2_X1 i_257_76_15738 (.A1(n_257_76_15518), .A2(n_257_76_15710), .ZN(
      n_257_76_15711));
   NAND2_X1 i_257_76_15739 (.A1(n_257_76_15401), .A2(n_257_76_15711), .ZN(n_27));
   NAND2_X1 i_257_76_15740 (.A1(n_257_1055), .A2(n_257_443), .ZN(n_257_76_15712));
   NAND2_X1 i_257_76_15741 (.A1(n_257_1023), .A2(n_257_444), .ZN(n_257_76_15713));
   NAND2_X1 i_257_76_15742 (.A1(n_257_441), .A2(n_257_991), .ZN(n_257_76_15714));
   NAND2_X1 i_257_76_15743 (.A1(n_257_959), .A2(n_257_442), .ZN(n_257_76_15715));
   NOR2_X1 i_257_76_15744 (.A1(n_257_1087), .A2(n_257_76_15715), .ZN(
      n_257_76_15716));
   NAND2_X1 i_257_76_15745 (.A1(n_257_440), .A2(n_257_76_15716), .ZN(
      n_257_76_15717));
   INV_X1 i_257_76_15746 (.A(n_257_76_15717), .ZN(n_257_76_15718));
   NAND2_X1 i_257_76_15747 (.A1(n_257_76_15714), .A2(n_257_76_15718), .ZN(
      n_257_76_15719));
   INV_X1 i_257_76_15748 (.A(n_257_76_15719), .ZN(n_257_76_15720));
   NAND2_X1 i_257_76_15749 (.A1(n_257_76_15713), .A2(n_257_76_15720), .ZN(
      n_257_76_15721));
   INV_X1 i_257_76_15750 (.A(n_257_76_15721), .ZN(n_257_76_15722));
   NAND2_X1 i_257_76_15751 (.A1(n_257_76_15712), .A2(n_257_76_15722), .ZN(
      n_257_76_15723));
   INV_X1 i_257_76_15752 (.A(n_257_76_15723), .ZN(n_257_76_15724));
   NAND2_X1 i_257_76_15753 (.A1(n_257_17), .A2(n_257_76_15724), .ZN(
      n_257_76_15725));
   NOR2_X1 i_257_76_15754 (.A1(n_257_1087), .A2(n_257_76_17412), .ZN(
      n_257_76_15726));
   NAND2_X1 i_257_76_15755 (.A1(n_257_443), .A2(n_257_76_15726), .ZN(
      n_257_76_15727));
   INV_X1 i_257_76_15756 (.A(n_257_76_15727), .ZN(n_257_76_15728));
   NAND2_X1 i_257_76_15757 (.A1(n_257_1055), .A2(n_257_76_15728), .ZN(
      n_257_76_15729));
   INV_X1 i_257_76_15758 (.A(n_257_76_15729), .ZN(n_257_76_15730));
   NAND2_X1 i_257_76_15759 (.A1(n_257_76_18072), .A2(n_257_76_15730), .ZN(
      n_257_76_15731));
   NAND2_X1 i_257_76_15760 (.A1(n_257_761), .A2(n_257_436), .ZN(n_257_76_15732));
   NAND2_X1 i_257_76_15761 (.A1(n_257_446), .A2(n_257_857), .ZN(n_257_76_15733));
   NAND2_X1 i_257_76_15762 (.A1(n_257_449), .A2(n_257_665), .ZN(n_257_76_15734));
   NAND3_X1 i_257_76_15763 (.A1(n_257_76_15732), .A2(n_257_76_15733), .A3(
      n_257_76_15734), .ZN(n_257_76_15735));
   INV_X1 i_257_76_15764 (.A(n_257_76_15714), .ZN(n_257_76_15736));
   NOR2_X1 i_257_76_15765 (.A1(n_257_76_15735), .A2(n_257_76_15736), .ZN(
      n_257_76_15737));
   NAND2_X1 i_257_76_15766 (.A1(n_257_447), .A2(n_257_793), .ZN(n_257_76_15738));
   NAND2_X1 i_257_76_15767 (.A1(n_257_927), .A2(n_257_439), .ZN(n_257_76_15739));
   NAND2_X1 i_257_76_15768 (.A1(n_257_825), .A2(n_257_437), .ZN(n_257_76_15740));
   NAND3_X1 i_257_76_15769 (.A1(n_257_76_15738), .A2(n_257_76_15739), .A3(
      n_257_76_15740), .ZN(n_257_76_15741));
   NAND2_X1 i_257_76_15770 (.A1(n_257_450), .A2(n_257_76_15726), .ZN(
      n_257_76_15742));
   INV_X1 i_257_76_15771 (.A(n_257_76_15742), .ZN(n_257_76_15743));
   NAND2_X1 i_257_76_15772 (.A1(n_257_729), .A2(n_257_435), .ZN(n_257_76_15744));
   NAND3_X1 i_257_76_15773 (.A1(n_257_76_15743), .A2(n_257_657), .A3(
      n_257_76_15744), .ZN(n_257_76_15745));
   INV_X1 i_257_76_15774 (.A(n_257_76_15745), .ZN(n_257_76_15746));
   NAND2_X1 i_257_76_15775 (.A1(n_257_889), .A2(n_257_445), .ZN(n_257_76_15747));
   NAND2_X1 i_257_76_15776 (.A1(n_257_440), .A2(n_257_959), .ZN(n_257_76_15748));
   NAND2_X1 i_257_76_15777 (.A1(n_257_438), .A2(n_257_895), .ZN(n_257_76_15749));
   NAND4_X1 i_257_76_15778 (.A1(n_257_76_15746), .A2(n_257_76_15747), .A3(
      n_257_76_15748), .A4(n_257_76_15749), .ZN(n_257_76_15750));
   NOR2_X1 i_257_76_15779 (.A1(n_257_76_15741), .A2(n_257_76_15750), .ZN(
      n_257_76_15751));
   NAND3_X1 i_257_76_15780 (.A1(n_257_76_15713), .A2(n_257_76_15737), .A3(
      n_257_76_15751), .ZN(n_257_76_15752));
   INV_X1 i_257_76_15781 (.A(n_257_76_15752), .ZN(n_257_76_15753));
   NAND2_X1 i_257_76_15782 (.A1(n_257_697), .A2(n_257_448), .ZN(n_257_76_15754));
   NAND3_X1 i_257_76_15783 (.A1(n_257_76_15753), .A2(n_257_76_15754), .A3(
      n_257_76_15712), .ZN(n_257_76_15755));
   INV_X1 i_257_76_15784 (.A(n_257_76_15755), .ZN(n_257_76_15756));
   NAND2_X1 i_257_76_15785 (.A1(n_257_28), .A2(n_257_76_15756), .ZN(
      n_257_76_15757));
   NAND3_X1 i_257_76_15786 (.A1(n_257_76_15725), .A2(n_257_76_15731), .A3(
      n_257_76_15757), .ZN(n_257_76_15758));
   INV_X1 i_257_76_15787 (.A(n_257_76_15712), .ZN(n_257_76_15759));
   INV_X1 i_257_76_15788 (.A(n_257_76_15726), .ZN(n_257_76_15760));
   INV_X1 i_257_76_15789 (.A(n_257_857), .ZN(n_257_76_15761));
   NOR2_X1 i_257_76_15790 (.A1(n_257_76_15760), .A2(n_257_76_15761), .ZN(
      n_257_76_15762));
   NAND4_X1 i_257_76_15791 (.A1(n_257_446), .A2(n_257_76_15748), .A3(
      n_257_76_15749), .A4(n_257_76_15762), .ZN(n_257_76_15763));
   INV_X1 i_257_76_15792 (.A(n_257_76_15763), .ZN(n_257_76_15764));
   NAND2_X1 i_257_76_15793 (.A1(n_257_76_15739), .A2(n_257_76_15747), .ZN(
      n_257_76_15765));
   INV_X1 i_257_76_15794 (.A(n_257_76_15765), .ZN(n_257_76_15766));
   NAND3_X1 i_257_76_15795 (.A1(n_257_76_15764), .A2(n_257_76_15766), .A3(
      n_257_76_15714), .ZN(n_257_76_15767));
   INV_X1 i_257_76_15796 (.A(n_257_76_15767), .ZN(n_257_76_15768));
   NAND2_X1 i_257_76_15797 (.A1(n_257_76_15768), .A2(n_257_76_15713), .ZN(
      n_257_76_15769));
   NOR2_X1 i_257_76_15798 (.A1(n_257_76_15759), .A2(n_257_76_15769), .ZN(
      n_257_76_15770));
   NAND2_X1 i_257_76_15799 (.A1(n_257_76_18070), .A2(n_257_76_15770), .ZN(
      n_257_76_15771));
   NAND2_X1 i_257_76_15800 (.A1(n_257_439), .A2(n_257_76_15726), .ZN(
      n_257_76_15772));
   INV_X1 i_257_76_15801 (.A(n_257_76_15772), .ZN(n_257_76_15773));
   NAND3_X1 i_257_76_15802 (.A1(n_257_76_15773), .A2(n_257_927), .A3(
      n_257_76_15748), .ZN(n_257_76_15774));
   INV_X1 i_257_76_15803 (.A(n_257_76_15774), .ZN(n_257_76_15775));
   NAND2_X1 i_257_76_15804 (.A1(n_257_76_15714), .A2(n_257_76_15775), .ZN(
      n_257_76_15776));
   INV_X1 i_257_76_15805 (.A(n_257_76_15776), .ZN(n_257_76_15777));
   NAND2_X1 i_257_76_15806 (.A1(n_257_76_15713), .A2(n_257_76_15777), .ZN(
      n_257_76_15778));
   INV_X1 i_257_76_15807 (.A(n_257_76_15778), .ZN(n_257_76_15779));
   NAND2_X1 i_257_76_15808 (.A1(n_257_76_15712), .A2(n_257_76_15779), .ZN(
      n_257_76_15780));
   INV_X1 i_257_76_15809 (.A(n_257_76_15780), .ZN(n_257_76_15781));
   NAND2_X1 i_257_76_15810 (.A1(n_257_76_18084), .A2(n_257_76_15781), .ZN(
      n_257_76_15782));
   NAND3_X1 i_257_76_15811 (.A1(n_257_76_15733), .A2(n_257_76_15734), .A3(
      n_257_76_15738), .ZN(n_257_76_15783));
   INV_X1 i_257_76_15812 (.A(n_257_76_15783), .ZN(n_257_76_15784));
   NAND2_X1 i_257_76_15813 (.A1(n_257_451), .A2(n_257_480), .ZN(n_257_76_15785));
   NAND3_X1 i_257_76_15814 (.A1(n_257_76_15785), .A2(n_257_76_15739), .A3(
      n_257_76_15740), .ZN(n_257_76_15786));
   INV_X1 i_257_76_15815 (.A(n_257_76_15786), .ZN(n_257_76_15787));
   NAND2_X1 i_257_76_15816 (.A1(n_257_427), .A2(n_257_220), .ZN(n_257_76_15788));
   NAND4_X1 i_257_76_15817 (.A1(n_257_76_15747), .A2(n_257_76_15748), .A3(
      n_257_76_15749), .A4(n_257_76_15788), .ZN(n_257_76_15789));
   INV_X1 i_257_76_15818 (.A(n_257_76_15789), .ZN(n_257_76_15790));
   NAND3_X1 i_257_76_15819 (.A1(n_257_76_15784), .A2(n_257_76_15787), .A3(
      n_257_76_15790), .ZN(n_257_76_15791));
   NAND2_X1 i_257_76_15820 (.A1(n_257_260), .A2(n_257_425), .ZN(n_257_76_15792));
   NAND2_X1 i_257_76_15821 (.A1(n_257_103), .A2(n_257_431), .ZN(n_257_76_15793));
   NAND4_X1 i_257_76_15822 (.A1(n_257_76_15792), .A2(n_257_76_15714), .A3(
      n_257_76_15793), .A4(n_257_76_15732), .ZN(n_257_76_15794));
   NOR2_X1 i_257_76_15823 (.A1(n_257_76_15791), .A2(n_257_76_15794), .ZN(
      n_257_76_15795));
   NAND2_X1 i_257_76_15824 (.A1(n_257_657), .A2(n_257_450), .ZN(n_257_76_15796));
   INV_X1 i_257_76_15825 (.A(n_257_76_15796), .ZN(n_257_76_15797));
   NAND2_X1 i_257_76_15826 (.A1(n_257_529), .A2(n_257_424), .ZN(n_257_76_15798));
   NAND2_X1 i_257_76_15827 (.A1(n_257_63), .A2(n_257_433), .ZN(n_257_76_15799));
   NAND2_X1 i_257_76_15828 (.A1(n_257_76_15798), .A2(n_257_76_15799), .ZN(
      n_257_76_15800));
   NOR2_X1 i_257_76_15829 (.A1(n_257_76_15797), .A2(n_257_76_15800), .ZN(
      n_257_76_15801));
   NAND2_X1 i_257_76_15830 (.A1(n_257_300), .A2(n_257_76_15744), .ZN(
      n_257_76_15802));
   NAND2_X1 i_257_76_15831 (.A1(n_257_432), .A2(n_257_625), .ZN(n_257_76_15803));
   NOR2_X1 i_257_76_15832 (.A1(n_257_1087), .A2(n_257_76_17476), .ZN(
      n_257_76_15804));
   INV_X1 i_257_76_15833 (.A(n_257_593), .ZN(n_257_76_15805));
   NAND2_X1 i_257_76_15834 (.A1(n_257_76_15805), .A2(n_257_442), .ZN(
      n_257_76_15806));
   OAI21_X1 i_257_76_15835 (.A(n_257_76_15806), .B1(n_257_428), .B2(
      n_257_76_17412), .ZN(n_257_76_15807));
   NAND3_X1 i_257_76_15836 (.A1(n_257_76_15803), .A2(n_257_76_15804), .A3(
      n_257_76_15807), .ZN(n_257_76_15808));
   NOR2_X1 i_257_76_15837 (.A1(n_257_76_15802), .A2(n_257_76_15808), .ZN(
      n_257_76_15809));
   NAND2_X1 i_257_76_15838 (.A1(n_257_561), .A2(n_257_426), .ZN(n_257_76_15810));
   NAND2_X1 i_257_76_15839 (.A1(n_257_141), .A2(n_257_430), .ZN(n_257_76_15811));
   NAND4_X1 i_257_76_15840 (.A1(n_257_76_15801), .A2(n_257_76_15809), .A3(
      n_257_76_15810), .A4(n_257_76_15811), .ZN(n_257_76_15812));
   INV_X1 i_257_76_15841 (.A(n_257_76_15812), .ZN(n_257_76_15813));
   NAND2_X1 i_257_76_15842 (.A1(n_257_180), .A2(n_257_429), .ZN(n_257_76_15814));
   NAND3_X1 i_257_76_15843 (.A1(n_257_76_15713), .A2(n_257_76_15813), .A3(
      n_257_76_15814), .ZN(n_257_76_15815));
   INV_X1 i_257_76_15844 (.A(n_257_76_15815), .ZN(n_257_76_15816));
   NAND4_X1 i_257_76_15845 (.A1(n_257_76_15795), .A2(n_257_76_15754), .A3(
      n_257_76_15712), .A4(n_257_76_15816), .ZN(n_257_76_15817));
   INV_X1 i_257_76_15846 (.A(n_257_76_15817), .ZN(n_257_76_15818));
   NAND2_X1 i_257_76_15847 (.A1(n_257_76_18066), .A2(n_257_76_15818), .ZN(
      n_257_76_15819));
   NAND3_X1 i_257_76_15848 (.A1(n_257_76_15771), .A2(n_257_76_15782), .A3(
      n_257_76_15819), .ZN(n_257_76_15820));
   NOR2_X1 i_257_76_15849 (.A1(n_257_76_15758), .A2(n_257_76_15820), .ZN(
      n_257_76_15821));
   NAND2_X1 i_257_76_15850 (.A1(n_257_991), .A2(n_257_76_15726), .ZN(
      n_257_76_15822));
   INV_X1 i_257_76_15851 (.A(n_257_76_15822), .ZN(n_257_76_15823));
   NAND2_X1 i_257_76_15852 (.A1(n_257_441), .A2(n_257_76_15823), .ZN(
      n_257_76_15824));
   INV_X1 i_257_76_15853 (.A(n_257_76_15824), .ZN(n_257_76_15825));
   NAND2_X1 i_257_76_15854 (.A1(n_257_76_15713), .A2(n_257_76_15825), .ZN(
      n_257_76_15826));
   INV_X1 i_257_76_15855 (.A(n_257_76_15826), .ZN(n_257_76_15827));
   NAND2_X1 i_257_76_15856 (.A1(n_257_76_15712), .A2(n_257_76_15827), .ZN(
      n_257_76_15828));
   INV_X1 i_257_76_15857 (.A(n_257_76_15828), .ZN(n_257_76_15829));
   NAND2_X1 i_257_76_15858 (.A1(n_257_76_18071), .A2(n_257_76_15829), .ZN(
      n_257_76_15830));
   NAND2_X1 i_257_76_15859 (.A1(n_257_76_15732), .A2(n_257_76_15733), .ZN(
      n_257_76_15831));
   NOR2_X1 i_257_76_15860 (.A1(n_257_76_15736), .A2(n_257_76_15831), .ZN(
      n_257_76_15832));
   NAND3_X1 i_257_76_15861 (.A1(n_257_76_15726), .A2(n_257_729), .A3(n_257_435), 
      .ZN(n_257_76_15833));
   INV_X1 i_257_76_15862 (.A(n_257_76_15833), .ZN(n_257_76_15834));
   NAND4_X1 i_257_76_15863 (.A1(n_257_76_15747), .A2(n_257_76_15748), .A3(
      n_257_76_15749), .A4(n_257_76_15834), .ZN(n_257_76_15835));
   NOR2_X1 i_257_76_15864 (.A1(n_257_76_15741), .A2(n_257_76_15835), .ZN(
      n_257_76_15836));
   NAND3_X1 i_257_76_15865 (.A1(n_257_76_15713), .A2(n_257_76_15832), .A3(
      n_257_76_15836), .ZN(n_257_76_15837));
   NOR2_X1 i_257_76_15866 (.A1(n_257_76_15837), .A2(n_257_76_15759), .ZN(
      n_257_76_15838));
   NAND2_X1 i_257_76_15867 (.A1(n_257_76_18078), .A2(n_257_76_15838), .ZN(
      n_257_76_15839));
   NAND4_X1 i_257_76_15868 (.A1(n_257_76_15738), .A2(n_257_76_15785), .A3(
      n_257_76_15739), .A4(n_257_76_15740), .ZN(n_257_76_15840));
   INV_X1 i_257_76_15869 (.A(n_257_76_15840), .ZN(n_257_76_15841));
   INV_X1 i_257_76_15870 (.A(n_257_76_15735), .ZN(n_257_76_15842));
   NAND2_X1 i_257_76_15871 (.A1(n_257_593), .A2(n_257_442), .ZN(n_257_76_15843));
   INV_X1 i_257_76_15872 (.A(n_257_76_15843), .ZN(n_257_76_15844));
   NAND2_X1 i_257_76_15873 (.A1(n_257_428), .A2(n_257_76_15844), .ZN(
      n_257_76_15845));
   NOR2_X1 i_257_76_15874 (.A1(n_257_76_15845), .A2(n_257_1087), .ZN(
      n_257_76_15846));
   NAND3_X1 i_257_76_15875 (.A1(n_257_76_15744), .A2(n_257_76_15846), .A3(
      n_257_76_15803), .ZN(n_257_76_15847));
   INV_X1 i_257_76_15876 (.A(n_257_76_15847), .ZN(n_257_76_15848));
   NAND4_X1 i_257_76_15877 (.A1(n_257_76_15749), .A2(n_257_76_15848), .A3(
      n_257_76_15796), .A4(n_257_76_15799), .ZN(n_257_76_15849));
   NAND3_X1 i_257_76_15878 (.A1(n_257_76_15747), .A2(n_257_76_15811), .A3(
      n_257_76_15748), .ZN(n_257_76_15850));
   NOR2_X1 i_257_76_15879 (.A1(n_257_76_15849), .A2(n_257_76_15850), .ZN(
      n_257_76_15851));
   NAND3_X1 i_257_76_15880 (.A1(n_257_76_15841), .A2(n_257_76_15842), .A3(
      n_257_76_15851), .ZN(n_257_76_15852));
   INV_X1 i_257_76_15881 (.A(n_257_76_15852), .ZN(n_257_76_15853));
   NAND2_X1 i_257_76_15882 (.A1(n_257_76_15714), .A2(n_257_76_15793), .ZN(
      n_257_76_15854));
   INV_X1 i_257_76_15883 (.A(n_257_76_15854), .ZN(n_257_76_15855));
   NAND3_X1 i_257_76_15884 (.A1(n_257_76_15713), .A2(n_257_76_15855), .A3(
      n_257_76_15814), .ZN(n_257_76_15856));
   INV_X1 i_257_76_15885 (.A(n_257_76_15856), .ZN(n_257_76_15857));
   NAND4_X1 i_257_76_15886 (.A1(n_257_76_15754), .A2(n_257_76_15853), .A3(
      n_257_76_15857), .A4(n_257_76_15712), .ZN(n_257_76_15858));
   INV_X1 i_257_76_15887 (.A(n_257_76_15858), .ZN(n_257_76_15859));
   NAND2_X1 i_257_76_15888 (.A1(n_257_76_18074), .A2(n_257_76_15859), .ZN(
      n_257_76_15860));
   NAND3_X1 i_257_76_15889 (.A1(n_257_76_15830), .A2(n_257_76_15839), .A3(
      n_257_76_15860), .ZN(n_257_76_15861));
   NAND2_X1 i_257_76_15890 (.A1(n_257_1087), .A2(n_257_442), .ZN(n_257_76_15862));
   INV_X1 i_257_76_15891 (.A(n_257_76_15862), .ZN(n_257_76_15863));
   NAND2_X1 i_257_76_15892 (.A1(n_257_13), .A2(n_257_76_15863), .ZN(
      n_257_76_15864));
   NAND2_X1 i_257_76_15893 (.A1(n_257_445), .A2(n_257_76_15726), .ZN(
      n_257_76_15865));
   INV_X1 i_257_76_15894 (.A(n_257_76_15865), .ZN(n_257_76_15866));
   NAND4_X1 i_257_76_15895 (.A1(n_257_76_15748), .A2(n_257_76_15749), .A3(
      n_257_889), .A4(n_257_76_15866), .ZN(n_257_76_15867));
   INV_X1 i_257_76_15896 (.A(n_257_76_15867), .ZN(n_257_76_15868));
   NAND3_X1 i_257_76_15897 (.A1(n_257_76_15868), .A2(n_257_76_15714), .A3(
      n_257_76_15739), .ZN(n_257_76_15869));
   INV_X1 i_257_76_15898 (.A(n_257_76_15869), .ZN(n_257_76_15870));
   NAND2_X1 i_257_76_15899 (.A1(n_257_76_15870), .A2(n_257_76_15713), .ZN(
      n_257_76_15871));
   NOR2_X1 i_257_76_15900 (.A1(n_257_76_15759), .A2(n_257_76_15871), .ZN(
      n_257_76_15872));
   NAND2_X1 i_257_76_15901 (.A1(n_257_76_18077), .A2(n_257_76_15872), .ZN(
      n_257_76_15873));
   NAND2_X1 i_257_76_15902 (.A1(n_257_76_15864), .A2(n_257_76_15873), .ZN(
      n_257_76_15874));
   NOR2_X1 i_257_76_15903 (.A1(n_257_76_15861), .A2(n_257_76_15874), .ZN(
      n_257_76_15875));
   NOR2_X1 i_257_76_15904 (.A1(n_257_1087), .A2(n_257_76_17564), .ZN(
      n_257_76_15876));
   NAND2_X1 i_257_76_15905 (.A1(n_257_76_15876), .A2(n_257_76_15807), .ZN(
      n_257_76_15877));
   INV_X1 i_257_76_15906 (.A(n_257_76_15877), .ZN(n_257_76_15878));
   NAND4_X1 i_257_76_15907 (.A1(n_257_76_15878), .A2(n_257_76_15799), .A3(
      n_257_76_15744), .A4(n_257_76_15803), .ZN(n_257_76_15879));
   INV_X1 i_257_76_15908 (.A(n_257_76_15879), .ZN(n_257_76_15880));
   NAND4_X1 i_257_76_15909 (.A1(n_257_76_15880), .A2(n_257_76_15811), .A3(
      n_257_561), .A4(n_257_76_15796), .ZN(n_257_76_15881));
   INV_X1 i_257_76_15910 (.A(n_257_76_15881), .ZN(n_257_76_15882));
   NAND3_X1 i_257_76_15911 (.A1(n_257_76_15882), .A2(n_257_76_15814), .A3(
      n_257_76_15714), .ZN(n_257_76_15883));
   INV_X1 i_257_76_15912 (.A(n_257_76_15713), .ZN(n_257_76_15884));
   NOR2_X1 i_257_76_15913 (.A1(n_257_76_15883), .A2(n_257_76_15884), .ZN(
      n_257_76_15885));
   NAND2_X1 i_257_76_15914 (.A1(n_257_76_15738), .A2(n_257_76_15785), .ZN(
      n_257_76_15886));
   INV_X1 i_257_76_15915 (.A(n_257_76_15886), .ZN(n_257_76_15887));
   NAND2_X1 i_257_76_15916 (.A1(n_257_76_15739), .A2(n_257_76_15740), .ZN(
      n_257_76_15888));
   INV_X1 i_257_76_15917 (.A(n_257_76_15888), .ZN(n_257_76_15889));
   NAND3_X1 i_257_76_15918 (.A1(n_257_76_15887), .A2(n_257_76_15889), .A3(
      n_257_76_15790), .ZN(n_257_76_15890));
   NAND4_X1 i_257_76_15919 (.A1(n_257_76_15793), .A2(n_257_76_15732), .A3(
      n_257_76_15733), .A4(n_257_76_15734), .ZN(n_257_76_15891));
   NOR2_X1 i_257_76_15920 (.A1(n_257_76_15890), .A2(n_257_76_15891), .ZN(
      n_257_76_15892));
   NAND4_X1 i_257_76_15921 (.A1(n_257_76_15885), .A2(n_257_76_15754), .A3(
      n_257_76_15712), .A4(n_257_76_15892), .ZN(n_257_76_15893));
   INV_X1 i_257_76_15922 (.A(n_257_76_15893), .ZN(n_257_76_15894));
   NAND2_X1 i_257_76_15923 (.A1(n_257_76_18076), .A2(n_257_76_15894), .ZN(
      n_257_76_15895));
   NAND2_X1 i_257_76_15924 (.A1(n_257_76_15733), .A2(n_257_76_15738), .ZN(
      n_257_76_15896));
   NOR2_X1 i_257_76_15925 (.A1(n_257_76_15736), .A2(n_257_76_15896), .ZN(
      n_257_76_15897));
   NAND3_X1 i_257_76_15926 (.A1(n_257_76_15739), .A2(n_257_76_15740), .A3(
      n_257_76_15747), .ZN(n_257_76_15898));
   NAND2_X1 i_257_76_15927 (.A1(n_257_436), .A2(n_257_76_15726), .ZN(
      n_257_76_15899));
   INV_X1 i_257_76_15928 (.A(n_257_76_15899), .ZN(n_257_76_15900));
   NAND4_X1 i_257_76_15929 (.A1(n_257_761), .A2(n_257_76_15748), .A3(
      n_257_76_15749), .A4(n_257_76_15900), .ZN(n_257_76_15901));
   NOR2_X1 i_257_76_15930 (.A1(n_257_76_15898), .A2(n_257_76_15901), .ZN(
      n_257_76_15902));
   NAND3_X1 i_257_76_15931 (.A1(n_257_76_15713), .A2(n_257_76_15897), .A3(
      n_257_76_15902), .ZN(n_257_76_15903));
   NOR2_X1 i_257_76_15932 (.A1(n_257_76_15903), .A2(n_257_76_15759), .ZN(
      n_257_76_15904));
   NAND2_X1 i_257_76_15933 (.A1(n_257_76_18069), .A2(n_257_76_15904), .ZN(
      n_257_76_15905));
   INV_X1 i_257_76_15934 (.A(n_257_1087), .ZN(n_257_76_15906));
   NAND2_X1 i_257_76_15935 (.A1(n_257_442), .A2(n_257_625), .ZN(n_257_76_15907));
   INV_X1 i_257_76_15936 (.A(n_257_76_15907), .ZN(n_257_76_15908));
   NAND3_X1 i_257_76_15937 (.A1(n_257_432), .A2(n_257_76_15906), .A3(
      n_257_76_15908), .ZN(n_257_76_15909));
   INV_X1 i_257_76_15938 (.A(n_257_76_15909), .ZN(n_257_76_15910));
   NAND3_X1 i_257_76_15939 (.A1(n_257_76_15799), .A2(n_257_76_15910), .A3(
      n_257_76_15744), .ZN(n_257_76_15911));
   INV_X1 i_257_76_15940 (.A(n_257_76_15911), .ZN(n_257_76_15912));
   NAND4_X1 i_257_76_15941 (.A1(n_257_76_15912), .A2(n_257_76_15748), .A3(
      n_257_76_15749), .A4(n_257_76_15796), .ZN(n_257_76_15913));
   NAND2_X1 i_257_76_15942 (.A1(n_257_76_15740), .A2(n_257_76_15747), .ZN(
      n_257_76_15914));
   NOR2_X1 i_257_76_15943 (.A1(n_257_76_15913), .A2(n_257_76_15914), .ZN(
      n_257_76_15915));
   NAND4_X1 i_257_76_15944 (.A1(n_257_76_15734), .A2(n_257_76_15738), .A3(
      n_257_76_15785), .A4(n_257_76_15739), .ZN(n_257_76_15916));
   INV_X1 i_257_76_15945 (.A(n_257_76_15916), .ZN(n_257_76_15917));
   NAND4_X1 i_257_76_15946 (.A1(n_257_76_15832), .A2(n_257_76_15713), .A3(
      n_257_76_15915), .A4(n_257_76_15917), .ZN(n_257_76_15918));
   INV_X1 i_257_76_15947 (.A(n_257_76_15918), .ZN(n_257_76_15919));
   NAND3_X1 i_257_76_15948 (.A1(n_257_76_15919), .A2(n_257_76_15754), .A3(
      n_257_76_15712), .ZN(n_257_76_15920));
   INV_X1 i_257_76_15949 (.A(n_257_76_15920), .ZN(n_257_76_15921));
   NAND2_X1 i_257_76_15950 (.A1(n_257_68), .A2(n_257_76_15921), .ZN(
      n_257_76_15922));
   NAND3_X1 i_257_76_15951 (.A1(n_257_76_15895), .A2(n_257_76_15905), .A3(
      n_257_76_15922), .ZN(n_257_76_15923));
   INV_X1 i_257_76_15952 (.A(n_257_437), .ZN(n_257_76_15924));
   NOR2_X1 i_257_76_15953 (.A1(n_257_76_15760), .A2(n_257_76_15924), .ZN(
      n_257_76_15925));
   NAND4_X1 i_257_76_15954 (.A1(n_257_76_15748), .A2(n_257_76_15749), .A3(
      n_257_825), .A4(n_257_76_15925), .ZN(n_257_76_15926));
   NOR2_X1 i_257_76_15955 (.A1(n_257_76_15765), .A2(n_257_76_15926), .ZN(
      n_257_76_15927));
   NAND2_X1 i_257_76_15956 (.A1(n_257_76_15714), .A2(n_257_76_15733), .ZN(
      n_257_76_15928));
   INV_X1 i_257_76_15957 (.A(n_257_76_15928), .ZN(n_257_76_15929));
   NAND3_X1 i_257_76_15958 (.A1(n_257_76_15927), .A2(n_257_76_15713), .A3(
      n_257_76_15929), .ZN(n_257_76_15930));
   NOR2_X1 i_257_76_15959 (.A1(n_257_76_15759), .A2(n_257_76_15930), .ZN(
      n_257_76_15931));
   NAND2_X1 i_257_76_15960 (.A1(n_257_22), .A2(n_257_76_15931), .ZN(
      n_257_76_15932));
   NAND2_X1 i_257_76_15961 (.A1(n_257_444), .A2(n_257_76_15726), .ZN(
      n_257_76_15933));
   INV_X1 i_257_76_15962 (.A(n_257_76_15933), .ZN(n_257_76_15934));
   NAND2_X1 i_257_76_15963 (.A1(n_257_1023), .A2(n_257_76_15934), .ZN(
      n_257_76_15935));
   INV_X1 i_257_76_15964 (.A(n_257_76_15935), .ZN(n_257_76_15936));
   NAND2_X1 i_257_76_15965 (.A1(n_257_76_15712), .A2(n_257_76_15936), .ZN(
      n_257_76_15937));
   INV_X1 i_257_76_15966 (.A(n_257_76_15937), .ZN(n_257_76_15938));
   NAND2_X1 i_257_76_15967 (.A1(n_257_76_18075), .A2(n_257_76_15938), .ZN(
      n_257_76_15939));
   NAND2_X1 i_257_76_15968 (.A1(n_257_76_15932), .A2(n_257_76_15939), .ZN(
      n_257_76_15940));
   NOR2_X1 i_257_76_15969 (.A1(n_257_76_15923), .A2(n_257_76_15940), .ZN(
      n_257_76_15941));
   NAND3_X1 i_257_76_15970 (.A1(n_257_76_15821), .A2(n_257_76_15875), .A3(
      n_257_76_15941), .ZN(n_257_76_15942));
   INV_X1 i_257_76_15971 (.A(n_257_76_15942), .ZN(n_257_76_15943));
   NAND4_X1 i_257_76_15972 (.A1(n_257_76_15744), .A2(n_257_76_15726), .A3(
      n_257_63), .A4(n_257_433), .ZN(n_257_76_15944));
   INV_X1 i_257_76_15973 (.A(n_257_76_15944), .ZN(n_257_76_15945));
   NAND4_X1 i_257_76_15974 (.A1(n_257_76_15748), .A2(n_257_76_15749), .A3(
      n_257_76_15945), .A4(n_257_76_15796), .ZN(n_257_76_15946));
   NOR2_X1 i_257_76_15975 (.A1(n_257_76_15946), .A2(n_257_76_15914), .ZN(
      n_257_76_15947));
   NAND4_X1 i_257_76_15976 (.A1(n_257_76_15832), .A2(n_257_76_15713), .A3(
      n_257_76_15947), .A4(n_257_76_15917), .ZN(n_257_76_15948));
   INV_X1 i_257_76_15977 (.A(n_257_76_15948), .ZN(n_257_76_15949));
   NAND3_X1 i_257_76_15978 (.A1(n_257_76_15949), .A2(n_257_76_15754), .A3(
      n_257_76_15712), .ZN(n_257_76_15950));
   INV_X1 i_257_76_15979 (.A(n_257_76_15950), .ZN(n_257_76_15951));
   NAND2_X1 i_257_76_15980 (.A1(n_257_76_18081), .A2(n_257_76_15951), .ZN(
      n_257_76_15952));
   NAND3_X1 i_257_76_15981 (.A1(n_257_76_15732), .A2(n_257_76_15733), .A3(
      n_257_76_15738), .ZN(n_257_76_15953));
   NOR2_X1 i_257_76_15982 (.A1(n_257_76_15953), .A2(n_257_76_15736), .ZN(
      n_257_76_15954));
   NAND2_X1 i_257_76_15983 (.A1(n_257_442), .A2(n_257_665), .ZN(n_257_76_15955));
   NOR2_X1 i_257_76_15984 (.A1(n_257_1087), .A2(n_257_76_15955), .ZN(
      n_257_76_15956));
   NAND2_X1 i_257_76_15985 (.A1(n_257_76_15744), .A2(n_257_76_15956), .ZN(
      n_257_76_15957));
   INV_X1 i_257_76_15986 (.A(n_257_76_15957), .ZN(n_257_76_15958));
   NAND4_X1 i_257_76_15987 (.A1(n_257_449), .A2(n_257_76_15748), .A3(
      n_257_76_15749), .A4(n_257_76_15958), .ZN(n_257_76_15959));
   NOR2_X1 i_257_76_15988 (.A1(n_257_76_15898), .A2(n_257_76_15959), .ZN(
      n_257_76_15960));
   NAND3_X1 i_257_76_15989 (.A1(n_257_76_15954), .A2(n_257_76_15713), .A3(
      n_257_76_15960), .ZN(n_257_76_15961));
   INV_X1 i_257_76_15990 (.A(n_257_76_15961), .ZN(n_257_76_15962));
   NAND3_X1 i_257_76_15991 (.A1(n_257_76_15962), .A2(n_257_76_15754), .A3(
      n_257_76_15712), .ZN(n_257_76_15963));
   INV_X1 i_257_76_15992 (.A(n_257_76_15963), .ZN(n_257_76_15964));
   NAND2_X1 i_257_76_15993 (.A1(n_257_76_18083), .A2(n_257_76_15964), .ZN(
      n_257_76_15965));
   NAND3_X1 i_257_76_15994 (.A1(n_257_180), .A2(n_257_76_15732), .A3(
      n_257_76_15733), .ZN(n_257_76_15966));
   INV_X1 i_257_76_15995 (.A(n_257_76_15966), .ZN(n_257_76_15967));
   NAND3_X1 i_257_76_15996 (.A1(n_257_76_15713), .A2(n_257_76_15855), .A3(
      n_257_76_15967), .ZN(n_257_76_15968));
   INV_X1 i_257_76_15997 (.A(n_257_76_15968), .ZN(n_257_76_15969));
   INV_X1 i_257_76_15998 (.A(n_257_76_15914), .ZN(n_257_76_15970));
   NAND3_X1 i_257_76_15999 (.A1(n_257_76_15811), .A2(n_257_76_15748), .A3(
      n_257_76_15749), .ZN(n_257_76_15971));
   INV_X1 i_257_76_16000 (.A(n_257_76_15971), .ZN(n_257_76_15972));
   NAND2_X1 i_257_76_16001 (.A1(n_257_76_15799), .A2(n_257_76_15744), .ZN(
      n_257_76_15973));
   INV_X1 i_257_76_16002 (.A(n_257_76_15973), .ZN(n_257_76_15974));
   NAND3_X1 i_257_76_16003 (.A1(n_257_76_15803), .A2(n_257_76_15726), .A3(
      n_257_429), .ZN(n_257_76_15975));
   INV_X1 i_257_76_16004 (.A(n_257_76_15975), .ZN(n_257_76_15976));
   NAND3_X1 i_257_76_16005 (.A1(n_257_76_15974), .A2(n_257_76_15796), .A3(
      n_257_76_15976), .ZN(n_257_76_15977));
   INV_X1 i_257_76_16006 (.A(n_257_76_15977), .ZN(n_257_76_15978));
   NAND3_X1 i_257_76_16007 (.A1(n_257_76_15970), .A2(n_257_76_15972), .A3(
      n_257_76_15978), .ZN(n_257_76_15979));
   NOR2_X1 i_257_76_16008 (.A1(n_257_76_15979), .A2(n_257_76_15916), .ZN(
      n_257_76_15980));
   NAND4_X1 i_257_76_16009 (.A1(n_257_76_15754), .A2(n_257_76_15969), .A3(
      n_257_76_15980), .A4(n_257_76_15712), .ZN(n_257_76_15981));
   INV_X1 i_257_76_16010 (.A(n_257_76_15981), .ZN(n_257_76_15982));
   NAND2_X1 i_257_76_16011 (.A1(n_257_76_18061), .A2(n_257_76_15982), .ZN(
      n_257_76_15983));
   NAND3_X1 i_257_76_16012 (.A1(n_257_76_15952), .A2(n_257_76_15965), .A3(
      n_257_76_15983), .ZN(n_257_76_15984));
   INV_X1 i_257_76_16013 (.A(n_257_76_15984), .ZN(n_257_76_15985));
   NAND2_X1 i_257_76_16014 (.A1(n_257_442), .A2(n_257_895), .ZN(n_257_76_15986));
   NOR2_X1 i_257_76_16015 (.A1(n_257_1087), .A2(n_257_76_15986), .ZN(
      n_257_76_15987));
   NAND2_X1 i_257_76_16016 (.A1(n_257_438), .A2(n_257_76_15987), .ZN(
      n_257_76_15988));
   INV_X1 i_257_76_16017 (.A(n_257_76_15988), .ZN(n_257_76_15989));
   NAND3_X1 i_257_76_16018 (.A1(n_257_76_15739), .A2(n_257_76_15748), .A3(
      n_257_76_15989), .ZN(n_257_76_15990));
   INV_X1 i_257_76_16019 (.A(n_257_76_15990), .ZN(n_257_76_15991));
   NAND2_X1 i_257_76_16020 (.A1(n_257_76_15991), .A2(n_257_76_15714), .ZN(
      n_257_76_15992));
   NOR2_X1 i_257_76_16021 (.A1(n_257_76_15884), .A2(n_257_76_15992), .ZN(
      n_257_76_15993));
   NAND2_X1 i_257_76_16022 (.A1(n_257_76_15712), .A2(n_257_76_15993), .ZN(
      n_257_76_15994));
   INV_X1 i_257_76_16023 (.A(n_257_76_15994), .ZN(n_257_76_15995));
   NAND2_X1 i_257_76_16024 (.A1(n_257_76_18067), .A2(n_257_76_15995), .ZN(
      n_257_76_15996));
   NAND2_X1 i_257_76_16025 (.A1(n_257_338), .A2(n_257_422), .ZN(n_257_76_15997));
   NAND2_X1 i_257_76_16026 (.A1(n_257_428), .A2(n_257_593), .ZN(n_257_76_15998));
   NAND2_X1 i_257_76_16027 (.A1(n_257_76_15998), .A2(n_257_76_15906), .ZN(
      n_257_76_15999));
   INV_X1 i_257_76_16028 (.A(n_257_76_15999), .ZN(n_257_76_16000));
   NAND2_X1 i_257_76_16029 (.A1(n_257_442), .A2(n_257_497), .ZN(n_257_76_16001));
   INV_X1 i_257_76_16030 (.A(n_257_76_16001), .ZN(n_257_76_16002));
   NAND2_X1 i_257_76_16031 (.A1(n_257_420), .A2(n_257_76_16002), .ZN(
      n_257_76_16003));
   INV_X1 i_257_76_16032 (.A(n_257_76_16003), .ZN(n_257_76_16004));
   NAND4_X1 i_257_76_16033 (.A1(n_257_76_15997), .A2(n_257_76_16000), .A3(
      n_257_76_15803), .A4(n_257_76_16004), .ZN(n_257_76_16005));
   NOR2_X1 i_257_76_16034 (.A1(n_257_76_16005), .A2(n_257_76_15973), .ZN(
      n_257_76_16006));
   NAND2_X1 i_257_76_16035 (.A1(n_257_76_15749), .A2(n_257_76_15796), .ZN(
      n_257_76_16007));
   INV_X1 i_257_76_16036 (.A(n_257_76_16007), .ZN(n_257_76_16008));
   NAND2_X1 i_257_76_16037 (.A1(n_257_300), .A2(n_257_423), .ZN(n_257_76_16009));
   NAND3_X1 i_257_76_16038 (.A1(n_257_76_15788), .A2(n_257_76_16009), .A3(
      n_257_76_15798), .ZN(n_257_76_16010));
   INV_X1 i_257_76_16039 (.A(n_257_76_16010), .ZN(n_257_76_16011));
   NAND3_X1 i_257_76_16040 (.A1(n_257_76_16006), .A2(n_257_76_16008), .A3(
      n_257_76_16011), .ZN(n_257_76_16012));
   NAND4_X1 i_257_76_16041 (.A1(n_257_76_15810), .A2(n_257_76_15747), .A3(
      n_257_76_15811), .A4(n_257_76_15748), .ZN(n_257_76_16013));
   NOR2_X1 i_257_76_16042 (.A1(n_257_76_16012), .A2(n_257_76_16013), .ZN(
      n_257_76_16014));
   NAND3_X1 i_257_76_16043 (.A1(n_257_76_16014), .A2(n_257_76_15713), .A3(
      n_257_76_15814), .ZN(n_257_76_16015));
   INV_X1 i_257_76_16044 (.A(n_257_76_16015), .ZN(n_257_76_16016));
   INV_X1 i_257_76_16045 (.A(n_257_76_15831), .ZN(n_257_76_16017));
   NAND2_X1 i_257_76_16046 (.A1(n_257_76_15734), .A2(n_257_76_15738), .ZN(
      n_257_76_16018));
   INV_X1 i_257_76_16047 (.A(n_257_76_16018), .ZN(n_257_76_16019));
   NAND3_X1 i_257_76_16048 (.A1(n_257_76_15787), .A2(n_257_76_16017), .A3(
      n_257_76_16019), .ZN(n_257_76_16020));
   NAND2_X1 i_257_76_16049 (.A1(n_257_377), .A2(n_257_421), .ZN(n_257_76_16021));
   NAND4_X1 i_257_76_16050 (.A1(n_257_76_15792), .A2(n_257_76_15714), .A3(
      n_257_76_15793), .A4(n_257_76_16021), .ZN(n_257_76_16022));
   NOR2_X1 i_257_76_16051 (.A1(n_257_76_16020), .A2(n_257_76_16022), .ZN(
      n_257_76_16023));
   NAND4_X1 i_257_76_16052 (.A1(n_257_76_15754), .A2(n_257_76_16016), .A3(
      n_257_76_16023), .A4(n_257_76_15712), .ZN(n_257_76_16024));
   INV_X1 i_257_76_16053 (.A(n_257_76_16024), .ZN(n_257_76_16025));
   NAND2_X1 i_257_76_16054 (.A1(n_257_76_18073), .A2(n_257_76_16025), .ZN(
      n_257_76_16026));
   NAND3_X1 i_257_76_16055 (.A1(n_257_76_15738), .A2(n_257_76_15785), .A3(
      n_257_76_15739), .ZN(n_257_76_16027));
   NOR2_X1 i_257_76_16056 (.A1(n_257_76_15735), .A2(n_257_76_16027), .ZN(
      n_257_76_16028));
   NAND2_X1 i_257_76_16057 (.A1(n_257_141), .A2(n_257_76_15799), .ZN(
      n_257_76_16029));
   INV_X1 i_257_76_16058 (.A(n_257_76_16029), .ZN(n_257_76_16030));
   NAND4_X1 i_257_76_16059 (.A1(n_257_76_15744), .A2(n_257_76_15803), .A3(
      n_257_76_15726), .A4(n_257_430), .ZN(n_257_76_16031));
   INV_X1 i_257_76_16060 (.A(n_257_76_16031), .ZN(n_257_76_16032));
   NAND4_X1 i_257_76_16061 (.A1(n_257_76_16030), .A2(n_257_76_16032), .A3(
      n_257_76_15749), .A4(n_257_76_15796), .ZN(n_257_76_16033));
   NAND3_X1 i_257_76_16062 (.A1(n_257_76_15740), .A2(n_257_76_15747), .A3(
      n_257_76_15748), .ZN(n_257_76_16034));
   NOR2_X1 i_257_76_16063 (.A1(n_257_76_16033), .A2(n_257_76_16034), .ZN(
      n_257_76_16035));
   NAND4_X1 i_257_76_16064 (.A1(n_257_76_16028), .A2(n_257_76_15713), .A3(
      n_257_76_15855), .A4(n_257_76_16035), .ZN(n_257_76_16036));
   INV_X1 i_257_76_16065 (.A(n_257_76_16036), .ZN(n_257_76_16037));
   NAND3_X1 i_257_76_16066 (.A1(n_257_76_16037), .A2(n_257_76_15754), .A3(
      n_257_76_15712), .ZN(n_257_76_16038));
   INV_X1 i_257_76_16067 (.A(n_257_76_16038), .ZN(n_257_76_16039));
   NAND2_X1 i_257_76_16068 (.A1(n_257_76_18068), .A2(n_257_76_16039), .ZN(
      n_257_76_16040));
   NAND3_X1 i_257_76_16069 (.A1(n_257_76_15996), .A2(n_257_76_16026), .A3(
      n_257_76_16040), .ZN(n_257_76_16041));
   INV_X1 i_257_76_16070 (.A(n_257_76_16041), .ZN(n_257_76_16042));
   NAND2_X1 i_257_76_16071 (.A1(n_257_793), .A2(n_257_442), .ZN(n_257_76_16043));
   NOR2_X1 i_257_76_16072 (.A1(n_257_1087), .A2(n_257_76_16043), .ZN(
      n_257_76_16044));
   NAND4_X1 i_257_76_16073 (.A1(n_257_447), .A2(n_257_76_15748), .A3(
      n_257_76_15749), .A4(n_257_76_16044), .ZN(n_257_76_16045));
   NOR2_X1 i_257_76_16074 (.A1(n_257_76_15898), .A2(n_257_76_16045), .ZN(
      n_257_76_16046));
   NAND3_X1 i_257_76_16075 (.A1(n_257_76_16046), .A2(n_257_76_15713), .A3(
      n_257_76_15929), .ZN(n_257_76_16047));
   NOR2_X1 i_257_76_16076 (.A1(n_257_76_15759), .A2(n_257_76_16047), .ZN(
      n_257_76_16048));
   NAND3_X1 i_257_76_16077 (.A1(n_257_76_15785), .A2(n_257_76_15739), .A3(
      n_257_103), .ZN(n_257_76_16049));
   NOR2_X1 i_257_76_16078 (.A1(n_257_76_15783), .A2(n_257_76_16049), .ZN(
      n_257_76_16050));
   NAND2_X1 i_257_76_16079 (.A1(n_257_76_15714), .A2(n_257_76_15732), .ZN(
      n_257_76_16051));
   INV_X1 i_257_76_16080 (.A(n_257_76_16051), .ZN(n_257_76_16052));
   NAND3_X1 i_257_76_16081 (.A1(n_257_76_15803), .A2(n_257_76_15726), .A3(
      n_257_431), .ZN(n_257_76_16053));
   INV_X1 i_257_76_16082 (.A(n_257_76_16053), .ZN(n_257_76_16054));
   NAND4_X1 i_257_76_16083 (.A1(n_257_76_15749), .A2(n_257_76_15974), .A3(
      n_257_76_15796), .A4(n_257_76_16054), .ZN(n_257_76_16055));
   NOR2_X1 i_257_76_16084 (.A1(n_257_76_16034), .A2(n_257_76_16055), .ZN(
      n_257_76_16056));
   NAND4_X1 i_257_76_16085 (.A1(n_257_76_16050), .A2(n_257_76_15713), .A3(
      n_257_76_16052), .A4(n_257_76_16056), .ZN(n_257_76_16057));
   INV_X1 i_257_76_16086 (.A(n_257_76_16057), .ZN(n_257_76_16058));
   NAND3_X1 i_257_76_16087 (.A1(n_257_76_16058), .A2(n_257_76_15754), .A3(
      n_257_76_15712), .ZN(n_257_76_16059));
   INV_X1 i_257_76_16088 (.A(n_257_76_16059), .ZN(n_257_76_16060));
   AOI22_X1 i_257_76_16089 (.A1(n_257_76_18085), .A2(n_257_76_16048), .B1(
      n_257_76_18080), .B2(n_257_76_16060), .ZN(n_257_76_16061));
   NAND3_X1 i_257_76_16090 (.A1(n_257_76_15985), .A2(n_257_76_16042), .A3(
      n_257_76_16061), .ZN(n_257_76_16062));
   NAND4_X1 i_257_76_16091 (.A1(n_257_76_15714), .A2(n_257_76_15732), .A3(
      n_257_76_15733), .A4(n_257_76_15738), .ZN(n_257_76_16063));
   NAND4_X1 i_257_76_16092 (.A1(n_257_76_15748), .A2(n_257_76_17980), .A3(
      n_257_76_15749), .A4(n_257_448), .ZN(n_257_76_16064));
   INV_X1 i_257_76_16093 (.A(n_257_76_16064), .ZN(n_257_76_16065));
   NAND3_X1 i_257_76_16094 (.A1(n_257_76_16065), .A2(n_257_76_15970), .A3(
      n_257_76_15739), .ZN(n_257_76_16066));
   NOR2_X1 i_257_76_16095 (.A1(n_257_76_16063), .A2(n_257_76_16066), .ZN(
      n_257_76_16067));
   NAND4_X1 i_257_76_16096 (.A1(n_257_76_16067), .A2(n_257_76_15712), .A3(
      n_257_697), .A4(n_257_76_15713), .ZN(n_257_76_16068));
   INV_X1 i_257_76_16097 (.A(n_257_76_16068), .ZN(n_257_76_16069));
   NAND2_X1 i_257_76_16098 (.A1(n_257_76_18079), .A2(n_257_76_16069), .ZN(
      n_257_76_16070));
   NAND2_X1 i_257_76_16099 (.A1(n_257_76_15814), .A2(n_257_76_15714), .ZN(
      n_257_76_16071));
   INV_X1 i_257_76_16100 (.A(n_257_76_16071), .ZN(n_257_76_16072));
   NAND4_X1 i_257_76_16101 (.A1(n_257_76_15733), .A2(n_257_76_15734), .A3(
      n_257_76_15738), .A4(n_257_76_15785), .ZN(n_257_76_16073));
   INV_X1 i_257_76_16102 (.A(n_257_76_16073), .ZN(n_257_76_16074));
   NAND3_X1 i_257_76_16103 (.A1(n_257_76_16072), .A2(n_257_76_15713), .A3(
      n_257_76_16074), .ZN(n_257_76_16075));
   INV_X1 i_257_76_16104 (.A(n_257_76_16075), .ZN(n_257_76_16076));
   NAND4_X1 i_257_76_16105 (.A1(n_257_76_15747), .A2(n_257_76_15811), .A3(
      n_257_76_15748), .A4(n_257_76_15749), .ZN(n_257_76_16077));
   NOR2_X1 i_257_76_16106 (.A1(n_257_1087), .A2(n_257_76_17778), .ZN(
      n_257_76_16078));
   NAND3_X1 i_257_76_16107 (.A1(n_257_76_15803), .A2(n_257_76_16078), .A3(
      n_257_76_15807), .ZN(n_257_76_16079));
   INV_X1 i_257_76_16108 (.A(n_257_76_16079), .ZN(n_257_76_16080));
   NAND4_X1 i_257_76_16109 (.A1(n_257_76_15974), .A2(n_257_76_16080), .A3(
      n_257_76_15796), .A4(n_257_76_15788), .ZN(n_257_76_16081));
   NOR2_X1 i_257_76_16110 (.A1(n_257_76_16077), .A2(n_257_76_16081), .ZN(
      n_257_76_16082));
   NAND2_X1 i_257_76_16111 (.A1(n_257_76_15793), .A2(n_257_260), .ZN(
      n_257_76_16083));
   INV_X1 i_257_76_16112 (.A(n_257_76_16083), .ZN(n_257_76_16084));
   NAND4_X1 i_257_76_16113 (.A1(n_257_76_15732), .A2(n_257_76_15739), .A3(
      n_257_76_15740), .A4(n_257_76_15810), .ZN(n_257_76_16085));
   INV_X1 i_257_76_16114 (.A(n_257_76_16085), .ZN(n_257_76_16086));
   NAND3_X1 i_257_76_16115 (.A1(n_257_76_16082), .A2(n_257_76_16084), .A3(
      n_257_76_16086), .ZN(n_257_76_16087));
   INV_X1 i_257_76_16116 (.A(n_257_76_16087), .ZN(n_257_76_16088));
   NAND4_X1 i_257_76_16117 (.A1(n_257_76_15754), .A2(n_257_76_16076), .A3(
      n_257_76_16088), .A4(n_257_76_15712), .ZN(n_257_76_16089));
   INV_X1 i_257_76_16118 (.A(n_257_76_16089), .ZN(n_257_76_16090));
   NAND2_X1 i_257_76_16119 (.A1(n_257_76_18064), .A2(n_257_76_16090), .ZN(
      n_257_76_16091));
   NAND3_X1 i_257_76_16120 (.A1(n_257_76_15796), .A2(n_257_76_15788), .A3(
      n_257_76_16009), .ZN(n_257_76_16092));
   INV_X1 i_257_76_16121 (.A(n_257_76_16092), .ZN(n_257_76_16093));
   NAND3_X1 i_257_76_16122 (.A1(n_257_76_15798), .A2(n_257_76_15799), .A3(
      n_257_76_15744), .ZN(n_257_76_16094));
   NOR2_X1 i_257_76_16123 (.A1(n_257_76_17792), .A2(n_257_1087), .ZN(
      n_257_76_16095));
   NAND4_X1 i_257_76_16124 (.A1(n_257_76_15997), .A2(n_257_76_16095), .A3(
      n_257_76_15803), .A4(n_257_76_15807), .ZN(n_257_76_16096));
   NOR2_X1 i_257_76_16125 (.A1(n_257_76_16094), .A2(n_257_76_16096), .ZN(
      n_257_76_16097));
   NAND2_X1 i_257_76_16126 (.A1(n_257_76_16093), .A2(n_257_76_16097), .ZN(
      n_257_76_16098));
   NOR2_X1 i_257_76_16127 (.A1(n_257_76_16098), .A2(n_257_76_16077), .ZN(
      n_257_76_16099));
   NAND2_X1 i_257_76_16128 (.A1(n_257_76_15792), .A2(n_257_76_15793), .ZN(
      n_257_76_16100));
   INV_X1 i_257_76_16129 (.A(n_257_76_16100), .ZN(n_257_76_16101));
   NAND2_X1 i_257_76_16130 (.A1(n_257_76_15732), .A2(n_257_76_15739), .ZN(
      n_257_76_16102));
   NAND3_X1 i_257_76_16131 (.A1(n_257_76_15740), .A2(n_257_377), .A3(
      n_257_76_15810), .ZN(n_257_76_16103));
   NOR2_X1 i_257_76_16132 (.A1(n_257_76_16102), .A2(n_257_76_16103), .ZN(
      n_257_76_16104));
   NAND3_X1 i_257_76_16133 (.A1(n_257_76_16099), .A2(n_257_76_16101), .A3(
      n_257_76_16104), .ZN(n_257_76_16105));
   INV_X1 i_257_76_16134 (.A(n_257_76_16105), .ZN(n_257_76_16106));
   NAND4_X1 i_257_76_16135 (.A1(n_257_76_16106), .A2(n_257_76_15754), .A3(
      n_257_76_16076), .A4(n_257_76_15712), .ZN(n_257_76_16107));
   INV_X1 i_257_76_16136 (.A(n_257_76_16107), .ZN(n_257_76_16108));
   NAND2_X1 i_257_76_16137 (.A1(n_257_76_18082), .A2(n_257_76_16108), .ZN(
      n_257_76_16109));
   NAND3_X1 i_257_76_16138 (.A1(n_257_76_16070), .A2(n_257_76_16091), .A3(
      n_257_76_16109), .ZN(n_257_76_16110));
   INV_X1 i_257_76_16139 (.A(n_257_76_16110), .ZN(n_257_76_16111));
   NAND2_X1 i_257_76_16140 (.A1(n_257_220), .A2(n_257_76_15906), .ZN(
      n_257_76_16112));
   INV_X1 i_257_76_16141 (.A(n_257_76_16112), .ZN(n_257_76_16113));
   NAND4_X1 i_257_76_16142 (.A1(n_257_76_15744), .A2(n_257_76_16113), .A3(
      n_257_76_15803), .A4(n_257_76_15807), .ZN(n_257_76_16114));
   INV_X1 i_257_76_16143 (.A(n_257_76_16114), .ZN(n_257_76_16115));
   NAND2_X1 i_257_76_16144 (.A1(n_257_76_15799), .A2(n_257_427), .ZN(
      n_257_76_16116));
   INV_X1 i_257_76_16145 (.A(n_257_76_16116), .ZN(n_257_76_16117));
   NAND4_X1 i_257_76_16146 (.A1(n_257_76_15811), .A2(n_257_76_16115), .A3(
      n_257_76_16117), .A4(n_257_76_15796), .ZN(n_257_76_16118));
   INV_X1 i_257_76_16147 (.A(n_257_76_16118), .ZN(n_257_76_16119));
   NAND3_X1 i_257_76_16148 (.A1(n_257_76_15814), .A2(n_257_76_16119), .A3(
      n_257_76_15714), .ZN(n_257_76_16120));
   NOR2_X1 i_257_76_16149 (.A1(n_257_76_16120), .A2(n_257_76_15884), .ZN(
      n_257_76_16121));
   NAND3_X1 i_257_76_16150 (.A1(n_257_76_15747), .A2(n_257_76_15748), .A3(
      n_257_76_15749), .ZN(n_257_76_16122));
   INV_X1 i_257_76_16151 (.A(n_257_76_16122), .ZN(n_257_76_16123));
   NAND3_X1 i_257_76_16152 (.A1(n_257_76_15887), .A2(n_257_76_15889), .A3(
      n_257_76_16123), .ZN(n_257_76_16124));
   NOR2_X1 i_257_76_16153 (.A1(n_257_76_16124), .A2(n_257_76_15891), .ZN(
      n_257_76_16125));
   NAND4_X1 i_257_76_16154 (.A1(n_257_76_16121), .A2(n_257_76_15754), .A3(
      n_257_76_16125), .A4(n_257_76_15712), .ZN(n_257_76_16126));
   INV_X1 i_257_76_16155 (.A(n_257_76_16126), .ZN(n_257_76_16127));
   NAND2_X1 i_257_76_16156 (.A1(n_257_76_18065), .A2(n_257_76_16127), .ZN(
      n_257_76_16128));
   NAND4_X1 i_257_76_16157 (.A1(n_257_76_15738), .A2(n_257_76_15739), .A3(
      n_257_76_15740), .A4(n_257_76_15747), .ZN(n_257_76_16129));
   NAND2_X1 i_257_76_16158 (.A1(n_257_451), .A2(n_257_76_15748), .ZN(
      n_257_76_16130));
   INV_X1 i_257_76_16159 (.A(n_257_76_16130), .ZN(n_257_76_16131));
   NAND2_X1 i_257_76_16160 (.A1(n_257_76_15749), .A2(n_257_76_17980), .ZN(
      n_257_76_16132));
   INV_X1 i_257_76_16161 (.A(n_257_76_16132), .ZN(n_257_76_16133));
   NAND2_X1 i_257_76_16162 (.A1(n_257_76_15796), .A2(n_257_480), .ZN(
      n_257_76_16134));
   INV_X1 i_257_76_16163 (.A(n_257_76_16134), .ZN(n_257_76_16135));
   NAND3_X1 i_257_76_16164 (.A1(n_257_76_16131), .A2(n_257_76_16133), .A3(
      n_257_76_16135), .ZN(n_257_76_16136));
   NOR2_X1 i_257_76_16165 (.A1(n_257_76_16129), .A2(n_257_76_16136), .ZN(
      n_257_76_16137));
   NAND3_X1 i_257_76_16166 (.A1(n_257_76_16137), .A2(n_257_76_15713), .A3(
      n_257_76_15737), .ZN(n_257_76_16138));
   INV_X1 i_257_76_16167 (.A(n_257_76_16138), .ZN(n_257_76_16139));
   NAND3_X1 i_257_76_16168 (.A1(n_257_76_16139), .A2(n_257_76_15754), .A3(
      n_257_76_15712), .ZN(n_257_76_16140));
   INV_X1 i_257_76_16169 (.A(n_257_76_16140), .ZN(n_257_76_16141));
   NAND2_X1 i_257_76_16170 (.A1(n_257_76_18063), .A2(n_257_76_16141), .ZN(
      n_257_76_16142));
   NAND4_X1 i_257_76_16171 (.A1(n_257_76_15814), .A2(n_257_76_15792), .A3(
      n_257_76_15714), .A4(n_257_76_15793), .ZN(n_257_76_16143));
   NOR2_X1 i_257_76_16172 (.A1(n_257_76_16143), .A2(n_257_76_15884), .ZN(
      n_257_76_16144));
   INV_X1 i_257_76_16173 (.A(n_257_424), .ZN(n_257_76_16145));
   NOR2_X1 i_257_76_16174 (.A1(n_257_76_16145), .A2(n_257_1087), .ZN(
      n_257_76_16146));
   NAND3_X1 i_257_76_16175 (.A1(n_257_76_16146), .A2(n_257_529), .A3(
      n_257_76_15807), .ZN(n_257_76_16147));
   INV_X1 i_257_76_16176 (.A(n_257_76_16147), .ZN(n_257_76_16148));
   NAND3_X1 i_257_76_16177 (.A1(n_257_76_15748), .A2(n_257_76_15749), .A3(
      n_257_76_16148), .ZN(n_257_76_16149));
   NAND2_X1 i_257_76_16178 (.A1(n_257_76_15744), .A2(n_257_76_15803), .ZN(
      n_257_76_16150));
   INV_X1 i_257_76_16179 (.A(n_257_76_16150), .ZN(n_257_76_16151));
   NAND4_X1 i_257_76_16180 (.A1(n_257_76_15796), .A2(n_257_76_16151), .A3(
      n_257_76_15788), .A4(n_257_76_15799), .ZN(n_257_76_16152));
   NOR2_X1 i_257_76_16181 (.A1(n_257_76_16149), .A2(n_257_76_16152), .ZN(
      n_257_76_16153));
   INV_X1 i_257_76_16182 (.A(n_257_76_16027), .ZN(n_257_76_16154));
   NAND4_X1 i_257_76_16183 (.A1(n_257_76_15740), .A2(n_257_76_15810), .A3(
      n_257_76_15747), .A4(n_257_76_15811), .ZN(n_257_76_16155));
   INV_X1 i_257_76_16184 (.A(n_257_76_16155), .ZN(n_257_76_16156));
   NAND4_X1 i_257_76_16185 (.A1(n_257_76_16153), .A2(n_257_76_15842), .A3(
      n_257_76_16154), .A4(n_257_76_16156), .ZN(n_257_76_16157));
   INV_X1 i_257_76_16186 (.A(n_257_76_16157), .ZN(n_257_76_16158));
   NAND4_X1 i_257_76_16187 (.A1(n_257_76_16144), .A2(n_257_76_15754), .A3(
      n_257_76_16158), .A4(n_257_76_15712), .ZN(n_257_76_16159));
   INV_X1 i_257_76_16188 (.A(n_257_76_16159), .ZN(n_257_76_16160));
   NAND2_X1 i_257_76_16189 (.A1(n_257_76_18062), .A2(n_257_76_16160), .ZN(
      n_257_76_16161));
   NAND3_X1 i_257_76_16190 (.A1(n_257_76_16128), .A2(n_257_76_16142), .A3(
      n_257_76_16161), .ZN(n_257_76_16162));
   INV_X1 i_257_76_16191 (.A(n_257_76_16162), .ZN(n_257_76_16163));
   NAND2_X1 i_257_76_16192 (.A1(n_257_338), .A2(n_257_76_15807), .ZN(
      n_257_76_16164));
   INV_X1 i_257_76_16193 (.A(n_257_76_16164), .ZN(n_257_76_16165));
   NAND2_X1 i_257_76_16194 (.A1(n_257_76_15906), .A2(n_257_422), .ZN(
      n_257_76_16166));
   INV_X1 i_257_76_16195 (.A(n_257_76_16166), .ZN(n_257_76_16167));
   NAND3_X1 i_257_76_16196 (.A1(n_257_76_16165), .A2(n_257_76_15798), .A3(
      n_257_76_16167), .ZN(n_257_76_16168));
   INV_X1 i_257_76_16197 (.A(n_257_76_16168), .ZN(n_257_76_16169));
   NAND3_X1 i_257_76_16198 (.A1(n_257_76_16169), .A2(n_257_76_15747), .A3(
      n_257_76_15811), .ZN(n_257_76_16170));
   NAND2_X1 i_257_76_16199 (.A1(n_257_76_15740), .A2(n_257_76_15810), .ZN(
      n_257_76_16171));
   NOR2_X1 i_257_76_16200 (.A1(n_257_76_16170), .A2(n_257_76_16171), .ZN(
      n_257_76_16172));
   NAND3_X1 i_257_76_16201 (.A1(n_257_76_15748), .A2(n_257_76_15749), .A3(
      n_257_76_15796), .ZN(n_257_76_16173));
   NAND4_X1 i_257_76_16202 (.A1(n_257_76_15788), .A2(n_257_76_16151), .A3(
      n_257_76_16009), .A4(n_257_76_15799), .ZN(n_257_76_16174));
   NOR2_X1 i_257_76_16203 (.A1(n_257_76_16173), .A2(n_257_76_16174), .ZN(
      n_257_76_16175));
   NAND4_X1 i_257_76_16204 (.A1(n_257_76_16172), .A2(n_257_76_16175), .A3(
      n_257_76_15842), .A4(n_257_76_16154), .ZN(n_257_76_16176));
   INV_X1 i_257_76_16205 (.A(n_257_76_16176), .ZN(n_257_76_16177));
   NAND4_X1 i_257_76_16206 (.A1(n_257_76_15754), .A2(n_257_76_16144), .A3(
      n_257_76_15712), .A4(n_257_76_16177), .ZN(n_257_76_16178));
   INV_X1 i_257_76_16207 (.A(n_257_76_16178), .ZN(n_257_76_16179));
   NAND2_X1 i_257_76_16208 (.A1(n_257_342), .A2(n_257_76_16179), .ZN(
      n_257_76_16180));
   NAND2_X1 i_257_76_16209 (.A1(n_257_442), .A2(n_257_416), .ZN(n_257_76_16181));
   INV_X1 i_257_76_16210 (.A(n_257_76_16181), .ZN(n_257_76_16182));
   NAND2_X1 i_257_76_16211 (.A1(n_257_484), .A2(n_257_76_16182), .ZN(
      n_257_76_16183));
   INV_X1 i_257_76_16212 (.A(n_257_76_16183), .ZN(n_257_76_16184));
   NAND3_X1 i_257_76_16213 (.A1(n_257_76_15998), .A2(n_257_76_15906), .A3(
      n_257_76_16184), .ZN(n_257_76_16185));
   INV_X1 i_257_76_16214 (.A(n_257_76_16185), .ZN(n_257_76_16186));
   NAND2_X1 i_257_76_16215 (.A1(n_257_420), .A2(n_257_497), .ZN(n_257_76_16187));
   NAND4_X1 i_257_76_16216 (.A1(n_257_76_16186), .A2(n_257_76_15997), .A3(
      n_257_76_15803), .A4(n_257_76_16187), .ZN(n_257_76_16188));
   NOR2_X1 i_257_76_16217 (.A1(n_257_76_16094), .A2(n_257_76_16188), .ZN(
      n_257_76_16189));
   NAND2_X1 i_257_76_16218 (.A1(n_257_76_16093), .A2(n_257_76_16189), .ZN(
      n_257_76_16190));
   NOR2_X1 i_257_76_16219 (.A1(n_257_76_16190), .A2(n_257_76_16077), .ZN(
      n_257_76_16191));
   NAND3_X1 i_257_76_16220 (.A1(n_257_76_16191), .A2(n_257_76_15713), .A3(
      n_257_76_15814), .ZN(n_257_76_16192));
   INV_X1 i_257_76_16221 (.A(n_257_76_16192), .ZN(n_257_76_16193));
   NAND3_X1 i_257_76_16222 (.A1(n_257_76_15734), .A2(n_257_76_15738), .A3(
      n_257_76_15785), .ZN(n_257_76_16194));
   INV_X1 i_257_76_16223 (.A(n_257_76_16194), .ZN(n_257_76_16195));
   NAND3_X1 i_257_76_16224 (.A1(n_257_76_15739), .A2(n_257_76_15740), .A3(
      n_257_76_15810), .ZN(n_257_76_16196));
   INV_X1 i_257_76_16225 (.A(n_257_76_16196), .ZN(n_257_76_16197));
   NAND3_X1 i_257_76_16226 (.A1(n_257_76_16195), .A2(n_257_76_16017), .A3(
      n_257_76_16197), .ZN(n_257_76_16198));
   NOR2_X1 i_257_76_16227 (.A1(n_257_76_16198), .A2(n_257_76_16022), .ZN(
      n_257_76_16199));
   NAND4_X1 i_257_76_16228 (.A1(n_257_76_15754), .A2(n_257_76_16193), .A3(
      n_257_76_15712), .A4(n_257_76_16199), .ZN(n_257_76_16200));
   INV_X1 i_257_76_16229 (.A(n_257_76_16200), .ZN(n_257_76_16201));
   NAND2_X1 i_257_76_16230 (.A1(n_257_76_18060), .A2(n_257_76_16201), .ZN(
      n_257_76_16202));
   NAND2_X1 i_257_76_16231 (.A1(n_257_697), .A2(n_257_76_17958), .ZN(
      n_257_76_16203));
   NAND2_X1 i_257_76_16232 (.A1(n_257_76_16105), .A2(n_257_76_16203), .ZN(
      n_257_76_16204));
   INV_X1 i_257_76_16233 (.A(n_257_76_16204), .ZN(n_257_76_16205));
   NAND2_X1 i_257_76_16234 (.A1(n_257_889), .A2(n_257_76_17903), .ZN(
      n_257_76_16206));
   NAND2_X1 i_257_76_16235 (.A1(n_257_141), .A2(n_257_76_17925), .ZN(
      n_257_76_16207));
   NAND3_X1 i_257_76_16236 (.A1(n_257_76_16206), .A2(n_257_76_16168), .A3(
      n_257_76_16207), .ZN(n_257_76_16208));
   INV_X1 i_257_76_16237 (.A(n_257_76_16208), .ZN(n_257_76_16209));
   NAND3_X1 i_257_76_16238 (.A1(n_257_729), .A2(n_257_435), .A3(n_257_442), 
      .ZN(n_257_76_16210));
   NAND2_X1 i_257_76_16239 (.A1(n_257_432), .A2(n_257_76_15908), .ZN(
      n_257_76_16211));
   NAND2_X1 i_257_76_16240 (.A1(n_257_76_16210), .A2(n_257_76_16211), .ZN(
      n_257_76_16212));
   INV_X1 i_257_76_16241 (.A(n_257_76_16212), .ZN(n_257_76_16213));
   NAND2_X1 i_257_76_16242 (.A1(n_257_657), .A2(n_257_76_17928), .ZN(
      n_257_76_16214));
   NAND2_X1 i_257_76_16243 (.A1(n_257_63), .A2(n_257_76_17918), .ZN(
      n_257_76_16215));
   NAND4_X1 i_257_76_16244 (.A1(n_257_76_16213), .A2(n_257_76_16214), .A3(
      n_257_76_16147), .A4(n_257_76_16215), .ZN(n_257_76_16216));
   INV_X1 i_257_76_16245 (.A(n_257_76_16216), .ZN(n_257_76_16217));
   INV_X1 i_257_76_16246 (.A(n_257_76_15715), .ZN(n_257_76_16218));
   NAND2_X1 i_257_76_16247 (.A1(n_257_440), .A2(n_257_76_16218), .ZN(
      n_257_76_16219));
   INV_X1 i_257_76_16248 (.A(n_257_76_15986), .ZN(n_257_76_16220));
   NAND2_X1 i_257_76_16249 (.A1(n_257_438), .A2(n_257_76_16220), .ZN(
      n_257_76_16221));
   INV_X1 i_257_76_16250 (.A(n_257_416), .ZN(n_257_76_16222));
   NAND2_X1 i_257_76_16251 (.A1(n_257_76_16222), .A2(Small_Packet_Data_Size[28]), 
      .ZN(n_257_76_16223));
   INV_X1 i_257_76_16252 (.A(Small_Packet_Data_Size[28]), .ZN(n_257_76_16224));
   OAI21_X1 i_257_76_16253 (.A(n_257_76_16223), .B1(n_257_484), .B2(
      n_257_76_16224), .ZN(n_257_76_16225));
   NAND4_X1 i_257_76_16254 (.A1(n_257_76_16187), .A2(n_257_76_16225), .A3(
      n_257_76_15998), .A4(n_257_76_15906), .ZN(n_257_76_16226));
   NAND2_X1 i_257_76_16255 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[28]), 
      .ZN(n_257_76_16227));
   NAND2_X1 i_257_76_16256 (.A1(n_257_76_16226), .A2(n_257_76_16227), .ZN(
      n_257_76_16228));
   NAND3_X1 i_257_76_16257 (.A1(n_257_76_16219), .A2(n_257_76_16221), .A3(
      n_257_76_16228), .ZN(n_257_76_16229));
   INV_X1 i_257_76_16258 (.A(n_257_76_16229), .ZN(n_257_76_16230));
   NAND3_X1 i_257_76_16259 (.A1(n_257_76_16209), .A2(n_257_76_16217), .A3(
      n_257_76_16230), .ZN(n_257_76_16231));
   NAND2_X1 i_257_76_16260 (.A1(n_257_480), .A2(n_257_442), .ZN(n_257_76_16232));
   INV_X1 i_257_76_16261 (.A(n_257_76_16232), .ZN(n_257_76_16233));
   NAND2_X1 i_257_76_16262 (.A1(n_257_451), .A2(n_257_76_16233), .ZN(
      n_257_76_16234));
   NAND2_X1 i_257_76_16263 (.A1(n_257_76_17940), .A2(n_257_927), .ZN(
      n_257_76_16235));
   INV_X1 i_257_76_16264 (.A(n_257_76_16043), .ZN(n_257_76_16236));
   NAND2_X1 i_257_76_16265 (.A1(n_257_447), .A2(n_257_76_16236), .ZN(
      n_257_76_16237));
   NAND2_X1 i_257_76_16266 (.A1(n_257_825), .A2(n_257_76_17952), .ZN(
      n_257_76_16238));
   NAND4_X1 i_257_76_16267 (.A1(n_257_76_16234), .A2(n_257_76_16235), .A3(
      n_257_76_16237), .A4(n_257_76_16238), .ZN(n_257_76_16239));
   NOR2_X1 i_257_76_16268 (.A1(n_257_76_16231), .A2(n_257_76_16239), .ZN(
      n_257_76_16240));
   NAND2_X1 i_257_76_16269 (.A1(n_257_180), .A2(n_257_76_17331), .ZN(
      n_257_76_16241));
   NAND3_X1 i_257_76_16270 (.A1(n_257_76_16241), .A2(n_257_76_15881), .A3(
      n_257_76_16118), .ZN(n_257_76_16242));
   INV_X1 i_257_76_16271 (.A(n_257_76_16242), .ZN(n_257_76_16243));
   NAND2_X1 i_257_76_16272 (.A1(n_257_991), .A2(n_257_442), .ZN(n_257_76_16244));
   INV_X1 i_257_76_16273 (.A(n_257_76_16244), .ZN(n_257_76_16245));
   NAND2_X1 i_257_76_16274 (.A1(n_257_441), .A2(n_257_76_16245), .ZN(
      n_257_76_16246));
   NAND2_X1 i_257_76_16275 (.A1(n_257_103), .A2(n_257_76_17932), .ZN(
      n_257_76_16247));
   NAND2_X1 i_257_76_16276 (.A1(n_257_76_16246), .A2(n_257_76_16247), .ZN(
      n_257_76_16248));
   NAND2_X1 i_257_76_16277 (.A1(n_257_761), .A2(n_257_76_17935), .ZN(
      n_257_76_16249));
   NAND2_X1 i_257_76_16278 (.A1(n_257_857), .A2(n_257_442), .ZN(n_257_76_16250));
   INV_X1 i_257_76_16279 (.A(n_257_76_16250), .ZN(n_257_76_16251));
   NAND2_X1 i_257_76_16280 (.A1(n_257_446), .A2(n_257_76_16251), .ZN(
      n_257_76_16252));
   INV_X1 i_257_76_16281 (.A(n_257_76_15955), .ZN(n_257_76_16253));
   NAND2_X1 i_257_76_16282 (.A1(n_257_449), .A2(n_257_76_16253), .ZN(
      n_257_76_16254));
   NAND3_X1 i_257_76_16283 (.A1(n_257_76_16249), .A2(n_257_76_16252), .A3(
      n_257_76_16254), .ZN(n_257_76_16255));
   NOR2_X1 i_257_76_16284 (.A1(n_257_76_16248), .A2(n_257_76_16255), .ZN(
      n_257_76_16256));
   NAND3_X1 i_257_76_16285 (.A1(n_257_76_16240), .A2(n_257_76_16243), .A3(
      n_257_76_16256), .ZN(n_257_76_16257));
   INV_X1 i_257_76_16286 (.A(n_257_76_16257), .ZN(n_257_76_16258));
   NAND2_X1 i_257_76_16287 (.A1(n_257_1055), .A2(n_257_76_17969), .ZN(
      n_257_76_16259));
   INV_X1 i_257_76_16288 (.A(n_257_1023), .ZN(n_257_76_16260));
   OAI21_X1 i_257_76_16289 (.A(n_257_76_15812), .B1(n_257_76_16260), .B2(
      n_257_76_17963), .ZN(n_257_76_16261));
   INV_X1 i_257_76_16290 (.A(n_257_76_16261), .ZN(n_257_76_16262));
   NAND3_X1 i_257_76_16291 (.A1(n_257_76_16259), .A2(n_257_76_16262), .A3(
      n_257_76_16087), .ZN(n_257_76_16263));
   INV_X1 i_257_76_16292 (.A(n_257_76_16263), .ZN(n_257_76_16264));
   NAND3_X1 i_257_76_16293 (.A1(n_257_76_16205), .A2(n_257_76_16258), .A3(
      n_257_76_16264), .ZN(n_257_76_16265));
   NAND3_X1 i_257_76_16294 (.A1(n_257_76_16180), .A2(n_257_76_16202), .A3(
      n_257_76_16265), .ZN(n_257_76_16266));
   INV_X1 i_257_76_16295 (.A(n_257_76_16266), .ZN(n_257_76_16267));
   NAND3_X1 i_257_76_16296 (.A1(n_257_76_16111), .A2(n_257_76_16163), .A3(
      n_257_76_16267), .ZN(n_257_76_16268));
   NOR2_X1 i_257_76_16297 (.A1(n_257_76_16062), .A2(n_257_76_16268), .ZN(
      n_257_76_16269));
   NAND2_X1 i_257_76_16298 (.A1(n_257_76_15943), .A2(n_257_76_16269), .ZN(n_28));
   NAND2_X1 i_257_76_16299 (.A1(n_257_1056), .A2(n_257_443), .ZN(n_257_76_16270));
   NAND2_X1 i_257_76_16300 (.A1(n_257_1024), .A2(n_257_444), .ZN(n_257_76_16271));
   NAND2_X1 i_257_76_16301 (.A1(n_257_441), .A2(n_257_992), .ZN(n_257_76_16272));
   NOR2_X1 i_257_76_16302 (.A1(n_257_1088), .A2(n_257_76_17412), .ZN(
      n_257_76_16273));
   INV_X1 i_257_76_16303 (.A(n_257_76_16273), .ZN(n_257_76_16274));
   INV_X1 i_257_76_16304 (.A(n_257_960), .ZN(n_257_76_16275));
   NOR2_X1 i_257_76_16305 (.A1(n_257_76_16274), .A2(n_257_76_16275), .ZN(
      n_257_76_16276));
   NAND2_X1 i_257_76_16306 (.A1(n_257_440), .A2(n_257_76_16276), .ZN(
      n_257_76_16277));
   INV_X1 i_257_76_16307 (.A(n_257_76_16277), .ZN(n_257_76_16278));
   NAND2_X1 i_257_76_16308 (.A1(n_257_76_16272), .A2(n_257_76_16278), .ZN(
      n_257_76_16279));
   INV_X1 i_257_76_16309 (.A(n_257_76_16279), .ZN(n_257_76_16280));
   NAND2_X1 i_257_76_16310 (.A1(n_257_76_16271), .A2(n_257_76_16280), .ZN(
      n_257_76_16281));
   INV_X1 i_257_76_16311 (.A(n_257_76_16281), .ZN(n_257_76_16282));
   NAND2_X1 i_257_76_16312 (.A1(n_257_76_16270), .A2(n_257_76_16282), .ZN(
      n_257_76_16283));
   INV_X1 i_257_76_16313 (.A(n_257_76_16283), .ZN(n_257_76_16284));
   NAND2_X1 i_257_76_16314 (.A1(n_257_17), .A2(n_257_76_16284), .ZN(
      n_257_76_16285));
   NAND2_X1 i_257_76_16315 (.A1(n_257_443), .A2(n_257_76_16273), .ZN(
      n_257_76_16286));
   INV_X1 i_257_76_16316 (.A(n_257_76_16286), .ZN(n_257_76_16287));
   NAND2_X1 i_257_76_16317 (.A1(n_257_1056), .A2(n_257_76_16287), .ZN(
      n_257_76_16288));
   INV_X1 i_257_76_16318 (.A(n_257_76_16288), .ZN(n_257_76_16289));
   NAND2_X1 i_257_76_16319 (.A1(n_257_76_18072), .A2(n_257_76_16289), .ZN(
      n_257_76_16290));
   NAND2_X1 i_257_76_16320 (.A1(n_257_698), .A2(n_257_448), .ZN(n_257_76_16291));
   NAND2_X1 i_257_76_16321 (.A1(n_257_762), .A2(n_257_436), .ZN(n_257_76_16292));
   NAND2_X1 i_257_76_16322 (.A1(n_257_446), .A2(n_257_858), .ZN(n_257_76_16293));
   NAND2_X1 i_257_76_16323 (.A1(n_257_449), .A2(n_257_666), .ZN(n_257_76_16294));
   NAND3_X1 i_257_76_16324 (.A1(n_257_76_16292), .A2(n_257_76_16293), .A3(
      n_257_76_16294), .ZN(n_257_76_16295));
   INV_X1 i_257_76_16325 (.A(n_257_76_16272), .ZN(n_257_76_16296));
   NOR2_X1 i_257_76_16326 (.A1(n_257_76_16295), .A2(n_257_76_16296), .ZN(
      n_257_76_16297));
   NAND2_X1 i_257_76_16327 (.A1(n_257_447), .A2(n_257_794), .ZN(n_257_76_16298));
   NAND2_X1 i_257_76_16328 (.A1(n_257_928), .A2(n_257_439), .ZN(n_257_76_16299));
   NAND2_X1 i_257_76_16329 (.A1(n_257_826), .A2(n_257_437), .ZN(n_257_76_16300));
   NAND3_X1 i_257_76_16330 (.A1(n_257_76_16298), .A2(n_257_76_16299), .A3(
      n_257_76_16300), .ZN(n_257_76_16301));
   NAND2_X1 i_257_76_16331 (.A1(n_257_890), .A2(n_257_445), .ZN(n_257_76_16302));
   NAND2_X1 i_257_76_16332 (.A1(n_257_450), .A2(n_257_76_16273), .ZN(
      n_257_76_16303));
   INV_X1 i_257_76_16333 (.A(n_257_76_16303), .ZN(n_257_76_16304));
   NAND2_X1 i_257_76_16334 (.A1(n_257_730), .A2(n_257_435), .ZN(n_257_76_16305));
   NAND3_X1 i_257_76_16335 (.A1(n_257_658), .A2(n_257_76_16304), .A3(
      n_257_76_16305), .ZN(n_257_76_16306));
   INV_X1 i_257_76_16336 (.A(n_257_76_16306), .ZN(n_257_76_16307));
   NAND2_X1 i_257_76_16337 (.A1(n_257_440), .A2(n_257_960), .ZN(n_257_76_16308));
   NAND2_X1 i_257_76_16338 (.A1(n_257_438), .A2(n_257_896), .ZN(n_257_76_16309));
   NAND4_X1 i_257_76_16339 (.A1(n_257_76_16302), .A2(n_257_76_16307), .A3(
      n_257_76_16308), .A4(n_257_76_16309), .ZN(n_257_76_16310));
   NOR2_X1 i_257_76_16340 (.A1(n_257_76_16301), .A2(n_257_76_16310), .ZN(
      n_257_76_16311));
   NAND4_X1 i_257_76_16341 (.A1(n_257_76_16291), .A2(n_257_76_16297), .A3(
      n_257_76_16311), .A4(n_257_76_16271), .ZN(n_257_76_16312));
   INV_X1 i_257_76_16342 (.A(n_257_76_16270), .ZN(n_257_76_16313));
   NOR2_X1 i_257_76_16343 (.A1(n_257_76_16312), .A2(n_257_76_16313), .ZN(
      n_257_76_16314));
   NAND2_X1 i_257_76_16344 (.A1(n_257_28), .A2(n_257_76_16314), .ZN(
      n_257_76_16315));
   NAND3_X1 i_257_76_16345 (.A1(n_257_76_16285), .A2(n_257_76_16290), .A3(
      n_257_76_16315), .ZN(n_257_76_16316));
   NAND2_X1 i_257_76_16346 (.A1(n_257_76_16299), .A2(n_257_76_16302), .ZN(
      n_257_76_16317));
   INV_X1 i_257_76_16347 (.A(n_257_76_16317), .ZN(n_257_76_16318));
   INV_X1 i_257_76_16348 (.A(n_257_858), .ZN(n_257_76_16319));
   NOR2_X1 i_257_76_16349 (.A1(n_257_76_16274), .A2(n_257_76_16319), .ZN(
      n_257_76_16320));
   NAND4_X1 i_257_76_16350 (.A1(n_257_446), .A2(n_257_76_16308), .A3(
      n_257_76_16309), .A4(n_257_76_16320), .ZN(n_257_76_16321));
   INV_X1 i_257_76_16351 (.A(n_257_76_16321), .ZN(n_257_76_16322));
   NAND3_X1 i_257_76_16352 (.A1(n_257_76_16318), .A2(n_257_76_16322), .A3(
      n_257_76_16272), .ZN(n_257_76_16323));
   INV_X1 i_257_76_16353 (.A(n_257_76_16323), .ZN(n_257_76_16324));
   NAND2_X1 i_257_76_16354 (.A1(n_257_76_16324), .A2(n_257_76_16271), .ZN(
      n_257_76_16325));
   NOR2_X1 i_257_76_16355 (.A1(n_257_76_16313), .A2(n_257_76_16325), .ZN(
      n_257_76_16326));
   NAND2_X1 i_257_76_16356 (.A1(n_257_76_18070), .A2(n_257_76_16326), .ZN(
      n_257_76_16327));
   NAND2_X1 i_257_76_16357 (.A1(n_257_439), .A2(n_257_76_16273), .ZN(
      n_257_76_16328));
   INV_X1 i_257_76_16358 (.A(n_257_76_16328), .ZN(n_257_76_16329));
   NAND3_X1 i_257_76_16359 (.A1(n_257_76_16329), .A2(n_257_928), .A3(
      n_257_76_16308), .ZN(n_257_76_16330));
   INV_X1 i_257_76_16360 (.A(n_257_76_16330), .ZN(n_257_76_16331));
   NAND2_X1 i_257_76_16361 (.A1(n_257_76_16272), .A2(n_257_76_16331), .ZN(
      n_257_76_16332));
   INV_X1 i_257_76_16362 (.A(n_257_76_16332), .ZN(n_257_76_16333));
   NAND2_X1 i_257_76_16363 (.A1(n_257_76_16271), .A2(n_257_76_16333), .ZN(
      n_257_76_16334));
   INV_X1 i_257_76_16364 (.A(n_257_76_16334), .ZN(n_257_76_16335));
   NAND2_X1 i_257_76_16365 (.A1(n_257_76_16270), .A2(n_257_76_16335), .ZN(
      n_257_76_16336));
   INV_X1 i_257_76_16366 (.A(n_257_76_16336), .ZN(n_257_76_16337));
   NAND2_X1 i_257_76_16367 (.A1(n_257_76_18084), .A2(n_257_76_16337), .ZN(
      n_257_76_16338));
   NAND2_X1 i_257_76_16368 (.A1(n_257_181), .A2(n_257_429), .ZN(n_257_76_16339));
   NAND2_X1 i_257_76_16369 (.A1(n_257_261), .A2(n_257_425), .ZN(n_257_76_16340));
   NAND2_X1 i_257_76_16370 (.A1(n_257_530), .A2(n_257_424), .ZN(n_257_76_16341));
   NAND2_X1 i_257_76_16371 (.A1(n_257_64), .A2(n_257_433), .ZN(n_257_76_16342));
   NAND2_X1 i_257_76_16372 (.A1(n_257_76_16341), .A2(n_257_76_16342), .ZN(
      n_257_76_16343));
   INV_X1 i_257_76_16373 (.A(n_257_76_16343), .ZN(n_257_76_16344));
   NAND2_X1 i_257_76_16374 (.A1(n_257_301), .A2(n_257_76_16305), .ZN(
      n_257_76_16345));
   INV_X1 i_257_76_16375 (.A(n_257_76_16345), .ZN(n_257_76_16346));
   NAND2_X1 i_257_76_16376 (.A1(n_257_658), .A2(n_257_450), .ZN(n_257_76_16347));
   NAND2_X1 i_257_76_16377 (.A1(n_257_432), .A2(n_257_626), .ZN(n_257_76_16348));
   INV_X1 i_257_76_16378 (.A(n_257_594), .ZN(n_257_76_16349));
   NAND2_X1 i_257_76_16379 (.A1(n_257_76_16349), .A2(n_257_442), .ZN(
      n_257_76_16350));
   OAI21_X1 i_257_76_16380 (.A(n_257_76_16350), .B1(n_257_428), .B2(
      n_257_76_17412), .ZN(n_257_76_16351));
   INV_X1 i_257_76_16381 (.A(n_257_1088), .ZN(n_257_76_16352));
   NAND2_X1 i_257_76_16382 (.A1(n_257_423), .A2(n_257_76_16352), .ZN(
      n_257_76_16353));
   INV_X1 i_257_76_16383 (.A(n_257_76_16353), .ZN(n_257_76_16354));
   NAND3_X1 i_257_76_16384 (.A1(n_257_76_16348), .A2(n_257_76_16351), .A3(
      n_257_76_16354), .ZN(n_257_76_16355));
   INV_X1 i_257_76_16385 (.A(n_257_76_16355), .ZN(n_257_76_16356));
   NAND4_X1 i_257_76_16386 (.A1(n_257_76_16344), .A2(n_257_76_16346), .A3(
      n_257_76_16347), .A4(n_257_76_16356), .ZN(n_257_76_16357));
   INV_X1 i_257_76_16387 (.A(n_257_76_16357), .ZN(n_257_76_16358));
   NAND4_X1 i_257_76_16388 (.A1(n_257_76_16339), .A2(n_257_76_16340), .A3(
      n_257_76_16272), .A4(n_257_76_16358), .ZN(n_257_76_16359));
   INV_X1 i_257_76_16389 (.A(n_257_76_16271), .ZN(n_257_76_16360));
   NOR2_X1 i_257_76_16390 (.A1(n_257_76_16359), .A2(n_257_76_16360), .ZN(
      n_257_76_16361));
   NAND2_X1 i_257_76_16391 (.A1(n_257_562), .A2(n_257_426), .ZN(n_257_76_16362));
   NAND2_X1 i_257_76_16392 (.A1(n_257_142), .A2(n_257_430), .ZN(n_257_76_16363));
   NAND3_X1 i_257_76_16393 (.A1(n_257_76_16300), .A2(n_257_76_16362), .A3(
      n_257_76_16363), .ZN(n_257_76_16364));
   NAND2_X1 i_257_76_16394 (.A1(n_257_427), .A2(n_257_221), .ZN(n_257_76_16365));
   NAND4_X1 i_257_76_16395 (.A1(n_257_76_16302), .A2(n_257_76_16308), .A3(
      n_257_76_16309), .A4(n_257_76_16365), .ZN(n_257_76_16366));
   NOR2_X1 i_257_76_16396 (.A1(n_257_76_16364), .A2(n_257_76_16366), .ZN(
      n_257_76_16367));
   NAND2_X1 i_257_76_16397 (.A1(n_257_104), .A2(n_257_431), .ZN(n_257_76_16368));
   NAND3_X1 i_257_76_16398 (.A1(n_257_76_16368), .A2(n_257_76_16292), .A3(
      n_257_76_16293), .ZN(n_257_76_16369));
   INV_X1 i_257_76_16399 (.A(n_257_76_16369), .ZN(n_257_76_16370));
   NAND2_X1 i_257_76_16400 (.A1(n_257_451), .A2(n_257_481), .ZN(n_257_76_16371));
   NAND4_X1 i_257_76_16401 (.A1(n_257_76_16294), .A2(n_257_76_16298), .A3(
      n_257_76_16371), .A4(n_257_76_16299), .ZN(n_257_76_16372));
   INV_X1 i_257_76_16402 (.A(n_257_76_16372), .ZN(n_257_76_16373));
   NAND3_X1 i_257_76_16403 (.A1(n_257_76_16367), .A2(n_257_76_16370), .A3(
      n_257_76_16373), .ZN(n_257_76_16374));
   INV_X1 i_257_76_16404 (.A(n_257_76_16374), .ZN(n_257_76_16375));
   NAND4_X1 i_257_76_16405 (.A1(n_257_76_16361), .A2(n_257_76_16375), .A3(
      n_257_76_16270), .A4(n_257_76_16291), .ZN(n_257_76_16376));
   INV_X1 i_257_76_16406 (.A(n_257_76_16376), .ZN(n_257_76_16377));
   NAND2_X1 i_257_76_16407 (.A1(n_257_76_18066), .A2(n_257_76_16377), .ZN(
      n_257_76_16378));
   NAND3_X1 i_257_76_16408 (.A1(n_257_76_16327), .A2(n_257_76_16338), .A3(
      n_257_76_16378), .ZN(n_257_76_16379));
   NOR2_X1 i_257_76_16409 (.A1(n_257_76_16316), .A2(n_257_76_16379), .ZN(
      n_257_76_16380));
   NAND2_X1 i_257_76_16410 (.A1(n_257_992), .A2(n_257_76_16273), .ZN(
      n_257_76_16381));
   INV_X1 i_257_76_16411 (.A(n_257_76_16381), .ZN(n_257_76_16382));
   NAND2_X1 i_257_76_16412 (.A1(n_257_441), .A2(n_257_76_16382), .ZN(
      n_257_76_16383));
   INV_X1 i_257_76_16413 (.A(n_257_76_16383), .ZN(n_257_76_16384));
   NAND2_X1 i_257_76_16414 (.A1(n_257_76_16271), .A2(n_257_76_16384), .ZN(
      n_257_76_16385));
   INV_X1 i_257_76_16415 (.A(n_257_76_16385), .ZN(n_257_76_16386));
   NAND2_X1 i_257_76_16416 (.A1(n_257_76_16270), .A2(n_257_76_16386), .ZN(
      n_257_76_16387));
   INV_X1 i_257_76_16417 (.A(n_257_76_16387), .ZN(n_257_76_16388));
   NAND2_X1 i_257_76_16418 (.A1(n_257_76_18071), .A2(n_257_76_16388), .ZN(
      n_257_76_16389));
   NAND2_X1 i_257_76_16419 (.A1(n_257_76_16292), .A2(n_257_76_16293), .ZN(
      n_257_76_16390));
   NOR2_X1 i_257_76_16420 (.A1(n_257_76_16296), .A2(n_257_76_16390), .ZN(
      n_257_76_16391));
   NAND3_X1 i_257_76_16421 (.A1(n_257_730), .A2(n_257_435), .A3(n_257_76_16273), 
      .ZN(n_257_76_16392));
   INV_X1 i_257_76_16422 (.A(n_257_76_16392), .ZN(n_257_76_16393));
   NAND4_X1 i_257_76_16423 (.A1(n_257_76_16302), .A2(n_257_76_16308), .A3(
      n_257_76_16309), .A4(n_257_76_16393), .ZN(n_257_76_16394));
   NOR2_X1 i_257_76_16424 (.A1(n_257_76_16301), .A2(n_257_76_16394), .ZN(
      n_257_76_16395));
   NAND3_X1 i_257_76_16425 (.A1(n_257_76_16271), .A2(n_257_76_16391), .A3(
      n_257_76_16395), .ZN(n_257_76_16396));
   NOR2_X1 i_257_76_16426 (.A1(n_257_76_16396), .A2(n_257_76_16313), .ZN(
      n_257_76_16397));
   NAND2_X1 i_257_76_16427 (.A1(n_257_76_18078), .A2(n_257_76_16397), .ZN(
      n_257_76_16398));
   NAND4_X1 i_257_76_16428 (.A1(n_257_76_16298), .A2(n_257_76_16371), .A3(
      n_257_76_16299), .A4(n_257_76_16300), .ZN(n_257_76_16399));
   INV_X1 i_257_76_16429 (.A(n_257_76_16399), .ZN(n_257_76_16400));
   INV_X1 i_257_76_16430 (.A(n_257_76_16295), .ZN(n_257_76_16401));
   NAND3_X1 i_257_76_16431 (.A1(n_257_76_16363), .A2(n_257_76_16302), .A3(
      n_257_76_16308), .ZN(n_257_76_16402));
   NAND2_X1 i_257_76_16432 (.A1(n_257_594), .A2(n_257_442), .ZN(n_257_76_16403));
   INV_X1 i_257_76_16433 (.A(n_257_76_16403), .ZN(n_257_76_16404));
   NAND3_X1 i_257_76_16434 (.A1(n_257_428), .A2(n_257_76_16352), .A3(
      n_257_76_16404), .ZN(n_257_76_16405));
   INV_X1 i_257_76_16435 (.A(n_257_76_16405), .ZN(n_257_76_16406));
   NAND3_X1 i_257_76_16436 (.A1(n_257_76_16305), .A2(n_257_76_16348), .A3(
      n_257_76_16406), .ZN(n_257_76_16407));
   INV_X1 i_257_76_16437 (.A(n_257_76_16407), .ZN(n_257_76_16408));
   NAND4_X1 i_257_76_16438 (.A1(n_257_76_16309), .A2(n_257_76_16408), .A3(
      n_257_76_16347), .A4(n_257_76_16342), .ZN(n_257_76_16409));
   NOR2_X1 i_257_76_16439 (.A1(n_257_76_16402), .A2(n_257_76_16409), .ZN(
      n_257_76_16410));
   NAND3_X1 i_257_76_16440 (.A1(n_257_76_16400), .A2(n_257_76_16401), .A3(
      n_257_76_16410), .ZN(n_257_76_16411));
   INV_X1 i_257_76_16441 (.A(n_257_76_16411), .ZN(n_257_76_16412));
   NAND2_X1 i_257_76_16442 (.A1(n_257_76_16272), .A2(n_257_76_16368), .ZN(
      n_257_76_16413));
   INV_X1 i_257_76_16443 (.A(n_257_76_16413), .ZN(n_257_76_16414));
   NAND3_X1 i_257_76_16444 (.A1(n_257_76_16271), .A2(n_257_76_16414), .A3(
      n_257_76_16339), .ZN(n_257_76_16415));
   INV_X1 i_257_76_16445 (.A(n_257_76_16415), .ZN(n_257_76_16416));
   NAND4_X1 i_257_76_16446 (.A1(n_257_76_16412), .A2(n_257_76_16416), .A3(
      n_257_76_16270), .A4(n_257_76_16291), .ZN(n_257_76_16417));
   INV_X1 i_257_76_16447 (.A(n_257_76_16417), .ZN(n_257_76_16418));
   NAND2_X1 i_257_76_16448 (.A1(n_257_76_18074), .A2(n_257_76_16418), .ZN(
      n_257_76_16419));
   NAND3_X1 i_257_76_16449 (.A1(n_257_76_16389), .A2(n_257_76_16398), .A3(
      n_257_76_16419), .ZN(n_257_76_16420));
   NAND2_X1 i_257_76_16450 (.A1(n_257_1088), .A2(n_257_442), .ZN(n_257_76_16421));
   INV_X1 i_257_76_16451 (.A(n_257_76_16421), .ZN(n_257_76_16422));
   NAND2_X1 i_257_76_16452 (.A1(n_257_13), .A2(n_257_76_16422), .ZN(
      n_257_76_16423));
   NAND2_X1 i_257_76_16453 (.A1(n_257_445), .A2(n_257_76_16273), .ZN(
      n_257_76_16424));
   INV_X1 i_257_76_16454 (.A(n_257_76_16424), .ZN(n_257_76_16425));
   NAND4_X1 i_257_76_16455 (.A1(n_257_76_16308), .A2(n_257_76_16309), .A3(
      n_257_890), .A4(n_257_76_16425), .ZN(n_257_76_16426));
   INV_X1 i_257_76_16456 (.A(n_257_76_16426), .ZN(n_257_76_16427));
   NAND3_X1 i_257_76_16457 (.A1(n_257_76_16427), .A2(n_257_76_16272), .A3(
      n_257_76_16299), .ZN(n_257_76_16428));
   INV_X1 i_257_76_16458 (.A(n_257_76_16428), .ZN(n_257_76_16429));
   NAND2_X1 i_257_76_16459 (.A1(n_257_76_16429), .A2(n_257_76_16271), .ZN(
      n_257_76_16430));
   NOR2_X1 i_257_76_16460 (.A1(n_257_76_16313), .A2(n_257_76_16430), .ZN(
      n_257_76_16431));
   NAND2_X1 i_257_76_16461 (.A1(n_257_76_18077), .A2(n_257_76_16431), .ZN(
      n_257_76_16432));
   NAND2_X1 i_257_76_16462 (.A1(n_257_76_16423), .A2(n_257_76_16432), .ZN(
      n_257_76_16433));
   NOR2_X1 i_257_76_16463 (.A1(n_257_76_16420), .A2(n_257_76_16433), .ZN(
      n_257_76_16434));
   NAND3_X1 i_257_76_16464 (.A1(n_257_76_16309), .A2(n_257_562), .A3(
      n_257_76_16347), .ZN(n_257_76_16435));
   NAND2_X1 i_257_76_16465 (.A1(n_257_76_16305), .A2(n_257_76_16348), .ZN(
      n_257_76_16436));
   INV_X1 i_257_76_16466 (.A(n_257_76_16436), .ZN(n_257_76_16437));
   NAND2_X1 i_257_76_16467 (.A1(n_257_426), .A2(n_257_76_16352), .ZN(
      n_257_76_16438));
   INV_X1 i_257_76_16468 (.A(n_257_76_16438), .ZN(n_257_76_16439));
   NAND2_X1 i_257_76_16469 (.A1(n_257_76_16439), .A2(n_257_76_16351), .ZN(
      n_257_76_16440));
   INV_X1 i_257_76_16470 (.A(n_257_76_16440), .ZN(n_257_76_16441));
   NAND4_X1 i_257_76_16471 (.A1(n_257_76_16437), .A2(n_257_76_16365), .A3(
      n_257_76_16342), .A4(n_257_76_16441), .ZN(n_257_76_16442));
   NOR2_X1 i_257_76_16472 (.A1(n_257_76_16435), .A2(n_257_76_16442), .ZN(
      n_257_76_16443));
   NAND2_X1 i_257_76_16473 (.A1(n_257_76_16292), .A2(n_257_76_16299), .ZN(
      n_257_76_16444));
   INV_X1 i_257_76_16474 (.A(n_257_76_16444), .ZN(n_257_76_16445));
   NAND3_X1 i_257_76_16475 (.A1(n_257_76_16300), .A2(n_257_76_16363), .A3(
      n_257_76_16302), .ZN(n_257_76_16446));
   INV_X1 i_257_76_16476 (.A(n_257_76_16446), .ZN(n_257_76_16447));
   NAND3_X1 i_257_76_16477 (.A1(n_257_76_16443), .A2(n_257_76_16445), .A3(
      n_257_76_16447), .ZN(n_257_76_16448));
   INV_X1 i_257_76_16478 (.A(n_257_76_16448), .ZN(n_257_76_16449));
   NAND2_X1 i_257_76_16479 (.A1(n_257_76_16270), .A2(n_257_76_16449), .ZN(
      n_257_76_16450));
   NAND3_X1 i_257_76_16480 (.A1(n_257_76_16339), .A2(n_257_76_16272), .A3(
      n_257_76_16368), .ZN(n_257_76_16451));
   INV_X1 i_257_76_16481 (.A(n_257_76_16451), .ZN(n_257_76_16452));
   NAND3_X1 i_257_76_16482 (.A1(n_257_76_16298), .A2(n_257_76_16371), .A3(
      n_257_76_16308), .ZN(n_257_76_16453));
   NAND2_X1 i_257_76_16483 (.A1(n_257_76_16293), .A2(n_257_76_16294), .ZN(
      n_257_76_16454));
   NOR2_X1 i_257_76_16484 (.A1(n_257_76_16453), .A2(n_257_76_16454), .ZN(
      n_257_76_16455));
   NAND4_X1 i_257_76_16485 (.A1(n_257_76_16452), .A2(n_257_76_16291), .A3(
      n_257_76_16455), .A4(n_257_76_16271), .ZN(n_257_76_16456));
   NOR2_X1 i_257_76_16486 (.A1(n_257_76_16450), .A2(n_257_76_16456), .ZN(
      n_257_76_16457));
   NAND2_X1 i_257_76_16487 (.A1(n_257_76_18076), .A2(n_257_76_16457), .ZN(
      n_257_76_16458));
   NAND2_X1 i_257_76_16488 (.A1(n_257_76_16293), .A2(n_257_76_16298), .ZN(
      n_257_76_16459));
   NOR2_X1 i_257_76_16489 (.A1(n_257_76_16296), .A2(n_257_76_16459), .ZN(
      n_257_76_16460));
   NAND3_X1 i_257_76_16490 (.A1(n_257_76_16299), .A2(n_257_76_16300), .A3(
      n_257_76_16302), .ZN(n_257_76_16461));
   NAND2_X1 i_257_76_16491 (.A1(n_257_436), .A2(n_257_76_16273), .ZN(
      n_257_76_16462));
   INV_X1 i_257_76_16492 (.A(n_257_76_16462), .ZN(n_257_76_16463));
   NAND4_X1 i_257_76_16493 (.A1(n_257_762), .A2(n_257_76_16308), .A3(
      n_257_76_16309), .A4(n_257_76_16463), .ZN(n_257_76_16464));
   NOR2_X1 i_257_76_16494 (.A1(n_257_76_16461), .A2(n_257_76_16464), .ZN(
      n_257_76_16465));
   NAND3_X1 i_257_76_16495 (.A1(n_257_76_16271), .A2(n_257_76_16460), .A3(
      n_257_76_16465), .ZN(n_257_76_16466));
   NOR2_X1 i_257_76_16496 (.A1(n_257_76_16466), .A2(n_257_76_16313), .ZN(
      n_257_76_16467));
   NAND2_X1 i_257_76_16497 (.A1(n_257_76_18069), .A2(n_257_76_16467), .ZN(
      n_257_76_16468));
   NAND2_X1 i_257_76_16498 (.A1(n_257_76_16272), .A2(n_257_76_16292), .ZN(
      n_257_76_16469));
   INV_X1 i_257_76_16499 (.A(n_257_76_16469), .ZN(n_257_76_16470));
   NAND2_X1 i_257_76_16500 (.A1(n_257_76_16271), .A2(n_257_76_16470), .ZN(
      n_257_76_16471));
   INV_X1 i_257_76_16501 (.A(n_257_76_16471), .ZN(n_257_76_16472));
   NAND2_X1 i_257_76_16502 (.A1(n_257_626), .A2(n_257_442), .ZN(n_257_76_16473));
   NOR2_X1 i_257_76_16503 (.A1(n_257_1088), .A2(n_257_76_16473), .ZN(
      n_257_76_16474));
   NAND2_X1 i_257_76_16504 (.A1(n_257_432), .A2(n_257_76_16474), .ZN(
      n_257_76_16475));
   INV_X1 i_257_76_16505 (.A(n_257_76_16475), .ZN(n_257_76_16476));
   NAND3_X1 i_257_76_16506 (.A1(n_257_76_16342), .A2(n_257_76_16305), .A3(
      n_257_76_16476), .ZN(n_257_76_16477));
   INV_X1 i_257_76_16507 (.A(n_257_76_16477), .ZN(n_257_76_16478));
   NAND3_X1 i_257_76_16508 (.A1(n_257_76_16478), .A2(n_257_76_16309), .A3(
      n_257_76_16347), .ZN(n_257_76_16479));
   NAND2_X1 i_257_76_16509 (.A1(n_257_76_16302), .A2(n_257_76_16308), .ZN(
      n_257_76_16480));
   NOR2_X1 i_257_76_16510 (.A1(n_257_76_16479), .A2(n_257_76_16480), .ZN(
      n_257_76_16481));
   NAND3_X1 i_257_76_16511 (.A1(n_257_76_16293), .A2(n_257_76_16294), .A3(
      n_257_76_16298), .ZN(n_257_76_16482));
   INV_X1 i_257_76_16512 (.A(n_257_76_16482), .ZN(n_257_76_16483));
   NAND3_X1 i_257_76_16513 (.A1(n_257_76_16371), .A2(n_257_76_16299), .A3(
      n_257_76_16300), .ZN(n_257_76_16484));
   INV_X1 i_257_76_16514 (.A(n_257_76_16484), .ZN(n_257_76_16485));
   NAND3_X1 i_257_76_16515 (.A1(n_257_76_16481), .A2(n_257_76_16483), .A3(
      n_257_76_16485), .ZN(n_257_76_16486));
   INV_X1 i_257_76_16516 (.A(n_257_76_16486), .ZN(n_257_76_16487));
   NAND4_X1 i_257_76_16517 (.A1(n_257_76_16270), .A2(n_257_76_16472), .A3(
      n_257_76_16487), .A4(n_257_76_16291), .ZN(n_257_76_16488));
   INV_X1 i_257_76_16518 (.A(n_257_76_16488), .ZN(n_257_76_16489));
   NAND2_X1 i_257_76_16519 (.A1(n_257_68), .A2(n_257_76_16489), .ZN(
      n_257_76_16490));
   NAND3_X1 i_257_76_16520 (.A1(n_257_76_16458), .A2(n_257_76_16468), .A3(
      n_257_76_16490), .ZN(n_257_76_16491));
   NAND2_X1 i_257_76_16521 (.A1(n_257_437), .A2(n_257_76_16273), .ZN(
      n_257_76_16492));
   INV_X1 i_257_76_16522 (.A(n_257_76_16492), .ZN(n_257_76_16493));
   NAND4_X1 i_257_76_16523 (.A1(n_257_76_16308), .A2(n_257_76_16309), .A3(
      n_257_826), .A4(n_257_76_16493), .ZN(n_257_76_16494));
   NOR2_X1 i_257_76_16524 (.A1(n_257_76_16317), .A2(n_257_76_16494), .ZN(
      n_257_76_16495));
   NAND2_X1 i_257_76_16525 (.A1(n_257_76_16272), .A2(n_257_76_16293), .ZN(
      n_257_76_16496));
   INV_X1 i_257_76_16526 (.A(n_257_76_16496), .ZN(n_257_76_16497));
   NAND3_X1 i_257_76_16527 (.A1(n_257_76_16495), .A2(n_257_76_16271), .A3(
      n_257_76_16497), .ZN(n_257_76_16498));
   NOR2_X1 i_257_76_16528 (.A1(n_257_76_16313), .A2(n_257_76_16498), .ZN(
      n_257_76_16499));
   NAND2_X1 i_257_76_16529 (.A1(n_257_22), .A2(n_257_76_16499), .ZN(
      n_257_76_16500));
   NAND2_X1 i_257_76_16530 (.A1(n_257_444), .A2(n_257_76_16273), .ZN(
      n_257_76_16501));
   INV_X1 i_257_76_16531 (.A(n_257_76_16501), .ZN(n_257_76_16502));
   NAND2_X1 i_257_76_16532 (.A1(n_257_1024), .A2(n_257_76_16502), .ZN(
      n_257_76_16503));
   INV_X1 i_257_76_16533 (.A(n_257_76_16503), .ZN(n_257_76_16504));
   NAND2_X1 i_257_76_16534 (.A1(n_257_76_16270), .A2(n_257_76_16504), .ZN(
      n_257_76_16505));
   INV_X1 i_257_76_16535 (.A(n_257_76_16505), .ZN(n_257_76_16506));
   NAND2_X1 i_257_76_16536 (.A1(n_257_76_18075), .A2(n_257_76_16506), .ZN(
      n_257_76_16507));
   NAND2_X1 i_257_76_16537 (.A1(n_257_76_16500), .A2(n_257_76_16507), .ZN(
      n_257_76_16508));
   NOR2_X1 i_257_76_16538 (.A1(n_257_76_16491), .A2(n_257_76_16508), .ZN(
      n_257_76_16509));
   NAND3_X1 i_257_76_16539 (.A1(n_257_76_16380), .A2(n_257_76_16434), .A3(
      n_257_76_16509), .ZN(n_257_76_16510));
   INV_X1 i_257_76_16540 (.A(n_257_76_16510), .ZN(n_257_76_16511));
   INV_X1 i_257_76_16541 (.A(n_257_76_16480), .ZN(n_257_76_16512));
   NOR2_X1 i_257_76_16542 (.A1(n_257_76_16274), .A2(n_257_76_17074), .ZN(
      n_257_76_16513));
   NAND3_X1 i_257_76_16543 (.A1(n_257_76_16305), .A2(n_257_76_16513), .A3(
      n_257_64), .ZN(n_257_76_16514));
   INV_X1 i_257_76_16544 (.A(n_257_76_16514), .ZN(n_257_76_16515));
   NAND3_X1 i_257_76_16545 (.A1(n_257_76_16309), .A2(n_257_76_16515), .A3(
      n_257_76_16347), .ZN(n_257_76_16516));
   INV_X1 i_257_76_16546 (.A(n_257_76_16516), .ZN(n_257_76_16517));
   NAND4_X1 i_257_76_16547 (.A1(n_257_76_16512), .A2(n_257_76_16517), .A3(
      n_257_76_16299), .A4(n_257_76_16300), .ZN(n_257_76_16518));
   NAND4_X1 i_257_76_16548 (.A1(n_257_76_16293), .A2(n_257_76_16294), .A3(
      n_257_76_16298), .A4(n_257_76_16371), .ZN(n_257_76_16519));
   NOR2_X1 i_257_76_16549 (.A1(n_257_76_16518), .A2(n_257_76_16519), .ZN(
      n_257_76_16520));
   NAND4_X1 i_257_76_16550 (.A1(n_257_76_16520), .A2(n_257_76_16270), .A3(
      n_257_76_16472), .A4(n_257_76_16291), .ZN(n_257_76_16521));
   INV_X1 i_257_76_16551 (.A(n_257_76_16521), .ZN(n_257_76_16522));
   NAND2_X1 i_257_76_16552 (.A1(n_257_76_18081), .A2(n_257_76_16522), .ZN(
      n_257_76_16523));
   NAND3_X1 i_257_76_16553 (.A1(n_257_76_16292), .A2(n_257_76_16293), .A3(
      n_257_76_16298), .ZN(n_257_76_16524));
   NOR2_X1 i_257_76_16554 (.A1(n_257_76_16524), .A2(n_257_76_16296), .ZN(
      n_257_76_16525));
   NAND2_X1 i_257_76_16555 (.A1(n_257_442), .A2(n_257_666), .ZN(n_257_76_16526));
   NOR2_X1 i_257_76_16556 (.A1(n_257_1088), .A2(n_257_76_16526), .ZN(
      n_257_76_16527));
   NAND2_X1 i_257_76_16557 (.A1(n_257_76_16305), .A2(n_257_76_16527), .ZN(
      n_257_76_16528));
   INV_X1 i_257_76_16558 (.A(n_257_76_16528), .ZN(n_257_76_16529));
   NAND4_X1 i_257_76_16559 (.A1(n_257_449), .A2(n_257_76_16308), .A3(
      n_257_76_16309), .A4(n_257_76_16529), .ZN(n_257_76_16530));
   NOR2_X1 i_257_76_16560 (.A1(n_257_76_16461), .A2(n_257_76_16530), .ZN(
      n_257_76_16531));
   NAND4_X1 i_257_76_16561 (.A1(n_257_76_16525), .A2(n_257_76_16291), .A3(
      n_257_76_16531), .A4(n_257_76_16271), .ZN(n_257_76_16532));
   NOR2_X1 i_257_76_16562 (.A1(n_257_76_16532), .A2(n_257_76_16313), .ZN(
      n_257_76_16533));
   NAND2_X1 i_257_76_16563 (.A1(n_257_76_18083), .A2(n_257_76_16533), .ZN(
      n_257_76_16534));
   NAND3_X1 i_257_76_16564 (.A1(n_257_181), .A2(n_257_76_16292), .A3(
      n_257_76_16293), .ZN(n_257_76_16535));
   INV_X1 i_257_76_16565 (.A(n_257_76_16535), .ZN(n_257_76_16536));
   NAND3_X1 i_257_76_16566 (.A1(n_257_76_16271), .A2(n_257_76_16414), .A3(
      n_257_76_16536), .ZN(n_257_76_16537));
   INV_X1 i_257_76_16567 (.A(n_257_76_16537), .ZN(n_257_76_16538));
   NOR2_X1 i_257_76_16568 (.A1(n_257_76_16274), .A2(n_257_76_17101), .ZN(
      n_257_76_16539));
   NAND3_X1 i_257_76_16569 (.A1(n_257_76_16305), .A2(n_257_76_16539), .A3(
      n_257_76_16348), .ZN(n_257_76_16540));
   INV_X1 i_257_76_16570 (.A(n_257_76_16540), .ZN(n_257_76_16541));
   NAND4_X1 i_257_76_16571 (.A1(n_257_76_16309), .A2(n_257_76_16541), .A3(
      n_257_76_16347), .A4(n_257_76_16342), .ZN(n_257_76_16542));
   INV_X1 i_257_76_16572 (.A(n_257_76_16542), .ZN(n_257_76_16543));
   NAND2_X1 i_257_76_16573 (.A1(n_257_76_16300), .A2(n_257_76_16363), .ZN(
      n_257_76_16544));
   INV_X1 i_257_76_16574 (.A(n_257_76_16544), .ZN(n_257_76_16545));
   NAND3_X1 i_257_76_16575 (.A1(n_257_76_16543), .A2(n_257_76_16545), .A3(
      n_257_76_16512), .ZN(n_257_76_16546));
   NOR2_X1 i_257_76_16576 (.A1(n_257_76_16546), .A2(n_257_76_16372), .ZN(
      n_257_76_16547));
   NAND4_X1 i_257_76_16577 (.A1(n_257_76_16538), .A2(n_257_76_16547), .A3(
      n_257_76_16270), .A4(n_257_76_16291), .ZN(n_257_76_16548));
   INV_X1 i_257_76_16578 (.A(n_257_76_16548), .ZN(n_257_76_16549));
   NAND2_X1 i_257_76_16579 (.A1(n_257_76_18061), .A2(n_257_76_16549), .ZN(
      n_257_76_16550));
   NAND3_X1 i_257_76_16580 (.A1(n_257_76_16523), .A2(n_257_76_16534), .A3(
      n_257_76_16550), .ZN(n_257_76_16551));
   INV_X1 i_257_76_16581 (.A(n_257_76_16551), .ZN(n_257_76_16552));
   NAND2_X1 i_257_76_16582 (.A1(n_257_442), .A2(n_257_896), .ZN(n_257_76_16553));
   NOR2_X1 i_257_76_16583 (.A1(n_257_1088), .A2(n_257_76_16553), .ZN(
      n_257_76_16554));
   NAND2_X1 i_257_76_16584 (.A1(n_257_438), .A2(n_257_76_16554), .ZN(
      n_257_76_16555));
   INV_X1 i_257_76_16585 (.A(n_257_76_16555), .ZN(n_257_76_16556));
   NAND3_X1 i_257_76_16586 (.A1(n_257_76_16299), .A2(n_257_76_16308), .A3(
      n_257_76_16556), .ZN(n_257_76_16557));
   INV_X1 i_257_76_16587 (.A(n_257_76_16557), .ZN(n_257_76_16558));
   NAND2_X1 i_257_76_16588 (.A1(n_257_76_16558), .A2(n_257_76_16272), .ZN(
      n_257_76_16559));
   NOR2_X1 i_257_76_16589 (.A1(n_257_76_16360), .A2(n_257_76_16559), .ZN(
      n_257_76_16560));
   NAND2_X1 i_257_76_16590 (.A1(n_257_76_16270), .A2(n_257_76_16560), .ZN(
      n_257_76_16561));
   INV_X1 i_257_76_16591 (.A(n_257_76_16561), .ZN(n_257_76_16562));
   NAND2_X1 i_257_76_16592 (.A1(n_257_76_18067), .A2(n_257_76_16562), .ZN(
      n_257_76_16563));
   NAND4_X1 i_257_76_16593 (.A1(n_257_76_16339), .A2(n_257_76_16340), .A3(
      n_257_76_16272), .A4(n_257_76_16368), .ZN(n_257_76_16564));
   NOR2_X1 i_257_76_16594 (.A1(n_257_76_16564), .A2(n_257_76_16360), .ZN(
      n_257_76_16565));
   NAND2_X1 i_257_76_16595 (.A1(n_257_378), .A2(n_257_421), .ZN(n_257_76_16566));
   NAND3_X1 i_257_76_16596 (.A1(n_257_76_16302), .A2(n_257_76_16566), .A3(
      n_257_76_16308), .ZN(n_257_76_16567));
   NOR2_X1 i_257_76_16597 (.A1(n_257_76_16364), .A2(n_257_76_16567), .ZN(
      n_257_76_16568));
   NAND2_X1 i_257_76_16598 (.A1(n_257_339), .A2(n_257_422), .ZN(n_257_76_16569));
   NAND3_X1 i_257_76_16599 (.A1(n_257_76_16305), .A2(n_257_76_16569), .A3(
      n_257_76_16348), .ZN(n_257_76_16570));
   INV_X1 i_257_76_16600 (.A(n_257_76_16570), .ZN(n_257_76_16571));
   NAND2_X1 i_257_76_16601 (.A1(n_257_301), .A2(n_257_423), .ZN(n_257_76_16572));
   NAND2_X1 i_257_76_16602 (.A1(n_257_420), .A2(n_257_76_16352), .ZN(
      n_257_76_16573));
   INV_X1 i_257_76_16603 (.A(n_257_76_16573), .ZN(n_257_76_16574));
   NAND2_X1 i_257_76_16604 (.A1(n_257_442), .A2(n_257_498), .ZN(n_257_76_16575));
   INV_X1 i_257_76_16605 (.A(n_257_76_16575), .ZN(n_257_76_16576));
   NAND2_X1 i_257_76_16606 (.A1(n_257_76_16576), .A2(n_257_76_16349), .ZN(
      n_257_76_16577));
   OAI21_X1 i_257_76_16607 (.A(n_257_76_16577), .B1(n_257_428), .B2(
      n_257_76_16575), .ZN(n_257_76_16578));
   NAND2_X1 i_257_76_16608 (.A1(n_257_76_16574), .A2(n_257_76_16578), .ZN(
      n_257_76_16579));
   INV_X1 i_257_76_16609 (.A(n_257_76_16579), .ZN(n_257_76_16580));
   NAND4_X1 i_257_76_16610 (.A1(n_257_76_16344), .A2(n_257_76_16571), .A3(
      n_257_76_16572), .A4(n_257_76_16580), .ZN(n_257_76_16581));
   NAND3_X1 i_257_76_16611 (.A1(n_257_76_16309), .A2(n_257_76_16347), .A3(
      n_257_76_16365), .ZN(n_257_76_16582));
   NOR2_X1 i_257_76_16612 (.A1(n_257_76_16581), .A2(n_257_76_16582), .ZN(
      n_257_76_16583));
   NAND3_X1 i_257_76_16613 (.A1(n_257_76_16298), .A2(n_257_76_16371), .A3(
      n_257_76_16299), .ZN(n_257_76_16584));
   INV_X1 i_257_76_16614 (.A(n_257_76_16584), .ZN(n_257_76_16585));
   NAND4_X1 i_257_76_16615 (.A1(n_257_76_16568), .A2(n_257_76_16583), .A3(
      n_257_76_16401), .A4(n_257_76_16585), .ZN(n_257_76_16586));
   INV_X1 i_257_76_16616 (.A(n_257_76_16586), .ZN(n_257_76_16587));
   NAND4_X1 i_257_76_16617 (.A1(n_257_76_16565), .A2(n_257_76_16587), .A3(
      n_257_76_16270), .A4(n_257_76_16291), .ZN(n_257_76_16588));
   INV_X1 i_257_76_16618 (.A(n_257_76_16588), .ZN(n_257_76_16589));
   NAND2_X1 i_257_76_16619 (.A1(n_257_76_18073), .A2(n_257_76_16589), .ZN(
      n_257_76_16590));
   NAND3_X1 i_257_76_16620 (.A1(n_257_76_16308), .A2(n_257_76_16309), .A3(
      n_257_76_16347), .ZN(n_257_76_16591));
   NOR2_X1 i_257_76_16621 (.A1(n_257_76_16274), .A2(n_257_76_17162), .ZN(
      n_257_76_16592));
   NAND3_X1 i_257_76_16622 (.A1(n_257_76_16305), .A2(n_257_76_16592), .A3(
      n_257_76_16348), .ZN(n_257_76_16593));
   INV_X1 i_257_76_16623 (.A(n_257_76_16593), .ZN(n_257_76_16594));
   NAND3_X1 i_257_76_16624 (.A1(n_257_76_16594), .A2(n_257_142), .A3(
      n_257_76_16342), .ZN(n_257_76_16595));
   NOR2_X1 i_257_76_16625 (.A1(n_257_76_16591), .A2(n_257_76_16595), .ZN(
      n_257_76_16596));
   INV_X1 i_257_76_16626 (.A(n_257_76_16461), .ZN(n_257_76_16597));
   NAND2_X1 i_257_76_16627 (.A1(n_257_76_16298), .A2(n_257_76_16371), .ZN(
      n_257_76_16598));
   INV_X1 i_257_76_16628 (.A(n_257_76_16598), .ZN(n_257_76_16599));
   NAND3_X1 i_257_76_16629 (.A1(n_257_76_16596), .A2(n_257_76_16597), .A3(
      n_257_76_16599), .ZN(n_257_76_16600));
   INV_X1 i_257_76_16630 (.A(n_257_76_16454), .ZN(n_257_76_16601));
   NAND4_X1 i_257_76_16631 (.A1(n_257_76_16601), .A2(n_257_76_16272), .A3(
      n_257_76_16368), .A4(n_257_76_16292), .ZN(n_257_76_16602));
   NOR2_X1 i_257_76_16632 (.A1(n_257_76_16600), .A2(n_257_76_16602), .ZN(
      n_257_76_16603));
   NAND2_X1 i_257_76_16633 (.A1(n_257_76_16291), .A2(n_257_76_16271), .ZN(
      n_257_76_16604));
   INV_X1 i_257_76_16634 (.A(n_257_76_16604), .ZN(n_257_76_16605));
   NAND3_X1 i_257_76_16635 (.A1(n_257_76_16603), .A2(n_257_76_16605), .A3(
      n_257_76_16270), .ZN(n_257_76_16606));
   INV_X1 i_257_76_16636 (.A(n_257_76_16606), .ZN(n_257_76_16607));
   NAND2_X1 i_257_76_16637 (.A1(n_257_76_18068), .A2(n_257_76_16607), .ZN(
      n_257_76_16608));
   NAND3_X1 i_257_76_16638 (.A1(n_257_76_16563), .A2(n_257_76_16590), .A3(
      n_257_76_16608), .ZN(n_257_76_16609));
   INV_X1 i_257_76_16639 (.A(n_257_76_16609), .ZN(n_257_76_16610));
   NAND2_X1 i_257_76_16640 (.A1(n_257_794), .A2(n_257_442), .ZN(n_257_76_16611));
   NOR2_X1 i_257_76_16641 (.A1(n_257_1088), .A2(n_257_76_16611), .ZN(
      n_257_76_16612));
   NAND4_X1 i_257_76_16642 (.A1(n_257_447), .A2(n_257_76_16308), .A3(
      n_257_76_16309), .A4(n_257_76_16612), .ZN(n_257_76_16613));
   NOR2_X1 i_257_76_16643 (.A1(n_257_76_16461), .A2(n_257_76_16613), .ZN(
      n_257_76_16614));
   NAND3_X1 i_257_76_16644 (.A1(n_257_76_16614), .A2(n_257_76_16271), .A3(
      n_257_76_16497), .ZN(n_257_76_16615));
   NOR2_X1 i_257_76_16645 (.A1(n_257_76_16313), .A2(n_257_76_16615), .ZN(
      n_257_76_16616));
   NAND3_X1 i_257_76_16646 (.A1(n_257_76_16300), .A2(n_257_76_16302), .A3(
      n_257_76_16308), .ZN(n_257_76_16617));
   NOR2_X1 i_257_76_16647 (.A1(n_257_76_16274), .A2(n_257_76_17183), .ZN(
      n_257_76_16618));
   NAND3_X1 i_257_76_16648 (.A1(n_257_76_16305), .A2(n_257_76_16618), .A3(
      n_257_76_16348), .ZN(n_257_76_16619));
   INV_X1 i_257_76_16649 (.A(n_257_76_16619), .ZN(n_257_76_16620));
   NAND4_X1 i_257_76_16650 (.A1(n_257_76_16309), .A2(n_257_76_16620), .A3(
      n_257_76_16347), .A4(n_257_76_16342), .ZN(n_257_76_16621));
   NOR2_X1 i_257_76_16651 (.A1(n_257_76_16617), .A2(n_257_76_16621), .ZN(
      n_257_76_16622));
   NAND3_X1 i_257_76_16652 (.A1(n_257_76_16371), .A2(n_257_76_16299), .A3(
      n_257_104), .ZN(n_257_76_16623));
   INV_X1 i_257_76_16653 (.A(n_257_76_16623), .ZN(n_257_76_16624));
   NAND3_X1 i_257_76_16654 (.A1(n_257_76_16622), .A2(n_257_76_16483), .A3(
      n_257_76_16624), .ZN(n_257_76_16625));
   INV_X1 i_257_76_16655 (.A(n_257_76_16625), .ZN(n_257_76_16626));
   NAND4_X1 i_257_76_16656 (.A1(n_257_76_16626), .A2(n_257_76_16270), .A3(
      n_257_76_16472), .A4(n_257_76_16291), .ZN(n_257_76_16627));
   INV_X1 i_257_76_16657 (.A(n_257_76_16627), .ZN(n_257_76_16628));
   AOI22_X1 i_257_76_16658 (.A1(n_257_76_18085), .A2(n_257_76_16616), .B1(
      n_257_76_18080), .B2(n_257_76_16628), .ZN(n_257_76_16629));
   NAND3_X1 i_257_76_16659 (.A1(n_257_76_16552), .A2(n_257_76_16610), .A3(
      n_257_76_16629), .ZN(n_257_76_16630));
   NAND4_X1 i_257_76_16660 (.A1(n_257_76_16272), .A2(n_257_76_16292), .A3(
      n_257_76_16293), .A4(n_257_76_16298), .ZN(n_257_76_16631));
   NAND4_X1 i_257_76_16661 (.A1(n_257_76_16308), .A2(n_257_76_16309), .A3(
      n_257_448), .A4(n_257_76_17979), .ZN(n_257_76_16632));
   INV_X1 i_257_76_16662 (.A(n_257_76_16632), .ZN(n_257_76_16633));
   NAND2_X1 i_257_76_16663 (.A1(n_257_76_16300), .A2(n_257_76_16302), .ZN(
      n_257_76_16634));
   INV_X1 i_257_76_16664 (.A(n_257_76_16634), .ZN(n_257_76_16635));
   NAND3_X1 i_257_76_16665 (.A1(n_257_76_16633), .A2(n_257_76_16635), .A3(
      n_257_76_16299), .ZN(n_257_76_16636));
   NOR2_X1 i_257_76_16666 (.A1(n_257_76_16631), .A2(n_257_76_16636), .ZN(
      n_257_76_16637));
   NAND2_X1 i_257_76_16667 (.A1(n_257_76_16271), .A2(n_257_698), .ZN(
      n_257_76_16638));
   INV_X1 i_257_76_16668 (.A(n_257_76_16638), .ZN(n_257_76_16639));
   NAND3_X1 i_257_76_16669 (.A1(n_257_76_16637), .A2(n_257_76_16270), .A3(
      n_257_76_16639), .ZN(n_257_76_16640));
   INV_X1 i_257_76_16670 (.A(n_257_76_16640), .ZN(n_257_76_16641));
   NAND2_X1 i_257_76_16671 (.A1(n_257_76_18079), .A2(n_257_76_16641), .ZN(
      n_257_76_16642));
   NAND2_X1 i_257_76_16672 (.A1(n_257_76_16271), .A2(n_257_76_16272), .ZN(
      n_257_76_16643));
   INV_X1 i_257_76_16673 (.A(n_257_76_16643), .ZN(n_257_76_16644));
   NAND3_X1 i_257_76_16674 (.A1(n_257_76_16270), .A2(n_257_76_16644), .A3(
      n_257_76_16291), .ZN(n_257_76_16645));
   NOR2_X1 i_257_76_16675 (.A1(n_257_76_16482), .A2(n_257_76_16484), .ZN(
      n_257_76_16646));
   NAND4_X1 i_257_76_16676 (.A1(n_257_76_16362), .A2(n_257_76_16363), .A3(
      n_257_76_16302), .A4(n_257_76_16308), .ZN(n_257_76_16647));
   NAND2_X1 i_257_76_16677 (.A1(n_257_76_16347), .A2(n_257_76_16365), .ZN(
      n_257_76_16648));
   INV_X1 i_257_76_16678 (.A(n_257_76_16648), .ZN(n_257_76_16649));
   NAND2_X1 i_257_76_16679 (.A1(n_257_425), .A2(n_257_76_16352), .ZN(
      n_257_76_16650));
   INV_X1 i_257_76_16680 (.A(n_257_76_16650), .ZN(n_257_76_16651));
   NAND2_X1 i_257_76_16681 (.A1(n_257_76_16651), .A2(n_257_76_16351), .ZN(
      n_257_76_16652));
   INV_X1 i_257_76_16682 (.A(n_257_76_16652), .ZN(n_257_76_16653));
   NAND4_X1 i_257_76_16683 (.A1(n_257_76_16653), .A2(n_257_76_16342), .A3(
      n_257_76_16305), .A4(n_257_76_16348), .ZN(n_257_76_16654));
   INV_X1 i_257_76_16684 (.A(n_257_76_16654), .ZN(n_257_76_16655));
   NAND3_X1 i_257_76_16685 (.A1(n_257_76_16649), .A2(n_257_76_16655), .A3(
      n_257_76_16309), .ZN(n_257_76_16656));
   NOR2_X1 i_257_76_16686 (.A1(n_257_76_16647), .A2(n_257_76_16656), .ZN(
      n_257_76_16657));
   NAND3_X1 i_257_76_16687 (.A1(n_257_76_16368), .A2(n_257_261), .A3(
      n_257_76_16292), .ZN(n_257_76_16658));
   INV_X1 i_257_76_16688 (.A(n_257_76_16658), .ZN(n_257_76_16659));
   NAND4_X1 i_257_76_16689 (.A1(n_257_76_16646), .A2(n_257_76_16657), .A3(
      n_257_76_16659), .A4(n_257_76_16339), .ZN(n_257_76_16660));
   NOR2_X1 i_257_76_16690 (.A1(n_257_76_16645), .A2(n_257_76_16660), .ZN(
      n_257_76_16661));
   NAND2_X1 i_257_76_16691 (.A1(n_257_76_18064), .A2(n_257_76_16661), .ZN(
      n_257_76_16662));
   NAND4_X1 i_257_76_16692 (.A1(n_257_76_16294), .A2(n_257_76_16298), .A3(
      n_257_76_16371), .A4(n_257_76_16308), .ZN(n_257_76_16663));
   NAND2_X1 i_257_76_16693 (.A1(n_257_76_16368), .A2(n_257_76_16293), .ZN(
      n_257_76_16664));
   NOR2_X1 i_257_76_16694 (.A1(n_257_76_16663), .A2(n_257_76_16664), .ZN(
      n_257_76_16665));
   NAND3_X1 i_257_76_16695 (.A1(n_257_76_16339), .A2(n_257_76_16340), .A3(
      n_257_76_16272), .ZN(n_257_76_16666));
   INV_X1 i_257_76_16696 (.A(n_257_76_16666), .ZN(n_257_76_16667));
   NAND4_X1 i_257_76_16697 (.A1(n_257_76_16665), .A2(n_257_76_16667), .A3(
      n_257_76_16291), .A4(n_257_76_16271), .ZN(n_257_76_16668));
   NAND4_X1 i_257_76_16698 (.A1(n_257_76_16347), .A2(n_257_76_16365), .A3(
      n_257_76_16572), .A4(n_257_378), .ZN(n_257_76_16669));
   NAND2_X1 i_257_76_16699 (.A1(n_257_76_16305), .A2(n_257_76_16569), .ZN(
      n_257_76_16670));
   INV_X1 i_257_76_16700 (.A(n_257_76_16670), .ZN(n_257_76_16671));
   NAND2_X1 i_257_76_16701 (.A1(n_257_421), .A2(n_257_76_16352), .ZN(
      n_257_76_16672));
   INV_X1 i_257_76_16702 (.A(n_257_76_16672), .ZN(n_257_76_16673));
   NAND3_X1 i_257_76_16703 (.A1(n_257_76_16348), .A2(n_257_76_16351), .A3(
      n_257_76_16673), .ZN(n_257_76_16674));
   INV_X1 i_257_76_16704 (.A(n_257_76_16674), .ZN(n_257_76_16675));
   NAND4_X1 i_257_76_16705 (.A1(n_257_76_16671), .A2(n_257_76_16675), .A3(
      n_257_76_16341), .A4(n_257_76_16342), .ZN(n_257_76_16676));
   NOR2_X1 i_257_76_16706 (.A1(n_257_76_16669), .A2(n_257_76_16676), .ZN(
      n_257_76_16677));
   NAND3_X1 i_257_76_16707 (.A1(n_257_76_16292), .A2(n_257_76_16299), .A3(
      n_257_76_16300), .ZN(n_257_76_16678));
   INV_X1 i_257_76_16708 (.A(n_257_76_16678), .ZN(n_257_76_16679));
   NAND4_X1 i_257_76_16709 (.A1(n_257_76_16362), .A2(n_257_76_16363), .A3(
      n_257_76_16302), .A4(n_257_76_16309), .ZN(n_257_76_16680));
   INV_X1 i_257_76_16710 (.A(n_257_76_16680), .ZN(n_257_76_16681));
   NAND3_X1 i_257_76_16711 (.A1(n_257_76_16677), .A2(n_257_76_16679), .A3(
      n_257_76_16681), .ZN(n_257_76_16682));
   INV_X1 i_257_76_16712 (.A(n_257_76_16682), .ZN(n_257_76_16683));
   NAND2_X1 i_257_76_16713 (.A1(n_257_76_16270), .A2(n_257_76_16683), .ZN(
      n_257_76_16684));
   NOR2_X1 i_257_76_16714 (.A1(n_257_76_16668), .A2(n_257_76_16684), .ZN(
      n_257_76_16685));
   NAND2_X1 i_257_76_16715 (.A1(n_257_76_18082), .A2(n_257_76_16685), .ZN(
      n_257_76_16686));
   NAND3_X1 i_257_76_16716 (.A1(n_257_76_16642), .A2(n_257_76_16662), .A3(
      n_257_76_16686), .ZN(n_257_76_16687));
   INV_X1 i_257_76_16717 (.A(n_257_76_16687), .ZN(n_257_76_16688));
   NAND3_X1 i_257_76_16718 (.A1(n_257_76_16302), .A2(n_257_76_16308), .A3(
      n_257_76_16309), .ZN(n_257_76_16689));
   NOR2_X1 i_257_76_16719 (.A1(n_257_76_16544), .A2(n_257_76_16689), .ZN(
      n_257_76_16690));
   NAND3_X1 i_257_76_16720 (.A1(n_257_76_16690), .A2(n_257_76_16401), .A3(
      n_257_76_16585), .ZN(n_257_76_16691));
   INV_X1 i_257_76_16721 (.A(n_257_76_16691), .ZN(n_257_76_16692));
   NAND2_X1 i_257_76_16722 (.A1(n_257_76_16351), .A2(n_257_76_16352), .ZN(
      n_257_76_16693));
   INV_X1 i_257_76_16723 (.A(n_257_76_16693), .ZN(n_257_76_16694));
   NAND3_X1 i_257_76_16724 (.A1(n_257_76_16694), .A2(n_257_76_16342), .A3(
      n_257_427), .ZN(n_257_76_16695));
   INV_X1 i_257_76_16725 (.A(n_257_76_16695), .ZN(n_257_76_16696));
   NAND3_X1 i_257_76_16726 (.A1(n_257_76_16305), .A2(n_257_76_16348), .A3(
      n_257_221), .ZN(n_257_76_16697));
   INV_X1 i_257_76_16727 (.A(n_257_76_16697), .ZN(n_257_76_16698));
   NAND3_X1 i_257_76_16728 (.A1(n_257_76_16696), .A2(n_257_76_16347), .A3(
      n_257_76_16698), .ZN(n_257_76_16699));
   INV_X1 i_257_76_16729 (.A(n_257_76_16699), .ZN(n_257_76_16700));
   NAND4_X1 i_257_76_16730 (.A1(n_257_76_16339), .A2(n_257_76_16700), .A3(
      n_257_76_16272), .A4(n_257_76_16368), .ZN(n_257_76_16701));
   INV_X1 i_257_76_16731 (.A(n_257_76_16701), .ZN(n_257_76_16702));
   NAND2_X1 i_257_76_16732 (.A1(n_257_76_16692), .A2(n_257_76_16702), .ZN(
      n_257_76_16703));
   NOR3_X1 i_257_76_16733 (.A1(n_257_76_16703), .A2(n_257_76_16313), .A3(
      n_257_76_16604), .ZN(n_257_76_16704));
   NAND2_X1 i_257_76_16734 (.A1(n_257_76_18065), .A2(n_257_76_16704), .ZN(
      n_257_76_16705));
   NAND4_X1 i_257_76_16735 (.A1(n_257_76_16298), .A2(n_257_76_16299), .A3(
      n_257_76_16300), .A4(n_257_76_16302), .ZN(n_257_76_16706));
   NAND2_X1 i_257_76_16736 (.A1(n_257_76_16308), .A2(n_257_76_16309), .ZN(
      n_257_76_16707));
   INV_X1 i_257_76_16737 (.A(n_257_76_16707), .ZN(n_257_76_16708));
   NAND3_X1 i_257_76_16738 (.A1(n_257_76_16347), .A2(n_257_76_17979), .A3(
      n_257_481), .ZN(n_257_76_16709));
   INV_X1 i_257_76_16739 (.A(n_257_76_16709), .ZN(n_257_76_16710));
   NAND3_X1 i_257_76_16740 (.A1(n_257_76_16708), .A2(n_257_76_16710), .A3(
      n_257_451), .ZN(n_257_76_16711));
   NOR2_X1 i_257_76_16741 (.A1(n_257_76_16706), .A2(n_257_76_16711), .ZN(
      n_257_76_16712));
   NAND4_X1 i_257_76_16742 (.A1(n_257_76_16712), .A2(n_257_76_16291), .A3(
      n_257_76_16297), .A4(n_257_76_16271), .ZN(n_257_76_16713));
   NOR2_X1 i_257_76_16743 (.A1(n_257_76_16713), .A2(n_257_76_16313), .ZN(
      n_257_76_16714));
   NAND2_X1 i_257_76_16744 (.A1(n_257_76_18063), .A2(n_257_76_16714), .ZN(
      n_257_76_16715));
   NAND2_X1 i_257_76_16745 (.A1(n_257_76_16342), .A2(n_257_76_16694), .ZN(
      n_257_76_16716));
   INV_X1 i_257_76_16746 (.A(n_257_76_16716), .ZN(n_257_76_16717));
   NAND4_X1 i_257_76_16747 (.A1(n_257_76_16305), .A2(n_257_76_16348), .A3(
      n_257_530), .A4(n_257_424), .ZN(n_257_76_16718));
   INV_X1 i_257_76_16748 (.A(n_257_76_16718), .ZN(n_257_76_16719));
   NAND3_X1 i_257_76_16749 (.A1(n_257_76_16717), .A2(n_257_76_16719), .A3(
      n_257_76_16347), .ZN(n_257_76_16720));
   INV_X1 i_257_76_16750 (.A(n_257_76_16720), .ZN(n_257_76_16721));
   NAND4_X1 i_257_76_16751 (.A1(n_257_76_16339), .A2(n_257_76_16340), .A3(
      n_257_76_16272), .A4(n_257_76_16721), .ZN(n_257_76_16722));
   NOR2_X1 i_257_76_16752 (.A1(n_257_76_16722), .A2(n_257_76_16360), .ZN(
      n_257_76_16723));
   NAND4_X1 i_257_76_16753 (.A1(n_257_76_16723), .A2(n_257_76_16375), .A3(
      n_257_76_16270), .A4(n_257_76_16291), .ZN(n_257_76_16724));
   INV_X1 i_257_76_16754 (.A(n_257_76_16724), .ZN(n_257_76_16725));
   NAND2_X1 i_257_76_16755 (.A1(n_257_76_18062), .A2(n_257_76_16725), .ZN(
      n_257_76_16726));
   NAND3_X1 i_257_76_16756 (.A1(n_257_76_16705), .A2(n_257_76_16715), .A3(
      n_257_76_16726), .ZN(n_257_76_16727));
   INV_X1 i_257_76_16757 (.A(n_257_76_16727), .ZN(n_257_76_16728));
   NAND2_X1 i_257_76_16758 (.A1(n_257_76_16300), .A2(n_257_76_16362), .ZN(
      n_257_76_16729));
   NOR2_X1 i_257_76_16759 (.A1(n_257_76_16402), .A2(n_257_76_16729), .ZN(
      n_257_76_16730));
   NAND4_X1 i_257_76_16760 (.A1(n_257_76_16344), .A2(n_257_76_16365), .A3(
      n_257_76_16572), .A4(n_257_76_16437), .ZN(n_257_76_16731));
   NOR2_X1 i_257_76_16761 (.A1(n_257_76_16693), .A2(n_257_76_16569), .ZN(
      n_257_76_16732));
   NAND3_X1 i_257_76_16762 (.A1(n_257_76_16309), .A2(n_257_76_16732), .A3(
      n_257_76_16347), .ZN(n_257_76_16733));
   NOR2_X1 i_257_76_16763 (.A1(n_257_76_16731), .A2(n_257_76_16733), .ZN(
      n_257_76_16734));
   NAND4_X1 i_257_76_16764 (.A1(n_257_76_16730), .A2(n_257_76_16734), .A3(
      n_257_76_16401), .A4(n_257_76_16585), .ZN(n_257_76_16735));
   INV_X1 i_257_76_16765 (.A(n_257_76_16735), .ZN(n_257_76_16736));
   NAND4_X1 i_257_76_16766 (.A1(n_257_76_16565), .A2(n_257_76_16736), .A3(
      n_257_76_16270), .A4(n_257_76_16291), .ZN(n_257_76_16737));
   INV_X1 i_257_76_16767 (.A(n_257_76_16737), .ZN(n_257_76_16738));
   NAND2_X1 i_257_76_16768 (.A1(n_257_342), .A2(n_257_76_16738), .ZN(
      n_257_76_16739));
   NAND3_X1 i_257_76_16769 (.A1(n_257_76_16347), .A2(n_257_76_16365), .A3(
      n_257_76_16572), .ZN(n_257_76_16740));
   INV_X1 i_257_76_16770 (.A(n_257_76_16740), .ZN(n_257_76_16741));
   NAND3_X1 i_257_76_16771 (.A1(n_257_76_16341), .A2(n_257_76_16342), .A3(
      n_257_76_16305), .ZN(n_257_76_16742));
   NAND2_X1 i_257_76_16772 (.A1(n_257_428), .A2(n_257_594), .ZN(n_257_76_16743));
   NAND2_X1 i_257_76_16773 (.A1(n_257_442), .A2(n_257_417), .ZN(n_257_76_16744));
   INV_X1 i_257_76_16774 (.A(n_257_76_16744), .ZN(n_257_76_16745));
   NAND2_X1 i_257_76_16775 (.A1(n_257_484), .A2(n_257_76_16745), .ZN(
      n_257_76_16746));
   INV_X1 i_257_76_16776 (.A(n_257_76_16746), .ZN(n_257_76_16747));
   NAND3_X1 i_257_76_16777 (.A1(n_257_76_16743), .A2(n_257_76_16352), .A3(
      n_257_76_16747), .ZN(n_257_76_16748));
   INV_X1 i_257_76_16778 (.A(n_257_76_16748), .ZN(n_257_76_16749));
   NAND2_X1 i_257_76_16779 (.A1(n_257_420), .A2(n_257_498), .ZN(n_257_76_16750));
   NAND4_X1 i_257_76_16780 (.A1(n_257_76_16749), .A2(n_257_76_16569), .A3(
      n_257_76_16348), .A4(n_257_76_16750), .ZN(n_257_76_16751));
   NOR2_X1 i_257_76_16781 (.A1(n_257_76_16742), .A2(n_257_76_16751), .ZN(
      n_257_76_16752));
   NAND2_X1 i_257_76_16782 (.A1(n_257_76_16741), .A2(n_257_76_16752), .ZN(
      n_257_76_16753));
   NAND4_X1 i_257_76_16783 (.A1(n_257_76_16302), .A2(n_257_76_16566), .A3(
      n_257_76_16308), .A4(n_257_76_16309), .ZN(n_257_76_16754));
   NOR2_X1 i_257_76_16784 (.A1(n_257_76_16753), .A2(n_257_76_16754), .ZN(
      n_257_76_16755));
   NAND3_X1 i_257_76_16785 (.A1(n_257_76_16755), .A2(n_257_76_16291), .A3(
      n_257_76_16271), .ZN(n_257_76_16756));
   INV_X1 i_257_76_16786 (.A(n_257_76_16756), .ZN(n_257_76_16757));
   INV_X1 i_257_76_16787 (.A(n_257_76_16364), .ZN(n_257_76_16758));
   NAND3_X1 i_257_76_16788 (.A1(n_257_76_16401), .A2(n_257_76_16585), .A3(
      n_257_76_16758), .ZN(n_257_76_16759));
   NOR2_X1 i_257_76_16789 (.A1(n_257_76_16759), .A2(n_257_76_16564), .ZN(
      n_257_76_16760));
   NAND3_X1 i_257_76_16790 (.A1(n_257_76_16757), .A2(n_257_76_16760), .A3(
      n_257_76_16270), .ZN(n_257_76_16761));
   INV_X1 i_257_76_16791 (.A(n_257_76_16761), .ZN(n_257_76_16762));
   NAND2_X1 i_257_76_16792 (.A1(n_257_76_18060), .A2(n_257_76_16762), .ZN(
      n_257_76_16763));
   NAND2_X1 i_257_76_16793 (.A1(n_257_698), .A2(n_257_76_17958), .ZN(
      n_257_76_16764));
   NAND2_X1 i_257_76_16794 (.A1(n_257_76_16448), .A2(n_257_76_16764), .ZN(
      n_257_76_16765));
   NAND2_X1 i_257_76_16795 (.A1(n_257_1024), .A2(n_257_76_17964), .ZN(
      n_257_76_16766));
   NAND2_X1 i_257_76_16796 (.A1(n_257_992), .A2(n_257_442), .ZN(n_257_76_16767));
   INV_X1 i_257_76_16797 (.A(n_257_76_16767), .ZN(n_257_76_16768));
   AOI22_X1 i_257_76_16798 (.A1(n_257_181), .A2(n_257_76_17331), .B1(n_257_441), 
      .B2(n_257_76_16768), .ZN(n_257_76_16769));
   NAND2_X1 i_257_76_16799 (.A1(n_257_76_16766), .A2(n_257_76_16769), .ZN(
      n_257_76_16770));
   NOR2_X1 i_257_76_16800 (.A1(n_257_76_16765), .A2(n_257_76_16770), .ZN(
      n_257_76_16771));
   NAND2_X1 i_257_76_16801 (.A1(n_257_104), .A2(n_257_76_17932), .ZN(
      n_257_76_16772));
   NAND2_X1 i_257_76_16802 (.A1(n_257_76_16772), .A2(n_257_76_16699), .ZN(
      n_257_76_16773));
   NAND2_X1 i_257_76_16803 (.A1(n_257_76_16357), .A2(n_257_76_16720), .ZN(
      n_257_76_16774));
   NOR2_X1 i_257_76_16804 (.A1(n_257_76_16773), .A2(n_257_76_16774), .ZN(
      n_257_76_16775));
   NAND2_X1 i_257_76_16805 (.A1(n_257_762), .A2(n_257_76_17935), .ZN(
      n_257_76_16776));
   NAND2_X1 i_257_76_16806 (.A1(n_257_858), .A2(n_257_442), .ZN(n_257_76_16777));
   INV_X1 i_257_76_16807 (.A(n_257_76_16777), .ZN(n_257_76_16778));
   NAND2_X1 i_257_76_16808 (.A1(n_257_446), .A2(n_257_76_16778), .ZN(
      n_257_76_16779));
   NAND2_X1 i_257_76_16809 (.A1(n_257_76_16776), .A2(n_257_76_16779), .ZN(
      n_257_76_16780));
   INV_X1 i_257_76_16810 (.A(n_257_76_16526), .ZN(n_257_76_16781));
   NAND2_X1 i_257_76_16811 (.A1(n_257_449), .A2(n_257_76_16781), .ZN(
      n_257_76_16782));
   NAND2_X1 i_257_76_16812 (.A1(n_257_481), .A2(n_257_442), .ZN(n_257_76_16783));
   INV_X1 i_257_76_16813 (.A(n_257_76_16783), .ZN(n_257_76_16784));
   NAND2_X1 i_257_76_16814 (.A1(n_257_451), .A2(n_257_76_16784), .ZN(
      n_257_76_16785));
   NAND2_X1 i_257_76_16815 (.A1(n_257_76_16782), .A2(n_257_76_16785), .ZN(
      n_257_76_16786));
   NOR2_X1 i_257_76_16816 (.A1(n_257_76_16780), .A2(n_257_76_16786), .ZN(
      n_257_76_16787));
   NAND2_X1 i_257_76_16817 (.A1(n_257_76_16775), .A2(n_257_76_16787), .ZN(
      n_257_76_16788));
   NAND2_X1 i_257_76_16818 (.A1(n_257_890), .A2(n_257_76_17903), .ZN(
      n_257_76_16789));
   NAND2_X1 i_257_76_16819 (.A1(n_257_960), .A2(n_257_442), .ZN(n_257_76_16790));
   INV_X1 i_257_76_16820 (.A(n_257_76_16790), .ZN(n_257_76_16791));
   NAND2_X1 i_257_76_16821 (.A1(n_257_440), .A2(n_257_76_16791), .ZN(
      n_257_76_16792));
   NAND2_X1 i_257_76_16822 (.A1(n_257_76_16789), .A2(n_257_76_16792), .ZN(
      n_257_76_16793));
   INV_X1 i_257_76_16823 (.A(n_257_76_16732), .ZN(n_257_76_16794));
   INV_X1 i_257_76_16824 (.A(n_257_438), .ZN(n_257_76_16795));
   OAI21_X1 i_257_76_16825 (.A(n_257_76_16794), .B1(n_257_76_16795), .B2(
      n_257_76_16553), .ZN(n_257_76_16796));
   NOR2_X1 i_257_76_16826 (.A1(n_257_76_16793), .A2(n_257_76_16796), .ZN(
      n_257_76_16797));
   NAND2_X1 i_257_76_16827 (.A1(n_257_64), .A2(n_257_76_17918), .ZN(
      n_257_76_16798));
   NAND2_X1 i_257_76_16828 (.A1(n_257_76_16798), .A2(n_257_76_16579), .ZN(
      n_257_76_16799));
   INV_X1 i_257_76_16829 (.A(n_257_76_16799), .ZN(n_257_76_16800));
   NAND2_X1 i_257_76_16830 (.A1(n_257_658), .A2(n_257_76_17928), .ZN(
      n_257_76_16801));
   NAND2_X1 i_257_76_16831 (.A1(n_257_76_16800), .A2(n_257_76_16801), .ZN(
      n_257_76_16802));
   NAND3_X1 i_257_76_16832 (.A1(n_257_730), .A2(n_257_435), .A3(n_257_442), 
      .ZN(n_257_76_16803));
   INV_X1 i_257_76_16833 (.A(n_257_76_16473), .ZN(n_257_76_16804));
   NAND2_X1 i_257_76_16834 (.A1(n_257_432), .A2(n_257_76_16804), .ZN(
      n_257_76_16805));
   NAND2_X1 i_257_76_16835 (.A1(n_257_76_16803), .A2(n_257_76_16805), .ZN(
      n_257_76_16806));
   INV_X1 i_257_76_16836 (.A(n_257_76_16806), .ZN(n_257_76_16807));
   NAND2_X1 i_257_76_16837 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[29]), 
      .ZN(n_257_76_16808));
   NAND2_X1 i_257_76_16838 (.A1(n_257_1088), .A2(n_257_76_16808), .ZN(
      n_257_76_16809));
   INV_X1 i_257_76_16839 (.A(n_257_428), .ZN(n_257_76_16810));
   NAND2_X1 i_257_76_16840 (.A1(n_257_76_16808), .A2(n_257_594), .ZN(
      n_257_76_16811));
   OAI21_X1 i_257_76_16841 (.A(n_257_76_16809), .B1(n_257_76_16810), .B2(
      n_257_76_16811), .ZN(n_257_76_16812));
   INV_X1 i_257_76_16842 (.A(Small_Packet_Data_Size[29]), .ZN(n_257_76_16813));
   NOR2_X1 i_257_76_16843 (.A1(n_257_484), .A2(n_257_76_16813), .ZN(
      n_257_76_16814));
   INV_X1 i_257_76_16844 (.A(n_257_417), .ZN(n_257_76_16815));
   NAND2_X1 i_257_76_16845 (.A1(n_257_76_16815), .A2(Small_Packet_Data_Size[29]), 
      .ZN(n_257_76_16816));
   NAND2_X1 i_257_76_16846 (.A1(n_257_76_16808), .A2(n_257_76_16816), .ZN(
      n_257_76_16817));
   NOR2_X1 i_257_76_16847 (.A1(n_257_76_16814), .A2(n_257_76_16817), .ZN(
      n_257_76_16818));
   NOR2_X1 i_257_76_16848 (.A1(n_257_76_16812), .A2(n_257_76_16818), .ZN(
      n_257_76_16819));
   NAND2_X1 i_257_76_16849 (.A1(n_257_76_16807), .A2(n_257_76_16819), .ZN(
      n_257_76_16820));
   NOR2_X1 i_257_76_16850 (.A1(n_257_76_16802), .A2(n_257_76_16820), .ZN(
      n_257_76_16821));
   NAND2_X1 i_257_76_16851 (.A1(n_257_76_16797), .A2(n_257_76_16821), .ZN(
      n_257_76_16822));
   INV_X1 i_257_76_16852 (.A(n_257_76_16822), .ZN(n_257_76_16823));
   NAND2_X1 i_257_76_16853 (.A1(n_257_76_17940), .A2(n_257_928), .ZN(
      n_257_76_16824));
   INV_X1 i_257_76_16854 (.A(n_257_76_16611), .ZN(n_257_76_16825));
   NAND2_X1 i_257_76_16855 (.A1(n_257_447), .A2(n_257_76_16825), .ZN(
      n_257_76_16826));
   NAND2_X1 i_257_76_16856 (.A1(n_257_76_16824), .A2(n_257_76_16826), .ZN(
      n_257_76_16827));
   NAND2_X1 i_257_76_16857 (.A1(n_257_826), .A2(n_257_76_17952), .ZN(
      n_257_76_16828));
   NAND2_X1 i_257_76_16858 (.A1(n_257_142), .A2(n_257_76_17925), .ZN(
      n_257_76_16829));
   NAND2_X1 i_257_76_16859 (.A1(n_257_76_16828), .A2(n_257_76_16829), .ZN(
      n_257_76_16830));
   NOR2_X1 i_257_76_16860 (.A1(n_257_76_16827), .A2(n_257_76_16830), .ZN(
      n_257_76_16831));
   NAND2_X1 i_257_76_16861 (.A1(n_257_76_16823), .A2(n_257_76_16831), .ZN(
      n_257_76_16832));
   NOR2_X1 i_257_76_16862 (.A1(n_257_76_16788), .A2(n_257_76_16832), .ZN(
      n_257_76_16833));
   NAND2_X1 i_257_76_16863 (.A1(n_257_76_16771), .A2(n_257_76_16833), .ZN(
      n_257_76_16834));
   INV_X1 i_257_76_16864 (.A(n_257_76_16834), .ZN(n_257_76_16835));
   INV_X1 i_257_76_16865 (.A(n_257_1056), .ZN(n_257_76_16836));
   OAI21_X1 i_257_76_16866 (.A(n_257_76_16682), .B1(n_257_76_16836), .B2(
      n_257_76_17968), .ZN(n_257_76_16837));
   INV_X1 i_257_76_16867 (.A(n_257_76_16660), .ZN(n_257_76_16838));
   NOR2_X1 i_257_76_16868 (.A1(n_257_76_16837), .A2(n_257_76_16838), .ZN(
      n_257_76_16839));
   NAND2_X1 i_257_76_16869 (.A1(n_257_76_16835), .A2(n_257_76_16839), .ZN(
      n_257_76_16840));
   NAND3_X1 i_257_76_16870 (.A1(n_257_76_16739), .A2(n_257_76_16763), .A3(
      n_257_76_16840), .ZN(n_257_76_16841));
   INV_X1 i_257_76_16871 (.A(n_257_76_16841), .ZN(n_257_76_16842));
   NAND3_X1 i_257_76_16872 (.A1(n_257_76_16688), .A2(n_257_76_16728), .A3(
      n_257_76_16842), .ZN(n_257_76_16843));
   NOR2_X1 i_257_76_16873 (.A1(n_257_76_16630), .A2(n_257_76_16843), .ZN(
      n_257_76_16844));
   NAND2_X1 i_257_76_16874 (.A1(n_257_76_16511), .A2(n_257_76_16844), .ZN(n_29));
   NAND2_X1 i_257_76_16875 (.A1(n_257_1057), .A2(n_257_443), .ZN(n_257_76_16845));
   NAND2_X1 i_257_76_16876 (.A1(n_257_1025), .A2(n_257_444), .ZN(n_257_76_16846));
   NAND2_X1 i_257_76_16877 (.A1(n_257_441), .A2(n_257_993), .ZN(n_257_76_16847));
   NOR2_X1 i_257_76_16878 (.A1(n_257_1089), .A2(n_257_76_17412), .ZN(
      n_257_76_16848));
   INV_X1 i_257_76_16879 (.A(n_257_76_16848), .ZN(n_257_76_16849));
   INV_X1 i_257_76_16880 (.A(n_257_961), .ZN(n_257_76_16850));
   NOR2_X1 i_257_76_16881 (.A1(n_257_76_16849), .A2(n_257_76_16850), .ZN(
      n_257_76_16851));
   NAND2_X1 i_257_76_16882 (.A1(n_257_440), .A2(n_257_76_16851), .ZN(
      n_257_76_16852));
   INV_X1 i_257_76_16883 (.A(n_257_76_16852), .ZN(n_257_76_16853));
   NAND2_X1 i_257_76_16884 (.A1(n_257_76_16847), .A2(n_257_76_16853), .ZN(
      n_257_76_16854));
   INV_X1 i_257_76_16885 (.A(n_257_76_16854), .ZN(n_257_76_16855));
   NAND2_X1 i_257_76_16886 (.A1(n_257_76_16846), .A2(n_257_76_16855), .ZN(
      n_257_76_16856));
   INV_X1 i_257_76_16887 (.A(n_257_76_16856), .ZN(n_257_76_16857));
   NAND2_X1 i_257_76_16888 (.A1(n_257_76_16845), .A2(n_257_76_16857), .ZN(
      n_257_76_16858));
   INV_X1 i_257_76_16889 (.A(n_257_76_16858), .ZN(n_257_76_16859));
   NAND2_X1 i_257_76_16890 (.A1(n_257_17), .A2(n_257_76_16859), .ZN(
      n_257_76_16860));
   NAND2_X1 i_257_76_16891 (.A1(n_257_443), .A2(n_257_76_16848), .ZN(
      n_257_76_16861));
   INV_X1 i_257_76_16892 (.A(n_257_76_16861), .ZN(n_257_76_16862));
   NAND2_X1 i_257_76_16893 (.A1(n_257_1057), .A2(n_257_76_16862), .ZN(
      n_257_76_16863));
   INV_X1 i_257_76_16894 (.A(n_257_76_16863), .ZN(n_257_76_16864));
   NAND2_X1 i_257_76_16895 (.A1(n_257_76_18072), .A2(n_257_76_16864), .ZN(
      n_257_76_16865));
   NAND2_X1 i_257_76_16896 (.A1(n_257_699), .A2(n_257_448), .ZN(n_257_76_16866));
   NAND2_X1 i_257_76_16897 (.A1(n_257_446), .A2(n_257_859), .ZN(n_257_76_16867));
   NAND2_X1 i_257_76_16898 (.A1(n_257_449), .A2(n_257_667), .ZN(n_257_76_16868));
   NAND2_X1 i_257_76_16899 (.A1(n_257_763), .A2(n_257_436), .ZN(n_257_76_16869));
   NAND3_X1 i_257_76_16900 (.A1(n_257_76_16867), .A2(n_257_76_16868), .A3(
      n_257_76_16869), .ZN(n_257_76_16870));
   INV_X1 i_257_76_16901 (.A(n_257_76_16847), .ZN(n_257_76_16871));
   NOR2_X1 i_257_76_16902 (.A1(n_257_76_16870), .A2(n_257_76_16871), .ZN(
      n_257_76_16872));
   NAND2_X1 i_257_76_16903 (.A1(n_257_447), .A2(n_257_795), .ZN(n_257_76_16873));
   NAND2_X1 i_257_76_16904 (.A1(n_257_929), .A2(n_257_439), .ZN(n_257_76_16874));
   NAND2_X1 i_257_76_16905 (.A1(n_257_827), .A2(n_257_437), .ZN(n_257_76_16875));
   NAND3_X1 i_257_76_16906 (.A1(n_257_76_16873), .A2(n_257_76_16874), .A3(
      n_257_76_16875), .ZN(n_257_76_16876));
   NAND2_X1 i_257_76_16907 (.A1(n_257_731), .A2(n_257_435), .ZN(n_257_76_16877));
   NAND2_X1 i_257_76_16908 (.A1(n_257_450), .A2(n_257_76_16848), .ZN(
      n_257_76_16878));
   INV_X1 i_257_76_16909 (.A(n_257_76_16878), .ZN(n_257_76_16879));
   NAND3_X1 i_257_76_16910 (.A1(n_257_659), .A2(n_257_76_16877), .A3(
      n_257_76_16879), .ZN(n_257_76_16880));
   INV_X1 i_257_76_16911 (.A(n_257_76_16880), .ZN(n_257_76_16881));
   NAND2_X1 i_257_76_16912 (.A1(n_257_891), .A2(n_257_445), .ZN(n_257_76_16882));
   NAND2_X1 i_257_76_16913 (.A1(n_257_440), .A2(n_257_961), .ZN(n_257_76_16883));
   NAND2_X1 i_257_76_16914 (.A1(n_257_438), .A2(n_257_897), .ZN(n_257_76_16884));
   NAND4_X1 i_257_76_16915 (.A1(n_257_76_16881), .A2(n_257_76_16882), .A3(
      n_257_76_16883), .A4(n_257_76_16884), .ZN(n_257_76_16885));
   NOR2_X1 i_257_76_16916 (.A1(n_257_76_16876), .A2(n_257_76_16885), .ZN(
      n_257_76_16886));
   NAND4_X1 i_257_76_16917 (.A1(n_257_76_16866), .A2(n_257_76_16872), .A3(
      n_257_76_16886), .A4(n_257_76_16846), .ZN(n_257_76_16887));
   INV_X1 i_257_76_16918 (.A(n_257_76_16845), .ZN(n_257_76_16888));
   NOR2_X1 i_257_76_16919 (.A1(n_257_76_16887), .A2(n_257_76_16888), .ZN(
      n_257_76_16889));
   NAND2_X1 i_257_76_16920 (.A1(n_257_28), .A2(n_257_76_16889), .ZN(
      n_257_76_16890));
   NAND3_X1 i_257_76_16921 (.A1(n_257_76_16860), .A2(n_257_76_16865), .A3(
      n_257_76_16890), .ZN(n_257_76_16891));
   INV_X1 i_257_76_16922 (.A(n_257_859), .ZN(n_257_76_16892));
   NOR2_X1 i_257_76_16923 (.A1(n_257_76_16849), .A2(n_257_76_16892), .ZN(
      n_257_76_16893));
   NAND4_X1 i_257_76_16924 (.A1(n_257_446), .A2(n_257_76_16883), .A3(
      n_257_76_16884), .A4(n_257_76_16893), .ZN(n_257_76_16894));
   INV_X1 i_257_76_16925 (.A(n_257_76_16894), .ZN(n_257_76_16895));
   NAND2_X1 i_257_76_16926 (.A1(n_257_76_16874), .A2(n_257_76_16882), .ZN(
      n_257_76_16896));
   INV_X1 i_257_76_16927 (.A(n_257_76_16896), .ZN(n_257_76_16897));
   NAND3_X1 i_257_76_16928 (.A1(n_257_76_16895), .A2(n_257_76_16897), .A3(
      n_257_76_16847), .ZN(n_257_76_16898));
   INV_X1 i_257_76_16929 (.A(n_257_76_16898), .ZN(n_257_76_16899));
   NAND2_X1 i_257_76_16930 (.A1(n_257_76_16899), .A2(n_257_76_16846), .ZN(
      n_257_76_16900));
   NOR2_X1 i_257_76_16931 (.A1(n_257_76_16888), .A2(n_257_76_16900), .ZN(
      n_257_76_16901));
   NAND2_X1 i_257_76_16932 (.A1(n_257_76_18070), .A2(n_257_76_16901), .ZN(
      n_257_76_16902));
   NAND2_X1 i_257_76_16933 (.A1(n_257_439), .A2(n_257_76_16848), .ZN(
      n_257_76_16903));
   INV_X1 i_257_76_16934 (.A(n_257_76_16903), .ZN(n_257_76_16904));
   NAND3_X1 i_257_76_16935 (.A1(n_257_76_16904), .A2(n_257_929), .A3(
      n_257_76_16883), .ZN(n_257_76_16905));
   INV_X1 i_257_76_16936 (.A(n_257_76_16905), .ZN(n_257_76_16906));
   NAND2_X1 i_257_76_16937 (.A1(n_257_76_16847), .A2(n_257_76_16906), .ZN(
      n_257_76_16907));
   INV_X1 i_257_76_16938 (.A(n_257_76_16907), .ZN(n_257_76_16908));
   NAND2_X1 i_257_76_16939 (.A1(n_257_76_16846), .A2(n_257_76_16908), .ZN(
      n_257_76_16909));
   INV_X1 i_257_76_16940 (.A(n_257_76_16909), .ZN(n_257_76_16910));
   NAND2_X1 i_257_76_16941 (.A1(n_257_76_16845), .A2(n_257_76_16910), .ZN(
      n_257_76_16911));
   INV_X1 i_257_76_16942 (.A(n_257_76_16911), .ZN(n_257_76_16912));
   NAND2_X1 i_257_76_16943 (.A1(n_257_76_18084), .A2(n_257_76_16912), .ZN(
      n_257_76_16913));
   NAND2_X1 i_257_76_16944 (.A1(n_257_182), .A2(n_257_429), .ZN(n_257_76_16914));
   NAND2_X1 i_257_76_16945 (.A1(n_257_262), .A2(n_257_425), .ZN(n_257_76_16915));
   NAND2_X1 i_257_76_16946 (.A1(n_257_65), .A2(n_257_433), .ZN(n_257_76_16916));
   NAND2_X1 i_257_76_16947 (.A1(n_257_531), .A2(n_257_424), .ZN(n_257_76_16917));
   NAND3_X1 i_257_76_16948 (.A1(n_257_76_16916), .A2(n_257_302), .A3(
      n_257_76_16917), .ZN(n_257_76_16918));
   INV_X1 i_257_76_16949 (.A(n_257_76_16918), .ZN(n_257_76_16919));
   NAND2_X1 i_257_76_16950 (.A1(n_257_659), .A2(n_257_450), .ZN(n_257_76_16920));
   NAND2_X1 i_257_76_16951 (.A1(n_257_432), .A2(n_257_627), .ZN(n_257_76_16921));
   INV_X1 i_257_76_16952 (.A(n_257_595), .ZN(n_257_76_16922));
   NAND2_X1 i_257_76_16953 (.A1(n_257_76_16922), .A2(n_257_442), .ZN(
      n_257_76_16923));
   OAI21_X1 i_257_76_16954 (.A(n_257_76_16923), .B1(n_257_428), .B2(
      n_257_76_17412), .ZN(n_257_76_16924));
   INV_X1 i_257_76_16955 (.A(n_257_1089), .ZN(n_257_76_16925));
   NAND2_X1 i_257_76_16956 (.A1(n_257_76_16925), .A2(n_257_423), .ZN(
      n_257_76_16926));
   INV_X1 i_257_76_16957 (.A(n_257_76_16926), .ZN(n_257_76_16927));
   NAND4_X1 i_257_76_16958 (.A1(n_257_76_16877), .A2(n_257_76_16921), .A3(
      n_257_76_16924), .A4(n_257_76_16927), .ZN(n_257_76_16928));
   INV_X1 i_257_76_16959 (.A(n_257_76_16928), .ZN(n_257_76_16929));
   NAND3_X1 i_257_76_16960 (.A1(n_257_76_16919), .A2(n_257_76_16920), .A3(
      n_257_76_16929), .ZN(n_257_76_16930));
   INV_X1 i_257_76_16961 (.A(n_257_76_16930), .ZN(n_257_76_16931));
   NAND4_X1 i_257_76_16962 (.A1(n_257_76_16914), .A2(n_257_76_16915), .A3(
      n_257_76_16931), .A4(n_257_76_16847), .ZN(n_257_76_16932));
   INV_X1 i_257_76_16963 (.A(n_257_76_16846), .ZN(n_257_76_16933));
   NOR2_X1 i_257_76_16964 (.A1(n_257_76_16932), .A2(n_257_76_16933), .ZN(
      n_257_76_16934));
   NAND2_X1 i_257_76_16965 (.A1(n_257_563), .A2(n_257_426), .ZN(n_257_76_16935));
   NAND2_X1 i_257_76_16966 (.A1(n_257_143), .A2(n_257_430), .ZN(n_257_76_16936));
   NAND3_X1 i_257_76_16967 (.A1(n_257_76_16875), .A2(n_257_76_16935), .A3(
      n_257_76_16936), .ZN(n_257_76_16937));
   NAND2_X1 i_257_76_16968 (.A1(n_257_427), .A2(n_257_222), .ZN(n_257_76_16938));
   NAND4_X1 i_257_76_16969 (.A1(n_257_76_16882), .A2(n_257_76_16883), .A3(
      n_257_76_16884), .A4(n_257_76_16938), .ZN(n_257_76_16939));
   NOR2_X1 i_257_76_16970 (.A1(n_257_76_16937), .A2(n_257_76_16939), .ZN(
      n_257_76_16940));
   NAND2_X1 i_257_76_16971 (.A1(n_257_105), .A2(n_257_431), .ZN(n_257_76_16941));
   NAND3_X1 i_257_76_16972 (.A1(n_257_76_16941), .A2(n_257_76_16867), .A3(
      n_257_76_16868), .ZN(n_257_76_16942));
   INV_X1 i_257_76_16973 (.A(n_257_76_16942), .ZN(n_257_76_16943));
   NAND2_X1 i_257_76_16974 (.A1(n_257_451), .A2(n_257_482), .ZN(n_257_76_16944));
   NAND4_X1 i_257_76_16975 (.A1(n_257_76_16869), .A2(n_257_76_16873), .A3(
      n_257_76_16944), .A4(n_257_76_16874), .ZN(n_257_76_16945));
   INV_X1 i_257_76_16976 (.A(n_257_76_16945), .ZN(n_257_76_16946));
   NAND3_X1 i_257_76_16977 (.A1(n_257_76_16940), .A2(n_257_76_16943), .A3(
      n_257_76_16946), .ZN(n_257_76_16947));
   INV_X1 i_257_76_16978 (.A(n_257_76_16947), .ZN(n_257_76_16948));
   NAND4_X1 i_257_76_16979 (.A1(n_257_76_16934), .A2(n_257_76_16948), .A3(
      n_257_76_16845), .A4(n_257_76_16866), .ZN(n_257_76_16949));
   INV_X1 i_257_76_16980 (.A(n_257_76_16949), .ZN(n_257_76_16950));
   NAND2_X1 i_257_76_16981 (.A1(n_257_76_18066), .A2(n_257_76_16950), .ZN(
      n_257_76_16951));
   NAND3_X1 i_257_76_16982 (.A1(n_257_76_16902), .A2(n_257_76_16913), .A3(
      n_257_76_16951), .ZN(n_257_76_16952));
   NOR2_X1 i_257_76_16983 (.A1(n_257_76_16891), .A2(n_257_76_16952), .ZN(
      n_257_76_16953));
   NAND2_X1 i_257_76_16984 (.A1(n_257_993), .A2(n_257_76_16848), .ZN(
      n_257_76_16954));
   INV_X1 i_257_76_16985 (.A(n_257_76_16954), .ZN(n_257_76_16955));
   NAND2_X1 i_257_76_16986 (.A1(n_257_441), .A2(n_257_76_16955), .ZN(
      n_257_76_16956));
   INV_X1 i_257_76_16987 (.A(n_257_76_16956), .ZN(n_257_76_16957));
   NAND2_X1 i_257_76_16988 (.A1(n_257_76_16846), .A2(n_257_76_16957), .ZN(
      n_257_76_16958));
   INV_X1 i_257_76_16989 (.A(n_257_76_16958), .ZN(n_257_76_16959));
   NAND2_X1 i_257_76_16990 (.A1(n_257_76_16845), .A2(n_257_76_16959), .ZN(
      n_257_76_16960));
   INV_X1 i_257_76_16991 (.A(n_257_76_16960), .ZN(n_257_76_16961));
   NAND2_X1 i_257_76_16992 (.A1(n_257_76_18071), .A2(n_257_76_16961), .ZN(
      n_257_76_16962));
   NAND3_X1 i_257_76_16993 (.A1(n_257_76_16848), .A2(n_257_731), .A3(n_257_435), 
      .ZN(n_257_76_16963));
   INV_X1 i_257_76_16994 (.A(n_257_76_16963), .ZN(n_257_76_16964));
   NAND4_X1 i_257_76_16995 (.A1(n_257_76_16882), .A2(n_257_76_16883), .A3(
      n_257_76_16884), .A4(n_257_76_16964), .ZN(n_257_76_16965));
   NOR2_X1 i_257_76_16996 (.A1(n_257_76_16876), .A2(n_257_76_16965), .ZN(
      n_257_76_16966));
   NAND2_X1 i_257_76_16997 (.A1(n_257_76_16867), .A2(n_257_76_16869), .ZN(
      n_257_76_16967));
   NOR2_X1 i_257_76_16998 (.A1(n_257_76_16871), .A2(n_257_76_16967), .ZN(
      n_257_76_16968));
   NAND3_X1 i_257_76_16999 (.A1(n_257_76_16846), .A2(n_257_76_16966), .A3(
      n_257_76_16968), .ZN(n_257_76_16969));
   NOR2_X1 i_257_76_17000 (.A1(n_257_76_16969), .A2(n_257_76_16888), .ZN(
      n_257_76_16970));
   NAND2_X1 i_257_76_17001 (.A1(n_257_76_18078), .A2(n_257_76_16970), .ZN(
      n_257_76_16971));
   NAND3_X1 i_257_76_17002 (.A1(n_257_76_16914), .A2(n_257_76_16847), .A3(
      n_257_76_16941), .ZN(n_257_76_16972));
   INV_X1 i_257_76_17003 (.A(n_257_76_16972), .ZN(n_257_76_16973));
   NAND3_X1 i_257_76_17004 (.A1(n_257_76_16873), .A2(n_257_76_16944), .A3(
      n_257_76_16874), .ZN(n_257_76_16974));
   NOR2_X1 i_257_76_17005 (.A1(n_257_76_16870), .A2(n_257_76_16974), .ZN(
      n_257_76_16975));
   NAND2_X1 i_257_76_17006 (.A1(n_257_595), .A2(n_257_442), .ZN(n_257_76_16976));
   INV_X1 i_257_76_17007 (.A(n_257_76_16976), .ZN(n_257_76_16977));
   NAND3_X1 i_257_76_17008 (.A1(n_257_76_16925), .A2(n_257_428), .A3(
      n_257_76_16977), .ZN(n_257_76_16978));
   INV_X1 i_257_76_17009 (.A(n_257_76_16978), .ZN(n_257_76_16979));
   NAND3_X1 i_257_76_17010 (.A1(n_257_76_16877), .A2(n_257_76_16921), .A3(
      n_257_76_16979), .ZN(n_257_76_16980));
   INV_X1 i_257_76_17011 (.A(n_257_76_16916), .ZN(n_257_76_16981));
   NOR2_X1 i_257_76_17012 (.A1(n_257_76_16980), .A2(n_257_76_16981), .ZN(
      n_257_76_16982));
   NAND4_X1 i_257_76_17013 (.A1(n_257_76_16982), .A2(n_257_76_16883), .A3(
      n_257_76_16884), .A4(n_257_76_16920), .ZN(n_257_76_16983));
   NAND3_X1 i_257_76_17014 (.A1(n_257_76_16875), .A2(n_257_76_16936), .A3(
      n_257_76_16882), .ZN(n_257_76_16984));
   NOR2_X1 i_257_76_17015 (.A1(n_257_76_16983), .A2(n_257_76_16984), .ZN(
      n_257_76_16985));
   NAND4_X1 i_257_76_17016 (.A1(n_257_76_16973), .A2(n_257_76_16975), .A3(
      n_257_76_16985), .A4(n_257_76_16846), .ZN(n_257_76_16986));
   NAND2_X1 i_257_76_17017 (.A1(n_257_76_16845), .A2(n_257_76_16866), .ZN(
      n_257_76_16987));
   NOR2_X1 i_257_76_17018 (.A1(n_257_76_16986), .A2(n_257_76_16987), .ZN(
      n_257_76_16988));
   NAND2_X1 i_257_76_17019 (.A1(n_257_76_18074), .A2(n_257_76_16988), .ZN(
      n_257_76_16989));
   NAND3_X1 i_257_76_17020 (.A1(n_257_76_16962), .A2(n_257_76_16971), .A3(
      n_257_76_16989), .ZN(n_257_76_16990));
   NAND2_X1 i_257_76_17021 (.A1(n_257_1089), .A2(n_257_442), .ZN(n_257_76_16991));
   INV_X1 i_257_76_17022 (.A(n_257_76_16991), .ZN(n_257_76_16992));
   NAND2_X1 i_257_76_17023 (.A1(n_257_13), .A2(n_257_76_16992), .ZN(
      n_257_76_16993));
   NAND2_X1 i_257_76_17024 (.A1(n_257_445), .A2(n_257_76_16848), .ZN(
      n_257_76_16994));
   INV_X1 i_257_76_17025 (.A(n_257_76_16994), .ZN(n_257_76_16995));
   NAND4_X1 i_257_76_17026 (.A1(n_257_76_16883), .A2(n_257_76_16884), .A3(
      n_257_891), .A4(n_257_76_16995), .ZN(n_257_76_16996));
   INV_X1 i_257_76_17027 (.A(n_257_76_16996), .ZN(n_257_76_16997));
   NAND3_X1 i_257_76_17028 (.A1(n_257_76_16997), .A2(n_257_76_16847), .A3(
      n_257_76_16874), .ZN(n_257_76_16998));
   INV_X1 i_257_76_17029 (.A(n_257_76_16998), .ZN(n_257_76_16999));
   NAND2_X1 i_257_76_17030 (.A1(n_257_76_16999), .A2(n_257_76_16846), .ZN(
      n_257_76_17000));
   NOR2_X1 i_257_76_17031 (.A1(n_257_76_16888), .A2(n_257_76_17000), .ZN(
      n_257_76_17001));
   NAND2_X1 i_257_76_17032 (.A1(n_257_76_18077), .A2(n_257_76_17001), .ZN(
      n_257_76_17002));
   NAND2_X1 i_257_76_17033 (.A1(n_257_76_16993), .A2(n_257_76_17002), .ZN(
      n_257_76_17003));
   NOR2_X1 i_257_76_17034 (.A1(n_257_76_16990), .A2(n_257_76_17003), .ZN(
      n_257_76_17004));
   NOR2_X1 i_257_76_17035 (.A1(n_257_76_17564), .A2(n_257_1089), .ZN(
      n_257_76_17005));
   NAND4_X1 i_257_76_17036 (.A1(n_257_76_16877), .A2(n_257_76_16921), .A3(
      n_257_76_16924), .A4(n_257_76_17005), .ZN(n_257_76_17006));
   INV_X1 i_257_76_17037 (.A(n_257_76_17006), .ZN(n_257_76_17007));
   NAND4_X1 i_257_76_17038 (.A1(n_257_76_17007), .A2(n_257_563), .A3(
      n_257_76_16938), .A4(n_257_76_16916), .ZN(n_257_76_17008));
   NAND3_X1 i_257_76_17039 (.A1(n_257_76_16883), .A2(n_257_76_16884), .A3(
      n_257_76_16920), .ZN(n_257_76_17009));
   NOR2_X1 i_257_76_17040 (.A1(n_257_76_17008), .A2(n_257_76_17009), .ZN(
      n_257_76_17010));
   NAND2_X1 i_257_76_17041 (.A1(n_257_76_16869), .A2(n_257_76_16874), .ZN(
      n_257_76_17011));
   INV_X1 i_257_76_17042 (.A(n_257_76_17011), .ZN(n_257_76_17012));
   INV_X1 i_257_76_17043 (.A(n_257_76_16984), .ZN(n_257_76_17013));
   NAND4_X1 i_257_76_17044 (.A1(n_257_76_17010), .A2(n_257_76_17012), .A3(
      n_257_76_16941), .A4(n_257_76_17013), .ZN(n_257_76_17014));
   INV_X1 i_257_76_17045 (.A(n_257_76_17014), .ZN(n_257_76_17015));
   NAND2_X1 i_257_76_17046 (.A1(n_257_76_16845), .A2(n_257_76_17015), .ZN(
      n_257_76_17016));
   NAND2_X1 i_257_76_17047 (.A1(n_257_76_16914), .A2(n_257_76_16847), .ZN(
      n_257_76_17017));
   INV_X1 i_257_76_17048 (.A(n_257_76_17017), .ZN(n_257_76_17018));
   NAND4_X1 i_257_76_17049 (.A1(n_257_76_16867), .A2(n_257_76_16868), .A3(
      n_257_76_16873), .A4(n_257_76_16944), .ZN(n_257_76_17019));
   INV_X1 i_257_76_17050 (.A(n_257_76_17019), .ZN(n_257_76_17020));
   NAND4_X1 i_257_76_17051 (.A1(n_257_76_16866), .A2(n_257_76_17018), .A3(
      n_257_76_16846), .A4(n_257_76_17020), .ZN(n_257_76_17021));
   NOR2_X1 i_257_76_17052 (.A1(n_257_76_17016), .A2(n_257_76_17021), .ZN(
      n_257_76_17022));
   NAND2_X1 i_257_76_17053 (.A1(n_257_76_18076), .A2(n_257_76_17022), .ZN(
      n_257_76_17023));
   NAND2_X1 i_257_76_17054 (.A1(n_257_76_16867), .A2(n_257_76_16873), .ZN(
      n_257_76_17024));
   NOR2_X1 i_257_76_17055 (.A1(n_257_76_16871), .A2(n_257_76_17024), .ZN(
      n_257_76_17025));
   NAND3_X1 i_257_76_17056 (.A1(n_257_76_16874), .A2(n_257_76_16875), .A3(
      n_257_76_16882), .ZN(n_257_76_17026));
   NAND2_X1 i_257_76_17057 (.A1(n_257_436), .A2(n_257_76_16848), .ZN(
      n_257_76_17027));
   INV_X1 i_257_76_17058 (.A(n_257_76_17027), .ZN(n_257_76_17028));
   NAND4_X1 i_257_76_17059 (.A1(n_257_763), .A2(n_257_76_16883), .A3(
      n_257_76_16884), .A4(n_257_76_17028), .ZN(n_257_76_17029));
   NOR2_X1 i_257_76_17060 (.A1(n_257_76_17026), .A2(n_257_76_17029), .ZN(
      n_257_76_17030));
   NAND3_X1 i_257_76_17061 (.A1(n_257_76_16846), .A2(n_257_76_17025), .A3(
      n_257_76_17030), .ZN(n_257_76_17031));
   NOR2_X1 i_257_76_17062 (.A1(n_257_76_17031), .A2(n_257_76_16888), .ZN(
      n_257_76_17032));
   NAND2_X1 i_257_76_17063 (.A1(n_257_76_18069), .A2(n_257_76_17032), .ZN(
      n_257_76_17033));
   INV_X1 i_257_76_17064 (.A(n_257_76_17026), .ZN(n_257_76_17034));
   NAND2_X1 i_257_76_17065 (.A1(n_257_76_16873), .A2(n_257_76_16944), .ZN(
      n_257_76_17035));
   INV_X1 i_257_76_17066 (.A(n_257_76_17035), .ZN(n_257_76_17036));
   NAND2_X1 i_257_76_17067 (.A1(n_257_442), .A2(n_257_627), .ZN(n_257_76_17037));
   NOR2_X1 i_257_76_17068 (.A1(n_257_1089), .A2(n_257_76_17037), .ZN(
      n_257_76_17038));
   NAND2_X1 i_257_76_17069 (.A1(n_257_432), .A2(n_257_76_17038), .ZN(
      n_257_76_17039));
   INV_X1 i_257_76_17070 (.A(n_257_76_17039), .ZN(n_257_76_17040));
   NAND3_X1 i_257_76_17071 (.A1(n_257_76_16916), .A2(n_257_76_16877), .A3(
      n_257_76_17040), .ZN(n_257_76_17041));
   INV_X1 i_257_76_17072 (.A(n_257_76_17041), .ZN(n_257_76_17042));
   NAND4_X1 i_257_76_17073 (.A1(n_257_76_17042), .A2(n_257_76_16883), .A3(
      n_257_76_16884), .A4(n_257_76_16920), .ZN(n_257_76_17043));
   INV_X1 i_257_76_17074 (.A(n_257_76_17043), .ZN(n_257_76_17044));
   NAND3_X1 i_257_76_17075 (.A1(n_257_76_17034), .A2(n_257_76_17036), .A3(
      n_257_76_17044), .ZN(n_257_76_17045));
   NAND4_X1 i_257_76_17076 (.A1(n_257_76_16847), .A2(n_257_76_16867), .A3(
      n_257_76_16868), .A4(n_257_76_16869), .ZN(n_257_76_17046));
   NOR2_X1 i_257_76_17077 (.A1(n_257_76_17045), .A2(n_257_76_17046), .ZN(
      n_257_76_17047));
   NAND2_X1 i_257_76_17078 (.A1(n_257_76_16866), .A2(n_257_76_16846), .ZN(
      n_257_76_17048));
   INV_X1 i_257_76_17079 (.A(n_257_76_17048), .ZN(n_257_76_17049));
   NAND3_X1 i_257_76_17080 (.A1(n_257_76_17047), .A2(n_257_76_17049), .A3(
      n_257_76_16845), .ZN(n_257_76_17050));
   INV_X1 i_257_76_17081 (.A(n_257_76_17050), .ZN(n_257_76_17051));
   NAND2_X1 i_257_76_17082 (.A1(n_257_68), .A2(n_257_76_17051), .ZN(
      n_257_76_17052));
   NAND3_X1 i_257_76_17083 (.A1(n_257_76_17023), .A2(n_257_76_17033), .A3(
      n_257_76_17052), .ZN(n_257_76_17053));
   NAND2_X1 i_257_76_17084 (.A1(n_257_437), .A2(n_257_76_16848), .ZN(
      n_257_76_17054));
   INV_X1 i_257_76_17085 (.A(n_257_76_17054), .ZN(n_257_76_17055));
   NAND4_X1 i_257_76_17086 (.A1(n_257_76_16883), .A2(n_257_76_16884), .A3(
      n_257_827), .A4(n_257_76_17055), .ZN(n_257_76_17056));
   NOR2_X1 i_257_76_17087 (.A1(n_257_76_16896), .A2(n_257_76_17056), .ZN(
      n_257_76_17057));
   NAND2_X1 i_257_76_17088 (.A1(n_257_76_16847), .A2(n_257_76_16867), .ZN(
      n_257_76_17058));
   INV_X1 i_257_76_17089 (.A(n_257_76_17058), .ZN(n_257_76_17059));
   NAND3_X1 i_257_76_17090 (.A1(n_257_76_17057), .A2(n_257_76_16846), .A3(
      n_257_76_17059), .ZN(n_257_76_17060));
   NOR2_X1 i_257_76_17091 (.A1(n_257_76_16888), .A2(n_257_76_17060), .ZN(
      n_257_76_17061));
   NAND2_X1 i_257_76_17092 (.A1(n_257_22), .A2(n_257_76_17061), .ZN(
      n_257_76_17062));
   NAND2_X1 i_257_76_17093 (.A1(n_257_444), .A2(n_257_76_16848), .ZN(
      n_257_76_17063));
   INV_X1 i_257_76_17094 (.A(n_257_76_17063), .ZN(n_257_76_17064));
   NAND2_X1 i_257_76_17095 (.A1(n_257_1025), .A2(n_257_76_17064), .ZN(
      n_257_76_17065));
   INV_X1 i_257_76_17096 (.A(n_257_76_17065), .ZN(n_257_76_17066));
   NAND2_X1 i_257_76_17097 (.A1(n_257_76_16845), .A2(n_257_76_17066), .ZN(
      n_257_76_17067));
   INV_X1 i_257_76_17098 (.A(n_257_76_17067), .ZN(n_257_76_17068));
   NAND2_X1 i_257_76_17099 (.A1(n_257_76_18075), .A2(n_257_76_17068), .ZN(
      n_257_76_17069));
   NAND2_X1 i_257_76_17100 (.A1(n_257_76_17062), .A2(n_257_76_17069), .ZN(
      n_257_76_17070));
   NOR2_X1 i_257_76_17101 (.A1(n_257_76_17053), .A2(n_257_76_17070), .ZN(
      n_257_76_17071));
   NAND3_X1 i_257_76_17102 (.A1(n_257_76_16953), .A2(n_257_76_17004), .A3(
      n_257_76_17071), .ZN(n_257_76_17072));
   INV_X1 i_257_76_17103 (.A(n_257_76_17072), .ZN(n_257_76_17073));
   INV_X1 i_257_76_17104 (.A(n_257_433), .ZN(n_257_76_17074));
   NOR2_X1 i_257_76_17105 (.A1(n_257_76_16849), .A2(n_257_76_17074), .ZN(
      n_257_76_17075));
   NAND3_X1 i_257_76_17106 (.A1(n_257_76_17075), .A2(n_257_76_16877), .A3(
      n_257_65), .ZN(n_257_76_17076));
   INV_X1 i_257_76_17107 (.A(n_257_76_17076), .ZN(n_257_76_17077));
   NAND3_X1 i_257_76_17108 (.A1(n_257_76_17077), .A2(n_257_76_16884), .A3(
      n_257_76_16920), .ZN(n_257_76_17078));
   NAND2_X1 i_257_76_17109 (.A1(n_257_76_16882), .A2(n_257_76_16883), .ZN(
      n_257_76_17079));
   NOR2_X1 i_257_76_17110 (.A1(n_257_76_17078), .A2(n_257_76_17079), .ZN(
      n_257_76_17080));
   NAND2_X1 i_257_76_17111 (.A1(n_257_76_16874), .A2(n_257_76_16875), .ZN(
      n_257_76_17081));
   INV_X1 i_257_76_17112 (.A(n_257_76_17081), .ZN(n_257_76_17082));
   NAND3_X1 i_257_76_17113 (.A1(n_257_76_17080), .A2(n_257_76_17036), .A3(
      n_257_76_17082), .ZN(n_257_76_17083));
   NOR2_X1 i_257_76_17114 (.A1(n_257_76_17083), .A2(n_257_76_17046), .ZN(
      n_257_76_17084));
   NAND3_X1 i_257_76_17115 (.A1(n_257_76_17084), .A2(n_257_76_17049), .A3(
      n_257_76_16845), .ZN(n_257_76_17085));
   INV_X1 i_257_76_17116 (.A(n_257_76_17085), .ZN(n_257_76_17086));
   NAND2_X1 i_257_76_17117 (.A1(n_257_76_18081), .A2(n_257_76_17086), .ZN(
      n_257_76_17087));
   NAND3_X1 i_257_76_17118 (.A1(n_257_76_16867), .A2(n_257_76_16869), .A3(
      n_257_76_16873), .ZN(n_257_76_17088));
   NOR2_X1 i_257_76_17119 (.A1(n_257_76_17088), .A2(n_257_76_16871), .ZN(
      n_257_76_17089));
   NAND2_X1 i_257_76_17120 (.A1(n_257_442), .A2(n_257_667), .ZN(n_257_76_17090));
   NOR2_X1 i_257_76_17121 (.A1(n_257_1089), .A2(n_257_76_17090), .ZN(
      n_257_76_17091));
   NAND2_X1 i_257_76_17122 (.A1(n_257_76_16877), .A2(n_257_76_17091), .ZN(
      n_257_76_17092));
   INV_X1 i_257_76_17123 (.A(n_257_76_17092), .ZN(n_257_76_17093));
   NAND4_X1 i_257_76_17124 (.A1(n_257_449), .A2(n_257_76_16883), .A3(
      n_257_76_16884), .A4(n_257_76_17093), .ZN(n_257_76_17094));
   NOR2_X1 i_257_76_17125 (.A1(n_257_76_17026), .A2(n_257_76_17094), .ZN(
      n_257_76_17095));
   NAND4_X1 i_257_76_17126 (.A1(n_257_76_17089), .A2(n_257_76_16866), .A3(
      n_257_76_17095), .A4(n_257_76_16846), .ZN(n_257_76_17096));
   NOR2_X1 i_257_76_17127 (.A1(n_257_76_17096), .A2(n_257_76_16888), .ZN(
      n_257_76_17097));
   NAND2_X1 i_257_76_17128 (.A1(n_257_76_18083), .A2(n_257_76_17097), .ZN(
      n_257_76_17098));
   NAND4_X1 i_257_76_17129 (.A1(n_257_76_16847), .A2(n_257_76_16941), .A3(
      n_257_182), .A4(n_257_76_16867), .ZN(n_257_76_17099));
   NOR2_X1 i_257_76_17130 (.A1(n_257_76_16933), .A2(n_257_76_17099), .ZN(
      n_257_76_17100));
   INV_X1 i_257_76_17131 (.A(n_257_429), .ZN(n_257_76_17101));
   NOR2_X1 i_257_76_17132 (.A1(n_257_76_16849), .A2(n_257_76_17101), .ZN(
      n_257_76_17102));
   NAND3_X1 i_257_76_17133 (.A1(n_257_76_17102), .A2(n_257_76_16877), .A3(
      n_257_76_16921), .ZN(n_257_76_17103));
   INV_X1 i_257_76_17134 (.A(n_257_76_17103), .ZN(n_257_76_17104));
   NAND4_X1 i_257_76_17135 (.A1(n_257_76_17104), .A2(n_257_76_16884), .A3(
      n_257_76_16920), .A4(n_257_76_16916), .ZN(n_257_76_17105));
   NAND3_X1 i_257_76_17136 (.A1(n_257_76_16936), .A2(n_257_76_16882), .A3(
      n_257_76_16883), .ZN(n_257_76_17106));
   NOR2_X1 i_257_76_17137 (.A1(n_257_76_17105), .A2(n_257_76_17106), .ZN(
      n_257_76_17107));
   NAND3_X1 i_257_76_17138 (.A1(n_257_76_16868), .A2(n_257_76_16869), .A3(
      n_257_76_16873), .ZN(n_257_76_17108));
   INV_X1 i_257_76_17139 (.A(n_257_76_17108), .ZN(n_257_76_17109));
   NAND3_X1 i_257_76_17140 (.A1(n_257_76_16944), .A2(n_257_76_16874), .A3(
      n_257_76_16875), .ZN(n_257_76_17110));
   INV_X1 i_257_76_17141 (.A(n_257_76_17110), .ZN(n_257_76_17111));
   NAND3_X1 i_257_76_17142 (.A1(n_257_76_17107), .A2(n_257_76_17109), .A3(
      n_257_76_17111), .ZN(n_257_76_17112));
   INV_X1 i_257_76_17143 (.A(n_257_76_17112), .ZN(n_257_76_17113));
   NAND4_X1 i_257_76_17144 (.A1(n_257_76_17100), .A2(n_257_76_16845), .A3(
      n_257_76_17113), .A4(n_257_76_16866), .ZN(n_257_76_17114));
   INV_X1 i_257_76_17145 (.A(n_257_76_17114), .ZN(n_257_76_17115));
   NAND2_X1 i_257_76_17146 (.A1(n_257_76_18061), .A2(n_257_76_17115), .ZN(
      n_257_76_17116));
   NAND3_X1 i_257_76_17147 (.A1(n_257_76_17087), .A2(n_257_76_17098), .A3(
      n_257_76_17116), .ZN(n_257_76_17117));
   INV_X1 i_257_76_17148 (.A(n_257_76_17117), .ZN(n_257_76_17118));
   NAND2_X1 i_257_76_17149 (.A1(n_257_442), .A2(n_257_897), .ZN(n_257_76_17119));
   NOR2_X1 i_257_76_17150 (.A1(n_257_1089), .A2(n_257_76_17119), .ZN(
      n_257_76_17120));
   NAND2_X1 i_257_76_17151 (.A1(n_257_438), .A2(n_257_76_17120), .ZN(
      n_257_76_17121));
   INV_X1 i_257_76_17152 (.A(n_257_76_17121), .ZN(n_257_76_17122));
   NAND3_X1 i_257_76_17153 (.A1(n_257_76_16874), .A2(n_257_76_16883), .A3(
      n_257_76_17122), .ZN(n_257_76_17123));
   INV_X1 i_257_76_17154 (.A(n_257_76_17123), .ZN(n_257_76_17124));
   NAND2_X1 i_257_76_17155 (.A1(n_257_76_17124), .A2(n_257_76_16847), .ZN(
      n_257_76_17125));
   NOR2_X1 i_257_76_17156 (.A1(n_257_76_16933), .A2(n_257_76_17125), .ZN(
      n_257_76_17126));
   NAND2_X1 i_257_76_17157 (.A1(n_257_76_16845), .A2(n_257_76_17126), .ZN(
      n_257_76_17127));
   INV_X1 i_257_76_17158 (.A(n_257_76_17127), .ZN(n_257_76_17128));
   NAND2_X1 i_257_76_17159 (.A1(n_257_76_18067), .A2(n_257_76_17128), .ZN(
      n_257_76_17129));
   NAND4_X1 i_257_76_17160 (.A1(n_257_76_16867), .A2(n_257_76_16868), .A3(
      n_257_76_16869), .A4(n_257_76_16873), .ZN(n_257_76_17130));
   NAND4_X1 i_257_76_17161 (.A1(n_257_76_16944), .A2(n_257_76_16874), .A3(
      n_257_76_16875), .A4(n_257_76_16935), .ZN(n_257_76_17131));
   NOR2_X1 i_257_76_17162 (.A1(n_257_76_17130), .A2(n_257_76_17131), .ZN(
      n_257_76_17132));
   NAND4_X1 i_257_76_17163 (.A1(n_257_76_16914), .A2(n_257_76_16915), .A3(
      n_257_76_16847), .A4(n_257_76_16941), .ZN(n_257_76_17133));
   INV_X1 i_257_76_17164 (.A(n_257_76_17133), .ZN(n_257_76_17134));
   NAND4_X1 i_257_76_17165 (.A1(n_257_76_17132), .A2(n_257_76_17134), .A3(
      n_257_76_16866), .A4(n_257_76_16846), .ZN(n_257_76_17135));
   NAND2_X1 i_257_76_17166 (.A1(n_257_442), .A2(n_257_499), .ZN(n_257_76_17136));
   NOR2_X1 i_257_76_17167 (.A1(n_257_1089), .A2(n_257_76_17136), .ZN(
      n_257_76_17137));
   NAND2_X1 i_257_76_17168 (.A1(n_257_428), .A2(n_257_595), .ZN(n_257_76_17138));
   NAND3_X1 i_257_76_17169 (.A1(n_257_76_17137), .A2(n_257_76_17138), .A3(
      n_257_420), .ZN(n_257_76_17139));
   INV_X1 i_257_76_17170 (.A(n_257_76_17139), .ZN(n_257_76_17140));
   NAND2_X1 i_257_76_17171 (.A1(n_257_340), .A2(n_257_422), .ZN(n_257_76_17141));
   NAND4_X1 i_257_76_17172 (.A1(n_257_76_17140), .A2(n_257_76_16877), .A3(
      n_257_76_16921), .A4(n_257_76_17141), .ZN(n_257_76_17142));
   NAND2_X1 i_257_76_17173 (.A1(n_257_76_16916), .A2(n_257_76_16917), .ZN(
      n_257_76_17143));
   NOR2_X1 i_257_76_17174 (.A1(n_257_76_17142), .A2(n_257_76_17143), .ZN(
      n_257_76_17144));
   NAND2_X1 i_257_76_17175 (.A1(n_257_76_16884), .A2(n_257_76_16920), .ZN(
      n_257_76_17145));
   INV_X1 i_257_76_17176 (.A(n_257_76_17145), .ZN(n_257_76_17146));
   NAND2_X1 i_257_76_17177 (.A1(n_257_302), .A2(n_257_423), .ZN(n_257_76_17147));
   NAND2_X1 i_257_76_17178 (.A1(n_257_76_17147), .A2(n_257_76_16938), .ZN(
      n_257_76_17148));
   INV_X1 i_257_76_17179 (.A(n_257_76_17148), .ZN(n_257_76_17149));
   NAND3_X1 i_257_76_17180 (.A1(n_257_76_17144), .A2(n_257_76_17146), .A3(
      n_257_76_17149), .ZN(n_257_76_17150));
   NAND2_X1 i_257_76_17181 (.A1(n_257_379), .A2(n_257_421), .ZN(n_257_76_17151));
   NAND4_X1 i_257_76_17182 (.A1(n_257_76_16936), .A2(n_257_76_16882), .A3(
      n_257_76_16883), .A4(n_257_76_17151), .ZN(n_257_76_17152));
   NOR2_X1 i_257_76_17183 (.A1(n_257_76_17150), .A2(n_257_76_17152), .ZN(
      n_257_76_17153));
   NAND2_X1 i_257_76_17184 (.A1(n_257_76_16845), .A2(n_257_76_17153), .ZN(
      n_257_76_17154));
   NOR2_X1 i_257_76_17185 (.A1(n_257_76_17135), .A2(n_257_76_17154), .ZN(
      n_257_76_17155));
   NAND2_X1 i_257_76_17186 (.A1(n_257_76_18073), .A2(n_257_76_17155), .ZN(
      n_257_76_17156));
   NAND4_X1 i_257_76_17187 (.A1(n_257_76_16847), .A2(n_257_76_16941), .A3(
      n_257_76_16867), .A4(n_257_76_16868), .ZN(n_257_76_17157));
   NOR2_X1 i_257_76_17188 (.A1(n_257_76_16933), .A2(n_257_76_17157), .ZN(
      n_257_76_17158));
   NAND2_X1 i_257_76_17189 (.A1(n_257_76_16875), .A2(n_257_76_16882), .ZN(
      n_257_76_17159));
   INV_X1 i_257_76_17190 (.A(n_257_76_17159), .ZN(n_257_76_17160));
   INV_X1 i_257_76_17191 (.A(n_257_76_17009), .ZN(n_257_76_17161));
   INV_X1 i_257_76_17192 (.A(n_257_430), .ZN(n_257_76_17162));
   NOR2_X1 i_257_76_17193 (.A1(n_257_76_16849), .A2(n_257_76_17162), .ZN(
      n_257_76_17163));
   NAND3_X1 i_257_76_17194 (.A1(n_257_76_17163), .A2(n_257_76_16877), .A3(
      n_257_76_16921), .ZN(n_257_76_17164));
   INV_X1 i_257_76_17195 (.A(n_257_76_17164), .ZN(n_257_76_17165));
   NAND3_X1 i_257_76_17196 (.A1(n_257_76_17165), .A2(n_257_143), .A3(
      n_257_76_16916), .ZN(n_257_76_17166));
   INV_X1 i_257_76_17197 (.A(n_257_76_17166), .ZN(n_257_76_17167));
   NAND3_X1 i_257_76_17198 (.A1(n_257_76_17160), .A2(n_257_76_17161), .A3(
      n_257_76_17167), .ZN(n_257_76_17168));
   NOR2_X1 i_257_76_17199 (.A1(n_257_76_17168), .A2(n_257_76_16945), .ZN(
      n_257_76_17169));
   NAND4_X1 i_257_76_17200 (.A1(n_257_76_17158), .A2(n_257_76_16845), .A3(
      n_257_76_16866), .A4(n_257_76_17169), .ZN(n_257_76_17170));
   INV_X1 i_257_76_17201 (.A(n_257_76_17170), .ZN(n_257_76_17171));
   NAND2_X1 i_257_76_17202 (.A1(n_257_76_18068), .A2(n_257_76_17171), .ZN(
      n_257_76_17172));
   NAND3_X1 i_257_76_17203 (.A1(n_257_76_17129), .A2(n_257_76_17156), .A3(
      n_257_76_17172), .ZN(n_257_76_17173));
   INV_X1 i_257_76_17204 (.A(n_257_76_17173), .ZN(n_257_76_17174));
   NAND2_X1 i_257_76_17205 (.A1(n_257_795), .A2(n_257_442), .ZN(n_257_76_17175));
   NOR2_X1 i_257_76_17206 (.A1(n_257_1089), .A2(n_257_76_17175), .ZN(
      n_257_76_17176));
   NAND4_X1 i_257_76_17207 (.A1(n_257_447), .A2(n_257_76_16883), .A3(
      n_257_76_16884), .A4(n_257_76_17176), .ZN(n_257_76_17177));
   NOR2_X1 i_257_76_17208 (.A1(n_257_76_17026), .A2(n_257_76_17177), .ZN(
      n_257_76_17178));
   NAND3_X1 i_257_76_17209 (.A1(n_257_76_17178), .A2(n_257_76_16846), .A3(
      n_257_76_17059), .ZN(n_257_76_17179));
   NOR2_X1 i_257_76_17210 (.A1(n_257_76_16888), .A2(n_257_76_17179), .ZN(
      n_257_76_17180));
   NAND3_X1 i_257_76_17211 (.A1(n_257_76_16875), .A2(n_257_76_16882), .A3(
      n_257_76_16883), .ZN(n_257_76_17181));
   INV_X1 i_257_76_17212 (.A(n_257_76_17181), .ZN(n_257_76_17182));
   INV_X1 i_257_76_17213 (.A(n_257_431), .ZN(n_257_76_17183));
   NOR2_X1 i_257_76_17214 (.A1(n_257_76_16849), .A2(n_257_76_17183), .ZN(
      n_257_76_17184));
   NAND3_X1 i_257_76_17215 (.A1(n_257_76_17184), .A2(n_257_76_16877), .A3(
      n_257_76_16921), .ZN(n_257_76_17185));
   INV_X1 i_257_76_17216 (.A(n_257_76_17185), .ZN(n_257_76_17186));
   NAND4_X1 i_257_76_17217 (.A1(n_257_76_17186), .A2(n_257_76_16884), .A3(
      n_257_76_16920), .A4(n_257_76_16916), .ZN(n_257_76_17187));
   INV_X1 i_257_76_17218 (.A(n_257_76_17187), .ZN(n_257_76_17188));
   NAND2_X1 i_257_76_17219 (.A1(n_257_76_17182), .A2(n_257_76_17188), .ZN(
      n_257_76_17189));
   NAND3_X1 i_257_76_17220 (.A1(n_257_76_16944), .A2(n_257_76_16874), .A3(
      n_257_105), .ZN(n_257_76_17190));
   NOR3_X1 i_257_76_17221 (.A1(n_257_76_17189), .A2(n_257_76_17108), .A3(
      n_257_76_17190), .ZN(n_257_76_17191));
   NAND2_X1 i_257_76_17222 (.A1(n_257_76_16846), .A2(n_257_76_17059), .ZN(
      n_257_76_17192));
   INV_X1 i_257_76_17223 (.A(n_257_76_17192), .ZN(n_257_76_17193));
   NAND4_X1 i_257_76_17224 (.A1(n_257_76_17191), .A2(n_257_76_16845), .A3(
      n_257_76_17193), .A4(n_257_76_16866), .ZN(n_257_76_17194));
   INV_X1 i_257_76_17225 (.A(n_257_76_17194), .ZN(n_257_76_17195));
   AOI22_X1 i_257_76_17226 (.A1(n_257_76_18085), .A2(n_257_76_17180), .B1(
      n_257_76_18080), .B2(n_257_76_17195), .ZN(n_257_76_17196));
   NAND3_X1 i_257_76_17227 (.A1(n_257_76_17118), .A2(n_257_76_17174), .A3(
      n_257_76_17196), .ZN(n_257_76_17197));
   NAND3_X1 i_257_76_17228 (.A1(n_257_76_16884), .A2(n_257_448), .A3(
      n_257_76_17978), .ZN(n_257_76_17198));
   NOR2_X1 i_257_76_17229 (.A1(n_257_76_17198), .A2(n_257_76_17079), .ZN(
      n_257_76_17199));
   INV_X1 i_257_76_17230 (.A(n_257_76_16876), .ZN(n_257_76_17200));
   INV_X1 i_257_76_17231 (.A(n_257_76_16967), .ZN(n_257_76_17201));
   NAND4_X1 i_257_76_17232 (.A1(n_257_76_17199), .A2(n_257_76_17200), .A3(
      n_257_76_17201), .A4(n_257_76_16847), .ZN(n_257_76_17202));
   INV_X1 i_257_76_17233 (.A(n_257_76_17202), .ZN(n_257_76_17203));
   NAND2_X1 i_257_76_17234 (.A1(n_257_76_16846), .A2(n_257_699), .ZN(
      n_257_76_17204));
   INV_X1 i_257_76_17235 (.A(n_257_76_17204), .ZN(n_257_76_17205));
   NAND3_X1 i_257_76_17236 (.A1(n_257_76_17203), .A2(n_257_76_16845), .A3(
      n_257_76_17205), .ZN(n_257_76_17206));
   INV_X1 i_257_76_17237 (.A(n_257_76_17206), .ZN(n_257_76_17207));
   NAND2_X1 i_257_76_17238 (.A1(n_257_76_18079), .A2(n_257_76_17207), .ZN(
      n_257_76_17208));
   NAND2_X1 i_257_76_17239 (.A1(n_257_76_16846), .A2(n_257_76_16847), .ZN(
      n_257_76_17209));
   INV_X1 i_257_76_17240 (.A(n_257_76_17209), .ZN(n_257_76_17210));
   NAND3_X1 i_257_76_17241 (.A1(n_257_76_16845), .A2(n_257_76_17210), .A3(
      n_257_76_16866), .ZN(n_257_76_17211));
   INV_X1 i_257_76_17242 (.A(n_257_76_17079), .ZN(n_257_76_17212));
   NAND2_X1 i_257_76_17243 (.A1(n_257_76_16877), .A2(n_257_76_16921), .ZN(
      n_257_76_17213));
   INV_X1 i_257_76_17244 (.A(n_257_76_17213), .ZN(n_257_76_17214));
   NAND2_X1 i_257_76_17245 (.A1(n_257_76_16925), .A2(n_257_425), .ZN(
      n_257_76_17215));
   INV_X1 i_257_76_17246 (.A(n_257_76_17215), .ZN(n_257_76_17216));
   NAND2_X1 i_257_76_17247 (.A1(n_257_76_17216), .A2(n_257_76_16924), .ZN(
      n_257_76_17217));
   INV_X1 i_257_76_17248 (.A(n_257_76_17217), .ZN(n_257_76_17218));
   NAND4_X1 i_257_76_17249 (.A1(n_257_76_16938), .A2(n_257_76_17214), .A3(
      n_257_76_16916), .A4(n_257_76_17218), .ZN(n_257_76_17219));
   INV_X1 i_257_76_17250 (.A(n_257_76_17219), .ZN(n_257_76_17220));
   NAND3_X1 i_257_76_17251 (.A1(n_257_76_17212), .A2(n_257_76_17220), .A3(
      n_257_76_17146), .ZN(n_257_76_17221));
   NAND4_X1 i_257_76_17252 (.A1(n_257_76_16874), .A2(n_257_76_16875), .A3(
      n_257_76_16935), .A4(n_257_76_16936), .ZN(n_257_76_17222));
   NOR2_X1 i_257_76_17253 (.A1(n_257_76_17221), .A2(n_257_76_17222), .ZN(
      n_257_76_17223));
   NAND2_X1 i_257_76_17254 (.A1(n_257_76_16914), .A2(n_257_76_16941), .ZN(
      n_257_76_17224));
   INV_X1 i_257_76_17255 (.A(n_257_76_17224), .ZN(n_257_76_17225));
   NAND3_X1 i_257_76_17256 (.A1(n_257_262), .A2(n_257_76_16867), .A3(
      n_257_76_16868), .ZN(n_257_76_17226));
   NAND3_X1 i_257_76_17257 (.A1(n_257_76_16869), .A2(n_257_76_16873), .A3(
      n_257_76_16944), .ZN(n_257_76_17227));
   NOR2_X1 i_257_76_17258 (.A1(n_257_76_17226), .A2(n_257_76_17227), .ZN(
      n_257_76_17228));
   NAND3_X1 i_257_76_17259 (.A1(n_257_76_17223), .A2(n_257_76_17225), .A3(
      n_257_76_17228), .ZN(n_257_76_17229));
   NOR2_X1 i_257_76_17260 (.A1(n_257_76_17211), .A2(n_257_76_17229), .ZN(
      n_257_76_17230));
   NAND2_X1 i_257_76_17261 (.A1(n_257_76_18064), .A2(n_257_76_17230), .ZN(
      n_257_76_17231));
   INV_X1 i_257_76_17262 (.A(n_257_76_16937), .ZN(n_257_76_17232));
   INV_X1 i_257_76_17263 (.A(n_257_76_16939), .ZN(n_257_76_17233));
   NAND2_X1 i_257_76_17264 (.A1(n_257_76_17232), .A2(n_257_76_17233), .ZN(
      n_257_76_17234));
   NOR3_X1 i_257_76_17265 (.A1(n_257_76_17234), .A2(n_257_76_16870), .A3(
      n_257_76_16974), .ZN(n_257_76_17235));
   NAND3_X1 i_257_76_17266 (.A1(n_257_379), .A2(n_257_76_16916), .A3(
      n_257_76_16917), .ZN(n_257_76_17236));
   INV_X1 i_257_76_17267 (.A(n_257_76_17236), .ZN(n_257_76_17237));
   NAND2_X1 i_257_76_17268 (.A1(n_257_76_16925), .A2(n_257_421), .ZN(
      n_257_76_17238));
   INV_X1 i_257_76_17269 (.A(n_257_76_17238), .ZN(n_257_76_17239));
   NAND3_X1 i_257_76_17270 (.A1(n_257_76_17141), .A2(n_257_76_16924), .A3(
      n_257_76_17239), .ZN(n_257_76_17240));
   NOR2_X1 i_257_76_17271 (.A1(n_257_76_17213), .A2(n_257_76_17240), .ZN(
      n_257_76_17241));
   NAND4_X1 i_257_76_17272 (.A1(n_257_76_17237), .A2(n_257_76_17241), .A3(
      n_257_76_16920), .A4(n_257_76_17147), .ZN(n_257_76_17242));
   INV_X1 i_257_76_17273 (.A(n_257_76_17242), .ZN(n_257_76_17243));
   NAND2_X1 i_257_76_17274 (.A1(n_257_76_16914), .A2(n_257_76_17243), .ZN(
      n_257_76_17244));
   NAND3_X1 i_257_76_17275 (.A1(n_257_76_16915), .A2(n_257_76_16847), .A3(
      n_257_76_16941), .ZN(n_257_76_17245));
   NOR2_X1 i_257_76_17276 (.A1(n_257_76_17244), .A2(n_257_76_17245), .ZN(
      n_257_76_17246));
   NAND4_X1 i_257_76_17277 (.A1(n_257_76_17049), .A2(n_257_76_17235), .A3(
      n_257_76_16845), .A4(n_257_76_17246), .ZN(n_257_76_17247));
   INV_X1 i_257_76_17278 (.A(n_257_76_17247), .ZN(n_257_76_17248));
   NAND2_X1 i_257_76_17279 (.A1(n_257_76_18082), .A2(n_257_76_17248), .ZN(
      n_257_76_17249));
   NAND3_X1 i_257_76_17280 (.A1(n_257_76_17208), .A2(n_257_76_17231), .A3(
      n_257_76_17249), .ZN(n_257_76_17250));
   INV_X1 i_257_76_17281 (.A(n_257_76_17250), .ZN(n_257_76_17251));
   NAND2_X1 i_257_76_17282 (.A1(n_257_76_16875), .A2(n_257_76_16936), .ZN(
      n_257_76_17252));
   NAND3_X1 i_257_76_17283 (.A1(n_257_76_16882), .A2(n_257_76_16883), .A3(
      n_257_76_16884), .ZN(n_257_76_17253));
   NOR2_X1 i_257_76_17284 (.A1(n_257_76_17252), .A2(n_257_76_17253), .ZN(
      n_257_76_17254));
   INV_X1 i_257_76_17285 (.A(n_257_76_16870), .ZN(n_257_76_17255));
   INV_X1 i_257_76_17286 (.A(n_257_76_16974), .ZN(n_257_76_17256));
   NAND3_X1 i_257_76_17287 (.A1(n_257_76_17254), .A2(n_257_76_17255), .A3(
      n_257_76_17256), .ZN(n_257_76_17257));
   INV_X1 i_257_76_17288 (.A(n_257_76_17257), .ZN(n_257_76_17258));
   NAND4_X1 i_257_76_17289 (.A1(n_257_427), .A2(n_257_76_16877), .A3(
      n_257_76_16921), .A4(n_257_222), .ZN(n_257_76_17259));
   INV_X1 i_257_76_17290 (.A(n_257_76_17259), .ZN(n_257_76_17260));
   NAND2_X1 i_257_76_17291 (.A1(n_257_76_16924), .A2(n_257_76_16925), .ZN(
      n_257_76_17261));
   INV_X1 i_257_76_17292 (.A(n_257_76_17261), .ZN(n_257_76_17262));
   NAND2_X1 i_257_76_17293 (.A1(n_257_76_16916), .A2(n_257_76_17262), .ZN(
      n_257_76_17263));
   INV_X1 i_257_76_17294 (.A(n_257_76_17263), .ZN(n_257_76_17264));
   NAND3_X1 i_257_76_17295 (.A1(n_257_76_17260), .A2(n_257_76_17264), .A3(
      n_257_76_16920), .ZN(n_257_76_17265));
   INV_X1 i_257_76_17296 (.A(n_257_76_17265), .ZN(n_257_76_17266));
   NAND4_X1 i_257_76_17297 (.A1(n_257_76_16914), .A2(n_257_76_16847), .A3(
      n_257_76_17266), .A4(n_257_76_16941), .ZN(n_257_76_17267));
   INV_X1 i_257_76_17298 (.A(n_257_76_17267), .ZN(n_257_76_17268));
   NAND2_X1 i_257_76_17299 (.A1(n_257_76_17258), .A2(n_257_76_17268), .ZN(
      n_257_76_17269));
   NOR3_X1 i_257_76_17300 (.A1(n_257_76_17269), .A2(n_257_76_16888), .A3(
      n_257_76_17048), .ZN(n_257_76_17270));
   NAND2_X1 i_257_76_17301 (.A1(n_257_76_18065), .A2(n_257_76_17270), .ZN(
      n_257_76_17271));
   NAND4_X1 i_257_76_17302 (.A1(n_257_76_16884), .A2(n_257_76_16920), .A3(
      n_257_76_17978), .A4(n_257_482), .ZN(n_257_76_17272));
   NAND3_X1 i_257_76_17303 (.A1(n_257_76_16882), .A2(n_257_451), .A3(
      n_257_76_16883), .ZN(n_257_76_17273));
   NOR2_X1 i_257_76_17304 (.A1(n_257_76_17272), .A2(n_257_76_17273), .ZN(
      n_257_76_17274));
   NAND3_X1 i_257_76_17305 (.A1(n_257_76_17274), .A2(n_257_76_17255), .A3(
      n_257_76_17200), .ZN(n_257_76_17275));
   INV_X1 i_257_76_17306 (.A(n_257_76_17275), .ZN(n_257_76_17276));
   NAND4_X1 i_257_76_17307 (.A1(n_257_76_17276), .A2(n_257_76_16845), .A3(
      n_257_76_17210), .A4(n_257_76_16866), .ZN(n_257_76_17277));
   INV_X1 i_257_76_17308 (.A(n_257_76_17277), .ZN(n_257_76_17278));
   NAND2_X1 i_257_76_17309 (.A1(n_257_76_18063), .A2(n_257_76_17278), .ZN(
      n_257_76_17279));
   NOR2_X1 i_257_76_17310 (.A1(n_257_76_17133), .A2(n_257_76_16933), .ZN(
      n_257_76_17280));
   NAND4_X1 i_257_76_17311 (.A1(n_257_76_16920), .A2(n_257_76_16938), .A3(
      n_257_76_16916), .A4(n_257_76_17214), .ZN(n_257_76_17281));
   NOR2_X1 i_257_76_17312 (.A1(n_257_76_17253), .A2(n_257_76_17281), .ZN(
      n_257_76_17282));
   INV_X1 i_257_76_17313 (.A(n_257_76_17222), .ZN(n_257_76_17283));
   NAND3_X1 i_257_76_17314 (.A1(n_257_76_17262), .A2(n_257_531), .A3(n_257_424), 
      .ZN(n_257_76_17284));
   INV_X1 i_257_76_17315 (.A(n_257_76_17284), .ZN(n_257_76_17285));
   NAND3_X1 i_257_76_17316 (.A1(n_257_76_16873), .A2(n_257_76_16944), .A3(
      n_257_76_17285), .ZN(n_257_76_17286));
   INV_X1 i_257_76_17317 (.A(n_257_76_17286), .ZN(n_257_76_17287));
   NAND4_X1 i_257_76_17318 (.A1(n_257_76_17282), .A2(n_257_76_17255), .A3(
      n_257_76_17283), .A4(n_257_76_17287), .ZN(n_257_76_17288));
   INV_X1 i_257_76_17319 (.A(n_257_76_17288), .ZN(n_257_76_17289));
   NAND4_X1 i_257_76_17320 (.A1(n_257_76_17280), .A2(n_257_76_17289), .A3(
      n_257_76_16845), .A4(n_257_76_16866), .ZN(n_257_76_17290));
   INV_X1 i_257_76_17321 (.A(n_257_76_17290), .ZN(n_257_76_17291));
   NAND2_X1 i_257_76_17322 (.A1(n_257_76_18062), .A2(n_257_76_17291), .ZN(
      n_257_76_17292));
   NAND3_X1 i_257_76_17323 (.A1(n_257_76_17271), .A2(n_257_76_17279), .A3(
      n_257_76_17292), .ZN(n_257_76_17293));
   INV_X1 i_257_76_17324 (.A(n_257_76_17293), .ZN(n_257_76_17294));
   NAND3_X1 i_257_76_17325 (.A1(n_257_76_16914), .A2(n_257_76_16915), .A3(
      n_257_76_16847), .ZN(n_257_76_17295));
   NAND4_X1 i_257_76_17326 (.A1(n_257_76_16941), .A2(n_257_76_16867), .A3(
      n_257_76_16868), .A4(n_257_76_16869), .ZN(n_257_76_17296));
   NOR2_X1 i_257_76_17327 (.A1(n_257_76_17295), .A2(n_257_76_17296), .ZN(
      n_257_76_17297));
   NOR2_X1 i_257_76_17328 (.A1(n_257_76_17261), .A2(n_257_76_17141), .ZN(
      n_257_76_17298));
   NAND4_X1 i_257_76_17329 (.A1(n_257_76_17298), .A2(n_257_76_16884), .A3(
      n_257_76_16920), .A4(n_257_76_17147), .ZN(n_257_76_17299));
   NAND4_X1 i_257_76_17330 (.A1(n_257_76_16938), .A2(n_257_76_17214), .A3(
      n_257_76_16916), .A4(n_257_76_16917), .ZN(n_257_76_17300));
   NOR2_X1 i_257_76_17331 (.A1(n_257_76_17299), .A2(n_257_76_17300), .ZN(
      n_257_76_17301));
   NAND2_X1 i_257_76_17332 (.A1(n_257_76_16875), .A2(n_257_76_16935), .ZN(
      n_257_76_17302));
   NOR2_X1 i_257_76_17333 (.A1(n_257_76_17106), .A2(n_257_76_17302), .ZN(
      n_257_76_17303));
   NAND3_X1 i_257_76_17334 (.A1(n_257_76_17256), .A2(n_257_76_17301), .A3(
      n_257_76_17303), .ZN(n_257_76_17304));
   INV_X1 i_257_76_17335 (.A(n_257_76_17304), .ZN(n_257_76_17305));
   NAND4_X1 i_257_76_17336 (.A1(n_257_76_17049), .A2(n_257_76_17297), .A3(
      n_257_76_17305), .A4(n_257_76_16845), .ZN(n_257_76_17306));
   INV_X1 i_257_76_17337 (.A(n_257_76_17306), .ZN(n_257_76_17307));
   NAND2_X1 i_257_76_17338 (.A1(n_257_342), .A2(n_257_76_17307), .ZN(
      n_257_76_17308));
   NAND3_X1 i_257_76_17339 (.A1(n_257_76_16938), .A2(n_257_76_16916), .A3(
      n_257_76_16917), .ZN(n_257_76_17309));
   INV_X1 i_257_76_17340 (.A(n_257_76_17309), .ZN(n_257_76_17310));
   NAND2_X1 i_257_76_17341 (.A1(n_257_442), .A2(n_257_418), .ZN(n_257_76_17311));
   INV_X1 i_257_76_17342 (.A(n_257_76_17311), .ZN(n_257_76_17312));
   NAND2_X1 i_257_76_17343 (.A1(n_257_484), .A2(n_257_76_17312), .ZN(
      n_257_76_17313));
   NOR2_X1 i_257_76_17344 (.A1(n_257_76_17313), .A2(n_257_1089), .ZN(
      n_257_76_17314));
   NAND2_X1 i_257_76_17345 (.A1(n_257_420), .A2(n_257_499), .ZN(n_257_76_17315));
   NAND3_X1 i_257_76_17346 (.A1(n_257_76_17314), .A2(n_257_76_17315), .A3(
      n_257_76_17138), .ZN(n_257_76_17316));
   INV_X1 i_257_76_17347 (.A(n_257_76_17316), .ZN(n_257_76_17317));
   NAND4_X1 i_257_76_17348 (.A1(n_257_76_17317), .A2(n_257_76_16877), .A3(
      n_257_76_16921), .A4(n_257_76_17141), .ZN(n_257_76_17318));
   INV_X1 i_257_76_17349 (.A(n_257_76_17318), .ZN(n_257_76_17319));
   NAND2_X1 i_257_76_17350 (.A1(n_257_76_17310), .A2(n_257_76_17319), .ZN(
      n_257_76_17320));
   NAND3_X1 i_257_76_17351 (.A1(n_257_76_16882), .A2(n_257_76_16883), .A3(
      n_257_76_17151), .ZN(n_257_76_17321));
   NAND3_X1 i_257_76_17352 (.A1(n_257_76_16884), .A2(n_257_76_16920), .A3(
      n_257_76_17147), .ZN(n_257_76_17322));
   NOR3_X1 i_257_76_17353 (.A1(n_257_76_17320), .A2(n_257_76_17321), .A3(
      n_257_76_17322), .ZN(n_257_76_17323));
   NAND3_X1 i_257_76_17354 (.A1(n_257_76_17323), .A2(n_257_76_16866), .A3(
      n_257_76_16846), .ZN(n_257_76_17324));
   INV_X1 i_257_76_17355 (.A(n_257_76_17324), .ZN(n_257_76_17325));
   NAND3_X1 i_257_76_17356 (.A1(n_257_76_17255), .A2(n_257_76_17256), .A3(
      n_257_76_17232), .ZN(n_257_76_17326));
   NOR2_X1 i_257_76_17357 (.A1(n_257_76_17326), .A2(n_257_76_17133), .ZN(
      n_257_76_17327));
   NAND3_X1 i_257_76_17358 (.A1(n_257_76_17325), .A2(n_257_76_16845), .A3(
      n_257_76_17327), .ZN(n_257_76_17328));
   INV_X1 i_257_76_17359 (.A(n_257_76_17328), .ZN(n_257_76_17329));
   NAND2_X1 i_257_76_17360 (.A1(n_257_76_18060), .A2(n_257_76_17329), .ZN(
      n_257_76_17330));
   INV_X1 i_257_76_17361 (.A(n_257_76_17660), .ZN(n_257_76_17331));
   NAND2_X1 i_257_76_17362 (.A1(n_257_182), .A2(n_257_76_17331), .ZN(
      n_257_76_17332));
   NAND2_X1 i_257_76_17363 (.A1(n_257_76_17242), .A2(n_257_76_17332), .ZN(
      n_257_76_17333));
   INV_X1 i_257_76_17364 (.A(n_257_76_17333), .ZN(n_257_76_17334));
   NAND2_X1 i_257_76_17365 (.A1(n_257_699), .A2(n_257_76_17958), .ZN(
      n_257_76_17335));
   NAND2_X1 i_257_76_17366 (.A1(n_257_1025), .A2(n_257_76_17964), .ZN(
      n_257_76_17336));
   NAND2_X1 i_257_76_17367 (.A1(n_257_993), .A2(n_257_442), .ZN(n_257_76_17337));
   INV_X1 i_257_76_17368 (.A(n_257_76_17337), .ZN(n_257_76_17338));
   NAND2_X1 i_257_76_17369 (.A1(n_257_441), .A2(n_257_76_17338), .ZN(
      n_257_76_17339));
   NAND2_X1 i_257_76_17370 (.A1(n_257_105), .A2(n_257_76_17932), .ZN(
      n_257_76_17340));
   NAND3_X1 i_257_76_17371 (.A1(n_257_76_17339), .A2(n_257_76_16930), .A3(
      n_257_76_17340), .ZN(n_257_76_17341));
   INV_X1 i_257_76_17372 (.A(n_257_76_17341), .ZN(n_257_76_17342));
   NAND4_X1 i_257_76_17373 (.A1(n_257_76_17334), .A2(n_257_76_17335), .A3(
      n_257_76_17336), .A4(n_257_76_17342), .ZN(n_257_76_17343));
   INV_X1 i_257_76_17374 (.A(n_257_76_17343), .ZN(n_257_76_17344));
   INV_X1 i_257_76_17375 (.A(n_257_1057), .ZN(n_257_76_17345));
   OAI21_X1 i_257_76_17376 (.A(n_257_76_17014), .B1(n_257_76_17345), .B2(
      n_257_76_17968), .ZN(n_257_76_17346));
   INV_X1 i_257_76_17377 (.A(n_257_76_17346), .ZN(n_257_76_17347));
   NAND2_X1 i_257_76_17378 (.A1(n_257_482), .A2(n_257_442), .ZN(n_257_76_17348));
   INV_X1 i_257_76_17379 (.A(n_257_76_17348), .ZN(n_257_76_17349));
   NAND2_X1 i_257_76_17380 (.A1(n_257_76_17349), .A2(n_257_451), .ZN(
      n_257_76_17350));
   NAND2_X1 i_257_76_17381 (.A1(n_257_859), .A2(n_257_442), .ZN(n_257_76_17351));
   INV_X1 i_257_76_17382 (.A(n_257_76_17351), .ZN(n_257_76_17352));
   NAND2_X1 i_257_76_17383 (.A1(n_257_446), .A2(n_257_76_17352), .ZN(
      n_257_76_17353));
   INV_X1 i_257_76_17384 (.A(n_257_76_17090), .ZN(n_257_76_17354));
   NAND2_X1 i_257_76_17385 (.A1(n_257_449), .A2(n_257_76_17354), .ZN(
      n_257_76_17355));
   NAND4_X1 i_257_76_17386 (.A1(n_257_76_17265), .A2(n_257_76_17350), .A3(
      n_257_76_17353), .A4(n_257_76_17355), .ZN(n_257_76_17356));
   INV_X1 i_257_76_17387 (.A(n_257_76_17356), .ZN(n_257_76_17357));
   INV_X1 i_257_76_17388 (.A(n_257_76_17175), .ZN(n_257_76_17358));
   NAND2_X1 i_257_76_17389 (.A1(n_257_447), .A2(n_257_76_17358), .ZN(
      n_257_76_17359));
   NAND2_X1 i_257_76_17390 (.A1(n_257_827), .A2(n_257_76_17952), .ZN(
      n_257_76_17360));
   NAND2_X1 i_257_76_17391 (.A1(n_257_143), .A2(n_257_76_17925), .ZN(
      n_257_76_17361));
   NAND3_X1 i_257_76_17392 (.A1(n_257_76_17359), .A2(n_257_76_17360), .A3(
      n_257_76_17361), .ZN(n_257_76_17362));
   NAND2_X1 i_257_76_17393 (.A1(n_257_763), .A2(n_257_76_17935), .ZN(
      n_257_76_17363));
   NAND2_X1 i_257_76_17394 (.A1(n_257_76_17940), .A2(n_257_929), .ZN(
      n_257_76_17364));
   NAND2_X1 i_257_76_17395 (.A1(n_257_76_17363), .A2(n_257_76_17364), .ZN(
      n_257_76_17365));
   NOR2_X1 i_257_76_17396 (.A1(n_257_76_17362), .A2(n_257_76_17365), .ZN(
      n_257_76_17366));
   NAND2_X1 i_257_76_17397 (.A1(n_257_65), .A2(n_257_76_17918), .ZN(
      n_257_76_17367));
   NAND3_X1 i_257_76_17398 (.A1(n_257_731), .A2(n_257_435), .A3(n_257_442), 
      .ZN(n_257_76_17368));
   INV_X1 i_257_76_17399 (.A(n_257_76_17037), .ZN(n_257_76_17369));
   NAND2_X1 i_257_76_17400 (.A1(n_257_432), .A2(n_257_76_17369), .ZN(
      n_257_76_17370));
   NAND3_X1 i_257_76_17401 (.A1(n_257_76_17367), .A2(n_257_76_17368), .A3(
      n_257_76_17370), .ZN(n_257_76_17371));
   INV_X1 i_257_76_17402 (.A(n_257_76_17371), .ZN(n_257_76_17372));
   NAND2_X1 i_257_76_17403 (.A1(n_257_659), .A2(n_257_76_17928), .ZN(
      n_257_76_17373));
   INV_X1 i_257_76_17404 (.A(n_257_418), .ZN(n_257_76_17374));
   NAND2_X1 i_257_76_17405 (.A1(n_257_76_17374), .A2(Small_Packet_Data_Size[30]), 
      .ZN(n_257_76_17375));
   INV_X1 i_257_76_17406 (.A(Small_Packet_Data_Size[30]), .ZN(n_257_76_17376));
   OAI21_X1 i_257_76_17407 (.A(n_257_76_17375), .B1(n_257_484), .B2(
      n_257_76_17376), .ZN(n_257_76_17377));
   NAND4_X1 i_257_76_17408 (.A1(n_257_76_17315), .A2(n_257_76_17377), .A3(
      n_257_76_17138), .A4(n_257_76_16925), .ZN(n_257_76_17378));
   NAND2_X1 i_257_76_17409 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[30]), 
      .ZN(n_257_76_17379));
   NAND2_X1 i_257_76_17410 (.A1(n_257_76_17378), .A2(n_257_76_17379), .ZN(
      n_257_76_17380));
   INV_X1 i_257_76_17411 (.A(n_257_76_17298), .ZN(n_257_76_17381));
   NAND4_X1 i_257_76_17412 (.A1(n_257_76_17372), .A2(n_257_76_17373), .A3(
      n_257_76_17380), .A4(n_257_76_17381), .ZN(n_257_76_17382));
   NAND2_X1 i_257_76_17413 (.A1(n_257_891), .A2(n_257_76_17903), .ZN(
      n_257_76_17383));
   NAND2_X1 i_257_76_17414 (.A1(n_257_961), .A2(n_257_442), .ZN(n_257_76_17384));
   INV_X1 i_257_76_17415 (.A(n_257_76_17384), .ZN(n_257_76_17385));
   NAND2_X1 i_257_76_17416 (.A1(n_257_440), .A2(n_257_76_17385), .ZN(
      n_257_76_17386));
   INV_X1 i_257_76_17417 (.A(n_257_76_17119), .ZN(n_257_76_17387));
   NAND2_X1 i_257_76_17418 (.A1(n_257_438), .A2(n_257_76_17387), .ZN(
      n_257_76_17388));
   NAND4_X1 i_257_76_17419 (.A1(n_257_76_17383), .A2(n_257_76_17284), .A3(
      n_257_76_17386), .A4(n_257_76_17388), .ZN(n_257_76_17389));
   NOR2_X1 i_257_76_17420 (.A1(n_257_76_17382), .A2(n_257_76_17389), .ZN(
      n_257_76_17390));
   NAND3_X1 i_257_76_17421 (.A1(n_257_76_17357), .A2(n_257_76_17366), .A3(
      n_257_76_17390), .ZN(n_257_76_17391));
   INV_X1 i_257_76_17422 (.A(n_257_76_17391), .ZN(n_257_76_17392));
   NAND4_X1 i_257_76_17423 (.A1(n_257_76_17344), .A2(n_257_76_17347), .A3(
      n_257_76_17392), .A4(n_257_76_17229), .ZN(n_257_76_17393));
   NAND3_X1 i_257_76_17424 (.A1(n_257_76_17308), .A2(n_257_76_17330), .A3(
      n_257_76_17393), .ZN(n_257_76_17394));
   INV_X1 i_257_76_17425 (.A(n_257_76_17394), .ZN(n_257_76_17395));
   NAND3_X1 i_257_76_17426 (.A1(n_257_76_17251), .A2(n_257_76_17294), .A3(
      n_257_76_17395), .ZN(n_257_76_17396));
   NOR2_X1 i_257_76_17427 (.A1(n_257_76_17197), .A2(n_257_76_17396), .ZN(
      n_257_76_17397));
   NAND2_X1 i_257_76_17428 (.A1(n_257_76_17073), .A2(n_257_76_17397), .ZN(n_30));
   NAND2_X1 i_257_76_17429 (.A1(n_257_1026), .A2(n_257_444), .ZN(n_257_76_17398));
   NAND2_X1 i_257_76_17430 (.A1(n_257_441), .A2(n_257_994), .ZN(n_257_76_17399));
   NAND2_X1 i_257_76_17431 (.A1(n_257_962), .A2(n_257_442), .ZN(n_257_76_17400));
   NOR2_X1 i_257_76_17432 (.A1(n_257_1090), .A2(n_257_76_17400), .ZN(
      n_257_76_17401));
   NAND2_X1 i_257_76_17433 (.A1(n_257_440), .A2(n_257_76_17401), .ZN(
      n_257_76_17402));
   INV_X1 i_257_76_17434 (.A(n_257_76_17402), .ZN(n_257_76_17403));
   NAND2_X1 i_257_76_17435 (.A1(n_257_76_17399), .A2(n_257_76_17403), .ZN(
      n_257_76_17404));
   INV_X1 i_257_76_17436 (.A(n_257_76_17404), .ZN(n_257_76_17405));
   NAND2_X1 i_257_76_17437 (.A1(n_257_76_17398), .A2(n_257_76_17405), .ZN(
      n_257_76_17406));
   INV_X1 i_257_76_17438 (.A(n_257_76_17406), .ZN(n_257_76_17407));
   NAND2_X1 i_257_76_17439 (.A1(n_257_1058), .A2(n_257_443), .ZN(n_257_76_17408));
   NAND2_X1 i_257_76_17440 (.A1(n_257_76_17407), .A2(n_257_76_17408), .ZN(
      n_257_76_17409));
   INV_X1 i_257_76_17441 (.A(n_257_76_17409), .ZN(n_257_76_17410));
   NAND2_X1 i_257_76_17442 (.A1(n_257_17), .A2(n_257_76_17410), .ZN(
      n_257_76_17411));
   INV_X1 i_257_76_17443 (.A(n_257_442), .ZN(n_257_76_17412));
   NOR2_X1 i_257_76_17444 (.A1(n_257_1090), .A2(n_257_76_17412), .ZN(
      n_257_76_17413));
   NAND2_X1 i_257_76_17445 (.A1(n_257_443), .A2(n_257_76_17413), .ZN(
      n_257_76_17414));
   INV_X1 i_257_76_17446 (.A(n_257_76_17414), .ZN(n_257_76_17415));
   NAND2_X1 i_257_76_17447 (.A1(n_257_1058), .A2(n_257_76_17415), .ZN(
      n_257_76_17416));
   INV_X1 i_257_76_17448 (.A(n_257_76_17416), .ZN(n_257_76_17417));
   NAND2_X1 i_257_76_17449 (.A1(n_257_76_18072), .A2(n_257_76_17417), .ZN(
      n_257_76_17418));
   NAND2_X1 i_257_76_17450 (.A1(n_257_764), .A2(n_257_436), .ZN(n_257_76_17419));
   NAND2_X1 i_257_76_17451 (.A1(n_257_446), .A2(n_257_860), .ZN(n_257_76_17420));
   NAND2_X1 i_257_76_17452 (.A1(n_257_449), .A2(n_257_668), .ZN(n_257_76_17421));
   NAND3_X1 i_257_76_17453 (.A1(n_257_76_17419), .A2(n_257_76_17420), .A3(
      n_257_76_17421), .ZN(n_257_76_17422));
   INV_X1 i_257_76_17454 (.A(n_257_76_17422), .ZN(n_257_76_17423));
   NAND2_X1 i_257_76_17455 (.A1(n_257_447), .A2(n_257_796), .ZN(n_257_76_17424));
   NAND2_X1 i_257_76_17456 (.A1(n_257_930), .A2(n_257_439), .ZN(n_257_76_17425));
   NAND2_X1 i_257_76_17457 (.A1(n_257_828), .A2(n_257_437), .ZN(n_257_76_17426));
   NAND3_X1 i_257_76_17458 (.A1(n_257_76_17424), .A2(n_257_76_17425), .A3(
      n_257_76_17426), .ZN(n_257_76_17427));
   INV_X1 i_257_76_17459 (.A(n_257_76_17427), .ZN(n_257_76_17428));
   NAND2_X1 i_257_76_17460 (.A1(n_257_892), .A2(n_257_445), .ZN(n_257_76_17429));
   NAND2_X1 i_257_76_17461 (.A1(n_257_450), .A2(n_257_76_17413), .ZN(
      n_257_76_17430));
   INV_X1 i_257_76_17462 (.A(n_257_76_17430), .ZN(n_257_76_17431));
   NAND2_X1 i_257_76_17463 (.A1(n_257_732), .A2(n_257_435), .ZN(n_257_76_17432));
   NAND3_X1 i_257_76_17464 (.A1(n_257_76_17431), .A2(n_257_660), .A3(
      n_257_76_17432), .ZN(n_257_76_17433));
   INV_X1 i_257_76_17465 (.A(n_257_76_17433), .ZN(n_257_76_17434));
   NAND2_X1 i_257_76_17466 (.A1(n_257_440), .A2(n_257_962), .ZN(n_257_76_17435));
   NAND2_X1 i_257_76_17467 (.A1(n_257_438), .A2(n_257_898), .ZN(n_257_76_17436));
   NAND4_X1 i_257_76_17468 (.A1(n_257_76_17429), .A2(n_257_76_17434), .A3(
      n_257_76_17435), .A4(n_257_76_17436), .ZN(n_257_76_17437));
   INV_X1 i_257_76_17469 (.A(n_257_76_17437), .ZN(n_257_76_17438));
   NAND4_X1 i_257_76_17470 (.A1(n_257_76_17423), .A2(n_257_76_17428), .A3(
      n_257_76_17438), .A4(n_257_76_17399), .ZN(n_257_76_17439));
   INV_X1 i_257_76_17471 (.A(n_257_76_17439), .ZN(n_257_76_17440));
   NAND2_X1 i_257_76_17472 (.A1(n_257_700), .A2(n_257_448), .ZN(n_257_76_17441));
   NAND2_X1 i_257_76_17473 (.A1(n_257_76_17441), .A2(n_257_76_17398), .ZN(
      n_257_76_17442));
   INV_X1 i_257_76_17474 (.A(n_257_76_17442), .ZN(n_257_76_17443));
   NAND3_X1 i_257_76_17475 (.A1(n_257_76_17440), .A2(n_257_76_17443), .A3(
      n_257_76_17408), .ZN(n_257_76_17444));
   INV_X1 i_257_76_17476 (.A(n_257_76_17444), .ZN(n_257_76_17445));
   NAND2_X1 i_257_76_17477 (.A1(n_257_28), .A2(n_257_76_17445), .ZN(
      n_257_76_17446));
   NAND3_X1 i_257_76_17478 (.A1(n_257_76_17411), .A2(n_257_76_17418), .A3(
      n_257_76_17446), .ZN(n_257_76_17447));
   NAND2_X1 i_257_76_17479 (.A1(n_257_76_17425), .A2(n_257_76_17429), .ZN(
      n_257_76_17448));
   NAND2_X1 i_257_76_17480 (.A1(n_257_860), .A2(n_257_442), .ZN(n_257_76_17449));
   NOR2_X1 i_257_76_17481 (.A1(n_257_76_17449), .A2(n_257_1090), .ZN(
      n_257_76_17450));
   NAND4_X1 i_257_76_17482 (.A1(n_257_446), .A2(n_257_76_17435), .A3(
      n_257_76_17436), .A4(n_257_76_17450), .ZN(n_257_76_17451));
   NOR2_X1 i_257_76_17483 (.A1(n_257_76_17448), .A2(n_257_76_17451), .ZN(
      n_257_76_17452));
   NAND3_X1 i_257_76_17484 (.A1(n_257_76_17452), .A2(n_257_76_17398), .A3(
      n_257_76_17399), .ZN(n_257_76_17453));
   INV_X1 i_257_76_17485 (.A(n_257_76_17408), .ZN(n_257_76_17454));
   NOR2_X1 i_257_76_17486 (.A1(n_257_76_17453), .A2(n_257_76_17454), .ZN(
      n_257_76_17455));
   NAND2_X1 i_257_76_17487 (.A1(n_257_76_18070), .A2(n_257_76_17455), .ZN(
      n_257_76_17456));
   NAND2_X1 i_257_76_17488 (.A1(n_257_439), .A2(n_257_76_17413), .ZN(
      n_257_76_17457));
   INV_X1 i_257_76_17489 (.A(n_257_76_17457), .ZN(n_257_76_17458));
   NAND3_X1 i_257_76_17490 (.A1(n_257_930), .A2(n_257_76_17458), .A3(
      n_257_76_17435), .ZN(n_257_76_17459));
   INV_X1 i_257_76_17491 (.A(n_257_76_17459), .ZN(n_257_76_17460));
   NAND2_X1 i_257_76_17492 (.A1(n_257_76_17399), .A2(n_257_76_17460), .ZN(
      n_257_76_17461));
   INV_X1 i_257_76_17493 (.A(n_257_76_17461), .ZN(n_257_76_17462));
   NAND2_X1 i_257_76_17494 (.A1(n_257_76_17398), .A2(n_257_76_17462), .ZN(
      n_257_76_17463));
   INV_X1 i_257_76_17495 (.A(n_257_76_17463), .ZN(n_257_76_17464));
   NAND2_X1 i_257_76_17496 (.A1(n_257_76_17464), .A2(n_257_76_17408), .ZN(
      n_257_76_17465));
   INV_X1 i_257_76_17497 (.A(n_257_76_17465), .ZN(n_257_76_17466));
   NAND2_X1 i_257_76_17498 (.A1(n_257_76_18084), .A2(n_257_76_17466), .ZN(
      n_257_76_17467));
   NAND2_X1 i_257_76_17499 (.A1(n_257_183), .A2(n_257_429), .ZN(n_257_76_17468));
   NAND2_X1 i_257_76_17500 (.A1(n_257_106), .A2(n_257_431), .ZN(n_257_76_17469));
   NAND3_X1 i_257_76_17501 (.A1(n_257_76_17468), .A2(n_257_76_17399), .A3(
      n_257_76_17469), .ZN(n_257_76_17470));
   NAND2_X1 i_257_76_17502 (.A1(n_257_263), .A2(n_257_425), .ZN(n_257_76_17471));
   NAND2_X1 i_257_76_17503 (.A1(n_257_532), .A2(n_257_424), .ZN(n_257_76_17472));
   NAND2_X1 i_257_76_17504 (.A1(n_257_66), .A2(n_257_433), .ZN(n_257_76_17473));
   NAND3_X1 i_257_76_17505 (.A1(n_257_76_17472), .A2(n_257_303), .A3(
      n_257_76_17473), .ZN(n_257_76_17474));
   INV_X1 i_257_76_17506 (.A(n_257_76_17474), .ZN(n_257_76_17475));
   INV_X1 i_257_76_17507 (.A(n_257_423), .ZN(n_257_76_17476));
   NOR2_X1 i_257_76_17508 (.A1(n_257_76_17476), .A2(n_257_1090), .ZN(
      n_257_76_17477));
   NAND2_X1 i_257_76_17509 (.A1(n_257_432), .A2(n_257_628), .ZN(n_257_76_17478));
   INV_X1 i_257_76_17510 (.A(n_257_596), .ZN(n_257_76_17479));
   NAND2_X1 i_257_76_17511 (.A1(n_257_76_17479), .A2(n_257_442), .ZN(
      n_257_76_17480));
   OAI21_X1 i_257_76_17512 (.A(n_257_76_17480), .B1(n_257_428), .B2(
      n_257_76_17412), .ZN(n_257_76_17481));
   NAND4_X1 i_257_76_17513 (.A1(n_257_76_17432), .A2(n_257_76_17477), .A3(
      n_257_76_17478), .A4(n_257_76_17481), .ZN(n_257_76_17482));
   INV_X1 i_257_76_17514 (.A(n_257_76_17482), .ZN(n_257_76_17483));
   NAND2_X1 i_257_76_17515 (.A1(n_257_144), .A2(n_257_430), .ZN(n_257_76_17484));
   NAND2_X1 i_257_76_17516 (.A1(n_257_660), .A2(n_257_450), .ZN(n_257_76_17485));
   NAND4_X1 i_257_76_17517 (.A1(n_257_76_17475), .A2(n_257_76_17483), .A3(
      n_257_76_17484), .A4(n_257_76_17485), .ZN(n_257_76_17486));
   INV_X1 i_257_76_17518 (.A(n_257_76_17486), .ZN(n_257_76_17487));
   NAND2_X1 i_257_76_17519 (.A1(n_257_76_17471), .A2(n_257_76_17487), .ZN(
      n_257_76_17488));
   NOR2_X1 i_257_76_17520 (.A1(n_257_76_17470), .A2(n_257_76_17488), .ZN(
      n_257_76_17489));
   NAND3_X1 i_257_76_17521 (.A1(n_257_76_17421), .A2(n_257_76_17424), .A3(
      n_257_76_17425), .ZN(n_257_76_17490));
   INV_X1 i_257_76_17522 (.A(n_257_76_17490), .ZN(n_257_76_17491));
   NAND2_X1 i_257_76_17523 (.A1(n_257_427), .A2(n_257_223), .ZN(n_257_76_17492));
   NAND3_X1 i_257_76_17524 (.A1(n_257_76_17435), .A2(n_257_76_17436), .A3(
      n_257_76_17492), .ZN(n_257_76_17493));
   NAND2_X1 i_257_76_17525 (.A1(n_257_564), .A2(n_257_426), .ZN(n_257_76_17494));
   INV_X1 i_257_76_17526 (.A(n_257_76_17494), .ZN(n_257_76_17495));
   NOR2_X1 i_257_76_17527 (.A1(n_257_76_17493), .A2(n_257_76_17495), .ZN(
      n_257_76_17496));
   NAND2_X1 i_257_76_17528 (.A1(n_257_451), .A2(n_257_483), .ZN(n_257_76_17497));
   NAND3_X1 i_257_76_17529 (.A1(n_257_76_17497), .A2(n_257_76_17426), .A3(
      n_257_76_17429), .ZN(n_257_76_17498));
   INV_X1 i_257_76_17530 (.A(n_257_76_17498), .ZN(n_257_76_17499));
   NAND2_X1 i_257_76_17531 (.A1(n_257_76_17419), .A2(n_257_76_17420), .ZN(
      n_257_76_17500));
   INV_X1 i_257_76_17532 (.A(n_257_76_17500), .ZN(n_257_76_17501));
   NAND4_X1 i_257_76_17533 (.A1(n_257_76_17491), .A2(n_257_76_17496), .A3(
      n_257_76_17499), .A4(n_257_76_17501), .ZN(n_257_76_17502));
   INV_X1 i_257_76_17534 (.A(n_257_76_17502), .ZN(n_257_76_17503));
   NAND4_X1 i_257_76_17535 (.A1(n_257_76_17443), .A2(n_257_76_17489), .A3(
      n_257_76_17503), .A4(n_257_76_17408), .ZN(n_257_76_17504));
   INV_X1 i_257_76_17536 (.A(n_257_76_17504), .ZN(n_257_76_17505));
   NAND2_X1 i_257_76_17537 (.A1(n_257_76_18066), .A2(n_257_76_17505), .ZN(
      n_257_76_17506));
   NAND3_X1 i_257_76_17538 (.A1(n_257_76_17456), .A2(n_257_76_17467), .A3(
      n_257_76_17506), .ZN(n_257_76_17507));
   NOR2_X1 i_257_76_17539 (.A1(n_257_76_17447), .A2(n_257_76_17507), .ZN(
      n_257_76_17508));
   NAND2_X1 i_257_76_17540 (.A1(n_257_994), .A2(n_257_76_17413), .ZN(
      n_257_76_17509));
   INV_X1 i_257_76_17541 (.A(n_257_76_17509), .ZN(n_257_76_17510));
   NAND2_X1 i_257_76_17542 (.A1(n_257_441), .A2(n_257_76_17510), .ZN(
      n_257_76_17511));
   INV_X1 i_257_76_17543 (.A(n_257_76_17511), .ZN(n_257_76_17512));
   NAND2_X1 i_257_76_17544 (.A1(n_257_76_17398), .A2(n_257_76_17512), .ZN(
      n_257_76_17513));
   INV_X1 i_257_76_17545 (.A(n_257_76_17513), .ZN(n_257_76_17514));
   NAND2_X1 i_257_76_17546 (.A1(n_257_76_17514), .A2(n_257_76_17408), .ZN(
      n_257_76_17515));
   INV_X1 i_257_76_17547 (.A(n_257_76_17515), .ZN(n_257_76_17516));
   NAND2_X1 i_257_76_17548 (.A1(n_257_76_18071), .A2(n_257_76_17516), .ZN(
      n_257_76_17517));
   NAND3_X1 i_257_76_17549 (.A1(n_257_76_17413), .A2(n_257_732), .A3(n_257_435), 
      .ZN(n_257_76_17518));
   INV_X1 i_257_76_17550 (.A(n_257_76_17518), .ZN(n_257_76_17519));
   NAND4_X1 i_257_76_17551 (.A1(n_257_76_17429), .A2(n_257_76_17435), .A3(
      n_257_76_17436), .A4(n_257_76_17519), .ZN(n_257_76_17520));
   NOR2_X1 i_257_76_17552 (.A1(n_257_76_17427), .A2(n_257_76_17520), .ZN(
      n_257_76_17521));
   INV_X1 i_257_76_17553 (.A(n_257_76_17399), .ZN(n_257_76_17522));
   NOR2_X1 i_257_76_17554 (.A1(n_257_76_17522), .A2(n_257_76_17500), .ZN(
      n_257_76_17523));
   NAND3_X1 i_257_76_17555 (.A1(n_257_76_17521), .A2(n_257_76_17398), .A3(
      n_257_76_17523), .ZN(n_257_76_17524));
   NOR2_X1 i_257_76_17556 (.A1(n_257_76_17524), .A2(n_257_76_17454), .ZN(
      n_257_76_17525));
   NAND2_X1 i_257_76_17557 (.A1(n_257_76_18078), .A2(n_257_76_17525), .ZN(
      n_257_76_17526));
   NAND4_X1 i_257_76_17558 (.A1(n_257_76_17419), .A2(n_257_76_17420), .A3(
      n_257_76_17421), .A4(n_257_76_17424), .ZN(n_257_76_17527));
   NOR2_X1 i_257_76_17559 (.A1(n_257_76_17470), .A2(n_257_76_17527), .ZN(
      n_257_76_17528));
   NAND4_X1 i_257_76_17560 (.A1(n_257_76_17425), .A2(n_257_76_17497), .A3(
      n_257_76_17426), .A4(n_257_76_17429), .ZN(n_257_76_17529));
   NAND2_X1 i_257_76_17561 (.A1(n_257_596), .A2(n_257_442), .ZN(n_257_76_17530));
   INV_X1 i_257_76_17562 (.A(n_257_76_17530), .ZN(n_257_76_17531));
   NAND2_X1 i_257_76_17563 (.A1(n_257_428), .A2(n_257_76_17531), .ZN(
      n_257_76_17532));
   NOR2_X1 i_257_76_17564 (.A1(n_257_76_17532), .A2(n_257_1090), .ZN(
      n_257_76_17533));
   NAND4_X1 i_257_76_17565 (.A1(n_257_76_17473), .A2(n_257_76_17533), .A3(
      n_257_76_17432), .A4(n_257_76_17478), .ZN(n_257_76_17534));
   INV_X1 i_257_76_17566 (.A(n_257_76_17485), .ZN(n_257_76_17535));
   NOR2_X1 i_257_76_17567 (.A1(n_257_76_17534), .A2(n_257_76_17535), .ZN(
      n_257_76_17536));
   NAND2_X1 i_257_76_17568 (.A1(n_257_76_17436), .A2(n_257_76_17484), .ZN(
      n_257_76_17537));
   INV_X1 i_257_76_17569 (.A(n_257_76_17537), .ZN(n_257_76_17538));
   NAND3_X1 i_257_76_17570 (.A1(n_257_76_17536), .A2(n_257_76_17538), .A3(
      n_257_76_17435), .ZN(n_257_76_17539));
   NOR2_X1 i_257_76_17571 (.A1(n_257_76_17529), .A2(n_257_76_17539), .ZN(
      n_257_76_17540));
   NAND4_X1 i_257_76_17572 (.A1(n_257_76_17443), .A2(n_257_76_17528), .A3(
      n_257_76_17408), .A4(n_257_76_17540), .ZN(n_257_76_17541));
   INV_X1 i_257_76_17573 (.A(n_257_76_17541), .ZN(n_257_76_17542));
   NAND2_X1 i_257_76_17574 (.A1(n_257_76_18074), .A2(n_257_76_17542), .ZN(
      n_257_76_17543));
   NAND3_X1 i_257_76_17575 (.A1(n_257_76_17517), .A2(n_257_76_17526), .A3(
      n_257_76_17543), .ZN(n_257_76_17544));
   NAND2_X1 i_257_76_17576 (.A1(n_257_1090), .A2(n_257_442), .ZN(n_257_76_17545));
   INV_X1 i_257_76_17577 (.A(n_257_76_17545), .ZN(n_257_76_17546));
   NAND2_X1 i_257_76_17578 (.A1(n_257_13), .A2(n_257_76_17546), .ZN(
      n_257_76_17547));
   NAND2_X1 i_257_76_17579 (.A1(n_257_76_17435), .A2(n_257_76_17436), .ZN(
      n_257_76_17548));
   INV_X1 i_257_76_17580 (.A(n_257_76_17548), .ZN(n_257_76_17549));
   NAND2_X1 i_257_76_17581 (.A1(n_257_445), .A2(n_257_76_17413), .ZN(
      n_257_76_17550));
   INV_X1 i_257_76_17582 (.A(n_257_76_17550), .ZN(n_257_76_17551));
   NAND2_X1 i_257_76_17583 (.A1(n_257_892), .A2(n_257_76_17551), .ZN(
      n_257_76_17552));
   INV_X1 i_257_76_17584 (.A(n_257_76_17552), .ZN(n_257_76_17553));
   NAND3_X1 i_257_76_17585 (.A1(n_257_76_17549), .A2(n_257_76_17425), .A3(
      n_257_76_17553), .ZN(n_257_76_17554));
   NOR2_X1 i_257_76_17586 (.A1(n_257_76_17554), .A2(n_257_76_17522), .ZN(
      n_257_76_17555));
   NAND2_X1 i_257_76_17587 (.A1(n_257_76_17398), .A2(n_257_76_17555), .ZN(
      n_257_76_17556));
   NOR2_X1 i_257_76_17588 (.A1(n_257_76_17556), .A2(n_257_76_17454), .ZN(
      n_257_76_17557));
   NAND2_X1 i_257_76_17589 (.A1(n_257_76_18077), .A2(n_257_76_17557), .ZN(
      n_257_76_17558));
   NAND2_X1 i_257_76_17590 (.A1(n_257_76_17547), .A2(n_257_76_17558), .ZN(
      n_257_76_17559));
   NOR2_X1 i_257_76_17591 (.A1(n_257_76_17544), .A2(n_257_76_17559), .ZN(
      n_257_76_17560));
   NAND4_X1 i_257_76_17592 (.A1(n_257_76_17435), .A2(n_257_76_17436), .A3(
      n_257_76_17484), .A4(n_257_564), .ZN(n_257_76_17561));
   NAND2_X1 i_257_76_17593 (.A1(n_257_76_17473), .A2(n_257_76_17432), .ZN(
      n_257_76_17562));
   INV_X1 i_257_76_17594 (.A(n_257_76_17562), .ZN(n_257_76_17563));
   INV_X1 i_257_76_17595 (.A(n_257_426), .ZN(n_257_76_17564));
   NOR2_X1 i_257_76_17596 (.A1(n_257_1090), .A2(n_257_76_17564), .ZN(
      n_257_76_17565));
   NAND3_X1 i_257_76_17597 (.A1(n_257_76_17478), .A2(n_257_76_17565), .A3(
      n_257_76_17481), .ZN(n_257_76_17566));
   INV_X1 i_257_76_17598 (.A(n_257_76_17566), .ZN(n_257_76_17567));
   NAND4_X1 i_257_76_17599 (.A1(n_257_76_17485), .A2(n_257_76_17563), .A3(
      n_257_76_17567), .A4(n_257_76_17492), .ZN(n_257_76_17568));
   NOR2_X1 i_257_76_17600 (.A1(n_257_76_17561), .A2(n_257_76_17568), .ZN(
      n_257_76_17569));
   NAND2_X1 i_257_76_17601 (.A1(n_257_76_17469), .A2(n_257_76_17419), .ZN(
      n_257_76_17570));
   INV_X1 i_257_76_17602 (.A(n_257_76_17570), .ZN(n_257_76_17571));
   NAND3_X1 i_257_76_17603 (.A1(n_257_76_17425), .A2(n_257_76_17426), .A3(
      n_257_76_17429), .ZN(n_257_76_17572));
   INV_X1 i_257_76_17604 (.A(n_257_76_17572), .ZN(n_257_76_17573));
   NAND3_X1 i_257_76_17605 (.A1(n_257_76_17569), .A2(n_257_76_17571), .A3(
      n_257_76_17573), .ZN(n_257_76_17574));
   INV_X1 i_257_76_17606 (.A(n_257_76_17574), .ZN(n_257_76_17575));
   NAND2_X1 i_257_76_17607 (.A1(n_257_76_17468), .A2(n_257_76_17399), .ZN(
      n_257_76_17576));
   NAND4_X1 i_257_76_17608 (.A1(n_257_76_17420), .A2(n_257_76_17421), .A3(
      n_257_76_17424), .A4(n_257_76_17497), .ZN(n_257_76_17577));
   NOR2_X1 i_257_76_17609 (.A1(n_257_76_17576), .A2(n_257_76_17577), .ZN(
      n_257_76_17578));
   NAND4_X1 i_257_76_17610 (.A1(n_257_76_17443), .A2(n_257_76_17575), .A3(
      n_257_76_17578), .A4(n_257_76_17408), .ZN(n_257_76_17579));
   INV_X1 i_257_76_17611 (.A(n_257_76_17579), .ZN(n_257_76_17580));
   NAND2_X1 i_257_76_17612 (.A1(n_257_76_18076), .A2(n_257_76_17580), .ZN(
      n_257_76_17581));
   NAND2_X1 i_257_76_17613 (.A1(n_257_436), .A2(n_257_76_17413), .ZN(
      n_257_76_17582));
   INV_X1 i_257_76_17614 (.A(n_257_76_17582), .ZN(n_257_76_17583));
   NAND4_X1 i_257_76_17615 (.A1(n_257_764), .A2(n_257_76_17435), .A3(
      n_257_76_17436), .A4(n_257_76_17583), .ZN(n_257_76_17584));
   NOR2_X1 i_257_76_17616 (.A1(n_257_76_17572), .A2(n_257_76_17584), .ZN(
      n_257_76_17585));
   NAND2_X1 i_257_76_17617 (.A1(n_257_76_17420), .A2(n_257_76_17424), .ZN(
      n_257_76_17586));
   NOR2_X1 i_257_76_17618 (.A1(n_257_76_17522), .A2(n_257_76_17586), .ZN(
      n_257_76_17587));
   NAND3_X1 i_257_76_17619 (.A1(n_257_76_17398), .A2(n_257_76_17585), .A3(
      n_257_76_17587), .ZN(n_257_76_17588));
   NOR2_X1 i_257_76_17620 (.A1(n_257_76_17588), .A2(n_257_76_17454), .ZN(
      n_257_76_17589));
   NAND2_X1 i_257_76_17621 (.A1(n_257_76_18069), .A2(n_257_76_17589), .ZN(
      n_257_76_17590));
   NAND2_X1 i_257_76_17622 (.A1(n_257_76_17421), .A2(n_257_76_17424), .ZN(
      n_257_76_17591));
   INV_X1 i_257_76_17623 (.A(n_257_76_17591), .ZN(n_257_76_17592));
   NAND3_X1 i_257_76_17624 (.A1(n_257_76_17501), .A2(n_257_76_17592), .A3(
      n_257_76_17399), .ZN(n_257_76_17593));
   NAND2_X1 i_257_76_17625 (.A1(n_257_76_17425), .A2(n_257_76_17497), .ZN(
      n_257_76_17594));
   INV_X1 i_257_76_17626 (.A(n_257_76_17594), .ZN(n_257_76_17595));
   NAND2_X1 i_257_76_17627 (.A1(n_257_76_17426), .A2(n_257_76_17429), .ZN(
      n_257_76_17596));
   INV_X1 i_257_76_17628 (.A(n_257_76_17596), .ZN(n_257_76_17597));
   INV_X1 i_257_76_17629 (.A(n_257_1090), .ZN(n_257_76_17598));
   NAND2_X1 i_257_76_17630 (.A1(n_257_628), .A2(n_257_442), .ZN(n_257_76_17599));
   INV_X1 i_257_76_17631 (.A(n_257_76_17599), .ZN(n_257_76_17600));
   NAND3_X1 i_257_76_17632 (.A1(n_257_432), .A2(n_257_76_17598), .A3(
      n_257_76_17600), .ZN(n_257_76_17601));
   INV_X1 i_257_76_17633 (.A(n_257_76_17601), .ZN(n_257_76_17602));
   NAND3_X1 i_257_76_17634 (.A1(n_257_76_17602), .A2(n_257_76_17473), .A3(
      n_257_76_17432), .ZN(n_257_76_17603));
   INV_X1 i_257_76_17635 (.A(n_257_76_17603), .ZN(n_257_76_17604));
   NAND4_X1 i_257_76_17636 (.A1(n_257_76_17604), .A2(n_257_76_17435), .A3(
      n_257_76_17436), .A4(n_257_76_17485), .ZN(n_257_76_17605));
   INV_X1 i_257_76_17637 (.A(n_257_76_17605), .ZN(n_257_76_17606));
   NAND3_X1 i_257_76_17638 (.A1(n_257_76_17595), .A2(n_257_76_17597), .A3(
      n_257_76_17606), .ZN(n_257_76_17607));
   NOR2_X1 i_257_76_17639 (.A1(n_257_76_17593), .A2(n_257_76_17607), .ZN(
      n_257_76_17608));
   NAND3_X1 i_257_76_17640 (.A1(n_257_76_17608), .A2(n_257_76_17443), .A3(
      n_257_76_17408), .ZN(n_257_76_17609));
   INV_X1 i_257_76_17641 (.A(n_257_76_17609), .ZN(n_257_76_17610));
   NAND2_X1 i_257_76_17642 (.A1(n_257_68), .A2(n_257_76_17610), .ZN(
      n_257_76_17611));
   NAND3_X1 i_257_76_17643 (.A1(n_257_76_17581), .A2(n_257_76_17590), .A3(
      n_257_76_17611), .ZN(n_257_76_17612));
   NAND2_X1 i_257_76_17644 (.A1(n_257_437), .A2(n_257_76_17413), .ZN(
      n_257_76_17613));
   INV_X1 i_257_76_17645 (.A(n_257_76_17613), .ZN(n_257_76_17614));
   NAND4_X1 i_257_76_17646 (.A1(n_257_828), .A2(n_257_76_17435), .A3(
      n_257_76_17436), .A4(n_257_76_17614), .ZN(n_257_76_17615));
   NOR2_X1 i_257_76_17647 (.A1(n_257_76_17448), .A2(n_257_76_17615), .ZN(
      n_257_76_17616));
   NAND2_X1 i_257_76_17648 (.A1(n_257_76_17399), .A2(n_257_76_17420), .ZN(
      n_257_76_17617));
   INV_X1 i_257_76_17649 (.A(n_257_76_17617), .ZN(n_257_76_17618));
   NAND3_X1 i_257_76_17650 (.A1(n_257_76_17616), .A2(n_257_76_17398), .A3(
      n_257_76_17618), .ZN(n_257_76_17619));
   NOR2_X1 i_257_76_17651 (.A1(n_257_76_17619), .A2(n_257_76_17454), .ZN(
      n_257_76_17620));
   NAND2_X1 i_257_76_17652 (.A1(n_257_22), .A2(n_257_76_17620), .ZN(
      n_257_76_17621));
   NAND2_X1 i_257_76_17653 (.A1(n_257_444), .A2(n_257_76_17413), .ZN(
      n_257_76_17622));
   INV_X1 i_257_76_17654 (.A(n_257_76_17622), .ZN(n_257_76_17623));
   NAND2_X1 i_257_76_17655 (.A1(n_257_1026), .A2(n_257_76_17623), .ZN(
      n_257_76_17624));
   INV_X1 i_257_76_17656 (.A(n_257_76_17624), .ZN(n_257_76_17625));
   NAND2_X1 i_257_76_17657 (.A1(n_257_76_17408), .A2(n_257_76_17625), .ZN(
      n_257_76_17626));
   INV_X1 i_257_76_17658 (.A(n_257_76_17626), .ZN(n_257_76_17627));
   NAND2_X1 i_257_76_17659 (.A1(n_257_76_18075), .A2(n_257_76_17627), .ZN(
      n_257_76_17628));
   NAND2_X1 i_257_76_17660 (.A1(n_257_76_17621), .A2(n_257_76_17628), .ZN(
      n_257_76_17629));
   NOR2_X1 i_257_76_17661 (.A1(n_257_76_17612), .A2(n_257_76_17629), .ZN(
      n_257_76_17630));
   NAND3_X1 i_257_76_17662 (.A1(n_257_76_17508), .A2(n_257_76_17560), .A3(
      n_257_76_17630), .ZN(n_257_76_17631));
   INV_X1 i_257_76_17663 (.A(n_257_76_17631), .ZN(n_257_76_17632));
   NAND2_X1 i_257_76_17664 (.A1(n_257_433), .A2(n_257_442), .ZN(n_257_76_17633));
   NOR2_X1 i_257_76_17665 (.A1(n_257_76_17633), .A2(n_257_1090), .ZN(
      n_257_76_17634));
   NAND3_X1 i_257_76_17666 (.A1(n_257_76_17634), .A2(n_257_76_17432), .A3(
      n_257_66), .ZN(n_257_76_17635));
   INV_X1 i_257_76_17667 (.A(n_257_76_17635), .ZN(n_257_76_17636));
   NAND4_X1 i_257_76_17668 (.A1(n_257_76_17435), .A2(n_257_76_17436), .A3(
      n_257_76_17636), .A4(n_257_76_17485), .ZN(n_257_76_17637));
   INV_X1 i_257_76_17669 (.A(n_257_76_17637), .ZN(n_257_76_17638));
   NAND3_X1 i_257_76_17670 (.A1(n_257_76_17595), .A2(n_257_76_17597), .A3(
      n_257_76_17638), .ZN(n_257_76_17639));
   NOR2_X1 i_257_76_17671 (.A1(n_257_76_17593), .A2(n_257_76_17639), .ZN(
      n_257_76_17640));
   NAND3_X1 i_257_76_17672 (.A1(n_257_76_17640), .A2(n_257_76_17443), .A3(
      n_257_76_17408), .ZN(n_257_76_17641));
   INV_X1 i_257_76_17673 (.A(n_257_76_17641), .ZN(n_257_76_17642));
   NAND2_X1 i_257_76_17674 (.A1(n_257_76_18081), .A2(n_257_76_17642), .ZN(
      n_257_76_17643));
   NAND3_X1 i_257_76_17675 (.A1(n_257_76_17419), .A2(n_257_76_17420), .A3(
      n_257_76_17424), .ZN(n_257_76_17644));
   INV_X1 i_257_76_17676 (.A(n_257_76_17644), .ZN(n_257_76_17645));
   NAND2_X1 i_257_76_17677 (.A1(n_257_442), .A2(n_257_668), .ZN(n_257_76_17646));
   NOR2_X1 i_257_76_17678 (.A1(n_257_1090), .A2(n_257_76_17646), .ZN(
      n_257_76_17647));
   NAND2_X1 i_257_76_17679 (.A1(n_257_76_17432), .A2(n_257_76_17647), .ZN(
      n_257_76_17648));
   INV_X1 i_257_76_17680 (.A(n_257_76_17648), .ZN(n_257_76_17649));
   NAND4_X1 i_257_76_17681 (.A1(n_257_449), .A2(n_257_76_17435), .A3(
      n_257_76_17436), .A4(n_257_76_17649), .ZN(n_257_76_17650));
   INV_X1 i_257_76_17682 (.A(n_257_76_17650), .ZN(n_257_76_17651));
   NAND4_X1 i_257_76_17683 (.A1(n_257_76_17645), .A2(n_257_76_17573), .A3(
      n_257_76_17399), .A4(n_257_76_17651), .ZN(n_257_76_17652));
   INV_X1 i_257_76_17684 (.A(n_257_76_17652), .ZN(n_257_76_17653));
   NAND3_X1 i_257_76_17685 (.A1(n_257_76_17653), .A2(n_257_76_17443), .A3(
      n_257_76_17408), .ZN(n_257_76_17654));
   INV_X1 i_257_76_17686 (.A(n_257_76_17654), .ZN(n_257_76_17655));
   NAND2_X1 i_257_76_17687 (.A1(n_257_76_18083), .A2(n_257_76_17655), .ZN(
      n_257_76_17656));
   NAND3_X1 i_257_76_17688 (.A1(n_257_76_17424), .A2(n_257_76_17425), .A3(
      n_257_76_17497), .ZN(n_257_76_17657));
   NOR2_X1 i_257_76_17689 (.A1(n_257_76_17422), .A2(n_257_76_17657), .ZN(
      n_257_76_17658));
   NAND3_X1 i_257_76_17690 (.A1(n_257_76_17426), .A2(n_257_76_17429), .A3(
      n_257_76_17435), .ZN(n_257_76_17659));
   NAND2_X1 i_257_76_17691 (.A1(n_257_429), .A2(n_257_442), .ZN(n_257_76_17660));
   NOR2_X1 i_257_76_17692 (.A1(n_257_76_17660), .A2(n_257_1090), .ZN(
      n_257_76_17661));
   NAND4_X1 i_257_76_17693 (.A1(n_257_76_17473), .A2(n_257_76_17661), .A3(
      n_257_76_17432), .A4(n_257_76_17478), .ZN(n_257_76_17662));
   INV_X1 i_257_76_17694 (.A(n_257_76_17662), .ZN(n_257_76_17663));
   NAND4_X1 i_257_76_17695 (.A1(n_257_76_17663), .A2(n_257_76_17436), .A3(
      n_257_76_17484), .A4(n_257_76_17485), .ZN(n_257_76_17664));
   NOR2_X1 i_257_76_17696 (.A1(n_257_76_17659), .A2(n_257_76_17664), .ZN(
      n_257_76_17665));
   NAND3_X1 i_257_76_17697 (.A1(n_257_76_17399), .A2(n_257_76_17469), .A3(
      n_257_183), .ZN(n_257_76_17666));
   INV_X1 i_257_76_17698 (.A(n_257_76_17666), .ZN(n_257_76_17667));
   NAND4_X1 i_257_76_17699 (.A1(n_257_76_17658), .A2(n_257_76_17665), .A3(
      n_257_76_17667), .A4(n_257_76_17398), .ZN(n_257_76_17668));
   NAND2_X1 i_257_76_17700 (.A1(n_257_76_17408), .A2(n_257_76_17441), .ZN(
      n_257_76_17669));
   NOR2_X1 i_257_76_17701 (.A1(n_257_76_17668), .A2(n_257_76_17669), .ZN(
      n_257_76_17670));
   NAND2_X1 i_257_76_17702 (.A1(n_257_76_18061), .A2(n_257_76_17670), .ZN(
      n_257_76_17671));
   NAND3_X1 i_257_76_17703 (.A1(n_257_76_17643), .A2(n_257_76_17656), .A3(
      n_257_76_17671), .ZN(n_257_76_17672));
   INV_X1 i_257_76_17704 (.A(n_257_76_17672), .ZN(n_257_76_17673));
   INV_X1 i_257_76_17705 (.A(n_257_76_17435), .ZN(n_257_76_17674));
   NAND2_X1 i_257_76_17706 (.A1(n_257_442), .A2(n_257_898), .ZN(n_257_76_17675));
   NOR2_X1 i_257_76_17707 (.A1(n_257_1090), .A2(n_257_76_17675), .ZN(
      n_257_76_17676));
   NAND2_X1 i_257_76_17708 (.A1(n_257_438), .A2(n_257_76_17676), .ZN(
      n_257_76_17677));
   NOR2_X1 i_257_76_17709 (.A1(n_257_76_17674), .A2(n_257_76_17677), .ZN(
      n_257_76_17678));
   NAND3_X1 i_257_76_17710 (.A1(n_257_76_17399), .A2(n_257_76_17678), .A3(
      n_257_76_17425), .ZN(n_257_76_17679));
   INV_X1 i_257_76_17711 (.A(n_257_76_17679), .ZN(n_257_76_17680));
   NAND2_X1 i_257_76_17712 (.A1(n_257_76_17680), .A2(n_257_76_17398), .ZN(
      n_257_76_17681));
   NOR2_X1 i_257_76_17713 (.A1(n_257_76_17454), .A2(n_257_76_17681), .ZN(
      n_257_76_17682));
   NAND2_X1 i_257_76_17714 (.A1(n_257_76_18067), .A2(n_257_76_17682), .ZN(
      n_257_76_17683));
   NAND2_X1 i_257_76_17715 (.A1(n_257_76_17472), .A2(n_257_76_17473), .ZN(
      n_257_76_17684));
   INV_X1 i_257_76_17716 (.A(n_257_76_17492), .ZN(n_257_76_17685));
   NOR2_X1 i_257_76_17717 (.A1(n_257_76_17684), .A2(n_257_76_17685), .ZN(
      n_257_76_17686));
   NAND2_X1 i_257_76_17718 (.A1(n_257_341), .A2(n_257_422), .ZN(n_257_76_17687));
   NAND2_X1 i_257_76_17719 (.A1(n_257_442), .A2(n_257_500), .ZN(n_257_76_17688));
   INV_X1 i_257_76_17720 (.A(n_257_76_17688), .ZN(n_257_76_17689));
   NAND2_X1 i_257_76_17721 (.A1(n_257_76_17689), .A2(n_257_76_17479), .ZN(
      n_257_76_17690));
   OAI21_X1 i_257_76_17722 (.A(n_257_76_17690), .B1(n_257_428), .B2(
      n_257_76_17688), .ZN(n_257_76_17691));
   NAND2_X1 i_257_76_17723 (.A1(n_257_76_17687), .A2(n_257_76_17691), .ZN(
      n_257_76_17692));
   INV_X1 i_257_76_17724 (.A(n_257_76_17692), .ZN(n_257_76_17693));
   INV_X1 i_257_76_17725 (.A(n_257_420), .ZN(n_257_76_17694));
   NOR2_X1 i_257_76_17726 (.A1(n_257_76_17694), .A2(n_257_1090), .ZN(
      n_257_76_17695));
   NAND2_X1 i_257_76_17727 (.A1(n_257_76_17693), .A2(n_257_76_17695), .ZN(
      n_257_76_17696));
   NAND2_X1 i_257_76_17728 (.A1(n_257_76_17432), .A2(n_257_76_17478), .ZN(
      n_257_76_17697));
   NOR2_X1 i_257_76_17729 (.A1(n_257_76_17696), .A2(n_257_76_17697), .ZN(
      n_257_76_17698));
   NAND2_X1 i_257_76_17730 (.A1(n_257_76_17686), .A2(n_257_76_17698), .ZN(
      n_257_76_17699));
   NAND2_X1 i_257_76_17731 (.A1(n_257_303), .A2(n_257_423), .ZN(n_257_76_17700));
   NAND2_X1 i_257_76_17732 (.A1(n_257_76_17485), .A2(n_257_76_17700), .ZN(
      n_257_76_17701));
   INV_X1 i_257_76_17733 (.A(n_257_76_17701), .ZN(n_257_76_17702));
   NAND2_X1 i_257_76_17734 (.A1(n_257_76_17702), .A2(n_257_76_17484), .ZN(
      n_257_76_17703));
   NOR2_X1 i_257_76_17735 (.A1(n_257_76_17699), .A2(n_257_76_17703), .ZN(
      n_257_76_17704));
   NAND2_X1 i_257_76_17736 (.A1(n_257_380), .A2(n_257_421), .ZN(n_257_76_17705));
   NAND2_X1 i_257_76_17737 (.A1(n_257_76_17494), .A2(n_257_76_17705), .ZN(
      n_257_76_17706));
   NOR2_X1 i_257_76_17738 (.A1(n_257_76_17706), .A2(n_257_76_17548), .ZN(
      n_257_76_17707));
   NAND2_X1 i_257_76_17739 (.A1(n_257_76_17704), .A2(n_257_76_17707), .ZN(
      n_257_76_17708));
   NOR2_X1 i_257_76_17740 (.A1(n_257_76_17594), .A2(n_257_76_17596), .ZN(
      n_257_76_17709));
   INV_X1 i_257_76_17741 (.A(n_257_76_17420), .ZN(n_257_76_17710));
   NOR2_X1 i_257_76_17742 (.A1(n_257_76_17591), .A2(n_257_76_17710), .ZN(
      n_257_76_17711));
   NAND2_X1 i_257_76_17743 (.A1(n_257_76_17709), .A2(n_257_76_17711), .ZN(
      n_257_76_17712));
   NOR2_X1 i_257_76_17744 (.A1(n_257_76_17708), .A2(n_257_76_17712), .ZN(
      n_257_76_17713));
   NAND2_X1 i_257_76_17745 (.A1(n_257_76_17571), .A2(n_257_76_17399), .ZN(
      n_257_76_17714));
   NAND2_X1 i_257_76_17746 (.A1(n_257_76_17471), .A2(n_257_76_17468), .ZN(
      n_257_76_17715));
   NOR2_X1 i_257_76_17747 (.A1(n_257_76_17714), .A2(n_257_76_17715), .ZN(
      n_257_76_17716));
   NAND2_X1 i_257_76_17748 (.A1(n_257_76_17713), .A2(n_257_76_17716), .ZN(
      n_257_76_17717));
   NAND2_X1 i_257_76_17749 (.A1(n_257_76_17443), .A2(n_257_76_17408), .ZN(
      n_257_76_17718));
   NOR2_X1 i_257_76_17750 (.A1(n_257_76_17717), .A2(n_257_76_17718), .ZN(
      n_257_76_17719));
   NAND2_X1 i_257_76_17751 (.A1(n_257_76_18073), .A2(n_257_76_17719), .ZN(
      n_257_76_17720));
   NAND2_X1 i_257_76_17752 (.A1(n_257_76_17399), .A2(n_257_76_17469), .ZN(
      n_257_76_17721));
   INV_X1 i_257_76_17753 (.A(n_257_76_17721), .ZN(n_257_76_17722));
   NAND2_X1 i_257_76_17754 (.A1(n_257_430), .A2(n_257_442), .ZN(n_257_76_17723));
   NOR2_X1 i_257_76_17755 (.A1(n_257_76_17723), .A2(n_257_1090), .ZN(
      n_257_76_17724));
   NAND4_X1 i_257_76_17756 (.A1(n_257_76_17473), .A2(n_257_76_17432), .A3(
      n_257_76_17724), .A4(n_257_76_17478), .ZN(n_257_76_17725));
   INV_X1 i_257_76_17757 (.A(n_257_76_17725), .ZN(n_257_76_17726));
   NAND4_X1 i_257_76_17758 (.A1(n_257_76_17726), .A2(n_257_76_17436), .A3(
      n_257_76_17485), .A4(n_257_144), .ZN(n_257_76_17727));
   NOR2_X1 i_257_76_17759 (.A1(n_257_76_17659), .A2(n_257_76_17727), .ZN(
      n_257_76_17728));
   NAND4_X1 i_257_76_17760 (.A1(n_257_76_17658), .A2(n_257_76_17398), .A3(
      n_257_76_17722), .A4(n_257_76_17728), .ZN(n_257_76_17729));
   NOR2_X1 i_257_76_17761 (.A1(n_257_76_17729), .A2(n_257_76_17669), .ZN(
      n_257_76_17730));
   NAND2_X1 i_257_76_17762 (.A1(n_257_76_18068), .A2(n_257_76_17730), .ZN(
      n_257_76_17731));
   NAND3_X1 i_257_76_17763 (.A1(n_257_76_17683), .A2(n_257_76_17720), .A3(
      n_257_76_17731), .ZN(n_257_76_17732));
   INV_X1 i_257_76_17764 (.A(n_257_76_17732), .ZN(n_257_76_17733));
   NAND2_X1 i_257_76_17765 (.A1(n_257_76_17420), .A2(n_257_76_17425), .ZN(
      n_257_76_17734));
   INV_X1 i_257_76_17766 (.A(n_257_76_17734), .ZN(n_257_76_17735));
   NAND2_X1 i_257_76_17767 (.A1(n_257_796), .A2(n_257_442), .ZN(n_257_76_17736));
   NOR2_X1 i_257_76_17768 (.A1(n_257_1090), .A2(n_257_76_17736), .ZN(
      n_257_76_17737));
   NAND4_X1 i_257_76_17769 (.A1(n_257_447), .A2(n_257_76_17435), .A3(
      n_257_76_17436), .A4(n_257_76_17737), .ZN(n_257_76_17738));
   INV_X1 i_257_76_17770 (.A(n_257_76_17738), .ZN(n_257_76_17739));
   NAND4_X1 i_257_76_17771 (.A1(n_257_76_17735), .A2(n_257_76_17739), .A3(
      n_257_76_17597), .A4(n_257_76_17399), .ZN(n_257_76_17740));
   INV_X1 i_257_76_17772 (.A(n_257_76_17740), .ZN(n_257_76_17741));
   NAND3_X1 i_257_76_17773 (.A1(n_257_76_17741), .A2(n_257_76_17408), .A3(
      n_257_76_17398), .ZN(n_257_76_17742));
   INV_X1 i_257_76_17774 (.A(n_257_76_17742), .ZN(n_257_76_17743));
   NOR2_X1 i_257_76_17775 (.A1(n_257_76_17422), .A2(n_257_76_17522), .ZN(
      n_257_76_17744));
   NAND4_X1 i_257_76_17776 (.A1(n_257_76_17424), .A2(n_257_76_17425), .A3(
      n_257_76_17497), .A4(n_257_76_17426), .ZN(n_257_76_17745));
   INV_X1 i_257_76_17777 (.A(n_257_76_17745), .ZN(n_257_76_17746));
   NAND2_X1 i_257_76_17778 (.A1(n_257_431), .A2(n_257_442), .ZN(n_257_76_17747));
   NOR2_X1 i_257_76_17779 (.A1(n_257_76_17747), .A2(n_257_1090), .ZN(
      n_257_76_17748));
   NAND4_X1 i_257_76_17780 (.A1(n_257_76_17473), .A2(n_257_76_17432), .A3(
      n_257_76_17748), .A4(n_257_76_17478), .ZN(n_257_76_17749));
   INV_X1 i_257_76_17781 (.A(n_257_76_17749), .ZN(n_257_76_17750));
   NAND4_X1 i_257_76_17782 (.A1(n_257_76_17750), .A2(n_257_76_17435), .A3(
      n_257_76_17436), .A4(n_257_76_17485), .ZN(n_257_76_17751));
   NAND2_X1 i_257_76_17783 (.A1(n_257_76_17429), .A2(n_257_106), .ZN(
      n_257_76_17752));
   NOR2_X1 i_257_76_17784 (.A1(n_257_76_17751), .A2(n_257_76_17752), .ZN(
      n_257_76_17753));
   NAND4_X1 i_257_76_17785 (.A1(n_257_76_17744), .A2(n_257_76_17398), .A3(
      n_257_76_17746), .A4(n_257_76_17753), .ZN(n_257_76_17754));
   NOR2_X1 i_257_76_17786 (.A1(n_257_76_17754), .A2(n_257_76_17669), .ZN(
      n_257_76_17755));
   AOI22_X1 i_257_76_17787 (.A1(n_257_76_18085), .A2(n_257_76_17743), .B1(
      n_257_76_18080), .B2(n_257_76_17755), .ZN(n_257_76_17756));
   NAND3_X1 i_257_76_17788 (.A1(n_257_76_17673), .A2(n_257_76_17733), .A3(
      n_257_76_17756), .ZN(n_257_76_17757));
   INV_X1 i_257_76_17789 (.A(n_257_732), .ZN(n_257_76_17758));
   NAND2_X1 i_257_76_17790 (.A1(n_257_76_17758), .A2(n_257_442), .ZN(
      n_257_76_17759));
   INV_X1 i_257_76_17791 (.A(n_257_435), .ZN(n_257_76_17760));
   NAND2_X1 i_257_76_17792 (.A1(n_257_76_17760), .A2(n_257_442), .ZN(
      n_257_76_17761));
   AOI21_X1 i_257_76_17793 (.A(n_257_1090), .B1(n_257_76_17759), .B2(
      n_257_76_17761), .ZN(n_257_76_17762));
   NAND4_X1 i_257_76_17794 (.A1(n_257_76_17762), .A2(n_257_76_17435), .A3(
      n_257_76_17436), .A4(n_257_448), .ZN(n_257_76_17763));
   INV_X1 i_257_76_17795 (.A(n_257_76_17763), .ZN(n_257_76_17764));
   NAND4_X1 i_257_76_17796 (.A1(n_257_76_17645), .A2(n_257_76_17573), .A3(
      n_257_76_17399), .A4(n_257_76_17764), .ZN(n_257_76_17765));
   INV_X1 i_257_76_17797 (.A(n_257_76_17765), .ZN(n_257_76_17766));
   NAND2_X1 i_257_76_17798 (.A1(n_257_76_17398), .A2(n_257_700), .ZN(
      n_257_76_17767));
   INV_X1 i_257_76_17799 (.A(n_257_76_17767), .ZN(n_257_76_17768));
   NAND3_X1 i_257_76_17800 (.A1(n_257_76_17766), .A2(n_257_76_17768), .A3(
      n_257_76_17408), .ZN(n_257_76_17769));
   INV_X1 i_257_76_17801 (.A(n_257_76_17769), .ZN(n_257_76_17770));
   NAND2_X1 i_257_76_17802 (.A1(n_257_76_18079), .A2(n_257_76_17770), .ZN(
      n_257_76_17771));
   NAND2_X1 i_257_76_17803 (.A1(n_257_76_17398), .A2(n_257_76_17399), .ZN(
      n_257_76_17772));
   INV_X1 i_257_76_17804 (.A(n_257_76_17772), .ZN(n_257_76_17773));
   NAND3_X1 i_257_76_17805 (.A1(n_257_76_17773), .A2(n_257_76_17408), .A3(
      n_257_76_17441), .ZN(n_257_76_17774));
   INV_X1 i_257_76_17806 (.A(n_257_76_17468), .ZN(n_257_76_17775));
   NAND2_X1 i_257_76_17807 (.A1(n_257_76_17469), .A2(n_257_263), .ZN(
      n_257_76_17776));
   NOR2_X1 i_257_76_17808 (.A1(n_257_76_17775), .A2(n_257_76_17776), .ZN(
      n_257_76_17777));
   INV_X1 i_257_76_17809 (.A(n_257_425), .ZN(n_257_76_17778));
   NOR2_X1 i_257_76_17810 (.A1(n_257_76_17778), .A2(n_257_1090), .ZN(
      n_257_76_17779));
   NAND3_X1 i_257_76_17811 (.A1(n_257_76_17478), .A2(n_257_76_17779), .A3(
      n_257_76_17481), .ZN(n_257_76_17780));
   INV_X1 i_257_76_17812 (.A(n_257_76_17780), .ZN(n_257_76_17781));
   NAND3_X1 i_257_76_17813 (.A1(n_257_76_17781), .A2(n_257_76_17563), .A3(
      n_257_76_17492), .ZN(n_257_76_17782));
   INV_X1 i_257_76_17814 (.A(n_257_76_17782), .ZN(n_257_76_17783));
   NAND2_X1 i_257_76_17815 (.A1(n_257_76_17484), .A2(n_257_76_17485), .ZN(
      n_257_76_17784));
   INV_X1 i_257_76_17816 (.A(n_257_76_17784), .ZN(n_257_76_17785));
   NAND3_X1 i_257_76_17817 (.A1(n_257_76_17549), .A2(n_257_76_17783), .A3(
      n_257_76_17785), .ZN(n_257_76_17786));
   NAND3_X1 i_257_76_17818 (.A1(n_257_76_17426), .A2(n_257_76_17429), .A3(
      n_257_76_17494), .ZN(n_257_76_17787));
   NOR2_X1 i_257_76_17819 (.A1(n_257_76_17786), .A2(n_257_76_17787), .ZN(
      n_257_76_17788));
   NAND3_X1 i_257_76_17820 (.A1(n_257_76_17777), .A2(n_257_76_17658), .A3(
      n_257_76_17788), .ZN(n_257_76_17789));
   NOR2_X1 i_257_76_17821 (.A1(n_257_76_17774), .A2(n_257_76_17789), .ZN(
      n_257_76_17790));
   NAND2_X1 i_257_76_17822 (.A1(n_257_76_18064), .A2(n_257_76_17790), .ZN(
      n_257_76_17791));
   INV_X1 i_257_76_17823 (.A(n_257_421), .ZN(n_257_76_17792));
   NOR2_X1 i_257_76_17824 (.A1(n_257_76_17792), .A2(n_257_1090), .ZN(
      n_257_76_17793));
   NAND3_X1 i_257_76_17825 (.A1(n_257_76_17793), .A2(n_257_76_17687), .A3(
      n_257_76_17481), .ZN(n_257_76_17794));
   NOR2_X1 i_257_76_17826 (.A1(n_257_76_17794), .A2(n_257_76_17697), .ZN(
      n_257_76_17795));
   INV_X1 i_257_76_17827 (.A(n_257_76_17684), .ZN(n_257_76_17796));
   NAND4_X1 i_257_76_17828 (.A1(n_257_76_17795), .A2(n_257_76_17796), .A3(
      n_257_76_17492), .A4(n_257_380), .ZN(n_257_76_17797));
   NAND4_X1 i_257_76_17829 (.A1(n_257_76_17436), .A2(n_257_76_17484), .A3(
      n_257_76_17485), .A4(n_257_76_17700), .ZN(n_257_76_17798));
   NOR2_X1 i_257_76_17830 (.A1(n_257_76_17797), .A2(n_257_76_17798), .ZN(
      n_257_76_17799));
   NAND3_X1 i_257_76_17831 (.A1(n_257_76_17469), .A2(n_257_76_17419), .A3(
      n_257_76_17425), .ZN(n_257_76_17800));
   INV_X1 i_257_76_17832 (.A(n_257_76_17800), .ZN(n_257_76_17801));
   NAND4_X1 i_257_76_17833 (.A1(n_257_76_17426), .A2(n_257_76_17429), .A3(
      n_257_76_17494), .A4(n_257_76_17435), .ZN(n_257_76_17802));
   INV_X1 i_257_76_17834 (.A(n_257_76_17802), .ZN(n_257_76_17803));
   NAND3_X1 i_257_76_17835 (.A1(n_257_76_17799), .A2(n_257_76_17801), .A3(
      n_257_76_17803), .ZN(n_257_76_17804));
   INV_X1 i_257_76_17836 (.A(n_257_76_17804), .ZN(n_257_76_17805));
   NAND2_X1 i_257_76_17837 (.A1(n_257_76_17408), .A2(n_257_76_17805), .ZN(
      n_257_76_17806));
   NAND3_X1 i_257_76_17838 (.A1(n_257_76_17471), .A2(n_257_76_17468), .A3(
      n_257_76_17399), .ZN(n_257_76_17807));
   INV_X1 i_257_76_17839 (.A(n_257_76_17807), .ZN(n_257_76_17808));
   INV_X1 i_257_76_17840 (.A(n_257_76_17577), .ZN(n_257_76_17809));
   NAND4_X1 i_257_76_17841 (.A1(n_257_76_17808), .A2(n_257_76_17441), .A3(
      n_257_76_17398), .A4(n_257_76_17809), .ZN(n_257_76_17810));
   NOR2_X1 i_257_76_17842 (.A1(n_257_76_17806), .A2(n_257_76_17810), .ZN(
      n_257_76_17811));
   NAND2_X1 i_257_76_17843 (.A1(n_257_76_18082), .A2(n_257_76_17811), .ZN(
      n_257_76_17812));
   NAND3_X1 i_257_76_17844 (.A1(n_257_76_17771), .A2(n_257_76_17791), .A3(
      n_257_76_17812), .ZN(n_257_76_17813));
   INV_X1 i_257_76_17845 (.A(n_257_76_17813), .ZN(n_257_76_17814));
   NAND3_X1 i_257_76_17846 (.A1(n_257_427), .A2(n_257_76_17473), .A3(
      n_257_76_17432), .ZN(n_257_76_17815));
   INV_X1 i_257_76_17847 (.A(n_257_76_17815), .ZN(n_257_76_17816));
   NAND2_X1 i_257_76_17848 (.A1(n_257_223), .A2(n_257_76_17598), .ZN(
      n_257_76_17817));
   INV_X1 i_257_76_17849 (.A(n_257_76_17817), .ZN(n_257_76_17818));
   NAND3_X1 i_257_76_17850 (.A1(n_257_76_17478), .A2(n_257_76_17818), .A3(
      n_257_76_17481), .ZN(n_257_76_17819));
   INV_X1 i_257_76_17851 (.A(n_257_76_17819), .ZN(n_257_76_17820));
   NAND4_X1 i_257_76_17852 (.A1(n_257_76_17816), .A2(n_257_76_17484), .A3(
      n_257_76_17485), .A4(n_257_76_17820), .ZN(n_257_76_17821));
   INV_X1 i_257_76_17853 (.A(n_257_76_17821), .ZN(n_257_76_17822));
   NAND3_X1 i_257_76_17854 (.A1(n_257_76_17468), .A2(n_257_76_17822), .A3(
      n_257_76_17399), .ZN(n_257_76_17823));
   NAND4_X1 i_257_76_17855 (.A1(n_257_76_17469), .A2(n_257_76_17419), .A3(
      n_257_76_17420), .A4(n_257_76_17421), .ZN(n_257_76_17824));
   NOR2_X1 i_257_76_17856 (.A1(n_257_76_17823), .A2(n_257_76_17824), .ZN(
      n_257_76_17825));
   NAND4_X1 i_257_76_17857 (.A1(n_257_76_17426), .A2(n_257_76_17429), .A3(
      n_257_76_17435), .A4(n_257_76_17436), .ZN(n_257_76_17826));
   NOR2_X1 i_257_76_17858 (.A1(n_257_76_17826), .A2(n_257_76_17657), .ZN(
      n_257_76_17827));
   NAND4_X1 i_257_76_17859 (.A1(n_257_76_17825), .A2(n_257_76_17443), .A3(
      n_257_76_17408), .A4(n_257_76_17827), .ZN(n_257_76_17828));
   INV_X1 i_257_76_17860 (.A(n_257_76_17828), .ZN(n_257_76_17829));
   NAND2_X1 i_257_76_17861 (.A1(n_257_76_18065), .A2(n_257_76_17829), .ZN(
      n_257_76_17830));
   NAND3_X1 i_257_76_17862 (.A1(n_257_76_17762), .A2(n_257_451), .A3(
      n_257_76_17435), .ZN(n_257_76_17831));
   NAND3_X1 i_257_76_17863 (.A1(n_257_76_17436), .A2(n_257_76_17485), .A3(
      n_257_483), .ZN(n_257_76_17832));
   NOR2_X1 i_257_76_17864 (.A1(n_257_76_17831), .A2(n_257_76_17832), .ZN(
      n_257_76_17833));
   NAND2_X1 i_257_76_17865 (.A1(n_257_76_17424), .A2(n_257_76_17425), .ZN(
      n_257_76_17834));
   INV_X1 i_257_76_17866 (.A(n_257_76_17834), .ZN(n_257_76_17835));
   NAND3_X1 i_257_76_17867 (.A1(n_257_76_17833), .A2(n_257_76_17835), .A3(
      n_257_76_17597), .ZN(n_257_76_17836));
   INV_X1 i_257_76_17868 (.A(n_257_76_17836), .ZN(n_257_76_17837));
   NAND4_X1 i_257_76_17869 (.A1(n_257_76_17399), .A2(n_257_76_17419), .A3(
      n_257_76_17420), .A4(n_257_76_17421), .ZN(n_257_76_17838));
   INV_X1 i_257_76_17870 (.A(n_257_76_17838), .ZN(n_257_76_17839));
   NAND2_X1 i_257_76_17871 (.A1(n_257_76_17837), .A2(n_257_76_17839), .ZN(
      n_257_76_17840));
   NOR3_X1 i_257_76_17872 (.A1(n_257_76_17840), .A2(n_257_76_17454), .A3(
      n_257_76_17442), .ZN(n_257_76_17841));
   NAND2_X1 i_257_76_17873 (.A1(n_257_76_18063), .A2(n_257_76_17841), .ZN(
      n_257_76_17842));
   NAND3_X1 i_257_76_17874 (.A1(n_257_76_17473), .A2(n_257_76_17432), .A3(
      n_257_76_17478), .ZN(n_257_76_17843));
   INV_X1 i_257_76_17875 (.A(n_257_76_17843), .ZN(n_257_76_17844));
   NAND2_X1 i_257_76_17876 (.A1(n_257_76_17598), .A2(n_257_424), .ZN(
      n_257_76_17845));
   INV_X1 i_257_76_17877 (.A(n_257_76_17845), .ZN(n_257_76_17846));
   NAND3_X1 i_257_76_17878 (.A1(n_257_532), .A2(n_257_76_17846), .A3(
      n_257_76_17481), .ZN(n_257_76_17847));
   INV_X1 i_257_76_17879 (.A(n_257_76_17847), .ZN(n_257_76_17848));
   NAND4_X1 i_257_76_17880 (.A1(n_257_76_17484), .A2(n_257_76_17844), .A3(
      n_257_76_17485), .A4(n_257_76_17848), .ZN(n_257_76_17849));
   INV_X1 i_257_76_17881 (.A(n_257_76_17849), .ZN(n_257_76_17850));
   NAND3_X1 i_257_76_17882 (.A1(n_257_76_17850), .A2(n_257_76_17399), .A3(
      n_257_76_17469), .ZN(n_257_76_17851));
   NOR2_X1 i_257_76_17883 (.A1(n_257_76_17851), .A2(n_257_76_17715), .ZN(
      n_257_76_17852));
   NAND4_X1 i_257_76_17884 (.A1(n_257_76_17443), .A2(n_257_76_17503), .A3(
      n_257_76_17852), .A4(n_257_76_17408), .ZN(n_257_76_17853));
   INV_X1 i_257_76_17885 (.A(n_257_76_17853), .ZN(n_257_76_17854));
   NAND2_X1 i_257_76_17886 (.A1(n_257_76_18062), .A2(n_257_76_17854), .ZN(
      n_257_76_17855));
   NAND3_X1 i_257_76_17887 (.A1(n_257_76_17830), .A2(n_257_76_17842), .A3(
      n_257_76_17855), .ZN(n_257_76_17856));
   INV_X1 i_257_76_17888 (.A(n_257_76_17856), .ZN(n_257_76_17857));
   NAND2_X1 i_257_76_17889 (.A1(n_257_76_17481), .A2(n_257_341), .ZN(
      n_257_76_17858));
   INV_X1 i_257_76_17890 (.A(n_257_76_17858), .ZN(n_257_76_17859));
   NAND2_X1 i_257_76_17891 (.A1(n_257_422), .A2(n_257_76_17598), .ZN(
      n_257_76_17860));
   INV_X1 i_257_76_17892 (.A(n_257_76_17860), .ZN(n_257_76_17861));
   NAND2_X1 i_257_76_17893 (.A1(n_257_76_17859), .A2(n_257_76_17861), .ZN(
      n_257_76_17862));
   NOR2_X1 i_257_76_17894 (.A1(n_257_76_17862), .A2(n_257_76_17697), .ZN(
      n_257_76_17863));
   NAND2_X1 i_257_76_17895 (.A1(n_257_76_17686), .A2(n_257_76_17863), .ZN(
      n_257_76_17864));
   NOR2_X1 i_257_76_17896 (.A1(n_257_76_17864), .A2(n_257_76_17703), .ZN(
      n_257_76_17865));
   NAND2_X1 i_257_76_17897 (.A1(n_257_76_17429), .A2(n_257_76_17494), .ZN(
      n_257_76_17866));
   NOR2_X1 i_257_76_17898 (.A1(n_257_76_17866), .A2(n_257_76_17548), .ZN(
      n_257_76_17867));
   NAND2_X1 i_257_76_17899 (.A1(n_257_76_17865), .A2(n_257_76_17867), .ZN(
      n_257_76_17868));
   NAND2_X1 i_257_76_17900 (.A1(n_257_76_17497), .A2(n_257_76_17426), .ZN(
      n_257_76_17869));
   INV_X1 i_257_76_17901 (.A(n_257_76_17425), .ZN(n_257_76_17870));
   NOR2_X1 i_257_76_17902 (.A1(n_257_76_17869), .A2(n_257_76_17870), .ZN(
      n_257_76_17871));
   NAND2_X1 i_257_76_17903 (.A1(n_257_76_17711), .A2(n_257_76_17871), .ZN(
      n_257_76_17872));
   NOR2_X1 i_257_76_17904 (.A1(n_257_76_17868), .A2(n_257_76_17872), .ZN(
      n_257_76_17873));
   NAND2_X1 i_257_76_17905 (.A1(n_257_76_17873), .A2(n_257_76_17716), .ZN(
      n_257_76_17874));
   NOR2_X1 i_257_76_17906 (.A1(n_257_76_17874), .A2(n_257_76_17718), .ZN(
      n_257_76_17875));
   NAND2_X1 i_257_76_17907 (.A1(n_257_342), .A2(n_257_76_17875), .ZN(
      n_257_76_17876));
   NAND3_X1 i_257_76_17908 (.A1(n_257_76_17420), .A2(n_257_76_17421), .A3(
      n_257_76_17424), .ZN(n_257_76_17877));
   NOR2_X1 i_257_76_17909 (.A1(n_257_76_17877), .A2(n_257_76_17570), .ZN(
      n_257_76_17878));
   NOR2_X1 i_257_76_17910 (.A1(n_257_76_17787), .A2(n_257_76_17594), .ZN(
      n_257_76_17879));
   NAND4_X1 i_257_76_17911 (.A1(n_257_76_17808), .A2(n_257_76_17878), .A3(
      n_257_76_17398), .A4(n_257_76_17879), .ZN(n_257_76_17880));
   NAND2_X1 i_257_76_17912 (.A1(n_257_442), .A2(n_257_419), .ZN(n_257_76_17881));
   INV_X1 i_257_76_17913 (.A(n_257_76_17881), .ZN(n_257_76_17882));
   NAND2_X1 i_257_76_17914 (.A1(n_257_484), .A2(n_257_76_17882), .ZN(
      n_257_76_17883));
   NOR2_X1 i_257_76_17915 (.A1(n_257_1090), .A2(n_257_76_17883), .ZN(
      n_257_76_17884));
   NAND2_X1 i_257_76_17916 (.A1(n_257_420), .A2(n_257_500), .ZN(n_257_76_17885));
   NAND2_X1 i_257_76_17917 (.A1(n_257_428), .A2(n_257_596), .ZN(n_257_76_17886));
   NAND4_X1 i_257_76_17918 (.A1(n_257_76_17884), .A2(n_257_76_17687), .A3(
      n_257_76_17885), .A4(n_257_76_17886), .ZN(n_257_76_17887));
   NOR2_X1 i_257_76_17919 (.A1(n_257_76_17843), .A2(n_257_76_17887), .ZN(
      n_257_76_17888));
   NAND2_X1 i_257_76_17920 (.A1(n_257_76_17492), .A2(n_257_76_17472), .ZN(
      n_257_76_17889));
   INV_X1 i_257_76_17921 (.A(n_257_76_17889), .ZN(n_257_76_17890));
   NAND3_X1 i_257_76_17922 (.A1(n_257_76_17888), .A2(n_257_76_17702), .A3(
      n_257_76_17890), .ZN(n_257_76_17891));
   NAND4_X1 i_257_76_17923 (.A1(n_257_76_17705), .A2(n_257_76_17435), .A3(
      n_257_76_17436), .A4(n_257_76_17484), .ZN(n_257_76_17892));
   NOR2_X1 i_257_76_17924 (.A1(n_257_76_17891), .A2(n_257_76_17892), .ZN(
      n_257_76_17893));
   NAND3_X1 i_257_76_17925 (.A1(n_257_76_17408), .A2(n_257_76_17893), .A3(
      n_257_76_17441), .ZN(n_257_76_17894));
   NOR2_X1 i_257_76_17926 (.A1(n_257_76_17880), .A2(n_257_76_17894), .ZN(
      n_257_76_17895));
   NAND2_X1 i_257_76_17927 (.A1(n_257_76_18060), .A2(n_257_76_17895), .ZN(
      n_257_76_17896));
   NAND2_X1 i_257_76_17928 (.A1(n_257_994), .A2(n_257_442), .ZN(n_257_76_17897));
   INV_X1 i_257_76_17929 (.A(n_257_76_17897), .ZN(n_257_76_17898));
   NAND2_X1 i_257_76_17930 (.A1(n_257_441), .A2(n_257_76_17898), .ZN(
      n_257_76_17899));
   NAND3_X1 i_257_76_17931 (.A1(n_257_76_17899), .A2(n_257_76_17849), .A3(
      n_257_76_17821), .ZN(n_257_76_17900));
   INV_X1 i_257_76_17932 (.A(n_257_76_17900), .ZN(n_257_76_17901));
   NAND2_X1 i_257_76_17933 (.A1(n_257_445), .A2(n_257_442), .ZN(n_257_76_17902));
   INV_X1 i_257_76_17934 (.A(n_257_76_17902), .ZN(n_257_76_17903));
   NAND2_X1 i_257_76_17935 (.A1(n_257_892), .A2(n_257_76_17903), .ZN(
      n_257_76_17904));
   NAND2_X1 i_257_76_17936 (.A1(n_257_76_17886), .A2(n_257_76_17598), .ZN(
      n_257_76_17905));
   INV_X1 i_257_76_17937 (.A(n_257_76_17905), .ZN(n_257_76_17906));
   INV_X1 i_257_76_17938 (.A(n_257_419), .ZN(n_257_76_17907));
   NAND2_X1 i_257_76_17939 (.A1(n_257_76_17907), .A2(Small_Packet_Data_Size[31]), 
      .ZN(n_257_76_17908));
   INV_X1 i_257_76_17940 (.A(Small_Packet_Data_Size[31]), .ZN(n_257_76_17909));
   OAI21_X1 i_257_76_17941 (.A(n_257_76_17908), .B1(n_257_484), .B2(
      n_257_76_17909), .ZN(n_257_76_17910));
   NAND4_X1 i_257_76_17942 (.A1(n_257_76_17906), .A2(n_257_76_17687), .A3(
      n_257_76_17885), .A4(n_257_76_17910), .ZN(n_257_76_17911));
   NAND2_X1 i_257_76_17943 (.A1(n_257_76_17412), .A2(Small_Packet_Data_Size[31]), 
      .ZN(n_257_76_17912));
   NAND2_X1 i_257_76_17944 (.A1(n_257_76_17911), .A2(n_257_76_17912), .ZN(
      n_257_76_17913));
   INV_X1 i_257_76_17945 (.A(n_257_76_17400), .ZN(n_257_76_17914));
   NAND2_X1 i_257_76_17946 (.A1(n_257_440), .A2(n_257_76_17914), .ZN(
      n_257_76_17915));
   NAND3_X1 i_257_76_17947 (.A1(n_257_76_17904), .A2(n_257_76_17913), .A3(
      n_257_76_17915), .ZN(n_257_76_17916));
   NAND3_X1 i_257_76_17948 (.A1(n_257_732), .A2(n_257_435), .A3(n_257_442), 
      .ZN(n_257_76_17917));
   INV_X1 i_257_76_17949 (.A(n_257_76_17633), .ZN(n_257_76_17918));
   NAND2_X1 i_257_76_17950 (.A1(n_257_66), .A2(n_257_76_17918), .ZN(
      n_257_76_17919));
   NAND2_X1 i_257_76_17951 (.A1(n_257_432), .A2(n_257_76_17600), .ZN(
      n_257_76_17920));
   NAND3_X1 i_257_76_17952 (.A1(n_257_76_17917), .A2(n_257_76_17919), .A3(
      n_257_76_17920), .ZN(n_257_76_17921));
   INV_X1 i_257_76_17953 (.A(n_257_76_17921), .ZN(n_257_76_17922));
   INV_X1 i_257_76_17954 (.A(n_257_76_17675), .ZN(n_257_76_17923));
   NAND2_X1 i_257_76_17955 (.A1(n_257_438), .A2(n_257_76_17923), .ZN(
      n_257_76_17924));
   INV_X1 i_257_76_17956 (.A(n_257_76_17723), .ZN(n_257_76_17925));
   NAND2_X1 i_257_76_17957 (.A1(n_257_144), .A2(n_257_76_17925), .ZN(
      n_257_76_17926));
   NAND2_X1 i_257_76_17958 (.A1(n_257_450), .A2(n_257_442), .ZN(n_257_76_17927));
   INV_X1 i_257_76_17959 (.A(n_257_76_17927), .ZN(n_257_76_17928));
   NAND2_X1 i_257_76_17960 (.A1(n_257_660), .A2(n_257_76_17928), .ZN(
      n_257_76_17929));
   NAND4_X1 i_257_76_17961 (.A1(n_257_76_17922), .A2(n_257_76_17924), .A3(
      n_257_76_17926), .A4(n_257_76_17929), .ZN(n_257_76_17930));
   NOR2_X1 i_257_76_17962 (.A1(n_257_76_17916), .A2(n_257_76_17930), .ZN(
      n_257_76_17931));
   INV_X1 i_257_76_17963 (.A(n_257_76_17747), .ZN(n_257_76_17932));
   NAND2_X1 i_257_76_17964 (.A1(n_257_106), .A2(n_257_76_17932), .ZN(
      n_257_76_17933));
   NAND2_X1 i_257_76_17965 (.A1(n_257_436), .A2(n_257_442), .ZN(n_257_76_17934));
   INV_X1 i_257_76_17966 (.A(n_257_76_17934), .ZN(n_257_76_17935));
   NAND2_X1 i_257_76_17967 (.A1(n_257_764), .A2(n_257_76_17935), .ZN(
      n_257_76_17936));
   INV_X1 i_257_76_17968 (.A(n_257_76_17449), .ZN(n_257_76_17937));
   NAND2_X1 i_257_76_17969 (.A1(n_257_446), .A2(n_257_76_17937), .ZN(
      n_257_76_17938));
   NAND2_X1 i_257_76_17970 (.A1(n_257_439), .A2(n_257_442), .ZN(n_257_76_17939));
   INV_X1 i_257_76_17971 (.A(n_257_76_17939), .ZN(n_257_76_17940));
   NAND2_X1 i_257_76_17972 (.A1(n_257_930), .A2(n_257_76_17940), .ZN(
      n_257_76_17941));
   NAND4_X1 i_257_76_17973 (.A1(n_257_76_17933), .A2(n_257_76_17936), .A3(
      n_257_76_17938), .A4(n_257_76_17941), .ZN(n_257_76_17942));
   INV_X1 i_257_76_17974 (.A(n_257_76_17942), .ZN(n_257_76_17943));
   INV_X1 i_257_76_17975 (.A(n_257_76_17646), .ZN(n_257_76_17944));
   NAND2_X1 i_257_76_17976 (.A1(n_257_449), .A2(n_257_76_17944), .ZN(
      n_257_76_17945));
   INV_X1 i_257_76_17977 (.A(n_257_76_17736), .ZN(n_257_76_17946));
   NAND2_X1 i_257_76_17978 (.A1(n_257_447), .A2(n_257_76_17946), .ZN(
      n_257_76_17947));
   NAND2_X1 i_257_76_17979 (.A1(n_257_483), .A2(n_257_442), .ZN(n_257_76_17948));
   INV_X1 i_257_76_17980 (.A(n_257_76_17948), .ZN(n_257_76_17949));
   NAND2_X1 i_257_76_17981 (.A1(n_257_451), .A2(n_257_76_17949), .ZN(
      n_257_76_17950));
   NAND2_X1 i_257_76_17982 (.A1(n_257_437), .A2(n_257_442), .ZN(n_257_76_17951));
   INV_X1 i_257_76_17983 (.A(n_257_76_17951), .ZN(n_257_76_17952));
   NAND2_X1 i_257_76_17984 (.A1(n_257_828), .A2(n_257_76_17952), .ZN(
      n_257_76_17953));
   NAND4_X1 i_257_76_17985 (.A1(n_257_76_17945), .A2(n_257_76_17947), .A3(
      n_257_76_17950), .A4(n_257_76_17953), .ZN(n_257_76_17954));
   INV_X1 i_257_76_17986 (.A(n_257_76_17954), .ZN(n_257_76_17955));
   NAND4_X1 i_257_76_17987 (.A1(n_257_76_17901), .A2(n_257_76_17931), .A3(
      n_257_76_17943), .A4(n_257_76_17955), .ZN(n_257_76_17956));
   NAND2_X1 i_257_76_17988 (.A1(n_257_448), .A2(n_257_442), .ZN(n_257_76_17957));
   INV_X1 i_257_76_17989 (.A(n_257_76_17957), .ZN(n_257_76_17958));
   NAND2_X1 i_257_76_17990 (.A1(n_257_700), .A2(n_257_76_17958), .ZN(
      n_257_76_17959));
   INV_X1 i_257_76_17991 (.A(n_257_183), .ZN(n_257_76_17960));
   OAI21_X1 i_257_76_17992 (.A(n_257_76_17486), .B1(n_257_76_17960), .B2(
      n_257_76_17660), .ZN(n_257_76_17961));
   INV_X1 i_257_76_17993 (.A(n_257_76_17961), .ZN(n_257_76_17962));
   NAND2_X1 i_257_76_17994 (.A1(n_257_444), .A2(n_257_442), .ZN(n_257_76_17963));
   INV_X1 i_257_76_17995 (.A(n_257_76_17963), .ZN(n_257_76_17964));
   NAND2_X1 i_257_76_17996 (.A1(n_257_1026), .A2(n_257_76_17964), .ZN(
      n_257_76_17965));
   NAND3_X1 i_257_76_17997 (.A1(n_257_76_17959), .A2(n_257_76_17962), .A3(
      n_257_76_17965), .ZN(n_257_76_17966));
   NOR2_X1 i_257_76_17998 (.A1(n_257_76_17956), .A2(n_257_76_17966), .ZN(
      n_257_76_17967));
   NAND2_X1 i_257_76_17999 (.A1(n_257_443), .A2(n_257_442), .ZN(n_257_76_17968));
   INV_X1 i_257_76_18000 (.A(n_257_76_17968), .ZN(n_257_76_17969));
   NAND2_X1 i_257_76_18001 (.A1(n_257_1058), .A2(n_257_76_17969), .ZN(
      n_257_76_17970));
   NAND3_X1 i_257_76_18002 (.A1(n_257_76_17970), .A2(n_257_76_17804), .A3(
      n_257_76_17574), .ZN(n_257_76_17971));
   INV_X1 i_257_76_18003 (.A(n_257_76_17971), .ZN(n_257_76_17972));
   NAND3_X1 i_257_76_18004 (.A1(n_257_76_17967), .A2(n_257_76_17972), .A3(
      n_257_76_17789), .ZN(n_257_76_17973));
   NAND3_X1 i_257_76_18005 (.A1(n_257_76_17876), .A2(n_257_76_17896), .A3(
      n_257_76_17973), .ZN(n_257_76_17974));
   INV_X1 i_257_76_18006 (.A(n_257_76_17974), .ZN(n_257_76_17975));
   NAND3_X1 i_257_76_18007 (.A1(n_257_76_17814), .A2(n_257_76_17857), .A3(
      n_257_76_17975), .ZN(n_257_76_17976));
   NOR2_X1 i_257_76_18008 (.A1(n_257_76_17757), .A2(n_257_76_17976), .ZN(
      n_257_76_17977));
   NAND2_X1 i_257_76_18009 (.A1(n_257_76_17632), .A2(n_257_76_17977), .ZN(n_31));
   AOI21_X1 i_257_76_18010 (.A(n_257_76_16849), .B1(n_257_731), .B2(n_257_435), 
      .ZN(n_257_76_17978));
   AOI21_X1 i_257_76_18011 (.A(n_257_76_16274), .B1(n_257_730), .B2(n_257_435), 
      .ZN(n_257_76_17979));
   AOI21_X1 i_257_76_18012 (.A(n_257_76_15760), .B1(n_257_729), .B2(n_257_435), 
      .ZN(n_257_76_17980));
   AOI21_X1 i_257_76_18013 (.A(n_257_76_15256), .B1(n_257_592), .B2(n_257_428), 
      .ZN(n_257_76_17981));
   AOI21_X1 i_257_76_18014 (.A(n_257_76_15335), .B1(n_257_592), .B2(n_257_428), 
      .ZN(n_257_76_17982));
   AOI21_X1 i_257_76_18015 (.A(n_257_76_17660), .B1(n_257_432), .B2(n_257_624), 
      .ZN(n_257_76_17983));
   AOI21_X1 i_257_76_18016 (.A(n_257_76_15456), .B1(n_257_592), .B2(n_257_428), 
      .ZN(n_257_76_17984));
   AOI21_X1 i_257_76_18017 (.A(n_257_76_15535), .B1(n_257_592), .B2(n_257_428), 
      .ZN(n_257_76_17985));
   AOI21_X1 i_257_76_18018 (.A(n_257_76_15546), .B1(n_257_592), .B2(n_257_428), 
      .ZN(n_257_76_17986));
   AOI21_X1 i_257_76_18019 (.A(n_257_76_17412), .B1(n_257_592), .B2(n_257_428), 
      .ZN(n_257_76_17987));
   AOI21_X1 i_257_76_18020 (.A(n_257_76_15640), .B1(n_257_592), .B2(n_257_428), 
      .ZN(n_257_76_17988));
   AOI21_X1 i_257_76_18021 (.A(n_257_76_15665), .B1(n_257_592), .B2(n_257_428), 
      .ZN(n_257_76_17989));
   AOI21_X1 i_257_76_18022 (.A(n_257_76_17412), .B1(n_257_591), .B2(n_257_428), 
      .ZN(n_257_76_17990));
   AOI21_X1 i_257_76_18023 (.A(n_257_76_14913), .B1(n_257_591), .B2(n_257_428), 
      .ZN(n_257_76_17991));
   AOI21_X1 i_257_76_18024 (.A(n_257_76_15113), .B1(n_257_414), .B2(n_257_484), 
      .ZN(n_257_76_17992));
   AOI21_X1 i_257_76_18025 (.A(n_257_76_17412), .B1(n_257_590), .B2(n_257_428), 
      .ZN(n_257_76_17993));
   AOI21_X1 i_257_76_18026 (.A(n_257_76_14406), .B1(n_257_590), .B2(n_257_428), 
      .ZN(n_257_76_17994));
   AOI21_X1 i_257_76_18027 (.A(n_257_76_17723), .B1(n_257_432), .B2(n_257_622), 
      .ZN(n_257_76_17995));
   AOI21_X1 i_257_76_18028 (.A(n_257_76_14594), .B1(n_257_413), .B2(n_257_484), 
      .ZN(n_257_76_17996));
   AOI21_X1 i_257_76_18029 (.A(n_257_76_17412), .B1(n_257_589), .B2(n_257_428), 
      .ZN(n_257_76_17997));
   AOI21_X1 i_257_76_18030 (.A(n_257_76_13868), .B1(n_257_589), .B2(n_257_428), 
      .ZN(n_257_76_17998));
   AOI21_X1 i_257_76_18031 (.A(n_257_76_17723), .B1(n_257_432), .B2(n_257_621), 
      .ZN(n_257_76_17999));
   AOI21_X1 i_257_76_18032 (.A(n_257_76_17747), .B1(n_257_432), .B2(n_257_621), 
      .ZN(n_257_76_18000));
   AOI21_X1 i_257_76_18033 (.A(n_257_76_14078), .B1(n_257_589), .B2(n_257_428), 
      .ZN(n_257_76_18001));
   AOI21_X1 i_257_76_18034 (.A(n_257_76_17412), .B1(n_257_588), .B2(n_257_428), 
      .ZN(n_257_76_18002));
   AOI21_X1 i_257_76_18035 (.A(n_257_76_17660), .B1(n_257_432), .B2(n_257_620), 
      .ZN(n_257_76_18003));
   AOI21_X1 i_257_76_18036 (.A(n_257_76_13332), .B1(n_257_588), .B2(n_257_428), 
      .ZN(n_257_76_18004));
   AOI21_X1 i_257_76_18037 (.A(n_257_76_17723), .B1(n_257_432), .B2(n_257_620), 
      .ZN(n_257_76_18005));
   AOI21_X1 i_257_76_18038 (.A(n_257_76_17747), .B1(n_257_432), .B2(n_257_620), 
      .ZN(n_257_76_18006));
   AOI21_X1 i_257_76_18039 (.A(n_257_76_13555), .B1(n_257_411), .B2(n_257_484), 
      .ZN(n_257_76_18007));
   AOI21_X1 i_257_76_18040 (.A(n_257_76_17412), .B1(n_257_587), .B2(n_257_428), 
      .ZN(n_257_76_18008));
   AOI21_X1 i_257_76_18041 (.A(n_257_76_12777), .B1(n_257_587), .B2(n_257_428), 
      .ZN(n_257_76_18009));
   AOI21_X1 i_257_76_18042 (.A(n_257_76_12997), .B1(n_257_484), .B2(n_257_410), 
      .ZN(n_257_76_18010));
   AOI21_X1 i_257_76_18043 (.A(n_257_76_17412), .B1(n_257_586), .B2(n_257_428), 
      .ZN(n_257_76_18011));
   AOI21_X1 i_257_76_18044 (.A(n_257_76_17747), .B1(n_257_432), .B2(n_257_618), 
      .ZN(n_257_76_18012));
   AOI21_X1 i_257_76_18045 (.A(n_257_76_17723), .B1(n_257_432), .B2(n_257_618), 
      .ZN(n_257_76_18013));
   AOI21_X1 i_257_76_18046 (.A(n_257_76_12292), .B1(n_257_586), .B2(n_257_428), 
      .ZN(n_257_76_18014));
   AOI21_X1 i_257_76_18047 (.A(n_257_76_12416), .B1(n_257_484), .B2(n_257_409), 
      .ZN(n_257_76_18015));
   AOI21_X1 i_257_76_18048 (.A(n_257_76_17412), .B1(n_257_585), .B2(n_257_428), 
      .ZN(n_257_76_18016));
   AOI21_X1 i_257_76_18049 (.A(n_257_76_17723), .B1(n_257_432), .B2(n_257_617), 
      .ZN(n_257_76_18017));
   AOI21_X1 i_257_76_18050 (.A(n_257_76_17747), .B1(n_257_432), .B2(n_257_617), 
      .ZN(n_257_76_18018));
   AOI21_X1 i_257_76_18051 (.A(n_257_76_11907), .B1(n_257_408), .B2(n_257_484), 
      .ZN(n_257_76_18019));
   AOI21_X1 i_257_76_18052 (.A(n_257_76_17412), .B1(n_257_584), .B2(n_257_428), 
      .ZN(n_257_76_18020));
   AOI21_X1 i_257_76_18053 (.A(n_257_76_11129), .B1(n_257_584), .B2(n_257_428), 
      .ZN(n_257_76_18021));
   AOI21_X1 i_257_76_18054 (.A(n_257_76_11365), .B1(n_257_484), .B2(n_257_407), 
      .ZN(n_257_76_18022));
   AOI21_X1 i_257_76_18055 (.A(n_257_76_17412), .B1(n_257_428), .B2(n_257_583), 
      .ZN(n_257_76_18023));
   AOI21_X1 i_257_76_18056 (.A(n_257_76_10568), .B1(n_257_428), .B2(n_257_583), 
      .ZN(n_257_76_18024));
   AOI21_X1 i_257_76_18057 (.A(n_257_76_17412), .B1(n_257_719), .B2(n_257_435), 
      .ZN(n_257_76_18025));
   AOI21_X1 i_257_76_18058 (.A(n_257_76_10771), .B1(n_257_484), .B2(n_257_406), 
      .ZN(n_257_76_18026));
   AOI21_X1 i_257_76_18059 (.A(n_257_76_17412), .B1(n_257_582), .B2(n_257_428), 
      .ZN(n_257_76_18027));
   AOI21_X1 i_257_76_18060 (.A(n_257_76_17412), .B1(n_257_432), .B2(n_257_614), 
      .ZN(n_257_76_18028));
   AOI21_X1 i_257_76_18061 (.A(n_257_76_10028), .B1(n_257_582), .B2(n_257_428), 
      .ZN(n_257_76_18029));
   AOI21_X1 i_257_76_18062 (.A(n_257_76_10228), .B1(n_257_405), .B2(n_257_484), 
      .ZN(n_257_76_18030));
   AOI21_X1 i_257_76_18063 (.A(n_257_76_17412), .B1(n_257_581), .B2(n_257_428), 
      .ZN(n_257_76_18031));
   AOI21_X1 i_257_76_18064 (.A(n_257_76_17747), .B1(n_257_432), .B2(n_257_613), 
      .ZN(n_257_76_18032));
   AOI21_X1 i_257_76_18065 (.A(n_257_76_17660), .B1(n_257_432), .B2(n_257_613), 
      .ZN(n_257_76_18033));
   AOI21_X1 i_257_76_18066 (.A(n_257_76_9487), .B1(n_257_581), .B2(n_257_428), 
      .ZN(n_257_76_18034));
   AOI21_X1 i_257_76_18067 (.A(n_257_76_17723), .B1(n_257_432), .B2(n_257_613), 
      .ZN(n_257_76_18035));
   AOI21_X1 i_257_76_18068 (.A(n_257_76_9683), .B1(n_257_404), .B2(n_257_484), 
      .ZN(n_257_76_18036));
   AOI21_X1 i_257_76_18069 (.A(n_257_76_17412), .B1(n_257_1080), .B2(n_257_438), 
      .ZN(n_257_76_18037));
   AOI21_X1 i_257_76_18070 (.A(n_257_76_9172), .B1(n_257_403), .B2(n_257_484), 
      .ZN(n_257_76_18038));
   AOI21_X1 i_257_76_18071 (.A(n_257_76_8623), .B1(n_257_484), .B2(n_257_402), 
      .ZN(n_257_76_18039));
   AOI21_X1 i_257_76_18072 (.A(n_257_76_8102), .B1(n_257_484), .B2(n_257_401), 
      .ZN(n_257_76_18040));
   AOI21_X1 i_257_76_18073 (.A(n_257_76_7467), .B1(n_257_400), .B2(n_257_484), 
      .ZN(n_257_76_18041));
   AOI21_X1 i_257_76_18074 (.A(n_257_76_17412), .B1(n_257_1077), .B2(n_257_438), 
      .ZN(n_257_76_18042));
   AOI21_X1 i_257_76_18075 (.A(n_257_76_6504), .B1(n_257_438), .B2(n_257_1076), 
      .ZN(n_257_76_18043));
   AOI21_X1 i_257_76_18076 (.A(n_257_76_6957), .B1(n_257_484), .B2(n_257_399), 
      .ZN(n_257_76_18044));
   AOI21_X1 i_257_76_18077 (.A(n_257_76_6371), .B1(n_257_398), .B2(n_257_484), 
      .ZN(n_257_76_18045));
   AOI21_X1 i_257_76_18078 (.A(n_257_76_17412), .B1(n_257_1075), .B2(n_257_438), 
      .ZN(n_257_76_18046));
   AOI21_X1 i_257_76_18079 (.A(n_257_76_17412), .B1(n_257_438), .B2(n_257_1074), 
      .ZN(n_257_76_18047));
   AOI21_X1 i_257_76_18080 (.A(n_257_76_5817), .B1(n_257_397), .B2(n_257_484), 
      .ZN(n_257_76_18048));
   AOI21_X1 i_257_76_18081 (.A(n_257_76_5289), .B1(n_257_396), .B2(n_257_484), 
      .ZN(n_257_76_18049));
   AOI21_X1 i_257_76_18082 (.A(n_257_76_4776), .B1(n_257_1066), .B2(n_257_442), 
      .ZN(n_257_76_18050));
   AOI21_X1 i_257_76_18083 (.A(n_257_76_4159), .B1(n_257_1065), .B2(n_257_442), 
      .ZN(n_257_76_18051));
   AOI21_X1 i_257_76_18084 (.A(n_257_76_3013), .B1(n_257_435), .B2(n_257_706), 
      .ZN(n_257_76_18052));
   AOI21_X1 i_257_76_18085 (.A(n_257_76_2415), .B1(n_257_435), .B2(n_257_705), 
      .ZN(n_257_76_18053));
   AOI21_X1 i_257_76_18086 (.A(n_257_76_1804), .B1(n_257_704), .B2(n_257_435), 
      .ZN(n_257_76_18054));
   AOI21_X1 i_257_76_18087 (.A(n_257_76_2378), .B1(n_257_442), .B2(n_257_1062), 
      .ZN(n_257_76_18055));
   AOI21_X1 i_257_76_18088 (.A(n_257_76_1216), .B1(n_257_703), .B2(n_257_435), 
      .ZN(n_257_76_18056));
   AOI21_X1 i_257_76_18089 (.A(n_257_76_1744), .B1(n_257_442), .B2(n_257_1061), 
      .ZN(n_257_76_18057));
   AOI21_X1 i_257_76_18090 (.A(n_257_76_1151), .B1(n_257_1060), .B2(n_257_442), 
      .ZN(n_257_76_18058));
   AOI21_X1 i_257_76_18091 (.A(n_257_76_521), .B1(n_257_1059), .B2(n_257_442), 
      .ZN(n_257_76_18059));
   BUF_X1 rt_shieldBuf__1 (.A(n_257_12), .Z(n_257_76_18060));
   BUF_X1 rt_shieldBuf__1__1__0 (.A(n_257_184), .Z(n_257_76_18061));
   BUF_X1 rt_shieldBuf__1__1__1 (.A(n_257_265), .Z(n_257_76_18062));
   BUF_X1 rt_shieldBuf__1__1__2 (.A(n_257_434), .Z(n_257_76_18063));
   BUF_X1 rt_shieldBuf__1__1__3 (.A(n_257_264), .Z(n_257_76_18064));
   BUF_X1 rt_shieldBuf__1__1__4 (.A(n_257_224), .Z(n_257_76_18065));
   BUF_X1 rt_shieldBuf__1__1__5 (.A(n_257_304), .Z(n_257_76_18066));
   BUF_X1 rt_shieldBuf__1__1__6 (.A(n_257_19), .Z(n_257_76_18067));
   BUF_X1 rt_shieldBuf__1__1__7 (.A(n_257_145), .Z(n_257_76_18068));
   BUF_X1 rt_shieldBuf__1__1__8 (.A(n_257_24), .Z(n_257_76_18069));
   BUF_X1 rt_shieldBuf__1__1__9 (.A(n_257_21), .Z(n_257_76_18070));
   BUF_X1 rt_shieldBuf__1__1__10 (.A(n_257_16), .Z(n_257_76_18071));
   BUF_X1 rt_shieldBuf__1__1__11 (.A(n_257_14), .Z(n_257_76_18072));
   BUF_X1 rt_shieldBuf__1__1__12 (.A(n_257_382), .Z(n_257_76_18073));
   BUF_X1 rt_shieldBuf__1__1__13 (.A(n_257_185), .Z(n_257_76_18074));
   BUF_X1 rt_shieldBuf__1__1__14 (.A(n_257_15), .Z(n_257_76_18075));
   BUF_X1 rt_shieldBuf__1__1__15 (.A(n_257_225), .Z(n_257_76_18076));
   BUF_X1 rt_shieldBuf__1__1__16 (.A(n_257_20), .Z(n_257_76_18077));
   BUF_X1 rt_shieldBuf__1__1__17 (.A(n_257_25), .Z(n_257_76_18078));
   BUF_X1 rt_shieldBuf__1__1__18 (.A(n_257_26), .Z(n_257_76_18079));
   BUF_X1 rt_shieldBuf__1__1__19 (.A(n_257_107), .Z(n_257_76_18080));
   BUF_X1 rt_shieldBuf__1__1__20 (.A(n_257_67), .Z(n_257_76_18081));
   BUF_X1 rt_shieldBuf__1__1__21 (.A(n_257_381), .Z(n_257_76_18082));
   BUF_X1 rt_shieldBuf__1__1__22 (.A(n_257_27), .Z(n_257_76_18083));
   BUF_X1 rt_shieldBuf__1__1__23 (.A(n_257_18), .Z(n_257_76_18084));
   BUF_X1 rt_shieldBuf__1__1__24 (.A(n_257_23), .Z(n_257_76_18085));
   datapath__0_22 i_2_3 (.PacketSize(PacketSize), .p_0({uc_617, uc_618, uc_619, 
      uc_620, uc_621, n_2_5, n_2_4, n_2_3, n_2_2, n_2_1, n_2_0, uc_622}));
   datapath__0_24 i_2_5 (.p_0({uc_623, uc_624, uc_625, uc_626, uc_627, n_2_206, 
      n_2_205, n_2_204, n_2_203, n_2_202, n_2_201, n_2_200}), 
      .Small_Packet_Indication_Bit_Location(Small_Packet_Indication_Bit_Location), 
      .p_1({n_2_11, n_2_10, n_2_9, n_2_8, n_2_7, n_2_6}));
   datapath__0_196 i_2_13 (.p_0({n_2_155, n_2_154, n_2_153, n_2_152, n_2_151, 
      n_2_150, n_2_149, n_2_148, n_2_147, n_2_146, n_2_145, n_2_144, n_2_143, 
      n_2_142, n_2_141, n_2_140, n_2_139, n_2_138, n_2_137, n_2_136, n_2_135, 
      n_2_134, n_2_133, n_2_132, n_2_131, n_2_130, n_2_129, n_2_128, n_2_127, 
      n_2_126, n_2_125, n_2_124}), .Data_Size({Data_Size[5], Data_Size[4], 
      Data_Size[3], Data_Size[2], Data_Size[1], Data_Size[0]}), .p_1({n_2_43, 
      n_2_42, n_2_41, n_2_40, n_2_39, n_2_38, n_2_37, n_2_36, n_2_35, n_2_34, 
      n_2_33, n_2_32, n_2_31, n_2_30, n_2_29, n_2_28, n_2_27, n_2_26, n_2_25, 
      n_2_24, n_2_23, n_2_22, n_2_21, n_2_20, n_2_19, n_2_18, n_2_17, n_2_16, 
      n_2_15, n_2_14, n_2_13, n_2_12}));
   datapath__0_197 i_2_14 (.Data_Size({Data_Size[31], Data_Size[30], 
      Data_Size[29], Data_Size[28], Data_Size[27], Data_Size[26], Data_Size[25], 
      Data_Size[24], Data_Size[23], Data_Size[22], Data_Size[21], Data_Size[20], 
      Data_Size[19], Data_Size[18], Data_Size[17], Data_Size[16], Data_Size[15], 
      Data_Size[14], Data_Size[13], Data_Size[12], Data_Size[11], Data_Size[10], 
      Data_Size[9], Data_Size[8], Data_Size[7], Data_Size[6], uc_628, uc_629, 
      uc_630, uc_631, uc_632, uc_633}), .p_0({n_2_68, n_2_67, n_2_66, n_2_65, 
      n_2_64, n_2_63, n_2_62, n_2_61, n_2_60, n_2_59, n_2_58, n_2_57, n_2_56, 
      n_2_55, n_2_54, n_2_53, n_2_52, n_2_51, n_2_50, n_2_49, n_2_48, n_2_47, 
      n_2_46, n_2_45, n_2_44, uc_634, uc_635, uc_636, uc_637, uc_638, uc_639, 
      uc_640}));
   datapath__0_393 i_2_207 (.p_0(n_2_69), .p_1({uc_641, uc_642, uc_643, uc_644, 
      uc_645, uc_646, uc_647, uc_648, uc_649, uc_650, uc_651, uc_652, uc_653, 
      uc_654, uc_655, uc_656, uc_657, uc_658, uc_659, uc_660, uc_661, uc_662, 
      uc_663, uc_664, uc_665, n_2_123, n_2_122, n_2_121, n_2_120, n_2_119, 
      n_2_118, n_2_117, n_2_116, n_2_115, n_2_114, n_2_113, n_2_112, uc_666}), 
      .RowsCount({RowsCount[15], RowsCount[14], RowsCount[13], RowsCount[12], 
      RowsCount[11], RowsCount[10], RowsCount[9], RowsCount[8], RowsCount[7], 
      RowsCount[6], RowsCount[5], RowsCount[4], RowsCount[3], RowsCount[2], 
      RowsCount[1], uc_667}));
   datapath i_2_0 (.PacketSize(PacketSize), .p_0({n_37, uc_668, uc_669, uc_670, 
      uc_671, uc_672, uc_673, uc_674, uc_675, uc_676, uc_677, uc_678, uc_679, 
      uc_680, uc_681, uc_682, uc_683, uc_684, uc_685, uc_686, uc_687, uc_688, 
      uc_689, uc_690, uc_691, uc_692, n_36, n_35, n_34, n_33, n_32, uc_693}));
   datapath__2_420 i_2_1 (.p_0({uc_694, uc_695, uc_696, uc_697, uc_698, uc_699, 
      uc_700, uc_701, uc_702, uc_703, uc_704, uc_705, uc_706, uc_707, uc_708, 
      uc_709, uc_710, uc_711, uc_712, uc_713, uc_714, uc_715, uc_716, uc_717, 
      uc_718, n_37, n_36, n_35, n_34, n_33, n_32, n_151}), 
      .Small_Packet_Indication_Bit_Location(Small_Packet_Indication_Bit_Location), 
      .p_1(n_2_70));
   AOI22_X1 i_2_2_0 (.A1(n_2_2_32), .A2(n_2_12), .B1(Data_Size[0]), .B2(n_2_214), 
      .ZN(n_2_2_0));
   INV_X1 i_2_2_1 (.A(n_2_2_0), .ZN(n_2_71));
   AOI22_X1 i_2_2_2 (.A1(n_2_2_32), .A2(n_2_13), .B1(n_2_214), .B2(Data_Size[1]), 
      .ZN(n_2_2_1));
   INV_X1 i_2_2_3 (.A(n_2_2_1), .ZN(n_2_72));
   AOI22_X1 i_2_2_4 (.A1(n_2_2_32), .A2(n_2_14), .B1(n_2_214), .B2(Data_Size[2]), 
      .ZN(n_2_2_2));
   INV_X1 i_2_2_5 (.A(n_2_2_2), .ZN(n_2_73));
   AOI22_X1 i_2_2_6 (.A1(n_2_2_32), .A2(n_2_15), .B1(n_2_214), .B2(Data_Size[3]), 
      .ZN(n_2_2_3));
   INV_X1 i_2_2_7 (.A(n_2_2_3), .ZN(n_2_74));
   AOI22_X1 i_2_2_8 (.A1(n_2_2_32), .A2(n_2_16), .B1(n_2_214), .B2(Data_Size[4]), 
      .ZN(n_2_2_4));
   INV_X1 i_2_2_9 (.A(n_2_2_4), .ZN(n_2_75));
   AOI22_X1 i_2_2_10 (.A1(n_2_2_32), .A2(n_2_17), .B1(n_2_214), .B2(Data_Size[5]), 
      .ZN(n_2_2_5));
   INV_X1 i_2_2_11 (.A(n_2_2_5), .ZN(n_2_76));
   AOI22_X1 i_2_2_12 (.A1(n_2_2_32), .A2(n_2_18), .B1(n_2_214), .B2(n_2_170), 
      .ZN(n_2_2_6));
   INV_X1 i_2_2_13 (.A(n_2_2_6), .ZN(n_2_77));
   AOI22_X1 i_2_2_14 (.A1(n_2_2_32), .A2(n_2_19), .B1(n_2_214), .B2(n_2_44), 
      .ZN(n_2_2_7));
   INV_X1 i_2_2_15 (.A(n_2_2_7), .ZN(n_2_78));
   AOI22_X1 i_2_2_16 (.A1(n_2_2_32), .A2(n_2_20), .B1(n_2_214), .B2(n_2_45), 
      .ZN(n_2_2_8));
   INV_X1 i_2_2_17 (.A(n_2_2_8), .ZN(n_2_79));
   AOI22_X1 i_2_2_18 (.A1(n_2_2_32), .A2(n_2_21), .B1(n_2_214), .B2(n_2_46), 
      .ZN(n_2_2_9));
   INV_X1 i_2_2_19 (.A(n_2_2_9), .ZN(n_2_80));
   AOI22_X1 i_2_2_20 (.A1(n_2_2_32), .A2(n_2_22), .B1(n_2_214), .B2(n_2_47), 
      .ZN(n_2_2_10));
   INV_X1 i_2_2_21 (.A(n_2_2_10), .ZN(n_2_81));
   AOI22_X1 i_2_2_22 (.A1(n_2_2_32), .A2(n_2_23), .B1(n_2_214), .B2(n_2_48), 
      .ZN(n_2_2_11));
   INV_X1 i_2_2_23 (.A(n_2_2_11), .ZN(n_2_82));
   AOI22_X1 i_2_2_24 (.A1(n_2_2_32), .A2(n_2_24), .B1(n_2_214), .B2(n_2_49), 
      .ZN(n_2_2_12));
   INV_X1 i_2_2_25 (.A(n_2_2_12), .ZN(n_2_83));
   AOI22_X1 i_2_2_26 (.A1(n_2_2_32), .A2(n_2_25), .B1(n_2_214), .B2(n_2_50), 
      .ZN(n_2_2_13));
   INV_X1 i_2_2_27 (.A(n_2_2_13), .ZN(n_2_84));
   AOI22_X1 i_2_2_28 (.A1(n_2_2_32), .A2(n_2_26), .B1(n_2_214), .B2(n_2_51), 
      .ZN(n_2_2_14));
   INV_X1 i_2_2_29 (.A(n_2_2_14), .ZN(n_2_85));
   AOI22_X1 i_2_2_30 (.A1(n_2_2_32), .A2(n_2_27), .B1(n_2_214), .B2(n_2_52), 
      .ZN(n_2_2_15));
   INV_X1 i_2_2_31 (.A(n_2_2_15), .ZN(n_2_86));
   AOI22_X1 i_2_2_32 (.A1(n_2_2_32), .A2(n_2_28), .B1(n_2_214), .B2(n_2_53), 
      .ZN(n_2_2_16));
   INV_X1 i_2_2_33 (.A(n_2_2_16), .ZN(n_2_87));
   AOI22_X1 i_2_2_34 (.A1(n_2_2_32), .A2(n_2_29), .B1(n_2_214), .B2(n_2_54), 
      .ZN(n_2_2_17));
   INV_X1 i_2_2_35 (.A(n_2_2_17), .ZN(n_2_88));
   AOI22_X1 i_2_2_36 (.A1(n_2_2_32), .A2(n_2_32), .B1(n_2_214), .B2(n_2_57), 
      .ZN(n_2_2_18));
   INV_X1 i_2_2_37 (.A(n_2_2_18), .ZN(n_2_91));
   AOI22_X1 i_2_2_38 (.A1(n_2_2_32), .A2(n_2_36), .B1(n_2_214), .B2(n_2_61), 
      .ZN(n_2_2_19));
   INV_X1 i_2_2_39 (.A(n_2_2_19), .ZN(n_2_95));
   AOI22_X1 i_2_2_40 (.A1(n_2_2_32), .A2(n_2_39), .B1(n_2_214), .B2(n_2_64), 
      .ZN(n_2_2_20));
   INV_X1 i_2_2_41 (.A(n_2_2_20), .ZN(n_2_98));
   MUX2_X1 i_2_2_42 (.A(n_2_30), .B(n_2_55), .S(n_2_214), .Z(n_2_89));
   MUX2_X1 i_2_2_43 (.A(n_2_31), .B(n_2_56), .S(n_2_214), .Z(n_2_90));
   AOI21_X1 i_2_2_44 (.A(n_2_2_21), .B1(n_2_2_22), .B2(n_2_2_32), .ZN(n_2_92));
   NOR2_X1 i_2_2_45 (.A1(n_2_58), .A2(n_2_2_32), .ZN(n_2_2_21));
   INV_X1 i_2_2_46 (.A(n_2_33), .ZN(n_2_2_22));
   AOI21_X1 i_2_2_47 (.A(n_2_2_23), .B1(n_2_2_24), .B2(n_2_2_32), .ZN(n_2_93));
   NOR2_X1 i_2_2_48 (.A1(n_2_59), .A2(n_2_2_32), .ZN(n_2_2_23));
   INV_X1 i_2_2_49 (.A(n_2_34), .ZN(n_2_2_24));
   MUX2_X1 i_2_2_50 (.A(n_2_35), .B(n_2_60), .S(n_2_214), .Z(n_2_94));
   AOI21_X1 i_2_2_51 (.A(n_2_2_25), .B1(n_2_2_26), .B2(n_2_2_32), .ZN(n_2_96));
   NOR2_X1 i_2_2_52 (.A1(n_2_62), .A2(n_2_2_32), .ZN(n_2_2_25));
   INV_X1 i_2_2_53 (.A(n_2_37), .ZN(n_2_2_26));
   MUX2_X1 i_2_2_54 (.A(n_2_38), .B(n_2_63), .S(n_2_214), .Z(n_2_97));
   AOI21_X1 i_2_2_55 (.A(n_2_2_27), .B1(n_2_2_28), .B2(n_2_2_32), .ZN(n_2_99));
   NOR2_X1 i_2_2_56 (.A1(n_2_65), .A2(n_2_2_32), .ZN(n_2_2_27));
   INV_X1 i_2_2_57 (.A(n_2_40), .ZN(n_2_2_28));
   AOI21_X1 i_2_2_58 (.A(n_2_2_29), .B1(n_2_2_30), .B2(n_2_2_32), .ZN(n_2_100));
   NOR2_X1 i_2_2_59 (.A1(n_2_66), .A2(n_2_2_32), .ZN(n_2_2_29));
   INV_X1 i_2_2_60 (.A(n_2_41), .ZN(n_2_2_30));
   AOI21_X1 i_2_2_61 (.A(n_2_2_31), .B1(n_2_2_33), .B2(n_2_2_32), .ZN(n_2_101));
   NOR2_X1 i_2_2_62 (.A1(n_2_67), .A2(n_2_2_32), .ZN(n_2_2_31));
   INV_X1 i_2_2_63 (.A(n_2_214), .ZN(n_2_2_32));
   INV_X1 i_2_2_64 (.A(n_2_42), .ZN(n_2_2_33));
   MUX2_X1 i_2_2_65 (.A(n_2_43), .B(n_2_68), .S(n_2_214), .Z(n_2_102));
   INV_X1 i_2_4_0 (.A(n_2_83), .ZN(n_2_4_0));
   INV_X1 i_2_4_1 (.A(n_2_84), .ZN(n_2_4_1));
   INV_X1 i_2_4_2 (.A(n_2_86), .ZN(n_2_4_2));
   NAND3_X1 i_2_4_3 (.A1(n_2_4_0), .A2(n_2_4_1), .A3(n_2_4_2), .ZN(n_2_4_3));
   INV_X1 i_2_4_4 (.A(n_2_4_3), .ZN(n_2_4_4));
   INV_X1 i_2_4_5 (.A(n_2_85), .ZN(n_2_4_5));
   INV_X1 i_2_4_6 (.A(n_2_82), .ZN(n_2_4_6));
   INV_X1 i_2_4_7 (.A(n_2_87), .ZN(n_2_4_7));
   INV_X1 i_2_4_8 (.A(n_2_80), .ZN(n_2_4_8));
   INV_X1 i_2_4_9 (.A(n_2_78), .ZN(n_2_4_9));
   INV_X1 i_2_4_10 (.A(n_2_77), .ZN(n_2_4_10));
   NAND2_X1 i_2_4_11 (.A1(n_2_4_9), .A2(n_2_4_10), .ZN(n_2_4_11));
   NOR2_X1 i_2_4_12 (.A1(n_2_79), .A2(n_2_4_11), .ZN(n_2_4_12));
   NAND2_X1 i_2_4_13 (.A1(n_2_4_8), .A2(n_2_4_12), .ZN(n_2_4_13));
   NOR2_X1 i_2_4_14 (.A1(n_2_4_13), .A2(n_2_81), .ZN(n_2_4_14));
   NAND4_X1 i_2_4_15 (.A1(n_2_4_5), .A2(n_2_4_6), .A3(n_2_4_7), .A4(n_2_4_14), 
      .ZN(n_2_4_15));
   INV_X1 i_2_4_16 (.A(n_2_4_15), .ZN(n_2_4_16));
   INV_X1 i_2_4_17 (.A(n_2_88), .ZN(n_2_4_17));
   INV_X1 i_2_4_18 (.A(n_2_98), .ZN(n_2_4_18));
   NAND4_X1 i_2_4_19 (.A1(n_2_4_4), .A2(n_2_4_16), .A3(n_2_4_17), .A4(n_2_4_18), 
      .ZN(n_2_4_19));
   INV_X1 i_2_4_20 (.A(n_2_89), .ZN(n_2_4_20));
   INV_X1 i_2_4_21 (.A(n_2_95), .ZN(n_2_4_21));
   INV_X1 i_2_4_22 (.A(n_2_97), .ZN(n_2_4_22));
   NAND3_X1 i_2_4_23 (.A1(n_2_4_20), .A2(n_2_4_21), .A3(n_2_4_22), .ZN(n_2_4_23));
   NOR2_X1 i_2_4_24 (.A1(n_2_4_19), .A2(n_2_4_23), .ZN(n_2_4_24));
   NOR2_X1 i_2_4_25 (.A1(n_2_99), .A2(n_2_91), .ZN(n_2_4_25));
   NOR2_X1 i_2_4_26 (.A1(n_2_102), .A2(n_2_96), .ZN(n_2_4_26));
   NAND3_X1 i_2_4_27 (.A1(n_2_4_24), .A2(n_2_4_25), .A3(n_2_4_26), .ZN(n_2_4_27));
   INV_X1 i_2_4_28 (.A(n_2_90), .ZN(n_2_4_28));
   INV_X1 i_2_4_29 (.A(n_2_94), .ZN(n_2_4_29));
   INV_X1 i_2_4_30 (.A(n_2_101), .ZN(n_2_4_30));
   NAND3_X1 i_2_4_31 (.A1(n_2_4_28), .A2(n_2_4_29), .A3(n_2_4_30), .ZN(n_2_4_31));
   NOR2_X1 i_2_4_32 (.A1(n_2_4_27), .A2(n_2_4_31), .ZN(n_2_4_32));
   INV_X1 i_2_4_33 (.A(n_2_92), .ZN(n_2_4_33));
   NOR2_X1 i_2_4_34 (.A1(n_2_100), .A2(n_2_93), .ZN(n_2_4_34));
   NAND3_X1 i_2_4_35 (.A1(n_2_4_32), .A2(n_2_4_33), .A3(n_2_4_34), .ZN(n_2_103));
   AND2_X1 i_2_6_0 (.A1(n_2_6_0), .A2(n_2_71), .ZN(n_2_104));
   AND2_X1 i_2_6_1 (.A1(n_2_6_0), .A2(n_2_209), .ZN(n_2_105));
   INV_X1 i_2_6_2 (.A(n_2_103), .ZN(n_2_6_0));
   NOR2_X1 i_2_6_3 (.A1(n_2_103), .A2(n_2_6_1), .ZN(n_2_106));
   INV_X1 i_2_6_4 (.A(n_2_210), .ZN(n_2_6_1));
   NOR2_X1 i_2_6_5 (.A1(n_2_103), .A2(n_2_6_2), .ZN(n_2_107));
   INV_X1 i_2_6_6 (.A(n_2_211), .ZN(n_2_6_2));
   NOR2_X1 i_2_6_7 (.A1(n_2_103), .A2(n_2_6_3), .ZN(n_2_108));
   INV_X1 i_2_6_8 (.A(n_2_212), .ZN(n_2_6_3));
   NOR2_X1 i_2_6_9 (.A1(n_2_103), .A2(n_2_6_4), .ZN(n_2_109));
   INV_X1 i_2_6_10 (.A(n_2_213), .ZN(n_2_6_4));
   NOR2_X1 i_2_7_0 (.A1(n_2_105), .A2(n_2_7_0), .ZN(n_2_110));
   NAND4_X1 i_2_7_1 (.A1(n_2_7_1), .A2(n_2_7_5), .A3(n_2_7_4), .A4(n_2_7_2), 
      .ZN(n_2_7_0));
   NOR2_X1 i_2_7_2 (.A1(n_2_107), .A2(n_2_106), .ZN(n_2_7_1));
   OR3_X1 i_2_7_3 (.A1(n_2_7_3), .A2(Writing_Start_Index[3]), .A3(
      Writing_Start_Index[2]), .ZN(n_2_7_2));
   OR4_X1 i_2_7_4 (.A1(Writing_Start_Index[5]), .A2(Writing_Start_Index[1]), 
      .A3(Writing_Start_Index[4]), .A4(Writing_Start_Index[0]), .ZN(n_2_7_3));
   INV_X1 i_2_7_5 (.A(n_2_108), .ZN(n_2_7_4));
   INV_X1 i_2_7_6 (.A(n_2_109), .ZN(n_2_7_5));
   INV_X1 i_2_8_0 (.A(n_2_8_0), .ZN(n_2_111));
   OAI21_X1 i_2_8_1 (.A(n_2_8_1), .B1(n_269), .B2(n_2_110), .ZN(n_2_8_0));
   NAND2_X1 i_2_8_2 (.A1(n_2_110), .A2(n_2_8_2), .ZN(n_2_8_1));
   INV_X1 i_2_8_3 (.A(n_2_215), .ZN(n_2_8_2));
   AOI22_X1 i_2_9_0 (.A1(n_2_9_13), .A2(N[5]), .B1(n_2_207), .B2(n_2_219), 
      .ZN(n_2_9_0));
   INV_X1 i_2_9_1 (.A(n_2_9_0), .ZN(n_2_117));
   AOI22_X1 i_2_9_2 (.A1(n_2_9_13), .A2(N[6]), .B1(n_2_207), .B2(n_2_220), 
      .ZN(n_2_9_1));
   INV_X1 i_2_9_3 (.A(n_2_9_1), .ZN(n_2_118));
   AOI22_X1 i_2_9_4 (.A1(n_2_9_13), .A2(N[7]), .B1(n_2_207), .B2(n_2_221), 
      .ZN(n_2_9_2));
   INV_X1 i_2_9_5 (.A(n_2_9_2), .ZN(n_2_119));
   AOI22_X1 i_2_9_6 (.A1(n_2_9_13), .A2(N[8]), .B1(n_2_207), .B2(n_2_222), 
      .ZN(n_2_9_3));
   INV_X1 i_2_9_7 (.A(n_2_9_3), .ZN(n_2_120));
   AOI22_X1 i_2_9_8 (.A1(n_2_9_13), .A2(N[9]), .B1(n_2_207), .B2(n_2_223), 
      .ZN(n_2_9_4));
   INV_X1 i_2_9_9 (.A(n_2_9_4), .ZN(n_2_121));
   AOI22_X1 i_2_9_10 (.A1(n_2_9_13), .A2(N[10]), .B1(n_2_207), .B2(n_2_224), 
      .ZN(n_2_9_5));
   INV_X1 i_2_9_11 (.A(n_2_9_5), .ZN(n_2_122));
   AOI22_X1 i_2_9_12 (.A1(n_2_9_13), .A2(N[11]), .B1(n_2_207), .B2(n_2_225), 
      .ZN(n_2_9_6));
   INV_X1 i_2_9_13 (.A(n_2_9_6), .ZN(n_2_123));
   INV_X1 i_2_9_14 (.A(n_2_207), .ZN(n_2_9_7));
   AOI22_X1 i_2_9_15 (.A1(n_2_208), .A2(n_2_207), .B1(n_2_9_7), .B2(N[0]), 
      .ZN(n_2_9_8));
   INV_X1 i_2_9_16 (.A(n_2_9_8), .ZN(n_2_112));
   AOI22_X1 i_2_9_17 (.A1(n_2_111), .A2(n_2_207), .B1(n_2_9_7), .B2(N[1]), 
      .ZN(n_2_9_9));
   INV_X1 i_2_9_18 (.A(n_2_9_9), .ZN(n_2_113));
   AOI22_X1 i_2_9_19 (.A1(n_2_216), .A2(n_2_207), .B1(n_2_9_7), .B2(N[2]), 
      .ZN(n_2_9_10));
   INV_X1 i_2_9_20 (.A(n_2_9_10), .ZN(n_2_114));
   AOI22_X1 i_2_9_21 (.A1(n_2_217), .A2(n_2_207), .B1(n_2_9_7), .B2(N[3]), 
      .ZN(n_2_9_11));
   INV_X1 i_2_9_22 (.A(n_2_9_11), .ZN(n_2_115));
   AOI22_X1 i_2_9_23 (.A1(n_2_218), .A2(n_2_207), .B1(n_2_9_7), .B2(N[4]), 
      .ZN(n_2_9_12));
   INV_X1 i_2_9_24 (.A(n_2_9_12), .ZN(n_2_116));
   BUF_X1 i_2_9_25 (.A(n_2_9_7), .Z(n_2_9_13));
   AOI22_X1 i_2_10_0 (.A1(n_2_10_42), .A2(n_0), .B1(Small_Packet_Data_Size[0]), 
      .B2(Done_Element), .ZN(n_2_10_0));
   INV_X1 i_2_10_1 (.A(n_2_10_0), .ZN(n_2_124));
   AOI22_X1 i_2_10_2 (.A1(n_2_10_42), .A2(n_3), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[3]), .ZN(n_2_10_1));
   INV_X1 i_2_10_3 (.A(n_2_10_1), .ZN(n_2_127));
   AOI22_X1 i_2_10_4 (.A1(n_2_10_42), .A2(n_4), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[4]), .ZN(n_2_10_2));
   INV_X1 i_2_10_5 (.A(n_2_10_2), .ZN(n_2_128));
   AOI22_X1 i_2_10_6 (.A1(n_2_10_42), .A2(n_8), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[8]), .ZN(n_2_10_3));
   INV_X1 i_2_10_7 (.A(n_2_10_3), .ZN(n_2_132));
   AOI22_X1 i_2_10_8 (.A1(n_2_10_42), .A2(n_11), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[11]), .ZN(n_2_10_4));
   INV_X1 i_2_10_9 (.A(n_2_10_4), .ZN(n_2_135));
   AOI22_X1 i_2_10_10 (.A1(n_2_10_42), .A2(n_13), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[13]), .ZN(n_2_10_5));
   INV_X1 i_2_10_11 (.A(n_2_10_5), .ZN(n_2_137));
   AOI22_X1 i_2_10_12 (.A1(n_2_10_42), .A2(n_14), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[14]), .ZN(n_2_10_6));
   INV_X1 i_2_10_13 (.A(n_2_10_6), .ZN(n_2_138));
   AOI22_X1 i_2_10_14 (.A1(n_2_10_42), .A2(n_16), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[16]), .ZN(n_2_10_7));
   INV_X1 i_2_10_15 (.A(n_2_10_7), .ZN(n_2_140));
   AOI22_X1 i_2_10_16 (.A1(n_2_10_42), .A2(n_17), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[17]), .ZN(n_2_10_8));
   INV_X1 i_2_10_17 (.A(n_2_10_8), .ZN(n_2_141));
   AOI22_X1 i_2_10_18 (.A1(n_2_10_42), .A2(n_18), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[18]), .ZN(n_2_10_9));
   INV_X1 i_2_10_19 (.A(n_2_10_9), .ZN(n_2_142));
   AOI22_X1 i_2_10_20 (.A1(n_2_10_42), .A2(n_19), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[19]), .ZN(n_2_10_10));
   INV_X1 i_2_10_21 (.A(n_2_10_10), .ZN(n_2_143));
   AOI22_X1 i_2_10_22 (.A1(n_2_10_42), .A2(n_20), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[20]), .ZN(n_2_10_11));
   INV_X1 i_2_10_23 (.A(n_2_10_11), .ZN(n_2_144));
   AOI22_X1 i_2_10_24 (.A1(n_2_10_42), .A2(n_21), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[21]), .ZN(n_2_10_12));
   INV_X1 i_2_10_25 (.A(n_2_10_12), .ZN(n_2_145));
   AOI22_X1 i_2_10_26 (.A1(n_2_10_42), .A2(n_22), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[22]), .ZN(n_2_10_13));
   INV_X1 i_2_10_27 (.A(n_2_10_13), .ZN(n_2_146));
   AOI22_X1 i_2_10_28 (.A1(n_2_10_42), .A2(n_23), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[23]), .ZN(n_2_10_14));
   INV_X1 i_2_10_29 (.A(n_2_10_14), .ZN(n_2_147));
   AOI22_X1 i_2_10_30 (.A1(n_2_10_42), .A2(n_24), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[24]), .ZN(n_2_10_15));
   INV_X1 i_2_10_31 (.A(n_2_10_15), .ZN(n_2_148));
   AOI22_X1 i_2_10_32 (.A1(n_2_10_42), .A2(n_26), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[26]), .ZN(n_2_10_16));
   INV_X1 i_2_10_33 (.A(n_2_10_16), .ZN(n_2_150));
   AOI22_X1 i_2_10_34 (.A1(n_2_10_42), .A2(n_28), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[28]), .ZN(n_2_10_17));
   INV_X1 i_2_10_35 (.A(n_2_10_17), .ZN(n_2_152));
   AOI22_X1 i_2_10_36 (.A1(n_2_10_42), .A2(n_29), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[29]), .ZN(n_2_10_18));
   INV_X1 i_2_10_37 (.A(n_2_10_18), .ZN(n_2_153));
   AOI22_X1 i_2_10_38 (.A1(n_2_10_42), .A2(n_30), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[30]), .ZN(n_2_10_19));
   INV_X1 i_2_10_39 (.A(n_2_10_19), .ZN(n_2_154));
   AOI22_X1 i_2_10_40 (.A1(n_2_10_42), .A2(n_31), .B1(Done_Element), .B2(
      Small_Packet_Data_Size[31]), .ZN(n_2_10_20));
   INV_X1 i_2_10_41 (.A(n_2_10_20), .ZN(n_2_155));
   NAND2_X1 i_2_10_42 (.A1(n_2_10_21), .A2(n_2_10_22), .ZN(n_2_125));
   NAND2_X1 i_2_10_43 (.A1(n_2_10_42), .A2(n_1), .ZN(n_2_10_21));
   NAND2_X1 i_2_10_44 (.A1(Small_Packet_Data_Size[1]), .A2(Done_Element), 
      .ZN(n_2_10_22));
   NAND2_X1 i_2_10_45 (.A1(n_2_10_23), .A2(n_2_10_24), .ZN(n_2_126));
   NAND2_X1 i_2_10_46 (.A1(n_2_10_42), .A2(n_2), .ZN(n_2_10_23));
   NAND2_X1 i_2_10_47 (.A1(Small_Packet_Data_Size[2]), .A2(Done_Element), 
      .ZN(n_2_10_24));
   NAND2_X1 i_2_10_48 (.A1(n_2_10_25), .A2(n_2_10_26), .ZN(n_2_129));
   NAND2_X1 i_2_10_49 (.A1(n_2_10_42), .A2(n_5), .ZN(n_2_10_25));
   NAND2_X1 i_2_10_50 (.A1(Small_Packet_Data_Size[5]), .A2(Done_Element), 
      .ZN(n_2_10_26));
   NAND2_X1 i_2_10_51 (.A1(n_2_10_27), .A2(n_2_10_28), .ZN(n_2_130));
   NAND2_X1 i_2_10_52 (.A1(n_2_10_42), .A2(n_6), .ZN(n_2_10_27));
   NAND2_X1 i_2_10_53 (.A1(Small_Packet_Data_Size[6]), .A2(Done_Element), 
      .ZN(n_2_10_28));
   NAND2_X1 i_2_10_54 (.A1(n_2_10_29), .A2(n_2_10_30), .ZN(n_2_131));
   NAND2_X1 i_2_10_55 (.A1(n_2_10_42), .A2(n_7), .ZN(n_2_10_29));
   NAND2_X1 i_2_10_56 (.A1(Small_Packet_Data_Size[7]), .A2(Done_Element), 
      .ZN(n_2_10_30));
   NAND2_X1 i_2_10_57 (.A1(n_2_10_31), .A2(n_2_10_32), .ZN(n_2_133));
   NAND2_X1 i_2_10_58 (.A1(n_2_10_42), .A2(n_9), .ZN(n_2_10_31));
   NAND2_X1 i_2_10_59 (.A1(Small_Packet_Data_Size[9]), .A2(Done_Element), 
      .ZN(n_2_10_32));
   NAND2_X1 i_2_10_60 (.A1(n_2_10_33), .A2(n_2_10_34), .ZN(n_2_134));
   NAND2_X1 i_2_10_61 (.A1(n_2_10_42), .A2(n_10), .ZN(n_2_10_33));
   NAND2_X1 i_2_10_62 (.A1(Small_Packet_Data_Size[10]), .A2(Done_Element), 
      .ZN(n_2_10_34));
   NAND2_X1 i_2_10_63 (.A1(n_2_10_35), .A2(n_2_10_36), .ZN(n_2_136));
   NAND2_X1 i_2_10_64 (.A1(n_2_10_42), .A2(n_12), .ZN(n_2_10_35));
   NAND2_X1 i_2_10_65 (.A1(Small_Packet_Data_Size[12]), .A2(Done_Element), 
      .ZN(n_2_10_36));
   NAND2_X1 i_2_10_66 (.A1(n_2_10_37), .A2(n_2_10_38), .ZN(n_2_139));
   NAND2_X1 i_2_10_67 (.A1(n_2_10_42), .A2(n_15), .ZN(n_2_10_37));
   NAND2_X1 i_2_10_68 (.A1(Small_Packet_Data_Size[15]), .A2(Done_Element), 
      .ZN(n_2_10_38));
   NAND2_X1 i_2_10_69 (.A1(n_2_10_39), .A2(n_2_10_40), .ZN(n_2_149));
   NAND2_X1 i_2_10_70 (.A1(n_2_10_42), .A2(n_25), .ZN(n_2_10_39));
   NAND2_X1 i_2_10_71 (.A1(Small_Packet_Data_Size[25]), .A2(Done_Element), 
      .ZN(n_2_10_40));
   NAND2_X1 i_2_10_72 (.A1(n_2_10_41), .A2(n_2_10_43), .ZN(n_2_151));
   NAND2_X1 i_2_10_73 (.A1(n_2_10_42), .A2(n_27), .ZN(n_2_10_41));
   INV_X1 i_2_10_74 (.A(Done_Element), .ZN(n_2_10_42));
   NAND2_X1 i_2_10_75 (.A1(Small_Packet_Data_Size[27]), .A2(Done_Element), 
      .ZN(n_2_10_43));
   datapath__2_568 i_2_11 (.p_0({n_2_123, n_2_122, n_2_121, n_2_120, n_2_119, 
      n_2_118, n_2_117, n_2_116, n_2_115, n_2_114, n_2_113, n_2_112}), .p_1({
      n_2_168, n_2_167, n_2_166, n_2_165, n_2_164, n_2_163, n_2_162, n_2_161, 
      n_2_160, n_2_159, n_2_158, n_2_157, n_2_156}));
   datapath__2_569 i_2_12 (.p_0({n_2_168, n_2_167, n_2_166, n_2_165, n_2_164, 
      n_2_163, n_2_162, n_2_161, n_2_160, n_2_159, n_2_158, n_2_157, n_2_156}), 
      .RowsCount(RowsCount), .p_1(n_2_169));
   OAI21_X1 i_2_15_0 (.A(n_2_15_4), .B1(n_2_169), .B2(n_2_15_0), .ZN(n_38));
   NAND3_X1 i_2_15_1 (.A1(n_2_15_3), .A2(n_2_69), .A3(n_2_15_1), .ZN(n_2_15_0));
   INV_X1 i_2_15_2 (.A(n_2_15_2), .ZN(n_2_15_1));
   NAND3_X1 i_2_15_3 (.A1(n_2_103), .A2(n_2_198), .A3(n_2_197), .ZN(n_2_15_2));
   INV_X1 i_2_15_4 (.A(n_2_196), .ZN(n_2_15_3));
   INV_X1 i_2_15_5 (.A(n_2_199), .ZN(n_2_15_4));
   AOI21_X1 i_2_16_0 (.A(n_2_16_0), .B1(n_2_16_4), .B2(n_2_16_2), .ZN(n_39));
   NAND2_X1 i_2_16_1 (.A1(n_2_16_1), .A2(n_2_197), .ZN(n_2_16_0));
   INV_X1 i_2_16_2 (.A(n_2_199), .ZN(n_2_16_1));
   INV_X1 i_2_16_3 (.A(n_2_16_3), .ZN(n_2_16_2));
   NAND2_X1 i_2_16_4 (.A1(n_2_103), .A2(n_2_198), .ZN(n_2_16_3));
   NAND3_X1 i_2_16_5 (.A1(n_2_16_7), .A2(n_2_16_6), .A3(n_2_16_5), .ZN(n_2_16_4));
   INV_X1 i_2_16_6 (.A(n_2_169), .ZN(n_2_16_5));
   INV_X1 i_2_16_7 (.A(n_2_196), .ZN(n_2_16_6));
   INV_X1 i_2_16_8 (.A(n_2_69), .ZN(n_2_16_7));
   NOR2_X1 i_2_17_0 (.A1(n_2_199), .A2(n_2_171), .ZN(n_2_17_0));
   NAND2_X1 i_2_17_1 (.A1(n_2_17_0), .A2(n_2_17_106), .ZN(n_2_17_1));
   INV_X1 i_2_17_2 (.A(n_2_17_0), .ZN(n_2_17_2));
   OAI21_X1 i_2_17_3 (.A(n_2_17_1), .B1(n_2_103), .B2(n_2_17_2), .ZN(n_2_17_3));
   NAND2_X1 i_2_17_4 (.A1(n_2_17_115), .A2(n_2_17_0), .ZN(n_2_17_4));
   NOR2_X1 i_2_17_5 (.A1(n_2_196), .A2(n_2_17_4), .ZN(n_2_17_5));
   AOI21_X1 i_2_17_6 (.A(n_2_17_3), .B1(n_2_17_99), .B2(n_2_17_5), .ZN(n_40));
   INV_X1 i_2_17_7 (.A(n_2_172), .ZN(n_2_17_6));
   INV_X1 i_2_17_8 (.A(n_2_184), .ZN(n_2_17_7));
   MUX2_X1 i_2_17_9 (.A(n_2_17_6), .B(n_2_17_7), .S(n_2_69), .Z(n_2_17_8));
   NAND3_X1 i_2_17_10 (.A1(n_2_17_99), .A2(n_2_17_8), .A3(n_2_17_68), .ZN(
      n_2_17_9));
   NAND2_X1 i_2_17_11 (.A1(n_2_17_6), .A2(n_2_17_106), .ZN(n_2_17_10));
   NOR2_X1 i_2_17_12 (.A1(n_2_199), .A2(n_2_17_10), .ZN(n_2_17_11));
   NOR2_X1 i_2_17_13 (.A1(n_2_199), .A2(n_2_172), .ZN(n_2_17_12));
   AOI21_X1 i_2_17_14 (.A(n_2_17_11), .B1(n_2_17_109), .B2(n_2_17_12), .ZN(
      n_2_17_13));
   NAND2_X1 i_2_17_15 (.A1(n_2_17_9), .A2(n_2_17_13), .ZN(n_2_17_14));
   INV_X1 i_2_17_16 (.A(n_2_17_14), .ZN(n_41));
   NAND2_X1 i_2_17_17 (.A1(n_2_173), .A2(n_2_17_106), .ZN(n_2_17_15));
   NAND2_X1 i_2_17_18 (.A1(n_2_17_96), .A2(n_2_17_15), .ZN(n_2_17_16));
   AOI21_X1 i_2_17_19 (.A(n_2_17_16), .B1(n_2_17_109), .B2(n_2_173), .ZN(
      n_2_17_17));
   NAND2_X1 i_2_17_20 (.A1(n_2_17_115), .A2(n_2_173), .ZN(n_2_17_18));
   NAND2_X1 i_2_17_21 (.A1(n_2_185), .A2(n_2_197), .ZN(n_2_17_19));
   INV_X1 i_2_17_22 (.A(n_2_17_19), .ZN(n_2_17_20));
   NAND3_X1 i_2_17_23 (.A1(n_2_69), .A2(n_2_103), .A3(n_2_17_20), .ZN(n_2_17_21));
   NAND2_X1 i_2_17_24 (.A1(n_2_17_18), .A2(n_2_17_21), .ZN(n_2_17_22));
   NOR2_X1 i_2_17_25 (.A1(n_2_17_114), .A2(n_2_17_22), .ZN(n_2_17_23));
   OAI21_X1 i_2_17_26 (.A(n_2_17_17), .B1(n_2_169), .B2(n_2_17_23), .ZN(n_42));
   INV_X1 i_2_17_27 (.A(n_2_174), .ZN(n_2_17_24));
   INV_X1 i_2_17_28 (.A(n_2_186), .ZN(n_2_17_25));
   MUX2_X1 i_2_17_29 (.A(n_2_17_24), .B(n_2_17_25), .S(n_2_69), .Z(n_2_17_26));
   NAND3_X1 i_2_17_30 (.A1(n_2_17_99), .A2(n_2_17_26), .A3(n_2_17_68), .ZN(
      n_2_17_27));
   NOR2_X1 i_2_17_31 (.A1(n_2_174), .A2(n_2_17_70), .ZN(n_2_17_28));
   NOR2_X1 i_2_17_32 (.A1(n_2_174), .A2(n_2_199), .ZN(n_2_17_29));
   AOI21_X1 i_2_17_33 (.A(n_2_17_28), .B1(n_2_17_109), .B2(n_2_17_29), .ZN(
      n_2_17_30));
   NAND2_X1 i_2_17_34 (.A1(n_2_17_27), .A2(n_2_17_30), .ZN(n_2_17_31));
   INV_X1 i_2_17_35 (.A(n_2_17_31), .ZN(n_43));
   NAND2_X1 i_2_17_36 (.A1(n_2_187), .A2(n_2_197), .ZN(n_2_17_32));
   INV_X1 i_2_17_37 (.A(n_2_17_32), .ZN(n_2_17_33));
   NAND2_X1 i_2_17_38 (.A1(n_2_103), .A2(n_2_17_33), .ZN(n_2_17_34));
   INV_X1 i_2_17_39 (.A(n_2_17_34), .ZN(n_2_17_35));
   MUX2_X1 i_2_17_40 (.A(n_2_175), .B(n_2_17_35), .S(n_2_69), .Z(n_2_17_36));
   NAND3_X1 i_2_17_41 (.A1(n_2_17_99), .A2(n_2_17_36), .A3(n_2_17_104), .ZN(
      n_2_17_37));
   AOI21_X1 i_2_17_42 (.A(n_2_199), .B1(n_2_175), .B2(n_2_17_106), .ZN(n_2_17_38));
   INV_X1 i_2_17_43 (.A(n_2_17_38), .ZN(n_2_17_39));
   AOI21_X1 i_2_17_44 (.A(n_2_17_39), .B1(n_2_17_109), .B2(n_2_175), .ZN(
      n_2_17_40));
   NAND2_X1 i_2_17_45 (.A1(n_2_17_37), .A2(n_2_17_40), .ZN(n_44));
   NAND2_X1 i_2_17_46 (.A1(n_2_188), .A2(n_2_197), .ZN(n_2_17_41));
   INV_X1 i_2_17_47 (.A(n_2_17_41), .ZN(n_2_17_42));
   NAND2_X1 i_2_17_48 (.A1(n_2_103), .A2(n_2_17_42), .ZN(n_2_17_43));
   INV_X1 i_2_17_49 (.A(n_2_17_43), .ZN(n_2_17_44));
   MUX2_X1 i_2_17_50 (.A(n_2_176), .B(n_2_17_44), .S(n_2_69), .Z(n_2_17_45));
   NAND3_X1 i_2_17_51 (.A1(n_2_17_99), .A2(n_2_17_45), .A3(n_2_17_104), .ZN(
      n_2_17_46));
   AOI21_X1 i_2_17_52 (.A(n_2_199), .B1(n_2_176), .B2(n_2_17_106), .ZN(n_2_17_47));
   INV_X1 i_2_17_53 (.A(n_2_17_47), .ZN(n_2_17_48));
   AOI21_X1 i_2_17_54 (.A(n_2_17_48), .B1(n_2_17_109), .B2(n_2_176), .ZN(
      n_2_17_49));
   NAND2_X1 i_2_17_55 (.A1(n_2_17_46), .A2(n_2_17_49), .ZN(n_45));
   INV_X1 i_2_17_56 (.A(n_2_177), .ZN(n_2_17_50));
   NAND2_X1 i_2_17_57 (.A1(n_2_17_50), .A2(n_2_17_94), .ZN(n_2_17_51));
   NAND2_X1 i_2_17_58 (.A1(n_2_17_50), .A2(n_2_17_96), .ZN(n_2_17_52));
   OAI21_X1 i_2_17_59 (.A(n_2_17_51), .B1(n_2_103), .B2(n_2_17_52), .ZN(
      n_2_17_53));
   INV_X1 i_2_17_60 (.A(n_2_189), .ZN(n_2_17_54));
   OAI22_X1 i_2_17_61 (.A1(n_2_17_115), .A2(n_2_17_54), .B1(n_2_69), .B2(
      n_2_17_50), .ZN(n_2_17_55));
   AOI21_X1 i_2_17_62 (.A(n_2_17_101), .B1(n_2_17_55), .B2(n_2_17_104), .ZN(
      n_2_17_56));
   AOI21_X1 i_2_17_63 (.A(n_2_17_53), .B1(n_2_17_99), .B2(n_2_17_56), .ZN(n_46));
   INV_X1 i_2_17_64 (.A(n_2_178), .ZN(n_2_17_57));
   INV_X1 i_2_17_65 (.A(n_2_190), .ZN(n_2_17_58));
   MUX2_X1 i_2_17_66 (.A(n_2_17_57), .B(n_2_17_58), .S(n_2_69), .Z(n_2_17_59));
   NAND3_X1 i_2_17_67 (.A1(n_2_17_99), .A2(n_2_17_59), .A3(n_2_17_68), .ZN(
      n_2_17_60));
   NOR2_X1 i_2_17_68 (.A1(n_2_178), .A2(n_2_17_70), .ZN(n_2_17_61));
   NOR2_X1 i_2_17_69 (.A1(n_2_178), .A2(n_2_199), .ZN(n_2_17_62));
   AOI21_X1 i_2_17_70 (.A(n_2_17_61), .B1(n_2_17_109), .B2(n_2_17_62), .ZN(
      n_2_17_63));
   NAND2_X1 i_2_17_71 (.A1(n_2_17_60), .A2(n_2_17_63), .ZN(n_2_17_64));
   INV_X1 i_2_17_72 (.A(n_2_17_64), .ZN(n_47));
   INV_X1 i_2_17_73 (.A(n_2_179), .ZN(n_2_17_65));
   INV_X1 i_2_17_74 (.A(n_2_191), .ZN(n_2_17_66));
   MUX2_X1 i_2_17_75 (.A(n_2_17_65), .B(n_2_17_66), .S(n_2_69), .Z(n_2_17_67));
   NOR2_X1 i_2_17_76 (.A1(n_2_196), .A2(n_2_17_101), .ZN(n_2_17_68));
   NAND3_X1 i_2_17_77 (.A1(n_2_17_99), .A2(n_2_17_67), .A3(n_2_17_68), .ZN(
      n_2_17_69));
   NAND2_X1 i_2_17_78 (.A1(n_2_17_96), .A2(n_2_17_106), .ZN(n_2_17_70));
   NOR2_X1 i_2_17_79 (.A1(n_2_179), .A2(n_2_17_70), .ZN(n_2_17_71));
   NOR2_X1 i_2_17_80 (.A1(n_2_179), .A2(n_2_199), .ZN(n_2_17_72));
   AOI21_X1 i_2_17_81 (.A(n_2_17_71), .B1(n_2_17_109), .B2(n_2_17_72), .ZN(
      n_2_17_73));
   NAND2_X1 i_2_17_82 (.A1(n_2_17_69), .A2(n_2_17_73), .ZN(n_2_17_74));
   INV_X1 i_2_17_83 (.A(n_2_17_74), .ZN(n_48));
   AOI21_X1 i_2_17_84 (.A(n_2_199), .B1(n_2_180), .B2(n_2_17_106), .ZN(n_2_17_75));
   INV_X1 i_2_17_85 (.A(n_2_17_75), .ZN(n_2_17_76));
   AOI21_X1 i_2_17_86 (.A(n_2_17_76), .B1(n_2_17_109), .B2(n_2_180), .ZN(
      n_2_17_77));
   NAND2_X1 i_2_17_87 (.A1(n_2_17_115), .A2(n_2_180), .ZN(n_2_17_78));
   NAND2_X1 i_2_17_88 (.A1(n_2_192), .A2(n_2_197), .ZN(n_2_17_79));
   INV_X1 i_2_17_89 (.A(n_2_17_79), .ZN(n_2_17_80));
   NAND3_X1 i_2_17_90 (.A1(n_2_69), .A2(n_2_103), .A3(n_2_17_80), .ZN(n_2_17_81));
   NAND2_X1 i_2_17_91 (.A1(n_2_17_78), .A2(n_2_17_81), .ZN(n_2_17_82));
   NOR2_X1 i_2_17_92 (.A1(n_2_17_114), .A2(n_2_17_82), .ZN(n_2_17_83));
   OAI21_X1 i_2_17_93 (.A(n_2_17_77), .B1(n_2_169), .B2(n_2_17_83), .ZN(n_49));
   NAND2_X1 i_2_17_94 (.A1(n_2_193), .A2(n_2_197), .ZN(n_2_17_84));
   INV_X1 i_2_17_95 (.A(n_2_17_84), .ZN(n_2_17_85));
   NAND2_X1 i_2_17_96 (.A1(n_2_103), .A2(n_2_17_85), .ZN(n_2_17_86));
   INV_X1 i_2_17_97 (.A(n_2_17_86), .ZN(n_2_17_87));
   MUX2_X1 i_2_17_98 (.A(n_2_181), .B(n_2_17_87), .S(n_2_69), .Z(n_2_17_88));
   NAND3_X1 i_2_17_99 (.A1(n_2_17_99), .A2(n_2_17_88), .A3(n_2_17_104), .ZN(
      n_2_17_89));
   AOI21_X1 i_2_17_100 (.A(n_2_199), .B1(n_2_181), .B2(n_2_17_106), .ZN(
      n_2_17_90));
   INV_X1 i_2_17_101 (.A(n_2_17_90), .ZN(n_2_17_91));
   AOI21_X1 i_2_17_102 (.A(n_2_17_91), .B1(n_2_17_109), .B2(n_2_181), .ZN(
      n_2_17_92));
   NAND2_X1 i_2_17_103 (.A1(n_2_17_89), .A2(n_2_17_92), .ZN(n_50));
   INV_X1 i_2_17_104 (.A(n_2_182), .ZN(n_2_17_93));
   NOR2_X1 i_2_17_105 (.A1(n_2_199), .A2(n_2_197), .ZN(n_2_17_94));
   NAND2_X1 i_2_17_106 (.A1(n_2_17_93), .A2(n_2_17_94), .ZN(n_2_17_95));
   INV_X1 i_2_17_107 (.A(n_2_199), .ZN(n_2_17_96));
   NAND2_X1 i_2_17_108 (.A1(n_2_17_93), .A2(n_2_17_96), .ZN(n_2_17_97));
   OAI21_X1 i_2_17_109 (.A(n_2_17_95), .B1(n_2_103), .B2(n_2_17_97), .ZN(
      n_2_17_98));
   INV_X1 i_2_17_110 (.A(n_2_169), .ZN(n_2_17_99));
   NOR2_X1 i_2_17_111 (.A1(n_2_199), .A2(n_2_17_106), .ZN(n_2_17_100));
   NAND2_X1 i_2_17_112 (.A1(n_2_103), .A2(n_2_17_100), .ZN(n_2_17_101));
   INV_X1 i_2_17_113 (.A(n_2_194), .ZN(n_2_17_102));
   OAI22_X1 i_2_17_114 (.A1(n_2_17_115), .A2(n_2_17_102), .B1(n_2_69), .B2(
      n_2_17_93), .ZN(n_2_17_103));
   INV_X1 i_2_17_115 (.A(n_2_196), .ZN(n_2_17_104));
   AOI21_X1 i_2_17_116 (.A(n_2_17_101), .B1(n_2_17_103), .B2(n_2_17_104), 
      .ZN(n_2_17_105));
   AOI21_X1 i_2_17_117 (.A(n_2_17_98), .B1(n_2_17_99), .B2(n_2_17_105), .ZN(n_51));
   INV_X1 i_2_17_118 (.A(n_2_197), .ZN(n_2_17_106));
   AOI21_X1 i_2_17_119 (.A(n_2_199), .B1(n_2_183), .B2(n_2_17_106), .ZN(
      n_2_17_107));
   INV_X1 i_2_17_120 (.A(n_2_17_107), .ZN(n_2_17_108));
   INV_X1 i_2_17_121 (.A(n_2_103), .ZN(n_2_17_109));
   AOI21_X1 i_2_17_122 (.A(n_2_17_108), .B1(n_2_17_109), .B2(n_2_183), .ZN(
      n_2_17_110));
   NAND2_X1 i_2_17_123 (.A1(n_2_103), .A2(n_2_197), .ZN(n_2_17_111));
   INV_X1 i_2_17_124 (.A(n_2_17_111), .ZN(n_2_17_112));
   NAND2_X1 i_2_17_125 (.A1(n_2_196), .A2(n_2_17_112), .ZN(n_2_17_113));
   INV_X1 i_2_17_126 (.A(n_2_17_113), .ZN(n_2_17_114));
   INV_X1 i_2_17_127 (.A(n_2_69), .ZN(n_2_17_115));
   NAND2_X1 i_2_17_128 (.A1(n_2_17_115), .A2(n_2_183), .ZN(n_2_17_116));
   NAND2_X1 i_2_17_129 (.A1(n_2_195), .A2(n_2_197), .ZN(n_2_17_117));
   INV_X1 i_2_17_130 (.A(n_2_17_117), .ZN(n_2_17_118));
   NAND3_X1 i_2_17_131 (.A1(n_2_69), .A2(n_2_103), .A3(n_2_17_118), .ZN(
      n_2_17_119));
   NAND2_X1 i_2_17_132 (.A1(n_2_17_116), .A2(n_2_17_119), .ZN(n_2_17_120));
   NOR2_X1 i_2_17_133 (.A1(n_2_17_114), .A2(n_2_17_120), .ZN(n_2_17_121));
   OAI21_X1 i_2_17_134 (.A(n_2_17_110), .B1(n_2_169), .B2(n_2_17_121), .ZN(n_52));
   HA_X1 i_2_18_0 (.A(n_2_18_79), .B(n_2_18_78), .CO(n_2_18_0), .S(n_2_209));
   HA_X1 i_2_18_1 (.A(n_2_18_80), .B(n_2_18_0), .CO(n_2_18_1), .S(n_2_210));
   HA_X1 i_2_18_2 (.A(n_2_18_81), .B(n_2_18_1), .CO(n_2_18_2), .S(n_2_211));
   HA_X1 i_2_18_3 (.A(n_2_18_82), .B(n_2_18_2), .CO(n_2_18_3), .S(n_2_212));
   HA_X1 i_2_18_4 (.A(Relative_Address[2]), .B(Relative_Address[1]), .CO(
      n_2_18_4), .S(n_2_185));
   HA_X1 i_2_18_5 (.A(Relative_Address[3]), .B(n_2_18_4), .CO(n_2_18_5), 
      .S(n_2_186));
   HA_X1 i_2_18_6 (.A(Relative_Address[6]), .B(n_2_18_154), .CO(n_2_18_6), 
      .S(n_2_189));
   HA_X1 i_2_18_7 (.A(Relative_Address[7]), .B(n_2_18_6), .CO(n_2_18_7), 
      .S(n_2_190));
   HA_X1 i_2_18_8 (.A(Relative_Address[8]), .B(n_2_18_7), .CO(n_2_18_8), 
      .S(n_2_191));
   HA_X1 i_2_18_9 (.A(Relative_Address[9]), .B(n_2_18_8), .CO(n_2_18_9), 
      .S(n_2_192));
   HA_X1 i_2_18_10 (.A(Relative_Address[10]), .B(n_2_18_9), .CO(n_2_18_10), 
      .S(n_2_193));
   HA_X1 i_2_18_11 (.A(Relative_Address[11]), .B(n_2_18_10), .CO(n_2_18_11), 
      .S(n_2_194));
   HA_X1 i_2_18_12 (.A(Relative_Address[12]), .B(n_2_18_11), .CO(n_2_18_12), 
      .S(n_2_195));
   HA_X1 i_2_18_13 (.A(Relative_Address[13]), .B(n_2_18_12), .CO(n_2_18_14), 
      .S(n_2_18_13));
   HA_X1 i_2_18_14 (.A(Relative_Address[14]), .B(n_2_18_14), .CO(n_2_18_16), 
      .S(n_2_18_15));
   HA_X1 i_2_18_15 (.A(RAM_Address[1]), .B(RAM_Address[0]), .CO(n_2_18_17), 
      .S(n_2_172));
   HA_X1 i_2_18_16 (.A(RAM_Address[2]), .B(n_2_18_17), .CO(n_2_18_18), .S(
      n_2_173));
   HA_X1 i_2_18_17 (.A(RAM_Address[3]), .B(n_2_18_18), .CO(n_2_18_19), .S(
      n_2_174));
   HA_X1 i_2_18_18 (.A(RAM_Address[4]), .B(n_2_18_19), .CO(n_2_18_20), .S(
      n_2_175));
   HA_X1 i_2_18_19 (.A(RAM_Address[5]), .B(n_2_18_20), .CO(n_2_18_21), .S(
      n_2_176));
   HA_X1 i_2_18_20 (.A(RAM_Address[6]), .B(n_2_18_21), .CO(n_2_18_22), .S(
      n_2_177));
   HA_X1 i_2_18_21 (.A(RAM_Address[7]), .B(n_2_18_22), .CO(n_2_18_23), .S(
      n_2_178));
   HA_X1 i_2_18_22 (.A(RAM_Address[8]), .B(n_2_18_23), .CO(n_2_18_24), .S(
      n_2_179));
   HA_X1 i_2_18_23 (.A(RAM_Address[9]), .B(n_2_18_24), .CO(n_2_18_25), .S(
      n_2_180));
   HA_X1 i_2_18_24 (.A(RAM_Address[10]), .B(n_2_18_25), .CO(n_2_18_26), .S(
      n_2_181));
   HA_X1 i_2_18_25 (.A(RAM_Address[11]), .B(n_2_18_26), .CO(n_2_18_27), .S(
      n_2_182));
   NOR2_X1 i_2_18_26 (.A1(Done_Loading), .A2(RST), .ZN(n_2_18_28));
   INV_X1 i_2_18_27 (.A(n_2_18_28), .ZN(n_2_199));
   INV_X1 i_2_18_28 (.A(InitCount[0]), .ZN(n_2_18_29));
   NAND2_X1 i_2_18_29 (.A1(n_2_18_29), .A2(InitCount[1]), .ZN(n_2_18_30));
   INV_X1 i_2_18_30 (.A(n_2_18_30), .ZN(n_2_198));
   NAND2_X1 i_2_18_31 (.A1(n_2_198), .A2(n_2_18_28), .ZN(n_2_18_31));
   INV_X1 i_2_18_32 (.A(n_2_18_31), .ZN(n_53));
   AND2_X1 i_2_18_33 (.A1(n_53), .A2(n_323), .ZN(n_54));
   INV_X1 i_2_18_34 (.A(n_2_227), .ZN(n_2_18_32));
   INV_X1 i_2_18_35 (.A(n_2_228), .ZN(n_2_18_33));
   AOI221_X1 i_2_18_36 (.A(n_2_18_32), .B1(CPU_Bus[27]), .B2(n_2_228), .C1(
      n_2_18_33), .C2(CPU_Bus[26]), .ZN(n_2_18_34));
   AOI221_X1 i_2_18_37 (.A(n_2_227), .B1(CPU_Bus[25]), .B2(n_2_228), .C1(
      CPU_Bus[24]), .C2(n_2_18_33), .ZN(n_2_18_35));
   AOI221_X1 i_2_18_38 (.A(n_2_18_32), .B1(CPU_Bus[31]), .B2(n_2_228), .C1(
      n_2_18_33), .C2(CPU_Bus[30]), .ZN(n_2_18_36));
   AOI221_X1 i_2_18_39 (.A(n_2_227), .B1(CPU_Bus[29]), .B2(n_2_228), .C1(
      CPU_Bus[28]), .C2(n_2_18_33), .ZN(n_2_18_37));
   INV_X1 i_2_18_40 (.A(n_2_226), .ZN(n_2_18_38));
   OAI33_X1 i_2_18_41 (.A1(n_2_18_34), .A2(n_2_18_35), .A3(n_2_226), .B1(
      n_2_18_36), .B2(n_2_18_37), .B3(n_2_18_38), .ZN(n_2_18_39));
   AOI221_X1 i_2_18_42 (.A(n_2_18_32), .B1(CPU_Bus[19]), .B2(n_2_228), .C1(
      n_2_18_33), .C2(CPU_Bus[18]), .ZN(n_2_18_40));
   AOI221_X1 i_2_18_43 (.A(n_2_227), .B1(CPU_Bus[17]), .B2(n_2_228), .C1(
      CPU_Bus[16]), .C2(n_2_18_33), .ZN(n_2_18_41));
   AOI221_X1 i_2_18_44 (.A(n_2_18_32), .B1(CPU_Bus[23]), .B2(n_2_228), .C1(
      n_2_18_33), .C2(CPU_Bus[22]), .ZN(n_2_18_42));
   AOI221_X1 i_2_18_45 (.A(n_2_227), .B1(CPU_Bus[21]), .B2(n_2_228), .C1(
      CPU_Bus[20]), .C2(n_2_18_33), .ZN(n_2_18_43));
   OAI33_X1 i_2_18_46 (.A1(n_2_18_40), .A2(n_2_18_41), .A3(n_2_226), .B1(
      n_2_18_42), .B2(n_2_18_43), .B3(n_2_18_38), .ZN(n_2_18_44));
   INV_X1 i_2_18_47 (.A(n_257), .ZN(n_2_18_45));
   AOI22_X1 i_2_18_48 (.A1(n_2_18_39), .A2(n_257), .B1(n_2_18_44), .B2(n_2_18_45), 
      .ZN(n_2_18_46));
   INV_X1 i_2_18_49 (.A(n_258), .ZN(n_2_18_47));
   INV_X1 i_2_18_50 (.A(CPU_Bus[7]), .ZN(n_2_18_48));
   INV_X1 i_2_18_51 (.A(CPU_Bus[6]), .ZN(n_2_18_49));
   AOI221_X1 i_2_18_52 (.A(n_2_18_32), .B1(n_2_18_48), .B2(n_2_228), .C1(
      n_2_18_49), .C2(n_2_18_33), .ZN(n_2_18_50));
   INV_X1 i_2_18_53 (.A(CPU_Bus[5]), .ZN(n_2_18_51));
   INV_X1 i_2_18_54 (.A(CPU_Bus[4]), .ZN(n_2_18_52));
   AOI221_X1 i_2_18_55 (.A(n_2_227), .B1(n_2_18_51), .B2(n_2_228), .C1(n_2_18_33), 
      .C2(n_2_18_52), .ZN(n_2_18_53));
   INV_X1 i_2_18_56 (.A(CPU_Bus[1]), .ZN(n_2_18_54));
   INV_X1 i_2_18_57 (.A(CPU_Bus[0]), .ZN(n_2_18_55));
   AOI221_X1 i_2_18_58 (.A(n_2_227), .B1(n_2_18_54), .B2(n_2_228), .C1(n_2_18_33), 
      .C2(n_2_18_55), .ZN(n_2_18_56));
   INV_X1 i_2_18_59 (.A(CPU_Bus[3]), .ZN(n_2_18_57));
   INV_X1 i_2_18_60 (.A(CPU_Bus[2]), .ZN(n_2_18_58));
   AOI221_X1 i_2_18_61 (.A(n_2_18_32), .B1(n_2_18_57), .B2(n_2_228), .C1(
      n_2_18_33), .C2(n_2_18_58), .ZN(n_2_18_59));
   OAI33_X1 i_2_18_62 (.A1(n_2_18_50), .A2(n_2_18_53), .A3(n_2_18_38), .B1(
      n_2_18_56), .B2(n_2_18_59), .B3(n_2_226), .ZN(n_2_18_60));
   AOI22_X1 i_2_18_63 (.A1(n_2_18_33), .A2(CPU_Bus[14]), .B1(CPU_Bus[15]), 
      .B2(n_2_228), .ZN(n_2_18_61));
   AOI22_X1 i_2_18_64 (.A1(n_2_18_33), .A2(CPU_Bus[12]), .B1(CPU_Bus[13]), 
      .B2(n_2_228), .ZN(n_2_18_62));
   OAI22_X1 i_2_18_65 (.A1(n_2_18_61), .A2(n_2_18_32), .B1(n_2_18_62), .B2(
      n_2_227), .ZN(n_2_18_63));
   AOI22_X1 i_2_18_66 (.A1(n_2_18_33), .A2(CPU_Bus[10]), .B1(CPU_Bus[11]), 
      .B2(n_2_228), .ZN(n_2_18_64));
   AOI22_X1 i_2_18_67 (.A1(n_2_18_33), .A2(CPU_Bus[8]), .B1(CPU_Bus[9]), 
      .B2(n_2_228), .ZN(n_2_18_65));
   OAI22_X1 i_2_18_68 (.A1(n_2_18_64), .A2(n_2_18_32), .B1(n_2_18_65), .B2(
      n_2_227), .ZN(n_2_18_66));
   AOI22_X1 i_2_18_69 (.A1(n_2_18_63), .A2(n_2_226), .B1(n_2_18_66), .B2(
      n_2_18_38), .ZN(n_2_18_67));
   OAI22_X1 i_2_18_70 (.A1(n_2_18_60), .A2(n_257), .B1(n_2_18_67), .B2(n_2_18_45), 
      .ZN(n_2_18_68));
   INV_X1 i_2_18_71 (.A(n_2_18_68), .ZN(n_2_18_69));
   OAI22_X1 i_2_18_72 (.A1(n_2_18_46), .A2(n_2_18_47), .B1(n_2_18_69), .B2(n_258), 
      .ZN(n_2_18_70));
   NAND2_X1 i_2_18_73 (.A1(n_2_18_70), .A2(Row_Done_Bit_Delayed), .ZN(n_2_18_71));
   INV_X1 i_2_18_74 (.A(n_2_18_71), .ZN(n_2_18_72));
   INV_X1 i_2_18_75 (.A(Row_Done_Bit_Delayed), .ZN(n_2_18_73));
   AOI21_X1 i_2_18_76 (.A(n_2_18_72), .B1(Row_Last_Bit), .B2(n_2_18_73), 
      .ZN(n_2_18_74));
   INV_X1 i_2_18_77 (.A(n_2_18_74), .ZN(n_2_18_75));
   INV_X1 i_2_18_78 (.A(n_2_18_70), .ZN(n_2_18_76));
   OAI22_X1 i_2_18_79 (.A1(n_2_18_70), .A2(n_2_18_75), .B1(n_2_18_74), .B2(
      n_2_18_76), .ZN(n_2_18_77));
   OAI33_X1 i_2_18_80 (.A1(n_2_18_77), .A2(Row_Done_Bit), .A3(n_2_18_31), 
      .B1(n_2_199), .B2(InitCount[0]), .B3(InitCount[1]), .ZN(n_55));
   INV_X1 i_2_18_81 (.A(n_2_71), .ZN(n_2_18_78));
   NOR2_X1 i_2_18_82 (.A1(n_2_199), .A2(n_2_18_78), .ZN(n_56));
   INV_X1 i_2_18_83 (.A(n_2_72), .ZN(n_2_18_79));
   NOR2_X1 i_2_18_84 (.A1(n_2_199), .A2(n_2_18_79), .ZN(n_57));
   INV_X1 i_2_18_85 (.A(n_2_73), .ZN(n_2_18_80));
   NOR2_X1 i_2_18_86 (.A1(n_2_199), .A2(n_2_18_80), .ZN(n_58));
   INV_X1 i_2_18_87 (.A(n_2_74), .ZN(n_2_18_81));
   NOR2_X1 i_2_18_88 (.A1(n_2_199), .A2(n_2_18_81), .ZN(n_59));
   INV_X1 i_2_18_89 (.A(n_2_75), .ZN(n_2_18_82));
   NOR2_X1 i_2_18_90 (.A1(n_2_199), .A2(n_2_18_82), .ZN(n_60));
   AND2_X1 i_2_18_91 (.A1(n_2_18_28), .A2(n_2_76), .ZN(n_61));
   AND2_X1 i_2_18_92 (.A1(n_2_18_28), .A2(n_2_77), .ZN(n_62));
   AND2_X1 i_2_18_93 (.A1(n_2_18_28), .A2(n_2_78), .ZN(n_63));
   AND2_X1 i_2_18_94 (.A1(n_2_18_28), .A2(n_2_79), .ZN(n_64));
   AND2_X1 i_2_18_95 (.A1(n_2_18_28), .A2(n_2_80), .ZN(n_65));
   AND2_X1 i_2_18_96 (.A1(n_2_18_28), .A2(n_2_81), .ZN(n_66));
   AND2_X1 i_2_18_97 (.A1(n_2_18_28), .A2(n_2_82), .ZN(n_67));
   AND2_X1 i_2_18_98 (.A1(n_2_18_28), .A2(n_2_83), .ZN(n_68));
   AND2_X1 i_2_18_99 (.A1(n_2_18_28), .A2(n_2_84), .ZN(n_69));
   AND2_X1 i_2_18_100 (.A1(n_2_18_28), .A2(n_2_85), .ZN(n_70));
   AND2_X1 i_2_18_101 (.A1(n_2_18_28), .A2(n_2_86), .ZN(n_71));
   AND2_X1 i_2_18_102 (.A1(n_2_18_28), .A2(n_2_87), .ZN(n_72));
   AND2_X1 i_2_18_103 (.A1(n_2_18_28), .A2(n_2_88), .ZN(n_73));
   AND2_X1 i_2_18_104 (.A1(n_2_18_28), .A2(n_2_89), .ZN(n_74));
   AND2_X1 i_2_18_105 (.A1(n_2_18_28), .A2(n_2_90), .ZN(n_75));
   AND2_X1 i_2_18_106 (.A1(n_2_18_28), .A2(n_2_91), .ZN(n_76));
   AND2_X1 i_2_18_107 (.A1(n_2_18_28), .A2(n_2_92), .ZN(n_77));
   AND2_X1 i_2_18_108 (.A1(n_2_18_28), .A2(n_2_93), .ZN(n_78));
   AND2_X1 i_2_18_109 (.A1(n_2_18_28), .A2(n_2_94), .ZN(n_79));
   AND2_X1 i_2_18_110 (.A1(n_2_18_28), .A2(n_2_95), .ZN(n_80));
   AND2_X1 i_2_18_111 (.A1(n_2_18_28), .A2(n_2_96), .ZN(n_81));
   AND2_X1 i_2_18_112 (.A1(n_2_18_28), .A2(n_2_97), .ZN(n_82));
   AND2_X1 i_2_18_113 (.A1(n_2_18_28), .A2(n_2_98), .ZN(n_83));
   AND2_X1 i_2_18_114 (.A1(n_2_18_28), .A2(n_2_99), .ZN(n_84));
   AND2_X1 i_2_18_115 (.A1(n_2_18_28), .A2(n_2_100), .ZN(n_85));
   AND2_X1 i_2_18_116 (.A1(n_2_18_28), .A2(n_2_101), .ZN(n_86));
   AND2_X1 i_2_18_117 (.A1(n_2_18_28), .A2(n_2_102), .ZN(n_87));
   NOR2_X1 i_2_18_118 (.A1(InitCount[0]), .A2(InitCount[1]), .ZN(n_2_18_83));
   INV_X1 i_2_18_119 (.A(n_2_18_83), .ZN(n_2_18_84));
   OAI22_X1 i_2_18_120 (.A1(n_2_18_84), .A2(CPU_Bus[0]), .B1(n_2_18_83), 
      .B2(PacketSize[0]), .ZN(n_2_18_85));
   NOR2_X1 i_2_18_121 (.A1(n_2_18_85), .A2(n_2_199), .ZN(n_88));
   OAI22_X1 i_2_18_122 (.A1(n_2_18_84), .A2(CPU_Bus[1]), .B1(n_2_18_83), 
      .B2(PacketSize[1]), .ZN(n_2_18_86));
   NOR2_X1 i_2_18_123 (.A1(n_2_18_86), .A2(n_2_199), .ZN(n_89));
   OAI22_X1 i_2_18_124 (.A1(n_2_18_84), .A2(CPU_Bus[2]), .B1(n_2_18_83), 
      .B2(PacketSize[2]), .ZN(n_2_18_87));
   NOR2_X1 i_2_18_125 (.A1(n_2_18_87), .A2(n_2_199), .ZN(n_90));
   OAI22_X1 i_2_18_126 (.A1(n_2_18_84), .A2(CPU_Bus[3]), .B1(n_2_18_83), 
      .B2(PacketSize[3]), .ZN(n_2_18_88));
   NOR2_X1 i_2_18_127 (.A1(n_2_18_88), .A2(n_2_199), .ZN(n_91));
   OAI22_X1 i_2_18_128 (.A1(n_2_18_84), .A2(CPU_Bus[4]), .B1(n_2_18_83), 
      .B2(PacketSize[4]), .ZN(n_2_18_89));
   NOR2_X1 i_2_18_129 (.A1(n_2_18_89), .A2(n_2_199), .ZN(n_92));
   OAI22_X1 i_2_18_130 (.A1(n_2_18_84), .A2(CPU_Bus[5]), .B1(n_2_18_83), 
      .B2(PacketSize[5]), .ZN(n_2_18_90));
   NOR2_X1 i_2_18_131 (.A1(n_2_18_90), .A2(n_2_199), .ZN(n_93));
   AND2_X1 i_2_18_132 (.A1(n_2_18_28), .A2(n_2_124), .ZN(n_94));
   AND2_X1 i_2_18_133 (.A1(n_2_18_28), .A2(n_2_125), .ZN(n_95));
   AND2_X1 i_2_18_134 (.A1(n_2_18_28), .A2(n_2_126), .ZN(n_96));
   AND2_X1 i_2_18_135 (.A1(n_2_18_28), .A2(n_2_127), .ZN(n_97));
   AND2_X1 i_2_18_136 (.A1(n_2_18_28), .A2(n_2_128), .ZN(n_98));
   AND2_X1 i_2_18_137 (.A1(n_2_18_28), .A2(n_2_129), .ZN(n_99));
   AND2_X1 i_2_18_138 (.A1(n_2_18_28), .A2(n_2_130), .ZN(n_100));
   AND2_X1 i_2_18_139 (.A1(n_2_18_28), .A2(n_2_131), .ZN(n_101));
   AND2_X1 i_2_18_140 (.A1(n_2_18_28), .A2(n_2_132), .ZN(n_102));
   AND2_X1 i_2_18_141 (.A1(n_2_18_28), .A2(n_2_133), .ZN(n_103));
   AND2_X1 i_2_18_142 (.A1(n_2_18_28), .A2(n_2_134), .ZN(n_104));
   AND2_X1 i_2_18_143 (.A1(n_2_18_28), .A2(n_2_135), .ZN(n_105));
   AND2_X1 i_2_18_144 (.A1(n_2_18_28), .A2(n_2_136), .ZN(n_106));
   AND2_X1 i_2_18_145 (.A1(n_2_18_28), .A2(n_2_137), .ZN(n_107));
   AND2_X1 i_2_18_146 (.A1(n_2_18_28), .A2(n_2_138), .ZN(n_108));
   AND2_X1 i_2_18_147 (.A1(n_2_18_28), .A2(n_2_139), .ZN(n_109));
   AND2_X1 i_2_18_148 (.A1(n_2_18_28), .A2(n_2_140), .ZN(n_110));
   AND2_X1 i_2_18_149 (.A1(n_2_18_28), .A2(n_2_141), .ZN(n_111));
   AND2_X1 i_2_18_150 (.A1(n_2_18_28), .A2(n_2_142), .ZN(n_112));
   AND2_X1 i_2_18_151 (.A1(n_2_18_28), .A2(n_2_143), .ZN(n_113));
   AND2_X1 i_2_18_152 (.A1(n_2_18_28), .A2(n_2_144), .ZN(n_114));
   AND2_X1 i_2_18_153 (.A1(n_2_18_28), .A2(n_2_145), .ZN(n_115));
   AND2_X1 i_2_18_154 (.A1(n_2_18_28), .A2(n_2_146), .ZN(n_116));
   AND2_X1 i_2_18_155 (.A1(n_2_18_28), .A2(n_2_147), .ZN(n_117));
   AND2_X1 i_2_18_156 (.A1(n_2_18_28), .A2(n_2_148), .ZN(n_118));
   AND2_X1 i_2_18_157 (.A1(n_2_18_28), .A2(n_2_149), .ZN(n_119));
   AND2_X1 i_2_18_158 (.A1(n_2_18_28), .A2(n_2_150), .ZN(n_120));
   AND2_X1 i_2_18_159 (.A1(n_2_18_28), .A2(n_2_151), .ZN(n_121));
   AND2_X1 i_2_18_160 (.A1(n_2_18_28), .A2(n_2_152), .ZN(n_122));
   AND2_X1 i_2_18_161 (.A1(n_2_18_28), .A2(n_2_153), .ZN(n_123));
   AND2_X1 i_2_18_162 (.A1(n_2_18_28), .A2(n_2_154), .ZN(n_124));
   AND2_X1 i_2_18_163 (.A1(n_2_18_28), .A2(n_2_155), .ZN(n_125));
   NAND2_X1 i_2_18_164 (.A1(n_2_18_30), .A2(n_2_18_28), .ZN(n_126));
   INV_X1 i_2_18_165 (.A(n_2_18_85), .ZN(n_2_18_91));
   OAI22_X1 i_2_18_166 (.A1(n_2_18_91), .A2(n_126), .B1(n_2_18_31), .B2(
      n_2_18_33), .ZN(n_127));
   NAND2_X1 i_2_18_167 (.A1(n_2_18_85), .A2(n_2_18_86), .ZN(n_2_18_92));
   OAI21_X1 i_2_18_168 (.A(n_2_18_92), .B1(n_2_18_85), .B2(n_2_18_86), .ZN(
      n_2_18_93));
   INV_X1 i_2_18_169 (.A(n_126), .ZN(n_2_18_94));
   AOI22_X1 i_2_18_170 (.A1(n_2_18_93), .A2(n_2_18_94), .B1(n_53), .B2(n_2_227), 
      .ZN(n_2_18_95));
   INV_X1 i_2_18_171 (.A(n_2_18_95), .ZN(n_128));
   INV_X1 i_2_18_172 (.A(n_2_18_92), .ZN(n_2_18_96));
   NAND2_X1 i_2_18_173 (.A1(n_2_18_96), .A2(n_2_18_87), .ZN(n_2_18_97));
   OAI21_X1 i_2_18_174 (.A(n_2_18_97), .B1(n_2_18_87), .B2(n_2_18_96), .ZN(
      n_2_18_98));
   AOI22_X1 i_2_18_175 (.A1(n_2_18_98), .A2(n_2_18_94), .B1(n_53), .B2(n_2_226), 
      .ZN(n_2_18_99));
   INV_X1 i_2_18_176 (.A(n_2_18_99), .ZN(n_129));
   INV_X1 i_2_18_177 (.A(n_2_18_97), .ZN(n_2_18_100));
   NAND2_X1 i_2_18_178 (.A1(n_2_18_100), .A2(n_2_18_88), .ZN(n_2_18_101));
   OAI21_X1 i_2_18_179 (.A(n_2_18_101), .B1(n_2_18_88), .B2(n_2_18_100), 
      .ZN(n_2_18_102));
   AOI22_X1 i_2_18_180 (.A1(n_2_18_102), .A2(n_2_18_94), .B1(n_53), .B2(n_257), 
      .ZN(n_2_18_103));
   INV_X1 i_2_18_181 (.A(n_2_18_103), .ZN(n_130));
   XNOR2_X1 i_2_18_182 (.A(n_2_18_101), .B(n_2_18_89), .ZN(n_2_18_104));
   OAI22_X1 i_2_18_183 (.A1(n_2_18_104), .A2(n_126), .B1(n_2_18_31), .B2(
      n_2_18_47), .ZN(n_131));
   INV_X1 i_2_18_184 (.A(n_2_18_101), .ZN(n_2_18_105));
   AND3_X1 i_2_18_185 (.A1(n_2_18_105), .A2(n_2_18_89), .A3(n_2_18_90), .ZN(
      n_2_18_106));
   AOI21_X1 i_2_18_186 (.A(n_2_18_90), .B1(n_2_18_105), .B2(n_2_18_89), .ZN(
      n_2_18_107));
   INV_X1 i_2_18_187 (.A(n_2_229), .ZN(n_2_18_108));
   OAI33_X1 i_2_18_188 (.A1(n_2_18_106), .A2(n_2_18_107), .A3(n_126), .B1(
      n_2_199), .B2(n_2_18_30), .B3(n_2_18_108), .ZN(n_132));
   NOR2_X1 i_2_18_189 (.A1(n_2_18_74), .A2(n_2_199), .ZN(n_133));
   INV_X1 i_2_18_190 (.A(InitCount[1]), .ZN(n_2_18_109));
   AOI21_X1 i_2_18_191 (.A(n_2_199), .B1(InitCount[0]), .B2(n_2_18_109), 
      .ZN(n_2_18_110));
   NOR3_X1 i_2_18_192 (.A1(n_2_199), .A2(n_2_18_29), .A3(InitCount[1]), .ZN(
      n_2_18_111));
   AOI22_X1 i_2_18_193 (.A1(n_2_18_110), .A2(RowsNum[0]), .B1(n_2_18_111), 
      .B2(CPU_Bus[0]), .ZN(n_2_18_112));
   INV_X1 i_2_18_194 (.A(n_2_18_112), .ZN(n_134));
   AOI22_X1 i_2_18_195 (.A1(n_2_18_110), .A2(RowsNum[1]), .B1(n_2_18_111), 
      .B2(CPU_Bus[1]), .ZN(n_2_18_113));
   INV_X1 i_2_18_196 (.A(n_2_18_113), .ZN(n_135));
   AOI22_X1 i_2_18_197 (.A1(n_2_18_110), .A2(RowsNum[2]), .B1(n_2_18_111), 
      .B2(CPU_Bus[2]), .ZN(n_2_18_114));
   INV_X1 i_2_18_198 (.A(n_2_18_114), .ZN(n_136));
   AOI22_X1 i_2_18_199 (.A1(n_2_18_110), .A2(RowsNum[3]), .B1(n_2_18_111), 
      .B2(CPU_Bus[3]), .ZN(n_2_18_115));
   INV_X1 i_2_18_200 (.A(n_2_18_115), .ZN(n_137));
   AOI22_X1 i_2_18_201 (.A1(n_2_18_110), .A2(RowsNum[4]), .B1(n_2_18_111), 
      .B2(CPU_Bus[4]), .ZN(n_2_18_116));
   INV_X1 i_2_18_202 (.A(n_2_18_116), .ZN(n_138));
   AOI22_X1 i_2_18_203 (.A1(n_2_18_110), .A2(RowsNum[5]), .B1(n_2_18_111), 
      .B2(CPU_Bus[5]), .ZN(n_2_18_117));
   INV_X1 i_2_18_204 (.A(n_2_18_117), .ZN(n_139));
   AOI22_X1 i_2_18_205 (.A1(n_2_18_110), .A2(RowsNum[6]), .B1(n_2_18_111), 
      .B2(CPU_Bus[6]), .ZN(n_2_18_118));
   INV_X1 i_2_18_206 (.A(n_2_18_118), .ZN(n_140));
   AOI22_X1 i_2_18_207 (.A1(n_2_18_110), .A2(RowsNum[7]), .B1(n_2_18_111), 
      .B2(CPU_Bus[7]), .ZN(n_2_18_119));
   INV_X1 i_2_18_208 (.A(n_2_18_119), .ZN(n_141));
   AOI22_X1 i_2_18_209 (.A1(n_2_18_110), .A2(RowsNum[8]), .B1(n_2_18_111), 
      .B2(CPU_Bus[8]), .ZN(n_2_18_120));
   INV_X1 i_2_18_210 (.A(n_2_18_120), .ZN(n_142));
   AOI22_X1 i_2_18_211 (.A1(n_2_18_110), .A2(RowsNum[9]), .B1(n_2_18_111), 
      .B2(CPU_Bus[9]), .ZN(n_2_18_121));
   INV_X1 i_2_18_212 (.A(n_2_18_121), .ZN(n_143));
   AOI22_X1 i_2_18_213 (.A1(n_2_18_110), .A2(RowsNum[10]), .B1(n_2_18_111), 
      .B2(CPU_Bus[10]), .ZN(n_2_18_122));
   INV_X1 i_2_18_214 (.A(n_2_18_122), .ZN(n_144));
   AOI22_X1 i_2_18_215 (.A1(n_2_18_110), .A2(RowsNum[11]), .B1(n_2_18_111), 
      .B2(CPU_Bus[11]), .ZN(n_2_18_123));
   INV_X1 i_2_18_216 (.A(n_2_18_123), .ZN(n_145));
   AOI22_X1 i_2_18_217 (.A1(n_2_18_110), .A2(RowsNum[12]), .B1(n_2_18_111), 
      .B2(CPU_Bus[12]), .ZN(n_2_18_124));
   INV_X1 i_2_18_218 (.A(n_2_18_124), .ZN(n_146));
   AOI22_X1 i_2_18_219 (.A1(n_2_18_110), .A2(RowsNum[13]), .B1(n_2_18_111), 
      .B2(CPU_Bus[13]), .ZN(n_2_18_125));
   INV_X1 i_2_18_220 (.A(n_2_18_125), .ZN(n_147));
   AOI22_X1 i_2_18_221 (.A1(n_2_18_110), .A2(RowsNum[14]), .B1(n_2_18_111), 
      .B2(CPU_Bus[14]), .ZN(n_2_18_126));
   INV_X1 i_2_18_222 (.A(n_2_18_126), .ZN(n_148));
   AOI22_X1 i_2_18_223 (.A1(n_2_18_110), .A2(RowsNum[15]), .B1(n_2_18_111), 
      .B2(CPU_Bus[15]), .ZN(n_2_18_127));
   INV_X1 i_2_18_224 (.A(n_2_18_127), .ZN(n_149));
   OR2_X1 i_2_18_225 (.A1(n_2_18_28), .A2(RST), .ZN(n_150));
   INV_X1 i_2_18_226 (.A(PacketSize[0]), .ZN(n_151));
   AOI22_X1 i_2_18_227 (.A1(n_2_18_32), .A2(n_32), .B1(n_2_18_108), .B2(n_36), 
      .ZN(n_2_18_128));
   OAI221_X1 i_2_18_228 (.A(n_2_18_128), .B1(n_2_18_108), .B2(n_36), .C1(
      n_2_18_33), .C2(n_151), .ZN(n_2_18_129));
   INV_X1 i_2_18_229 (.A(n_324), .ZN(n_2_18_130));
   NOR2_X1 i_2_18_230 (.A1(n_2_18_32), .A2(n_32), .ZN(n_2_18_131));
   NOR4_X1 i_2_18_231 (.A1(n_2_18_129), .A2(n_2_18_130), .A3(n_37), .A4(
      n_2_18_131), .ZN(n_2_18_132));
   AOI222_X1 i_2_18_232 (.A1(n_2_18_38), .A2(n_33), .B1(n_2_18_33), .B2(n_151), 
      .C1(n_2_18_47), .C2(n_35), .ZN(n_2_18_133));
   OAI22_X1 i_2_18_233 (.A1(n_2_18_38), .A2(n_33), .B1(n_2_18_45), .B2(n_34), 
      .ZN(n_2_18_134));
   INV_X1 i_2_18_234 (.A(n_35), .ZN(n_2_18_135));
   AOI221_X1 i_2_18_235 (.A(n_2_18_134), .B1(n_2_18_45), .B2(n_34), .C1(
      n_2_18_135), .C2(n_258), .ZN(n_2_18_136));
   NAND3_X1 i_2_18_236 (.A1(n_2_18_132), .A2(n_2_18_133), .A3(n_2_18_136), 
      .ZN(n_2_18_137));
   NAND2_X1 i_2_18_237 (.A1(n_2_18_137), .A2(n_2_18_28), .ZN(n_152));
   XOR2_X1 i_2_18_238 (.A(RAM_Address[12]), .B(n_2_18_27), .Z(n_2_183));
   INV_X1 i_2_18_239 (.A(n_2_103), .ZN(n_2_18_138));
   INV_X1 i_2_18_240 (.A(N_Indication_Bit), .ZN(n_2_18_139));
   AOI21_X1 i_2_18_241 (.A(n_2_199), .B1(n_2_18_138), .B2(n_2_18_139), .ZN(n_153));
   NOR2_X1 i_2_18_242 (.A1(n_2_199), .A2(n_2_18_138), .ZN(n_154));
   NAND3_X1 i_2_18_243 (.A1(n_53), .A2(n_2_18_138), .A3(n_2_71), .ZN(n_155));
   NAND3_X1 i_2_18_244 (.A1(n_53), .A2(n_2_18_138), .A3(n_2_72), .ZN(n_156));
   NAND3_X1 i_2_18_245 (.A1(n_53), .A2(n_2_18_138), .A3(n_2_73), .ZN(n_157));
   NAND3_X1 i_2_18_246 (.A1(n_53), .A2(n_2_18_138), .A3(n_2_74), .ZN(n_158));
   NAND3_X1 i_2_18_247 (.A1(n_53), .A2(n_2_18_138), .A3(n_2_75), .ZN(n_159));
   NAND3_X1 i_2_18_248 (.A1(n_53), .A2(n_2_18_138), .A3(n_2_76), .ZN(n_160));
   INV_X1 i_2_18_249 (.A(Done_Element), .ZN(n_2_18_140));
   OAI211_X1 i_2_18_250 (.A(n_2_18_71), .B(n_2_18_140), .C1(Data_Bit), .C2(
      Row_Done_Bit_Delayed), .ZN(n_2_18_141));
   OAI21_X1 i_2_18_251 (.A(n_2_18_141), .B1(n_2_18_140), .B2(Data_Bit), .ZN(
      n_2_18_142));
   NOR2_X1 i_2_18_252 (.A1(n_2_18_427), .A2(n_2_199), .ZN(n_161));
   INV_X1 i_2_18_253 (.A(n_2_112), .ZN(n_2_18_143));
   NOR2_X1 i_2_18_254 (.A1(n_2_199), .A2(n_2_18_143), .ZN(n_162));
   AND2_X1 i_2_18_255 (.A1(n_2_18_28), .A2(n_2_113), .ZN(n_163));
   AND2_X1 i_2_18_256 (.A1(n_2_18_28), .A2(n_2_114), .ZN(n_164));
   INV_X1 i_2_18_257 (.A(n_2_115), .ZN(n_2_18_144));
   NOR2_X1 i_2_18_258 (.A1(n_2_199), .A2(n_2_18_144), .ZN(n_165));
   AND2_X1 i_2_18_259 (.A1(n_2_18_28), .A2(n_2_116), .ZN(n_166));
   INV_X1 i_2_18_260 (.A(n_2_117), .ZN(n_2_18_145));
   NOR2_X1 i_2_18_261 (.A1(n_2_199), .A2(n_2_18_145), .ZN(n_167));
   INV_X1 i_2_18_262 (.A(n_2_118), .ZN(n_2_18_146));
   NOR2_X1 i_2_18_263 (.A1(n_2_199), .A2(n_2_18_146), .ZN(n_168));
   AND2_X1 i_2_18_264 (.A1(n_2_18_28), .A2(n_2_119), .ZN(n_169));
   AND2_X1 i_2_18_265 (.A1(n_2_18_28), .A2(n_2_120), .ZN(n_170));
   INV_X1 i_2_18_266 (.A(n_2_121), .ZN(n_2_18_147));
   NOR2_X1 i_2_18_267 (.A1(n_2_199), .A2(n_2_18_147), .ZN(n_171));
   INV_X1 i_2_18_268 (.A(n_2_122), .ZN(n_2_18_148));
   NOR2_X1 i_2_18_269 (.A1(n_2_199), .A2(n_2_18_148), .ZN(n_172));
   INV_X1 i_2_18_270 (.A(n_2_123), .ZN(n_2_18_149));
   NOR2_X1 i_2_18_271 (.A1(n_2_199), .A2(n_2_18_149), .ZN(n_173));
   NAND2_X1 i_2_18_272 (.A1(n_2_18_28), .A2(Relative_Address[1]), .ZN(n_174));
   OR2_X1 i_2_18_273 (.A1(n_2_199), .A2(n_2_185), .ZN(n_175));
   OR2_X1 i_2_18_274 (.A1(n_2_199), .A2(n_2_186), .ZN(n_176));
   NOR2_X1 i_2_18_275 (.A1(Relative_Address[4]), .A2(n_2_18_5), .ZN(n_2_18_150));
   AOI21_X1 i_2_18_276 (.A(n_2_18_150), .B1(Relative_Address[4]), .B2(n_2_18_5), 
      .ZN(n_2_18_151));
   NOR2_X1 i_2_18_277 (.A1(n_2_18_151), .A2(n_2_199), .ZN(n_177));
   INV_X1 i_2_18_278 (.A(n_2_18_150), .ZN(n_2_18_152));
   NOR2_X1 i_2_18_279 (.A1(n_2_18_152), .A2(Relative_Address[5]), .ZN(n_2_18_153));
   INV_X1 i_2_18_280 (.A(n_2_18_153), .ZN(n_2_18_154));
   AOI21_X1 i_2_18_281 (.A(n_2_18_153), .B1(Relative_Address[5]), .B2(n_2_18_152), 
      .ZN(n_2_18_155));
   INV_X1 i_2_18_282 (.A(n_2_18_155), .ZN(n_2_188));
   NOR2_X1 i_2_18_283 (.A1(n_2_18_155), .A2(n_2_199), .ZN(n_178));
   AND2_X1 i_2_18_284 (.A1(n_2_18_28), .A2(n_2_189), .ZN(n_179));
   OR2_X1 i_2_18_285 (.A1(n_2_199), .A2(n_2_190), .ZN(n_180));
   OR2_X1 i_2_18_286 (.A1(n_2_199), .A2(n_2_191), .ZN(n_181));
   OR2_X1 i_2_18_287 (.A1(n_2_199), .A2(n_2_192), .ZN(n_182));
   AND2_X1 i_2_18_288 (.A1(n_2_18_28), .A2(n_2_193), .ZN(n_183));
   AND2_X1 i_2_18_289 (.A1(n_2_18_28), .A2(n_2_194), .ZN(n_184));
   OR2_X1 i_2_18_290 (.A1(n_2_199), .A2(n_2_195), .ZN(n_185));
   AND2_X1 i_2_18_291 (.A1(n_2_18_28), .A2(n_2_18_13), .ZN(n_186));
   AND2_X1 i_2_18_292 (.A1(n_2_18_28), .A2(n_2_18_15), .ZN(n_187));
   INV_X1 i_2_18_293 (.A(Relative_Address[15]), .ZN(n_2_18_156));
   INV_X1 i_2_18_294 (.A(n_2_18_16), .ZN(n_2_18_157));
   AOI221_X1 i_2_18_295 (.A(n_2_199), .B1(n_2_18_156), .B2(n_2_18_157), .C1(
      Relative_Address[15]), .C2(n_2_18_16), .ZN(n_188));
   INV_X1 i_2_18_296 (.A(n_2_18_151), .ZN(n_2_187));
   XOR2_X1 i_2_18_297 (.A(n_2_114), .B(RowsCount[3]), .Z(n_2_18_158));
   INV_X1 i_2_18_298 (.A(RowsCount[11]), .ZN(n_2_18_159));
   AOI221_X1 i_2_18_299 (.A(n_2_18_158), .B1(n_2_18_159), .B2(n_2_122), .C1(
      RowsCount[11]), .C2(n_2_18_148), .ZN(n_2_18_160));
   XOR2_X1 i_2_18_300 (.A(n_2_116), .B(RowsCount[5]), .Z(n_2_18_161));
   INV_X1 i_2_18_301 (.A(RowsCount[7]), .ZN(n_2_18_162));
   AOI221_X1 i_2_18_302 (.A(n_2_18_161), .B1(n_2_18_162), .B2(n_2_118), .C1(
      RowsCount[7]), .C2(n_2_18_146), .ZN(n_2_18_163));
   XOR2_X1 i_2_18_303 (.A(n_2_113), .B(RowsCount[2]), .Z(n_2_18_164));
   INV_X1 i_2_18_304 (.A(RowsCount[10]), .ZN(n_2_18_165));
   AOI221_X1 i_2_18_305 (.A(n_2_18_164), .B1(n_2_18_165), .B2(n_2_121), .C1(
      RowsCount[10]), .C2(n_2_18_147), .ZN(n_2_18_166));
   INV_X1 i_2_18_306 (.A(RowsCount[0]), .ZN(n_2_18_167));
   NOR4_X1 i_2_18_307 (.A1(n_2_18_167), .A2(RowsCount[15]), .A3(RowsCount[14]), 
      .A4(RowsCount[13]), .ZN(n_2_18_168));
   NAND4_X1 i_2_18_308 (.A1(n_2_18_160), .A2(n_2_18_163), .A3(n_2_18_166), 
      .A4(n_2_18_168), .ZN(n_2_18_169));
   AOI22_X1 i_2_18_309 (.A1(n_2_18_145), .A2(RowsCount[6]), .B1(n_2_18_149), 
      .B2(RowsCount[12]), .ZN(n_2_18_170));
   OAI221_X1 i_2_18_310 (.A(n_2_18_170), .B1(n_2_18_149), .B2(RowsCount[12]), 
      .C1(n_2_18_145), .C2(RowsCount[6]), .ZN(n_2_18_171));
   XNOR2_X1 i_2_18_311 (.A(n_2_120), .B(RowsCount[9]), .ZN(n_2_18_172));
   INV_X1 i_2_18_312 (.A(RowsCount[1]), .ZN(n_2_18_173));
   OAI221_X1 i_2_18_313 (.A(n_2_18_172), .B1(n_2_18_143), .B2(RowsCount[1]), 
      .C1(n_2_18_173), .C2(n_2_112), .ZN(n_2_18_174));
   XNOR2_X1 i_2_18_314 (.A(n_2_119), .B(RowsCount[8]), .ZN(n_2_18_175));
   INV_X1 i_2_18_315 (.A(RowsCount[4]), .ZN(n_2_18_176));
   OAI221_X1 i_2_18_316 (.A(n_2_18_175), .B1(n_2_18_144), .B2(RowsCount[4]), 
      .C1(n_2_18_176), .C2(n_2_115), .ZN(n_2_18_177));
   NOR4_X1 i_2_18_317 (.A1(n_2_18_169), .A2(n_2_18_171), .A3(n_2_18_174), 
      .A4(n_2_18_177), .ZN(n_2_196));
   OR2_X1 i_2_18_318 (.A1(Row_Done_Bit_Delayed), .A2(
      Update_Address_Indication_Bit), .ZN(n_2_197));
   OAI21_X1 i_2_18_319 (.A(n_2_18_28), .B1(n_2_18_31), .B2(n_2_18_138), .ZN(
      n_189));
   NOR2_X1 i_2_18_320 (.A1(n_2_18_142), .A2(n_2_199), .ZN(n_190));
   AND2_X1 i_2_18_321 (.A1(n_2_18_28), .A2(n_2_111), .ZN(n_191));
   AND2_X1 i_2_18_322 (.A1(n_2_104), .A2(n_2_105), .ZN(n_2_18_178));
   NOR2_X1 i_2_18_323 (.A1(Writing_Start_Index[1]), .A2(Writing_Start_Index[2]), 
      .ZN(n_2_18_179));
   INV_X1 i_2_18_324 (.A(n_2_18_179), .ZN(n_2_18_180));
   NOR2_X1 i_2_18_325 (.A1(n_2_18_180), .A2(Writing_Start_Index[3]), .ZN(
      n_2_18_181));
   NOR2_X1 i_2_18_326 (.A1(Writing_Start_Index[4]), .A2(Writing_Start_Index[5]), 
      .ZN(n_2_18_182));
   NOR2_X1 i_2_18_327 (.A1(n_2_18_424), .A2(n_2_199), .ZN(n_192));
   OR2_X1 i_2_18_328 (.A1(Writing_Start_Index[3]), .A2(Writing_Start_Index[2]), 
      .ZN(n_2_18_183));
   NOR2_X1 i_2_18_329 (.A1(n_2_18_183), .A2(Writing_Start_Index[4]), .ZN(
      n_2_18_184));
   INV_X1 i_2_18_330 (.A(Writing_Start_Index[5]), .ZN(n_2_18_185));
   AND2_X1 i_2_18_331 (.A1(n_2_18_184), .A2(n_2_18_185), .ZN(n_2_18_186));
   NAND2_X1 i_2_18_332 (.A1(Writing_Start_Index[0]), .A2(Writing_Start_Index[1]), 
      .ZN(n_2_18_187));
   AOI211_X1 i_2_18_333 (.A(n_2_106), .B(n_2_18_439), .C1(n_2_18_186), .C2(
      n_2_18_187), .ZN(n_2_18_188));
   INV_X1 i_2_18_334 (.A(n_2_18_188), .ZN(n_2_18_189));
   OAI22_X1 i_2_18_335 (.A1(n_2_215), .A2(n_2_18_189), .B1(n_2_18_188), .B2(
      n_267), .ZN(n_2_18_190));
   INV_X1 i_2_18_336 (.A(n_2_18_190), .ZN(n_2_217));
   NOR2_X1 i_2_18_337 (.A1(n_2_18_190), .A2(n_2_199), .ZN(n_193));
   NOR2_X1 i_2_18_338 (.A1(n_2_18_431), .A2(n_2_18_432), .ZN(n_2_18_191));
   OR3_X1 i_2_18_339 (.A1(n_2_18_186), .A2(n_2_18_439), .A3(n_2_18_191), 
      .ZN(n_2_18_192));
   INV_X1 i_2_18_340 (.A(n_2_18_192), .ZN(n_2_18_193));
   OAI22_X1 i_2_18_341 (.A1(n_2_215), .A2(n_2_18_192), .B1(n_2_18_193), .B2(
      n_266), .ZN(n_2_18_194));
   INV_X1 i_2_18_342 (.A(n_2_18_194), .ZN(n_2_218));
   NOR2_X1 i_2_18_343 (.A1(n_2_18_194), .A2(n_2_199), .ZN(n_194));
   NAND2_X1 i_2_18_344 (.A1(n_2_105), .A2(n_2_106), .ZN(n_2_18_195));
   NOR2_X1 i_2_18_345 (.A1(Writing_Start_Index[3]), .A2(Writing_Start_Index[4]), 
      .ZN(n_2_18_196));
   NAND2_X1 i_2_18_346 (.A1(n_2_18_196), .A2(n_2_18_185), .ZN(n_2_18_197));
   NOR2_X1 i_2_18_347 (.A1(Writing_Start_Index[0]), .A2(Writing_Start_Index[1]), 
      .ZN(n_2_18_198));
   INV_X1 i_2_18_348 (.A(n_2_18_198), .ZN(n_2_18_199));
   NAND2_X1 i_2_18_349 (.A1(n_2_18_199), .A2(Writing_Start_Index[2]), .ZN(
      n_2_18_200));
   INV_X1 i_2_18_350 (.A(n_2_18_200), .ZN(n_2_18_201));
   OAI211_X1 i_2_18_351 (.A(n_2_18_434), .B(n_2_18_195), .C1(n_2_18_197), 
      .C2(n_2_18_201), .ZN(n_2_18_202));
   INV_X1 i_2_18_352 (.A(n_2_18_202), .ZN(n_2_18_203));
   AOI22_X1 i_2_18_353 (.A1(n_2_215), .A2(n_2_18_203), .B1(n_2_18_202), .B2(
      n_265), .ZN(n_2_18_204));
   INV_X1 i_2_18_354 (.A(n_2_18_204), .ZN(n_2_219));
   NOR2_X1 i_2_18_355 (.A1(n_2_18_204), .A2(n_2_199), .ZN(n_195));
   NAND2_X1 i_2_18_356 (.A1(n_2_18_178), .A2(n_2_106), .ZN(n_2_18_205));
   AND2_X1 i_2_18_357 (.A1(Writing_Start_Index[1]), .A2(Writing_Start_Index[2]), 
      .ZN(n_2_18_206));
   OAI211_X1 i_2_18_358 (.A(n_2_18_434), .B(n_2_18_205), .C1(n_2_18_197), 
      .C2(n_2_18_206), .ZN(n_2_18_207));
   INV_X1 i_2_18_359 (.A(n_2_18_207), .ZN(n_2_18_208));
   AOI22_X1 i_2_18_360 (.A1(n_2_215), .A2(n_2_18_208), .B1(n_2_18_207), .B2(
      n_264), .ZN(n_2_18_209));
   INV_X1 i_2_18_361 (.A(n_2_18_209), .ZN(n_2_220));
   NOR2_X1 i_2_18_362 (.A1(n_2_18_209), .A2(n_2_199), .ZN(n_196));
   INV_X1 i_2_18_363 (.A(n_2_18_187), .ZN(n_2_18_210));
   NAND2_X1 i_2_18_364 (.A1(n_2_18_210), .A2(Writing_Start_Index[2]), .ZN(
      n_2_18_211));
   INV_X1 i_2_18_365 (.A(n_2_18_211), .ZN(n_2_18_212));
   OAI21_X1 i_2_18_366 (.A(n_2_18_434), .B1(n_2_18_197), .B2(n_2_18_212), 
      .ZN(n_2_18_213));
   INV_X1 i_2_18_367 (.A(n_2_18_213), .ZN(n_2_18_214));
   AOI22_X1 i_2_18_368 (.A1(n_2_215), .A2(n_2_18_214), .B1(n_2_18_213), .B2(
      n_263), .ZN(n_2_18_215));
   INV_X1 i_2_18_369 (.A(n_2_18_215), .ZN(n_2_221));
   NOR2_X1 i_2_18_370 (.A1(n_2_18_215), .A2(n_2_199), .ZN(n_197));
   NAND2_X1 i_2_18_371 (.A1(n_2_18_428), .A2(n_2_107), .ZN(n_2_18_216));
   NOR2_X1 i_2_18_372 (.A1(n_2_108), .A2(n_2_109), .ZN(n_2_18_217));
   NAND3_X1 i_2_18_373 (.A1(n_2_18_216), .A2(n_2_18_197), .A3(n_2_18_217), 
      .ZN(n_2_18_218));
   INV_X1 i_2_18_374 (.A(n_2_18_218), .ZN(n_2_18_219));
   OAI22_X1 i_2_18_375 (.A1(n_2_215), .A2(n_2_18_218), .B1(n_2_18_219), .B2(
      n_262), .ZN(n_2_18_220));
   INV_X1 i_2_18_376 (.A(n_2_18_220), .ZN(n_2_222));
   NOR2_X1 i_2_18_377 (.A1(n_2_18_220), .A2(n_2_199), .ZN(n_198));
   OR2_X1 i_2_18_378 (.A1(n_2_105), .A2(n_2_106), .ZN(n_2_18_221));
   NAND2_X1 i_2_18_379 (.A1(n_2_18_221), .A2(n_2_107), .ZN(n_2_18_222));
   NOR2_X1 i_2_18_380 (.A1(n_2_18_199), .A2(Writing_Start_Index[2]), .ZN(
      n_2_18_223));
   INV_X1 i_2_18_381 (.A(Writing_Start_Index[3]), .ZN(n_2_18_224));
   NOR2_X1 i_2_18_382 (.A1(n_2_18_223), .A2(n_2_18_224), .ZN(n_2_18_225));
   OAI211_X1 i_2_18_383 (.A(n_2_18_217), .B(n_2_18_222), .C1(n_2_18_225), 
      .C2(n_2_18_425), .ZN(n_2_18_226));
   INV_X1 i_2_18_384 (.A(n_2_18_226), .ZN(n_2_18_227));
   AOI22_X1 i_2_18_385 (.A1(n_2_215), .A2(n_2_18_227), .B1(n_2_18_226), .B2(
      n_261), .ZN(n_2_18_228));
   INV_X1 i_2_18_386 (.A(n_2_18_228), .ZN(n_2_223));
   NOR2_X1 i_2_18_387 (.A1(n_2_18_228), .A2(n_2_199), .ZN(n_199));
   INV_X1 i_2_18_388 (.A(n_2_18_437), .ZN(n_2_18_229));
   AOI21_X1 i_2_18_389 (.A(n_2_108), .B1(n_2_18_229), .B2(n_2_107), .ZN(
      n_2_18_230));
   AOI21_X1 i_2_18_390 (.A(Writing_Start_Index[4]), .B1(n_2_18_180), .B2(
      Writing_Start_Index[3]), .ZN(n_2_18_231));
   INV_X1 i_2_18_391 (.A(n_2_18_231), .ZN(n_2_18_232));
   OAI211_X1 i_2_18_392 (.A(n_2_18_230), .B(n_2_18_444), .C1(n_2_18_232), 
      .C2(Writing_Start_Index[5]), .ZN(n_2_18_233));
   INV_X1 i_2_18_393 (.A(n_2_18_233), .ZN(n_2_18_234));
   AOI22_X1 i_2_18_394 (.A1(n_2_215), .A2(n_2_18_234), .B1(n_2_18_233), .B2(
      n_260), .ZN(n_2_18_235));
   INV_X1 i_2_18_395 (.A(n_2_18_235), .ZN(n_2_224));
   NOR2_X1 i_2_18_396 (.A1(n_2_18_235), .A2(n_2_199), .ZN(n_200));
   INV_X1 i_2_18_397 (.A(n_2_108), .ZN(n_2_18_236));
   INV_X1 i_2_18_398 (.A(n_2_107), .ZN(n_2_18_237));
   OAI21_X1 i_2_18_399 (.A(n_2_18_236), .B1(n_2_18_237), .B2(n_2_18_432), 
      .ZN(n_2_18_238));
   NOR2_X1 i_2_18_400 (.A1(n_2_18_210), .A2(Writing_Start_Index[2]), .ZN(
      n_2_18_239));
   INV_X1 i_2_18_401 (.A(n_2_18_239), .ZN(n_2_18_240));
   NAND2_X1 i_2_18_402 (.A1(n_2_18_240), .A2(Writing_Start_Index[3]), .ZN(
      n_2_18_241));
   AOI211_X1 i_2_18_403 (.A(n_2_109), .B(n_2_18_238), .C1(n_2_18_241), .C2(
      n_2_18_182), .ZN(n_2_18_242));
   INV_X1 i_2_18_404 (.A(n_2_18_242), .ZN(n_2_18_243));
   AOI22_X1 i_2_18_405 (.A1(n_2_215), .A2(n_2_18_242), .B1(n_2_18_243), .B2(
      n_259), .ZN(n_2_18_244));
   INV_X1 i_2_18_406 (.A(n_2_18_244), .ZN(n_2_225));
   NOR2_X1 i_2_18_407 (.A1(n_2_18_244), .A2(n_2_199), .ZN(n_201));
   INV_X1 i_2_18_408 (.A(n_2_18_217), .ZN(n_2_18_245));
   NOR3_X1 i_2_18_409 (.A1(n_2_18_431), .A2(n_2_18_237), .A3(n_2_18_432), 
      .ZN(n_2_18_246));
   NAND2_X1 i_2_18_410 (.A1(Writing_Start_Index[3]), .A2(Writing_Start_Index[2]), 
      .ZN(n_2_18_247));
   AOI211_X1 i_2_18_411 (.A(n_2_18_245), .B(n_2_18_246), .C1(n_2_18_182), 
      .C2(n_2_18_247), .ZN(n_2_18_248));
   OAI21_X1 i_2_18_412 (.A(n_2_18_28), .B1(n_2_18_248), .B2(n_322), .ZN(
      n_2_18_249));
   AOI21_X1 i_2_18_413 (.A(n_2_18_249), .B1(n_2_18_142), .B2(n_2_18_248), 
      .ZN(n_202));
   NOR2_X1 i_2_18_414 (.A1(n_2_18_195), .A2(n_2_18_237), .ZN(n_2_18_250));
   NAND2_X1 i_2_18_415 (.A1(n_2_18_201), .A2(Writing_Start_Index[3]), .ZN(
      n_2_18_251));
   AOI211_X1 i_2_18_416 (.A(n_2_18_245), .B(n_2_18_250), .C1(n_2_18_251), 
      .C2(n_2_18_182), .ZN(n_2_18_252));
   OAI21_X1 i_2_18_417 (.A(n_2_18_28), .B1(n_2_18_252), .B2(n_321), .ZN(
      n_2_18_253));
   AOI21_X1 i_2_18_418 (.A(n_2_18_253), .B1(n_2_18_142), .B2(n_2_18_252), 
      .ZN(n_203));
   OAI21_X1 i_2_18_419 (.A(n_2_18_236), .B1(n_2_18_205), .B2(n_2_18_237), 
      .ZN(n_2_18_254));
   NAND2_X1 i_2_18_420 (.A1(n_2_18_206), .A2(Writing_Start_Index[3]), .ZN(
      n_2_18_255));
   AOI211_X1 i_2_18_421 (.A(n_2_109), .B(n_2_18_254), .C1(n_2_18_182), .C2(
      n_2_18_255), .ZN(n_2_18_256));
   OAI21_X1 i_2_18_422 (.A(n_2_18_28), .B1(n_2_18_256), .B2(n_320), .ZN(
      n_2_18_257));
   AOI21_X1 i_2_18_423 (.A(n_2_18_257), .B1(n_2_18_142), .B2(n_2_18_256), 
      .ZN(n_204));
   NAND2_X1 i_2_18_424 (.A1(n_2_18_212), .A2(Writing_Start_Index[3]), .ZN(
      n_2_18_258));
   AOI21_X1 i_2_18_425 (.A(n_2_18_245), .B1(n_2_18_258), .B2(n_2_18_182), 
      .ZN(n_2_18_259));
   OAI21_X1 i_2_18_426 (.A(n_2_18_28), .B1(n_2_18_259), .B2(n_319), .ZN(
      n_2_18_260));
   AOI21_X1 i_2_18_427 (.A(n_2_18_260), .B1(n_2_18_142), .B2(n_2_18_259), 
      .ZN(n_205));
   NOR2_X1 i_2_18_428 (.A1(n_2_18_431), .A2(n_2_18_236), .ZN(n_2_18_261));
   OAI21_X1 i_2_18_429 (.A(n_2_18_445), .B1(n_2_18_446), .B2(n_2_106), .ZN(
      n_2_18_262));
   INV_X1 i_2_18_430 (.A(n_2_18_262), .ZN(n_2_18_263));
   NOR4_X1 i_2_18_431 (.A1(n_2_18_261), .A2(n_2_18_263), .A3(n_2_18_182), 
      .A4(n_2_109), .ZN(n_2_18_264));
   OAI21_X1 i_2_18_432 (.A(n_2_18_28), .B1(n_2_18_264), .B2(n_318), .ZN(
      n_2_18_265));
   AOI21_X1 i_2_18_433 (.A(n_2_18_265), .B1(n_2_18_142), .B2(n_2_18_264), 
      .ZN(n_206));
   NAND2_X1 i_2_18_434 (.A1(n_2_18_183), .A2(Writing_Start_Index[4]), .ZN(
      n_2_18_266));
   INV_X1 i_2_18_435 (.A(n_2_18_266), .ZN(n_2_18_267));
   AOI21_X1 i_2_18_436 (.A(n_2_18_267), .B1(n_2_18_199), .B2(
      Writing_Start_Index[4]), .ZN(n_2_18_268));
   INV_X1 i_2_18_437 (.A(n_2_18_268), .ZN(n_2_18_269));
   NOR2_X1 i_2_18_438 (.A1(n_2_18_221), .A2(n_2_18_446), .ZN(n_2_18_270));
   OAI22_X1 i_2_18_439 (.A1(n_2_18_269), .A2(Writing_Start_Index[5]), .B1(
      n_2_18_270), .B2(n_2_18_236), .ZN(n_2_18_271));
   NOR2_X1 i_2_18_440 (.A1(n_2_18_271), .A2(n_2_109), .ZN(n_2_18_272));
   OAI21_X1 i_2_18_441 (.A(n_2_18_28), .B1(n_2_18_272), .B2(n_317), .ZN(
      n_2_18_273));
   AOI21_X1 i_2_18_442 (.A(n_2_18_273), .B1(n_2_18_142), .B2(n_2_18_272), 
      .ZN(n_207));
   OAI21_X1 i_2_18_443 (.A(n_2_18_445), .B1(n_2_18_229), .B2(n_2_18_446), 
      .ZN(n_2_18_274));
   OAI211_X1 i_2_18_444 (.A(n_2_18_274), .B(n_2_18_425), .C1(n_2_18_426), 
      .C2(Writing_Start_Index[5]), .ZN(n_2_18_275));
   NOR2_X1 i_2_18_445 (.A1(n_2_18_275), .A2(n_2_109), .ZN(n_2_18_276));
   OAI21_X1 i_2_18_446 (.A(n_2_18_28), .B1(n_2_18_276), .B2(n_316), .ZN(
      n_2_18_277));
   AOI21_X1 i_2_18_447 (.A(n_2_18_277), .B1(n_2_18_142), .B2(n_2_18_276), 
      .ZN(n_208));
   NOR2_X1 i_2_18_448 (.A1(n_2_18_240), .A2(Writing_Start_Index[3]), .ZN(
      n_2_18_278));
   INV_X1 i_2_18_449 (.A(n_2_18_278), .ZN(n_2_18_279));
   AOI21_X1 i_2_18_450 (.A(Writing_Start_Index[5]), .B1(n_2_18_279), .B2(
      Writing_Start_Index[4]), .ZN(n_2_18_280));
   NOR3_X1 i_2_18_451 (.A1(n_2_18_280), .A2(n_2_109), .A3(n_2_18_263), .ZN(
      n_2_18_281));
   OAI21_X1 i_2_18_452 (.A(n_2_18_28), .B1(n_2_18_281), .B2(n_315), .ZN(
      n_2_18_282));
   AOI21_X1 i_2_18_453 (.A(n_2_18_282), .B1(n_2_18_142), .B2(n_2_18_281), 
      .ZN(n_209));
   OAI21_X1 i_2_18_454 (.A(n_2_18_445), .B1(n_2_18_191), .B2(n_2_18_446), 
      .ZN(n_2_18_283));
   OAI21_X1 i_2_18_455 (.A(n_2_18_283), .B1(Writing_Start_Index[5]), .B2(
      n_2_18_267), .ZN(n_2_18_284));
   NOR2_X1 i_2_18_456 (.A1(n_2_18_284), .A2(n_2_109), .ZN(n_2_18_285));
   OAI21_X1 i_2_18_457 (.A(n_2_18_28), .B1(n_2_18_285), .B2(n_314), .ZN(
      n_2_18_286));
   AOI21_X1 i_2_18_458 (.A(n_2_18_286), .B1(n_2_18_142), .B2(n_2_18_285), 
      .ZN(n_210));
   INV_X1 i_2_18_459 (.A(Writing_Start_Index[4]), .ZN(n_2_18_287));
   AOI21_X1 i_2_18_460 (.A(n_2_18_287), .B1(n_2_18_200), .B2(n_2_18_224), 
      .ZN(n_2_18_288));
   INV_X1 i_2_18_461 (.A(n_2_18_195), .ZN(n_2_18_289));
   NOR2_X1 i_2_18_462 (.A1(n_2_18_289), .A2(n_2_18_446), .ZN(n_2_18_290));
   OAI22_X1 i_2_18_463 (.A1(n_2_18_288), .A2(Writing_Start_Index[5]), .B1(
      n_2_18_290), .B2(n_2_18_236), .ZN(n_2_18_291));
   NOR2_X1 i_2_18_464 (.A1(n_2_18_291), .A2(n_2_109), .ZN(n_2_18_292));
   OAI21_X1 i_2_18_465 (.A(n_2_18_28), .B1(n_2_18_292), .B2(n_313), .ZN(
      n_2_18_293));
   AOI21_X1 i_2_18_466 (.A(n_2_18_293), .B1(n_2_18_142), .B2(n_2_18_292), 
      .ZN(n_211));
   NAND2_X1 i_2_18_467 (.A1(n_2_18_446), .A2(n_2_18_445), .ZN(n_2_18_294));
   NAND2_X1 i_2_18_468 (.A1(n_2_18_294), .A2(n_2_18_444), .ZN(n_2_18_295));
   INV_X1 i_2_18_469 (.A(n_2_18_205), .ZN(n_2_18_296));
   OAI21_X1 i_2_18_470 (.A(Writing_Start_Index[4]), .B1(n_2_18_206), .B2(
      Writing_Start_Index[3]), .ZN(n_2_18_297));
   AOI221_X1 i_2_18_471 (.A(n_2_18_295), .B1(n_2_18_296), .B2(n_2_18_445), 
      .C1(n_2_18_297), .C2(n_2_18_185), .ZN(n_2_18_298));
   OAI21_X1 i_2_18_472 (.A(n_2_18_28), .B1(n_2_18_298), .B2(n_312), .ZN(
      n_2_18_299));
   AOI21_X1 i_2_18_473 (.A(n_2_18_299), .B1(n_2_18_142), .B2(n_2_18_298), 
      .ZN(n_212));
   OAI21_X1 i_2_18_474 (.A(Writing_Start_Index[4]), .B1(n_2_18_212), .B2(
      Writing_Start_Index[3]), .ZN(n_2_18_300));
   AOI21_X1 i_2_18_475 (.A(n_2_18_295), .B1(n_2_18_300), .B2(n_2_18_185), 
      .ZN(n_2_18_301));
   OAI21_X1 i_2_18_476 (.A(n_2_18_28), .B1(n_2_18_301), .B2(n_311), .ZN(
      n_2_18_302));
   AOI21_X1 i_2_18_477 (.A(n_2_18_302), .B1(n_2_18_142), .B2(n_2_18_301), 
      .ZN(n_213));
   NOR2_X1 i_2_18_478 (.A1(n_2_18_216), .A2(n_2_18_236), .ZN(n_2_18_303));
   NOR2_X1 i_2_18_479 (.A1(n_2_18_224), .A2(n_2_18_287), .ZN(n_2_18_304));
   OAI21_X1 i_2_18_480 (.A(n_2_18_444), .B1(n_2_18_304), .B2(
      Writing_Start_Index[5]), .ZN(n_2_18_305));
   NOR2_X1 i_2_18_481 (.A1(n_2_18_303), .A2(n_2_18_305), .ZN(n_2_18_306));
   OAI21_X1 i_2_18_482 (.A(n_2_18_28), .B1(n_2_18_306), .B2(n_310), .ZN(
      n_2_18_307));
   AOI21_X1 i_2_18_483 (.A(n_2_18_307), .B1(n_2_18_142), .B2(n_2_18_306), 
      .ZN(n_214));
   NOR2_X1 i_2_18_484 (.A1(Writing_Start_Index[2]), .A2(Writing_Start_Index[5]), 
      .ZN(n_2_18_308));
   INV_X1 i_2_18_485 (.A(n_2_18_222), .ZN(n_2_18_309));
   AOI221_X1 i_2_18_486 (.A(n_2_18_305), .B1(n_2_18_198), .B2(n_2_18_308), 
      .C1(n_2_18_445), .C2(n_2_18_309), .ZN(n_2_18_310));
   OAI21_X1 i_2_18_487 (.A(n_2_18_28), .B1(n_2_18_310), .B2(n_309), .ZN(
      n_2_18_311));
   AOI21_X1 i_2_18_488 (.A(n_2_18_311), .B1(n_2_18_142), .B2(n_2_18_310), 
      .ZN(n_215));
   NOR2_X1 i_2_18_489 (.A1(n_2_18_437), .A2(n_2_18_294), .ZN(n_2_18_312));
   AOI21_X1 i_2_18_490 (.A(Writing_Start_Index[5]), .B1(n_2_18_180), .B2(
      n_2_18_304), .ZN(n_2_18_313));
   NOR3_X1 i_2_18_491 (.A1(n_2_18_312), .A2(n_2_18_313), .A3(n_2_109), .ZN(
      n_2_18_314));
   OAI21_X1 i_2_18_492 (.A(n_2_18_28), .B1(n_2_18_314), .B2(n_308), .ZN(
      n_2_18_315));
   AOI21_X1 i_2_18_493 (.A(n_2_18_315), .B1(n_2_18_142), .B2(n_2_18_314), 
      .ZN(n_216));
   NOR2_X1 i_2_18_494 (.A1(n_2_18_294), .A2(n_2_18_432), .ZN(n_2_18_316));
   AOI211_X1 i_2_18_495 (.A(n_2_18_316), .B(n_2_18_305), .C1(n_2_18_187), 
      .C2(n_2_18_308), .ZN(n_2_18_317));
   OAI21_X1 i_2_18_496 (.A(n_2_18_28), .B1(n_2_18_317), .B2(n_307), .ZN(
      n_2_18_318));
   AOI21_X1 i_2_18_497 (.A(n_2_18_318), .B1(n_2_18_142), .B2(n_2_18_317), 
      .ZN(n_217));
   AOI211_X1 i_2_18_498 (.A(n_2_18_308), .B(n_2_18_305), .C1(n_2_18_246), 
      .C2(n_2_18_445), .ZN(n_2_18_319));
   OAI21_X1 i_2_18_499 (.A(n_2_18_28), .B1(n_2_18_319), .B2(n_306), .ZN(
      n_2_18_320));
   AOI21_X1 i_2_18_500 (.A(n_2_18_320), .B1(n_2_18_142), .B2(n_2_18_319), 
      .ZN(n_218));
   AOI221_X1 i_2_18_501 (.A(n_2_18_305), .B1(n_2_18_185), .B2(n_2_18_200), 
      .C1(n_2_18_445), .C2(n_2_18_250), .ZN(n_2_18_321));
   OAI21_X1 i_2_18_502 (.A(n_2_18_28), .B1(n_2_18_321), .B2(n_305), .ZN(
      n_2_18_322));
   AOI21_X1 i_2_18_503 (.A(n_2_18_322), .B1(n_2_18_142), .B2(n_2_18_321), 
      .ZN(n_219));
   NOR2_X1 i_2_18_504 (.A1(n_2_18_255), .A2(n_2_18_287), .ZN(n_2_18_323));
   OAI22_X1 i_2_18_505 (.A1(n_2_18_323), .A2(Writing_Start_Index[5]), .B1(
      n_2_18_205), .B2(n_2_18_294), .ZN(n_2_18_324));
   NOR2_X1 i_2_18_506 (.A1(n_2_18_324), .A2(n_2_109), .ZN(n_2_18_325));
   OAI21_X1 i_2_18_507 (.A(n_2_18_28), .B1(n_2_18_325), .B2(n_304), .ZN(
      n_2_18_326));
   AOI21_X1 i_2_18_508 (.A(n_2_18_326), .B1(n_2_18_142), .B2(n_2_18_325), 
      .ZN(n_220));
   AOI21_X1 i_2_18_509 (.A(n_2_18_305), .B1(n_2_18_185), .B2(n_2_18_211), 
      .ZN(n_2_18_327));
   OAI21_X1 i_2_18_510 (.A(n_2_18_28), .B1(n_2_18_327), .B2(n_303), .ZN(
      n_2_18_328));
   AOI21_X1 i_2_18_511 (.A(n_2_18_328), .B1(n_2_18_142), .B2(n_2_18_327), 
      .ZN(n_221));
   OAI21_X1 i_2_18_512 (.A(Writing_Start_Index[5]), .B1(n_2_18_440), .B2(
      n_2_18_444), .ZN(n_2_18_329));
   AOI21_X1 i_2_18_513 (.A(n_2_18_329), .B1(n_2_109), .B2(n_2_18_428), .ZN(
      n_2_18_330));
   OAI21_X1 i_2_18_514 (.A(n_2_18_28), .B1(n_2_18_330), .B2(n_302), .ZN(
      n_2_18_331));
   AOI21_X1 i_2_18_515 (.A(n_2_18_331), .B1(n_2_18_142), .B2(n_2_18_330), 
      .ZN(n_222));
   AOI221_X1 i_2_18_516 (.A(n_2_18_329), .B1(n_2_109), .B2(n_2_18_221), .C1(
      n_2_18_184), .C2(n_2_18_198), .ZN(n_2_18_332));
   OAI21_X1 i_2_18_517 (.A(n_2_18_28), .B1(n_2_18_332), .B2(n_301), .ZN(
      n_2_18_333));
   AOI21_X1 i_2_18_518 (.A(n_2_18_333), .B1(n_2_18_142), .B2(n_2_18_332), 
      .ZN(n_223));
   AOI221_X1 i_2_18_519 (.A(n_2_18_329), .B1(n_2_109), .B2(n_2_18_229), .C1(
      n_2_18_181), .C2(n_2_18_287), .ZN(n_2_18_334));
   OAI21_X1 i_2_18_520 (.A(n_2_18_28), .B1(n_2_18_334), .B2(n_300), .ZN(
      n_2_18_335));
   AOI21_X1 i_2_18_521 (.A(n_2_18_335), .B1(n_2_18_142), .B2(n_2_18_334), 
      .ZN(n_224));
   AOI221_X1 i_2_18_522 (.A(n_2_18_329), .B1(n_2_106), .B2(n_2_109), .C1(
      n_2_18_184), .C2(n_2_18_187), .ZN(n_2_18_336));
   OAI21_X1 i_2_18_523 (.A(n_2_18_28), .B1(n_2_18_336), .B2(n_299), .ZN(
      n_2_18_337));
   AOI21_X1 i_2_18_524 (.A(n_2_18_337), .B1(n_2_18_142), .B2(n_2_18_336), 
      .ZN(n_225));
   AOI211_X1 i_2_18_525 (.A(n_2_18_184), .B(n_2_18_329), .C1(n_2_109), .C2(
      n_2_18_191), .ZN(n_2_18_338));
   OAI21_X1 i_2_18_526 (.A(n_2_18_28), .B1(n_2_18_338), .B2(n_298), .ZN(
      n_2_18_339));
   AOI21_X1 i_2_18_527 (.A(n_2_18_339), .B1(n_2_18_142), .B2(n_2_18_338), 
      .ZN(n_226));
   AOI221_X1 i_2_18_528 (.A(n_2_18_329), .B1(n_2_18_289), .B2(n_2_109), .C1(
      n_2_18_196), .C2(n_2_18_200), .ZN(n_2_18_340));
   OAI21_X1 i_2_18_529 (.A(n_2_18_28), .B1(n_2_18_340), .B2(n_297), .ZN(
      n_2_18_341));
   AOI21_X1 i_2_18_530 (.A(n_2_18_341), .B1(n_2_18_142), .B2(n_2_18_340), 
      .ZN(n_227));
   INV_X1 i_2_18_531 (.A(n_2_18_329), .ZN(n_2_18_342));
   INV_X1 i_2_18_532 (.A(n_2_18_196), .ZN(n_2_18_343));
   OAI21_X1 i_2_18_533 (.A(n_2_18_342), .B1(n_2_18_343), .B2(n_2_18_206), 
      .ZN(n_2_18_344));
   AOI21_X1 i_2_18_534 (.A(n_2_18_344), .B1(n_2_109), .B2(n_2_18_296), .ZN(
      n_2_18_345));
   OAI21_X1 i_2_18_535 (.A(n_2_18_28), .B1(n_2_18_345), .B2(n_296), .ZN(
      n_2_18_346));
   AOI21_X1 i_2_18_536 (.A(n_2_18_346), .B1(n_2_18_142), .B2(n_2_18_345), 
      .ZN(n_228));
   AOI21_X1 i_2_18_537 (.A(n_2_18_329), .B1(n_2_18_196), .B2(n_2_18_211), 
      .ZN(n_2_18_347));
   OAI21_X1 i_2_18_538 (.A(n_2_18_28), .B1(n_2_18_347), .B2(n_295), .ZN(
      n_2_18_348));
   AOI21_X1 i_2_18_539 (.A(n_2_18_348), .B1(n_2_18_142), .B2(n_2_18_347), 
      .ZN(n_229));
   NAND2_X1 i_2_18_540 (.A1(n_2_18_445), .A2(n_2_109), .ZN(n_2_18_349));
   NAND2_X1 i_2_18_541 (.A1(n_2_18_349), .A2(Writing_Start_Index[5]), .ZN(
      n_2_18_350));
   INV_X1 i_2_18_542 (.A(n_2_18_350), .ZN(n_2_18_351));
   NAND2_X1 i_2_18_543 (.A1(n_2_18_351), .A2(n_2_18_343), .ZN(n_2_18_352));
   INV_X1 i_2_18_544 (.A(n_2_18_216), .ZN(n_2_18_353));
   AOI21_X1 i_2_18_545 (.A(n_2_18_352), .B1(n_2_109), .B2(n_2_18_353), .ZN(
      n_2_18_354));
   OAI21_X1 i_2_18_546 (.A(n_2_18_28), .B1(n_2_18_354), .B2(n_294), .ZN(
      n_2_18_355));
   AOI21_X1 i_2_18_547 (.A(n_2_18_355), .B1(n_2_18_142), .B2(n_2_18_354), 
      .ZN(n_230));
   OAI21_X1 i_2_18_548 (.A(n_2_18_351), .B1(n_2_18_225), .B2(
      Writing_Start_Index[4]), .ZN(n_2_18_356));
   AOI21_X1 i_2_18_549 (.A(n_2_18_356), .B1(n_2_109), .B2(n_2_18_309), .ZN(
      n_2_18_357));
   OAI21_X1 i_2_18_550 (.A(n_2_18_28), .B1(n_2_18_357), .B2(n_293), .ZN(
      n_2_18_358));
   AOI21_X1 i_2_18_551 (.A(n_2_18_358), .B1(n_2_18_142), .B2(n_2_18_357), 
      .ZN(n_231));
   INV_X1 i_2_18_552 (.A(n_2_18_230), .ZN(n_2_18_359));
   AOI211_X1 i_2_18_553 (.A(n_2_18_185), .B(n_2_18_231), .C1(n_2_18_359), 
      .C2(n_2_109), .ZN(n_2_18_360));
   OAI21_X1 i_2_18_554 (.A(n_2_18_28), .B1(n_2_18_360), .B2(n_292), .ZN(
      n_2_18_361));
   AOI21_X1 i_2_18_555 (.A(n_2_18_361), .B1(n_2_18_142), .B2(n_2_18_360), 
      .ZN(n_232));
   AOI221_X1 i_2_18_556 (.A(n_2_18_185), .B1(n_2_18_238), .B2(n_2_109), .C1(
      n_2_18_241), .C2(n_2_18_287), .ZN(n_2_18_362));
   OAI21_X1 i_2_18_557 (.A(n_2_18_28), .B1(n_2_18_362), .B2(n_291), .ZN(
      n_2_18_363));
   AOI21_X1 i_2_18_558 (.A(n_2_18_363), .B1(n_2_18_142), .B2(n_2_18_362), 
      .ZN(n_233));
   INV_X1 i_2_18_559 (.A(n_2_18_349), .ZN(n_2_18_364));
   INV_X1 i_2_18_560 (.A(n_2_18_247), .ZN(n_2_18_365));
   OAI21_X1 i_2_18_561 (.A(Writing_Start_Index[5]), .B1(n_2_18_365), .B2(
      Writing_Start_Index[4]), .ZN(n_2_18_366));
   AOI211_X1 i_2_18_562 (.A(n_2_18_364), .B(n_2_18_366), .C1(n_2_18_246), 
      .C2(n_2_109), .ZN(n_2_18_367));
   OAI21_X1 i_2_18_563 (.A(n_2_18_28), .B1(n_2_18_367), .B2(n_290), .ZN(
      n_2_18_368));
   AOI21_X1 i_2_18_564 (.A(n_2_18_368), .B1(n_2_18_142), .B2(n_2_18_367), 
      .ZN(n_234));
   AOI221_X1 i_2_18_565 (.A(n_2_18_350), .B1(n_2_18_250), .B2(n_2_109), .C1(
      n_2_18_251), .C2(n_2_18_287), .ZN(n_2_18_369));
   OAI21_X1 i_2_18_566 (.A(n_2_18_28), .B1(n_2_18_369), .B2(n_289), .ZN(
      n_2_18_370));
   AOI21_X1 i_2_18_567 (.A(n_2_18_370), .B1(n_2_18_142), .B2(n_2_18_369), 
      .ZN(n_235));
   AOI221_X1 i_2_18_568 (.A(n_2_18_185), .B1(n_2_18_255), .B2(n_2_18_287), 
      .C1(n_2_18_254), .C2(n_2_109), .ZN(n_2_18_371));
   OAI21_X1 i_2_18_569 (.A(n_2_18_28), .B1(n_2_18_371), .B2(n_288), .ZN(
      n_2_18_372));
   AOI21_X1 i_2_18_570 (.A(n_2_18_372), .B1(n_2_18_142), .B2(n_2_18_371), 
      .ZN(n_236));
   AOI21_X1 i_2_18_571 (.A(n_2_18_350), .B1(n_2_18_258), .B2(n_2_18_287), 
      .ZN(n_2_18_373));
   OAI21_X1 i_2_18_572 (.A(n_2_18_28), .B1(n_2_18_373), .B2(n_287), .ZN(
      n_2_18_374));
   AOI21_X1 i_2_18_573 (.A(n_2_18_374), .B1(n_2_18_142), .B2(n_2_18_373), 
      .ZN(n_237));
   NAND2_X1 i_2_18_574 (.A1(Writing_Start_Index[4]), .A2(Writing_Start_Index[5]), 
      .ZN(n_2_18_375));
   NOR2_X1 i_2_18_575 (.A1(n_2_18_262), .A2(n_2_18_444), .ZN(n_2_18_376));
   AOI211_X1 i_2_18_576 (.A(n_2_18_375), .B(n_2_18_376), .C1(n_2_109), .C2(
      n_2_18_261), .ZN(n_2_18_377));
   OAI21_X1 i_2_18_577 (.A(n_2_18_28), .B1(n_2_18_377), .B2(n_286), .ZN(
      n_2_18_378));
   AOI21_X1 i_2_18_578 (.A(n_2_18_378), .B1(n_2_18_142), .B2(n_2_18_377), 
      .ZN(n_238));
   INV_X1 i_2_18_579 (.A(n_2_18_270), .ZN(n_2_18_379));
   AOI211_X1 i_2_18_580 (.A(n_2_18_185), .B(n_2_18_268), .C1(n_2_18_379), 
      .C2(n_2_18_364), .ZN(n_2_18_380));
   OAI21_X1 i_2_18_581 (.A(n_2_18_28), .B1(n_2_18_380), .B2(n_285), .ZN(
      n_2_18_381));
   AOI21_X1 i_2_18_582 (.A(n_2_18_381), .B1(n_2_18_142), .B2(n_2_18_380), 
      .ZN(n_239));
   INV_X1 i_2_18_583 (.A(n_2_18_274), .ZN(n_2_18_382));
   AOI211_X1 i_2_18_584 (.A(n_2_18_181), .B(n_2_18_375), .C1(n_2_18_382), 
      .C2(n_2_109), .ZN(n_2_18_383));
   OAI21_X1 i_2_18_585 (.A(n_2_18_28), .B1(n_2_18_383), .B2(n_284), .ZN(
      n_2_18_384));
   AOI21_X1 i_2_18_586 (.A(n_2_18_384), .B1(n_2_18_142), .B2(n_2_18_383), 
      .ZN(n_240));
   NOR3_X1 i_2_18_587 (.A1(n_2_18_376), .A2(n_2_18_278), .A3(n_2_18_375), 
      .ZN(n_2_18_385));
   OAI21_X1 i_2_18_588 (.A(n_2_18_28), .B1(n_2_18_385), .B2(n_283), .ZN(
      n_2_18_386));
   AOI21_X1 i_2_18_589 (.A(n_2_18_386), .B1(n_2_18_142), .B2(n_2_18_385), 
      .ZN(n_241));
   INV_X1 i_2_18_590 (.A(n_2_18_283), .ZN(n_2_18_387));
   AOI211_X1 i_2_18_591 (.A(n_2_18_185), .B(n_2_18_266), .C1(n_2_18_387), 
      .C2(n_2_109), .ZN(n_2_18_388));
   OAI21_X1 i_2_18_592 (.A(n_2_18_28), .B1(n_2_18_388), .B2(n_282), .ZN(
      n_2_18_389));
   AOI21_X1 i_2_18_593 (.A(n_2_18_389), .B1(n_2_18_142), .B2(n_2_18_388), 
      .ZN(n_242));
   OAI21_X1 i_2_18_594 (.A(n_2_18_288), .B1(n_2_18_290), .B2(n_2_18_349), 
      .ZN(n_2_18_390));
   NOR2_X1 i_2_18_595 (.A1(n_2_18_390), .A2(n_2_18_185), .ZN(n_2_18_391));
   OAI21_X1 i_2_18_596 (.A(n_2_18_28), .B1(n_2_18_391), .B2(n_281), .ZN(
      n_2_18_392));
   AOI21_X1 i_2_18_597 (.A(n_2_18_392), .B1(n_2_18_142), .B2(n_2_18_391), 
      .ZN(n_243));
   NOR2_X1 i_2_18_598 (.A1(n_2_18_205), .A2(n_2_18_349), .ZN(n_2_18_393));
   NOR2_X1 i_2_18_599 (.A1(n_2_18_294), .A2(n_2_18_444), .ZN(n_2_18_394));
   NOR4_X1 i_2_18_600 (.A1(n_2_18_297), .A2(n_2_18_393), .A3(n_2_18_185), 
      .A4(n_2_18_394), .ZN(n_2_18_395));
   OAI21_X1 i_2_18_601 (.A(n_2_18_28), .B1(n_2_18_395), .B2(n_280), .ZN(
      n_2_18_396));
   AOI21_X1 i_2_18_602 (.A(n_2_18_396), .B1(n_2_18_142), .B2(n_2_18_395), 
      .ZN(n_244));
   NOR3_X1 i_2_18_603 (.A1(n_2_18_300), .A2(n_2_18_185), .A3(n_2_18_394), 
      .ZN(n_2_18_397));
   OAI21_X1 i_2_18_604 (.A(n_2_18_28), .B1(n_2_18_397), .B2(n_279), .ZN(
      n_2_18_398));
   AOI21_X1 i_2_18_605 (.A(n_2_18_398), .B1(n_2_18_142), .B2(n_2_18_397), 
      .ZN(n_245));
   NAND2_X1 i_2_18_606 (.A1(n_2_18_304), .A2(Writing_Start_Index[5]), .ZN(
      n_2_18_399));
   AOI21_X1 i_2_18_607 (.A(n_2_18_399), .B1(n_2_18_303), .B2(n_2_109), .ZN(
      n_2_18_400));
   OAI21_X1 i_2_18_608 (.A(n_2_18_28), .B1(n_2_18_400), .B2(n_278), .ZN(
      n_2_18_401));
   AOI21_X1 i_2_18_609 (.A(n_2_18_401), .B1(n_2_18_142), .B2(n_2_18_400), 
      .ZN(n_246));
   AOI211_X1 i_2_18_610 (.A(n_2_18_223), .B(n_2_18_399), .C1(n_2_18_221), 
      .C2(n_2_18_394), .ZN(n_2_18_402));
   OAI21_X1 i_2_18_611 (.A(n_2_18_28), .B1(n_2_18_402), .B2(n_277), .ZN(
      n_2_18_403));
   AOI21_X1 i_2_18_612 (.A(n_2_18_403), .B1(n_2_18_142), .B2(n_2_18_402), 
      .ZN(n_247));
   AOI211_X1 i_2_18_613 (.A(n_2_18_179), .B(n_2_18_399), .C1(n_2_18_312), 
      .C2(n_2_109), .ZN(n_2_18_404));
   OAI21_X1 i_2_18_614 (.A(n_2_18_28), .B1(n_2_18_404), .B2(n_276), .ZN(
      n_2_18_405));
   AOI21_X1 i_2_18_615 (.A(n_2_18_405), .B1(n_2_18_142), .B2(n_2_18_404), 
      .ZN(n_248));
   AOI211_X1 i_2_18_616 (.A(n_2_18_239), .B(n_2_18_399), .C1(n_2_109), .C2(
      n_2_18_316), .ZN(n_2_18_406));
   OAI21_X1 i_2_18_617 (.A(n_2_18_28), .B1(n_2_18_406), .B2(n_275), .ZN(
      n_2_18_407));
   AOI21_X1 i_2_18_618 (.A(n_2_18_407), .B1(n_2_18_142), .B2(n_2_18_406), 
      .ZN(n_249));
   AOI211_X1 i_2_18_619 (.A(n_2_18_247), .B(n_2_18_375), .C1(n_2_18_246), 
      .C2(n_2_18_364), .ZN(n_2_18_408));
   OAI21_X1 i_2_18_620 (.A(n_2_18_28), .B1(n_2_18_408), .B2(n_274), .ZN(
      n_2_18_409));
   AOI21_X1 i_2_18_621 (.A(n_2_18_409), .B1(n_2_18_142), .B2(n_2_18_408), 
      .ZN(n_250));
   AOI211_X1 i_2_18_622 (.A(n_2_18_200), .B(n_2_18_399), .C1(n_2_18_250), 
      .C2(n_2_18_364), .ZN(n_2_18_410));
   OAI21_X1 i_2_18_623 (.A(n_2_18_28), .B1(n_2_18_410), .B2(n_273), .ZN(
      n_2_18_411));
   AOI21_X1 i_2_18_624 (.A(n_2_18_411), .B1(n_2_18_142), .B2(n_2_18_410), 
      .ZN(n_251));
   AOI211_X1 i_2_18_625 (.A(n_2_18_375), .B(n_2_18_255), .C1(n_2_18_296), 
      .C2(n_2_18_394), .ZN(n_2_18_412));
   OAI21_X1 i_2_18_626 (.A(n_2_18_28), .B1(n_2_18_412), .B2(n_272), .ZN(
      n_2_18_413));
   AOI21_X1 i_2_18_627 (.A(n_2_18_413), .B1(n_2_18_142), .B2(n_2_18_412), 
      .ZN(n_252));
   NOR2_X1 i_2_18_628 (.A1(n_2_18_211), .A2(n_2_18_399), .ZN(n_2_18_414));
   OAI21_X1 i_2_18_629 (.A(n_2_18_28), .B1(n_2_18_414), .B2(n_271), .ZN(
      n_2_18_415));
   AOI21_X1 i_2_18_630 (.A(n_2_18_415), .B1(n_2_18_142), .B2(n_2_18_414), 
      .ZN(n_253));
   INV_X1 i_2_18_631 (.A(Done_Element_Delayed), .ZN(n_2_200));
   AND2_X1 i_2_18_632 (.A1(n_2_200), .A2(n_2_0), .ZN(n_2_201));
   AND2_X1 i_2_18_633 (.A1(n_2_200), .A2(n_2_1), .ZN(n_2_202));
   AND2_X1 i_2_18_634 (.A1(n_2_200), .A2(n_2_2), .ZN(n_2_203));
   AND2_X1 i_2_18_635 (.A1(n_2_200), .A2(n_2_3), .ZN(n_2_204));
   AND2_X1 i_2_18_636 (.A1(n_2_200), .A2(n_2_4), .ZN(n_2_205));
   AND2_X1 i_2_18_637 (.A1(n_2_200), .A2(n_2_5), .ZN(n_2_206));
   NOR2_X1 i_2_18_638 (.A1(n_2_18_138), .A2(N_Indication_Bit), .ZN(n_2_207));
   XNOR2_X1 i_2_18_639 (.A(n_2_76), .B(n_2_18_3), .ZN(n_2_213));
   NOR4_X1 i_2_18_640 (.A1(Data_Size[17]), .A2(Data_Size[16]), .A3(Data_Size[18]), 
      .A4(Data_Size[19]), .ZN(n_2_18_416));
   NOR4_X1 i_2_18_641 (.A1(Data_Size[21]), .A2(Data_Size[20]), .A3(Data_Size[22]), 
      .A4(Data_Size[23]), .ZN(n_2_18_417));
   NOR4_X1 i_2_18_642 (.A1(Data_Size[25]), .A2(Data_Size[24]), .A3(Data_Size[26]), 
      .A4(Data_Size[27]), .ZN(n_2_18_418));
   NOR4_X1 i_2_18_643 (.A1(Data_Size[29]), .A2(Data_Size[28]), .A3(Data_Size[30]), 
      .A4(Data_Size[31]), .ZN(n_2_18_419));
   NAND4_X1 i_2_18_644 (.A1(n_2_18_416), .A2(n_2_18_417), .A3(n_2_18_418), 
      .A4(n_2_18_419), .ZN(n_2_18_420));
   NOR4_X1 i_2_18_645 (.A1(n_2_18_420), .A2(Data_Size[13]), .A3(Data_Size[14]), 
      .A4(Data_Size[15]), .ZN(n_2_18_421));
   NOR3_X1 i_2_18_646 (.A1(Data_Size[7]), .A2(Data_Size[8]), .A3(Data_Size[6]), 
      .ZN(n_2_18_422));
   NOR4_X1 i_2_18_647 (.A1(Data_Size[10]), .A2(Data_Size[9]), .A3(Data_Size[11]), 
      .A4(Data_Size[12]), .ZN(n_2_18_423));
   NAND3_X1 i_2_18_648 (.A1(n_2_18_421), .A2(n_2_18_422), .A3(n_2_18_423), 
      .ZN(n_2_214));
   INV_X1 i_2_18_649 (.A(RAM_Address[0]), .ZN(n_2_171));
   INV_X1 i_2_18_650 (.A(Relative_Address[1]), .ZN(n_2_184));
   INV_X1 i_2_18_651 (.A(Data_Size[6]), .ZN(n_2_170));
   INV_X1 i_2_18_652 (.A(n_2_216), .ZN(n_2_18_424));
   INV_X1 i_2_18_653 (.A(n_2_18_182), .ZN(n_2_18_425));
   INV_X1 i_2_18_654 (.A(n_2_18_181), .ZN(n_2_18_426));
   INV_X1 i_2_18_655 (.A(n_2_208), .ZN(n_2_18_427));
   NAND2_X1 i_2_18_656 (.A1(n_2_18_431), .A2(n_2_18_432), .ZN(n_2_18_428));
   OAI21_X1 i_2_18_657 (.A(n_2_18_429), .B1(n_2_18_430), .B2(n_2_18_142), 
      .ZN(n_2_208));
   NAND2_X1 i_2_18_658 (.A1(n_2_18_430), .A2(n_270), .ZN(n_2_18_429));
   NAND4_X1 i_2_18_659 (.A1(n_2_18_440), .A2(n_2_18_444), .A3(n_2_18_432), 
      .A4(n_2_18_431), .ZN(n_2_18_430));
   NOR2_X1 i_2_18_660 (.A1(n_2_105), .A2(n_2_104), .ZN(n_2_18_431));
   INV_X1 i_2_18_661 (.A(n_2_106), .ZN(n_2_18_432));
   NAND2_X1 i_2_18_662 (.A1(n_2_18_435), .A2(n_2_18_433), .ZN(n_2_216));
   NAND4_X1 i_2_18_663 (.A1(n_2_18_434), .A2(n_2_215), .A3(n_2_18_438), .A4(
      n_2_18_437), .ZN(n_2_18_433));
   INV_X1 i_2_18_664 (.A(n_2_18_439), .ZN(n_2_18_434));
   INV_X1 i_2_18_665 (.A(n_2_18_142), .ZN(n_2_215));
   OAI21_X1 i_2_18_666 (.A(n_268), .B1(n_2_18_436), .B2(n_2_18_439), .ZN(
      n_2_18_435));
   NAND2_X1 i_2_18_667 (.A1(n_2_18_437), .A2(n_2_18_438), .ZN(n_2_18_436));
   NOR2_X1 i_2_18_668 (.A1(n_2_18_178), .A2(n_2_106), .ZN(n_2_18_437));
   NAND2_X1 i_2_18_669 (.A1(n_2_18_181), .A2(n_2_18_182), .ZN(n_2_18_438));
   NAND2_X1 i_2_18_670 (.A1(n_2_18_440), .A2(n_2_18_444), .ZN(n_2_18_439));
   INV_X1 i_2_18_671 (.A(n_2_18_441), .ZN(n_2_18_440));
   NAND2_X1 i_2_18_672 (.A1(n_2_18_443), .A2(n_2_18_442), .ZN(n_2_18_441));
   INV_X1 i_2_18_673 (.A(n_2_107), .ZN(n_2_18_442));
   INV_X1 i_2_18_674 (.A(n_2_108), .ZN(n_2_18_443));
   INV_X1 i_2_18_675 (.A(n_2_109), .ZN(n_2_18_444));
   BUF_X1 rt_shieldBuf__2__2__2 (.A(n_2_108), .Z(n_2_18_445));
   BUF_X1 rt_shieldBuf__2__2__3 (.A(n_2_107), .Z(n_2_18_446));
   BUF_X1 rt_shieldBuf__2 (.A(n_256), .Z(n_2_226));
   BUF_X1 rt_shieldBuf__2__2__0 (.A(n_255), .Z(n_2_227));
   BUF_X1 rt_shieldBuf__2__2__1 (.A(n_254), .Z(n_2_228));
   AOI21_X1 i_2_19_0 (.A(n_2_6), .B1(n_2_70), .B2(n_2_19_5), .ZN(n_2_19_0));
   INV_X1 i_2_19_1 (.A(n_2_19_0), .ZN(n_254));
   AOI21_X1 i_2_19_2 (.A(n_2_7), .B1(n_2_70), .B2(n_2_19_5), .ZN(n_2_19_1));
   INV_X1 i_2_19_3 (.A(n_2_19_1), .ZN(n_255));
   AOI21_X1 i_2_19_4 (.A(n_2_8), .B1(n_2_70), .B2(n_2_19_5), .ZN(n_2_19_2));
   INV_X1 i_2_19_5 (.A(n_2_19_2), .ZN(n_256));
   AOI21_X1 i_2_19_6 (.A(n_2_9), .B1(n_2_19_8), .B2(n_2_19_5), .ZN(n_2_19_3));
   INV_X1 i_2_19_7 (.A(n_2_19_3), .ZN(n_257));
   AOI21_X1 i_2_19_8 (.A(n_2_10), .B1(n_2_19_8), .B2(n_2_19_5), .ZN(n_2_19_4));
   INV_X1 i_2_19_9 (.A(n_2_19_4), .ZN(n_258));
   INV_X1 i_2_19_10 (.A(Done_Element_Delayed), .ZN(n_2_19_5));
   NAND2_X1 i_2_19_11 (.A1(n_2_19_8), .A2(n_2_19_5), .ZN(n_2_19_6));
   NAND2_X1 i_2_19_12 (.A1(n_2_11), .A2(n_2_19_6), .ZN(n_2_19_7));
   INV_X1 i_2_19_13 (.A(n_2_19_7), .ZN(n_2_229));
   BUF_X1 rt_shieldBuf__2__2__4 (.A(n_2_70), .Z(n_2_19_8));
   DFF_X1 \RAM_Data_reg[63]  (.D(n_253), .CK(n_3_2), .Q(RAM_Data[63]), .QN());
   DFF_X1 \RAM_Data_reg[62]  (.D(n_252), .CK(n_3_2), .Q(RAM_Data[62]), .QN());
   DFF_X1 \RAM_Data_reg[61]  (.D(n_251), .CK(n_3_2), .Q(RAM_Data[61]), .QN());
   DFF_X1 \RAM_Data_reg[60]  (.D(n_250), .CK(n_3_2), .Q(RAM_Data[60]), .QN());
   DFF_X1 \RAM_Data_reg[59]  (.D(n_249), .CK(n_3_2), .Q(RAM_Data[59]), .QN());
   DFF_X1 \RAM_Data_reg[58]  (.D(n_248), .CK(n_3_2), .Q(RAM_Data[58]), .QN());
   DFF_X1 \RAM_Data_reg[57]  (.D(n_247), .CK(n_3_2), .Q(RAM_Data[57]), .QN());
   DFF_X1 \RAM_Data_reg[56]  (.D(n_246), .CK(n_3_2), .Q(RAM_Data[56]), .QN());
   DFF_X1 \RAM_Data_reg[55]  (.D(n_245), .CK(n_3_2), .Q(RAM_Data[55]), .QN());
   DFF_X1 \RAM_Data_reg[54]  (.D(n_244), .CK(n_3_2), .Q(RAM_Data[54]), .QN());
   DFF_X1 \RAM_Data_reg[53]  (.D(n_243), .CK(n_3_2), .Q(RAM_Data[53]), .QN());
   DFF_X1 \RAM_Data_reg[52]  (.D(n_242), .CK(n_3_2), .Q(RAM_Data[52]), .QN());
   DFF_X1 \RAM_Data_reg[51]  (.D(n_241), .CK(n_3_2), .Q(RAM_Data[51]), .QN());
   DFF_X1 \RAM_Data_reg[50]  (.D(n_240), .CK(n_3_2), .Q(RAM_Data[50]), .QN());
   DFF_X1 \RAM_Data_reg[49]  (.D(n_239), .CK(n_3_2), .Q(RAM_Data[49]), .QN());
   DFF_X1 \RAM_Data_reg[48]  (.D(n_238), .CK(n_3_2), .Q(RAM_Data[48]), .QN());
   DFF_X1 \RAM_Data_reg[47]  (.D(n_237), .CK(n_3_2), .Q(RAM_Data[47]), .QN());
   DFF_X1 \RAM_Data_reg[46]  (.D(n_236), .CK(n_3_2), .Q(RAM_Data[46]), .QN());
   DFF_X1 \RAM_Data_reg[45]  (.D(n_235), .CK(n_3_2), .Q(RAM_Data[45]), .QN());
   DFF_X1 \RAM_Data_reg[44]  (.D(n_234), .CK(n_3_2), .Q(RAM_Data[44]), .QN());
   DFF_X1 \RAM_Data_reg[43]  (.D(n_233), .CK(n_3_2), .Q(RAM_Data[43]), .QN());
   DFF_X1 \RAM_Data_reg[42]  (.D(n_232), .CK(n_3_2), .Q(RAM_Data[42]), .QN());
   DFF_X1 \RAM_Data_reg[41]  (.D(n_231), .CK(n_3_2), .Q(RAM_Data[41]), .QN());
   DFF_X1 \RAM_Data_reg[40]  (.D(n_230), .CK(n_3_2), .Q(RAM_Data[40]), .QN());
   DFF_X1 \RAM_Data_reg[39]  (.D(n_229), .CK(n_3_2), .Q(RAM_Data[39]), .QN());
   DFF_X1 \RAM_Data_reg[38]  (.D(n_228), .CK(n_3_2), .Q(RAM_Data[38]), .QN());
   DFF_X1 \RAM_Data_reg[37]  (.D(n_227), .CK(n_3_2), .Q(RAM_Data[37]), .QN());
   DFF_X1 \RAM_Data_reg[36]  (.D(n_226), .CK(n_3_2), .Q(RAM_Data[36]), .QN());
   DFF_X1 \RAM_Data_reg[35]  (.D(n_225), .CK(n_3_2), .Q(RAM_Data[35]), .QN());
   DFF_X1 \RAM_Data_reg[34]  (.D(n_224), .CK(n_3_2), .Q(RAM_Data[34]), .QN());
   DFF_X1 \RAM_Data_reg[33]  (.D(n_223), .CK(n_3_2), .Q(RAM_Data[33]), .QN());
   DFF_X1 \RAM_Data_reg[32]  (.D(n_222), .CK(n_3_2), .Q(RAM_Data[32]), .QN());
   DFF_X1 \RAM_Data_reg[31]  (.D(n_221), .CK(n_3_2), .Q(RAM_Data[31]), .QN());
   DFF_X1 \RAM_Data_reg[30]  (.D(n_220), .CK(n_3_2), .Q(RAM_Data[30]), .QN());
   DFF_X1 \RAM_Data_reg[29]  (.D(n_219), .CK(n_3_2), .Q(RAM_Data[29]), .QN());
   DFF_X1 \RAM_Data_reg[28]  (.D(n_218), .CK(n_3_2), .Q(RAM_Data[28]), .QN());
   DFF_X1 \RAM_Data_reg[27]  (.D(n_217), .CK(n_3_2), .Q(RAM_Data[27]), .QN());
   DFF_X1 \RAM_Data_reg[26]  (.D(n_216), .CK(n_3_2), .Q(RAM_Data[26]), .QN());
   DFF_X1 \RAM_Data_reg[25]  (.D(n_215), .CK(n_3_2), .Q(RAM_Data[25]), .QN());
   DFF_X1 \RAM_Data_reg[24]  (.D(n_214), .CK(n_3_2), .Q(RAM_Data[24]), .QN());
   DFF_X1 \RAM_Data_reg[23]  (.D(n_213), .CK(n_3_2), .Q(RAM_Data[23]), .QN());
   DFF_X1 \RAM_Data_reg[22]  (.D(n_212), .CK(n_3_2), .Q(RAM_Data[22]), .QN());
   DFF_X1 \RAM_Data_reg[21]  (.D(n_211), .CK(n_3_2), .Q(RAM_Data[21]), .QN());
   DFF_X1 \RAM_Data_reg[20]  (.D(n_210), .CK(n_3_2), .Q(RAM_Data[20]), .QN());
   DFF_X1 \RAM_Data_reg[19]  (.D(n_209), .CK(n_3_2), .Q(RAM_Data[19]), .QN());
   DFF_X1 \RAM_Data_reg[18]  (.D(n_208), .CK(n_3_2), .Q(RAM_Data[18]), .QN());
   DFF_X1 \RAM_Data_reg[17]  (.D(n_207), .CK(n_3_2), .Q(RAM_Data[17]), .QN());
   DFF_X1 \RAM_Data_reg[16]  (.D(n_206), .CK(n_3_2), .Q(RAM_Data[16]), .QN());
   DFF_X1 \RAM_Data_reg[15]  (.D(n_205), .CK(n_3_2), .Q(RAM_Data[15]), .QN());
   DFF_X1 \RAM_Data_reg[14]  (.D(n_204), .CK(n_3_2), .Q(RAM_Data[14]), .QN());
   DFF_X1 \RAM_Data_reg[13]  (.D(n_203), .CK(n_3_2), .Q(RAM_Data[13]), .QN());
   DFF_X1 \RAM_Data_reg[12]  (.D(n_202), .CK(n_3_2), .Q(RAM_Data[12]), .QN());
   DFF_X1 \RAM_Data_reg[11]  (.D(n_201), .CK(n_3_2), .Q(RAM_Data[11]), .QN());
   DFF_X1 \RAM_Data_reg[10]  (.D(n_200), .CK(n_3_2), .Q(RAM_Data[10]), .QN());
   DFF_X1 \RAM_Data_reg[9]  (.D(n_199), .CK(n_3_2), .Q(RAM_Data[9]), .QN());
   DFF_X1 \RAM_Data_reg[8]  (.D(n_198), .CK(n_3_2), .Q(RAM_Data[8]), .QN());
   DFF_X1 \RAM_Data_reg[7]  (.D(n_197), .CK(n_3_2), .Q(RAM_Data[7]), .QN());
   DFF_X1 \RAM_Data_reg[6]  (.D(n_196), .CK(n_3_2), .Q(RAM_Data[6]), .QN());
   DFF_X1 \RAM_Data_reg[5]  (.D(n_195), .CK(n_3_2), .Q(RAM_Data[5]), .QN());
   DFF_X1 \RAM_Data_reg[4]  (.D(n_194), .CK(n_3_2), .Q(RAM_Data[4]), .QN());
   DFF_X1 \RAM_Data_reg[3]  (.D(n_193), .CK(n_3_2), .Q(RAM_Data[3]), .QN());
   DFF_X1 \RAM_Data_reg[2]  (.D(n_192), .CK(n_3_2), .Q(RAM_Data[2]), .QN());
   DFF_X1 \RAM_Data_reg[1]  (.D(n_191), .CK(n_3_2), .Q(RAM_Data[1]), .QN());
   DFF_X1 \RAM_Data_reg[0]  (.D(n_190), .CK(n_3_2), .Q(RAM_Data[0]), .QN());
   DFF_X1 \RAM_Address_reg[12]  (.D(n_52), .CK(n_3_2), .Q(RAM_Address[12]), 
      .QN());
   DFF_X1 \RAM_Address_reg[11]  (.D(n_51), .CK(n_3_2), .Q(RAM_Address[11]), 
      .QN());
   DFF_X1 \RAM_Address_reg[10]  (.D(n_50), .CK(n_3_2), .Q(RAM_Address[10]), 
      .QN());
   DFF_X1 \RAM_Address_reg[9]  (.D(n_49), .CK(n_3_2), .Q(RAM_Address[9]), .QN());
   DFF_X1 \RAM_Address_reg[6]  (.D(n_46), .CK(n_3_2), .Q(RAM_Address[6]), .QN());
   DFF_X1 \RAM_Address_reg[5]  (.D(n_45), .CK(n_3_2), .Q(RAM_Address[5]), .QN());
   DFF_X1 \RAM_Address_reg[4]  (.D(n_44), .CK(n_3_2), .Q(RAM_Address[4]), .QN());
   DFF_X1 \RAM_Address_reg[2]  (.D(n_42), .CK(n_3_2), .Q(RAM_Address[2]), .QN());
   DFF_X1 \RAM_Address_reg[8]  (.D(n_48), .CK(n_3_2), .Q(RAM_Address[8]), .QN());
   DFF_X1 \RAM_Address_reg[7]  (.D(n_47), .CK(n_3_2), .Q(RAM_Address[7]), .QN());
   DFF_X1 \RAM_Address_reg[3]  (.D(n_43), .CK(n_3_2), .Q(RAM_Address[3]), .QN());
   DFF_X1 \RAM_Address_reg[1]  (.D(n_41), .CK(n_3_2), .Q(RAM_Address[1]), .QN());
   DFF_X1 \RAM_Address_reg[0]  (.D(n_40), .CK(n_3_2), .Q(RAM_Address[0]), .QN());
   DFF_X1 Done_Processing_Current_Packet_reg (.D(n_152), .CK(n_3_3), .Q(
      Done_Processing_Current_Packet), .QN());
   DFF_X1 Done_Loading_reg (.D(n_3_0), .CK(CLK), .Q(Done_Loading), .QN());
   MUX2_X1 Done_Loading_reg_enable_mux_0 (.A(Done_Loading), .B(n_54), .S(n_150), 
      .Z(n_3_0));
   DFF_X1 \RowsNum_reg[15]  (.D(n_149), .CK(CLK), .Q(RowsNum[15]), .QN());
   DFF_X1 \RowsNum_reg[14]  (.D(n_148), .CK(CLK), .Q(RowsNum[14]), .QN());
   DFF_X1 \RowsNum_reg[13]  (.D(n_147), .CK(CLK), .Q(RowsNum[13]), .QN());
   DFF_X1 \RowsNum_reg[12]  (.D(n_146), .CK(CLK), .Q(RowsNum[12]), .QN());
   DFF_X1 \RowsNum_reg[11]  (.D(n_145), .CK(CLK), .Q(RowsNum[11]), .QN());
   DFF_X1 \RowsNum_reg[10]  (.D(n_144), .CK(CLK), .Q(RowsNum[10]), .QN());
   DFF_X1 \RowsNum_reg[9]  (.D(n_143), .CK(CLK), .Q(RowsNum[9]), .QN());
   DFF_X1 \RowsNum_reg[8]  (.D(n_142), .CK(CLK), .Q(RowsNum[8]), .QN());
   DFF_X1 \RowsNum_reg[7]  (.D(n_141), .CK(CLK), .Q(RowsNum[7]), .QN());
   DFF_X1 \RowsNum_reg[6]  (.D(n_140), .CK(CLK), .Q(RowsNum[6]), .QN());
   DFF_X1 \RowsNum_reg[5]  (.D(n_139), .CK(CLK), .Q(RowsNum[5]), .QN());
   DFF_X1 \RowsNum_reg[4]  (.D(n_138), .CK(CLK), .Q(RowsNum[4]), .QN());
   DFF_X1 \RowsNum_reg[3]  (.D(n_137), .CK(CLK), .Q(RowsNum[3]), .QN());
   DFF_X1 \RowsNum_reg[2]  (.D(n_136), .CK(CLK), .Q(RowsNum[2]), .QN());
   DFF_X1 \RowsNum_reg[1]  (.D(n_135), .CK(CLK), .Q(RowsNum[1]), .QN());
   DFF_X1 \RowsNum_reg[0]  (.D(n_134), .CK(CLK), .Q(RowsNum[0]), .QN());
   DFF_X1 Start_Bit_reg (.D(n_53), .CK(CLK), .Q(Start_Bit), .QN());
   DFF_X1 Row_Done_Bit_reg (.D(n_55), .CK(CLK), .Q(Row_Done_Bit), .QN());
   DFF_X1 Done_Element_reg (.D(n_154), .CK(n_3_3), .Q(Done_Element), .QN());
   CLKGATETST_X1 clk_gate_Relative_Address_reg (.CK(CLK), .E(n_38), .SE(1'b0), 
      .GCK(n_3_1));
   DFF_X1 \Relative_Address_reg[15]  (.D(n_188), .CK(n_3_1), .Q(
      Relative_Address[15]), .QN());
   DFF_X1 \Relative_Address_reg[14]  (.D(n_187), .CK(n_3_1), .Q(
      Relative_Address[14]), .QN());
   DFF_X1 \Relative_Address_reg[13]  (.D(n_186), .CK(n_3_1), .Q(
      Relative_Address[13]), .QN());
   DFF_X1 \Relative_Address_reg[12]  (.D(n_185), .CK(n_3_1), .Q(
      Relative_Address[12]), .QN());
   DFF_X1 \Relative_Address_reg[11]  (.D(n_184), .CK(n_3_1), .Q(
      Relative_Address[11]), .QN());
   DFF_X1 \Relative_Address_reg[10]  (.D(n_183), .CK(n_3_1), .Q(
      Relative_Address[10]), .QN());
   DFF_X1 \Relative_Address_reg[9]  (.D(n_182), .CK(n_3_1), .Q(
      Relative_Address[9]), .QN());
   DFF_X1 \Relative_Address_reg[8]  (.D(n_181), .CK(n_3_1), .Q(
      Relative_Address[8]), .QN());
   DFF_X1 \Relative_Address_reg[7]  (.D(n_180), .CK(n_3_1), .Q(
      Relative_Address[7]), .QN());
   DFF_X1 \Relative_Address_reg[6]  (.D(n_179), .CK(n_3_1), .Q(
      Relative_Address[6]), .QN());
   DFF_X1 \Relative_Address_reg[5]  (.D(n_178), .CK(n_3_1), .Q(
      Relative_Address[5]), .QN());
   DFF_X1 \Relative_Address_reg[4]  (.D(n_177), .CK(n_3_1), .Q(
      Relative_Address[4]), .QN());
   DFF_X1 \Relative_Address_reg[3]  (.D(n_176), .CK(n_3_1), .Q(
      Relative_Address[3]), .QN());
   DFF_X1 \Relative_Address_reg[2]  (.D(n_175), .CK(n_3_1), .Q(
      Relative_Address[2]), .QN());
   DFF_X1 \Relative_Address_reg[1]  (.D(n_174), .CK(n_3_1), .Q(
      Relative_Address[1]), .QN());
   DFF_X1 Update_Address_Indication_Bit_reg (.D(n_39), .CK(n_3_3), .Q(
      Update_Address_Indication_Bit), .QN());
   DFF_X1 Data_Bit_reg (.D(n_190), .CK(n_3_3), .Q(Data_Bit), .QN());
   DFF_X1 \Decoded_Data_reg[11]  (.D(n_201), .CK(n_3_3), .Q(n_259), .QN());
   DFF_X1 \Decoded_Data_reg[10]  (.D(n_200), .CK(n_3_3), .Q(n_260), .QN());
   DFF_X1 \Decoded_Data_reg[9]  (.D(n_199), .CK(n_3_3), .Q(n_261), .QN());
   DFF_X1 \Decoded_Data_reg[8]  (.D(n_198), .CK(n_3_3), .Q(n_262), .QN());
   DFF_X1 \Decoded_Data_reg[7]  (.D(n_197), .CK(n_3_3), .Q(n_263), .QN());
   DFF_X1 \Decoded_Data_reg[6]  (.D(n_196), .CK(n_3_3), .Q(n_264), .QN());
   DFF_X1 \Decoded_Data_reg[5]  (.D(n_195), .CK(n_3_3), .Q(n_265), .QN());
   DFF_X1 \Decoded_Data_reg[4]  (.D(n_194), .CK(n_3_3), .Q(n_266), .QN());
   DFF_X1 \Decoded_Data_reg[3]  (.D(n_193), .CK(n_3_3), .Q(n_267), .QN());
   DFF_X1 \Decoded_Data_reg[2]  (.D(n_192), .CK(n_3_3), .Q(n_268), .QN());
   DFF_X1 \Decoded_Data_reg[1]  (.D(n_191), .CK(n_3_3), .Q(n_269), .QN());
   DFF_X1 \Decoded_Data_reg[0]  (.D(n_161), .CK(n_3_3), .Q(n_270), .QN());
   DFF_X1 \Decoded_Data_reg[63]  (.D(n_253), .CK(n_3_3), .Q(n_271), .QN());
   DFF_X1 \Decoded_Data_reg[62]  (.D(n_252), .CK(n_3_3), .Q(n_272), .QN());
   DFF_X1 \Decoded_Data_reg[61]  (.D(n_251), .CK(n_3_3), .Q(n_273), .QN());
   DFF_X1 \Decoded_Data_reg[60]  (.D(n_250), .CK(n_3_3), .Q(n_274), .QN());
   DFF_X1 \Decoded_Data_reg[59]  (.D(n_249), .CK(n_3_3), .Q(n_275), .QN());
   DFF_X1 \Decoded_Data_reg[58]  (.D(n_248), .CK(n_3_3), .Q(n_276), .QN());
   DFF_X1 \Decoded_Data_reg[57]  (.D(n_247), .CK(n_3_3), .Q(n_277), .QN());
   DFF_X1 \Decoded_Data_reg[56]  (.D(n_246), .CK(n_3_3), .Q(n_278), .QN());
   DFF_X1 \Decoded_Data_reg[55]  (.D(n_245), .CK(n_3_3), .Q(n_279), .QN());
   DFF_X1 \Decoded_Data_reg[54]  (.D(n_244), .CK(n_3_3), .Q(n_280), .QN());
   DFF_X1 \Decoded_Data_reg[53]  (.D(n_243), .CK(n_3_3), .Q(n_281), .QN());
   DFF_X1 \Decoded_Data_reg[52]  (.D(n_242), .CK(n_3_3), .Q(n_282), .QN());
   DFF_X1 \Decoded_Data_reg[51]  (.D(n_241), .CK(n_3_3), .Q(n_283), .QN());
   DFF_X1 \Decoded_Data_reg[50]  (.D(n_240), .CK(n_3_3), .Q(n_284), .QN());
   DFF_X1 \Decoded_Data_reg[49]  (.D(n_239), .CK(n_3_3), .Q(n_285), .QN());
   DFF_X1 \Decoded_Data_reg[48]  (.D(n_238), .CK(n_3_3), .Q(n_286), .QN());
   DFF_X1 \Decoded_Data_reg[47]  (.D(n_237), .CK(n_3_3), .Q(n_287), .QN());
   DFF_X1 \Decoded_Data_reg[46]  (.D(n_236), .CK(n_3_3), .Q(n_288), .QN());
   DFF_X1 \Decoded_Data_reg[45]  (.D(n_235), .CK(n_3_3), .Q(n_289), .QN());
   DFF_X1 \Decoded_Data_reg[44]  (.D(n_234), .CK(n_3_3), .Q(n_290), .QN());
   DFF_X1 \Decoded_Data_reg[43]  (.D(n_233), .CK(n_3_3), .Q(n_291), .QN());
   DFF_X1 \Decoded_Data_reg[42]  (.D(n_232), .CK(n_3_3), .Q(n_292), .QN());
   DFF_X1 \Decoded_Data_reg[41]  (.D(n_231), .CK(n_3_3), .Q(n_293), .QN());
   DFF_X1 \Decoded_Data_reg[40]  (.D(n_230), .CK(n_3_3), .Q(n_294), .QN());
   DFF_X1 \Decoded_Data_reg[39]  (.D(n_229), .CK(n_3_3), .Q(n_295), .QN());
   DFF_X1 \Decoded_Data_reg[38]  (.D(n_228), .CK(n_3_3), .Q(n_296), .QN());
   DFF_X1 \Decoded_Data_reg[37]  (.D(n_227), .CK(n_3_3), .Q(n_297), .QN());
   DFF_X1 \Decoded_Data_reg[36]  (.D(n_226), .CK(n_3_3), .Q(n_298), .QN());
   DFF_X1 \Decoded_Data_reg[35]  (.D(n_225), .CK(n_3_3), .Q(n_299), .QN());
   DFF_X1 \Decoded_Data_reg[34]  (.D(n_224), .CK(n_3_3), .Q(n_300), .QN());
   DFF_X1 \Decoded_Data_reg[33]  (.D(n_223), .CK(n_3_3), .Q(n_301), .QN());
   DFF_X1 \Decoded_Data_reg[32]  (.D(n_222), .CK(n_3_3), .Q(n_302), .QN());
   DFF_X1 \Decoded_Data_reg[31]  (.D(n_221), .CK(n_3_3), .Q(n_303), .QN());
   DFF_X1 \Decoded_Data_reg[30]  (.D(n_220), .CK(n_3_3), .Q(n_304), .QN());
   DFF_X1 \Decoded_Data_reg[29]  (.D(n_219), .CK(n_3_3), .Q(n_305), .QN());
   DFF_X1 \Decoded_Data_reg[28]  (.D(n_218), .CK(n_3_3), .Q(n_306), .QN());
   DFF_X1 \Decoded_Data_reg[27]  (.D(n_217), .CK(n_3_3), .Q(n_307), .QN());
   DFF_X1 \Decoded_Data_reg[26]  (.D(n_216), .CK(n_3_3), .Q(n_308), .QN());
   DFF_X1 \Decoded_Data_reg[25]  (.D(n_215), .CK(n_3_3), .Q(n_309), .QN());
   DFF_X1 \Decoded_Data_reg[24]  (.D(n_214), .CK(n_3_3), .Q(n_310), .QN());
   DFF_X1 \Decoded_Data_reg[23]  (.D(n_213), .CK(n_3_3), .Q(n_311), .QN());
   DFF_X1 \Decoded_Data_reg[22]  (.D(n_212), .CK(n_3_3), .Q(n_312), .QN());
   DFF_X1 \Decoded_Data_reg[21]  (.D(n_211), .CK(n_3_3), .Q(n_313), .QN());
   DFF_X1 \Decoded_Data_reg[20]  (.D(n_210), .CK(n_3_3), .Q(n_314), .QN());
   DFF_X1 \Decoded_Data_reg[19]  (.D(n_209), .CK(n_3_3), .Q(n_315), .QN());
   DFF_X1 \Decoded_Data_reg[18]  (.D(n_208), .CK(n_3_3), .Q(n_316), .QN());
   DFF_X1 \Decoded_Data_reg[17]  (.D(n_207), .CK(n_3_3), .Q(n_317), .QN());
   DFF_X1 \Decoded_Data_reg[16]  (.D(n_206), .CK(n_3_3), .Q(n_318), .QN());
   DFF_X1 \Decoded_Data_reg[15]  (.D(n_205), .CK(n_3_3), .Q(n_319), .QN());
   DFF_X1 \Decoded_Data_reg[14]  (.D(n_204), .CK(n_3_3), .Q(n_320), .QN());
   DFF_X1 \Decoded_Data_reg[13]  (.D(n_203), .CK(n_3_3), .Q(n_321), .QN());
   DFF_X1 \Writing_Start_Index_reg[5]  (.D(n_160), .CK(n_3_3), .Q(
      Writing_Start_Index[5]), .QN());
   DFF_X1 \Writing_Start_Index_reg[4]  (.D(n_159), .CK(n_3_3), .Q(
      Writing_Start_Index[4]), .QN());
   DFF_X1 \Writing_Start_Index_reg[3]  (.D(n_158), .CK(n_3_3), .Q(
      Writing_Start_Index[3]), .QN());
   DFF_X1 \Writing_Start_Index_reg[2]  (.D(n_157), .CK(n_3_3), .Q(
      Writing_Start_Index[2]), .QN());
   DFF_X1 \Writing_Start_Index_reg[1]  (.D(n_156), .CK(n_3_3), .Q(
      Writing_Start_Index[1]), .QN());
   DFF_X1 \Writing_Start_Index_reg[0]  (.D(n_155), .CK(n_3_3), .Q(
      Writing_Start_Index[0]), .QN());
   DFF_X1 \Decoded_Data_reg[12]  (.D(n_202), .CK(n_3_3), .Q(n_322), .QN());
   DFF_X1 \N_reg[11]  (.D(n_173), .CK(n_3_3), .Q(N[11]), .QN());
   DFF_X1 \N_reg[10]  (.D(n_172), .CK(n_3_3), .Q(N[10]), .QN());
   DFF_X1 \N_reg[9]  (.D(n_171), .CK(n_3_3), .Q(N[9]), .QN());
   DFF_X1 \N_reg[8]  (.D(n_170), .CK(n_3_3), .Q(N[8]), .QN());
   DFF_X1 \N_reg[7]  (.D(n_169), .CK(n_3_3), .Q(N[7]), .QN());
   DFF_X1 \N_reg[6]  (.D(n_168), .CK(n_3_3), .Q(N[6]), .QN());
   DFF_X1 \N_reg[5]  (.D(n_167), .CK(n_3_3), .Q(N[5]), .QN());
   DFF_X1 \N_reg[4]  (.D(n_166), .CK(n_3_3), .Q(N[4]), .QN());
   DFF_X1 \N_reg[3]  (.D(n_165), .CK(n_3_3), .Q(N[3]), .QN());
   DFF_X1 \N_reg[2]  (.D(n_164), .CK(n_3_3), .Q(N[2]), .QN());
   DFF_X1 \N_reg[1]  (.D(n_163), .CK(n_3_3), .Q(N[1]), .QN());
   DFF_X1 \N_reg[0]  (.D(n_162), .CK(n_3_3), .Q(N[0]), .QN());
   DFF_X1 N_Indication_Bit_reg (.D(n_153), .CK(n_3_3), .Q(N_Indication_Bit), 
      .QN());
   DFF_X1 Row_Last_Bit_reg (.D(n_133), .CK(n_3_3), .Q(Row_Last_Bit), .QN());
   DFF_X1 \Small_Packet_Indication_Bit_Location_reg[5]  (.D(n_132), .CK(CLK), 
      .Q(Small_Packet_Indication_Bit_Location[5]), .QN());
   DFF_X1 \Small_Packet_Indication_Bit_Location_reg[4]  (.D(n_131), .CK(CLK), 
      .Q(Small_Packet_Indication_Bit_Location[4]), .QN());
   DFF_X1 \Small_Packet_Indication_Bit_Location_reg[3]  (.D(n_130), .CK(CLK), 
      .Q(Small_Packet_Indication_Bit_Location[3]), .QN());
   DFF_X1 \Small_Packet_Indication_Bit_Location_reg[2]  (.D(n_129), .CK(CLK), 
      .Q(Small_Packet_Indication_Bit_Location[2]), .QN());
   DFF_X1 \Small_Packet_Indication_Bit_Location_reg[1]  (.D(n_128), .CK(CLK), 
      .Q(Small_Packet_Indication_Bit_Location[1]), .QN());
   DFF_X1 \Small_Packet_Indication_Bit_Location_reg[0]  (.D(n_127), .CK(CLK), 
      .Q(Small_Packet_Indication_Bit_Location[0]), .QN());
   DFF_X1 \PacketSize_reg[5]  (.D(n_93), .CK(CLK), .Q(PacketSize[5]), .QN());
   DFF_X1 \PacketSize_reg[4]  (.D(n_92), .CK(CLK), .Q(PacketSize[4]), .QN());
   DFF_X1 \PacketSize_reg[3]  (.D(n_91), .CK(CLK), .Q(PacketSize[3]), .QN());
   DFF_X1 \PacketSize_reg[2]  (.D(n_90), .CK(CLK), .Q(PacketSize[2]), .QN());
   DFF_X1 \PacketSize_reg[1]  (.D(n_89), .CK(CLK), .Q(PacketSize[1]), .QN());
   DFF_X1 \PacketSize_reg[0]  (.D(n_88), .CK(CLK), .Q(PacketSize[0]), .QN());
   DFF_X1 \Data_Size_reg[31]  (.D(n_87), .CK(n_3_3), .Q(Data_Size[31]), .QN());
   DFF_X1 \Data_Size_reg[30]  (.D(n_86), .CK(n_3_3), .Q(Data_Size[30]), .QN());
   DFF_X1 \Data_Size_reg[29]  (.D(n_85), .CK(n_3_3), .Q(Data_Size[29]), .QN());
   DFF_X1 \Data_Size_reg[28]  (.D(n_84), .CK(n_3_3), .Q(Data_Size[28]), .QN());
   DFF_X1 \Data_Size_reg[27]  (.D(n_83), .CK(n_3_3), .Q(Data_Size[27]), .QN());
   DFF_X1 \Data_Size_reg[26]  (.D(n_82), .CK(n_3_3), .Q(Data_Size[26]), .QN());
   DFF_X1 \Data_Size_reg[25]  (.D(n_81), .CK(n_3_3), .Q(Data_Size[25]), .QN());
   DFF_X1 \Data_Size_reg[24]  (.D(n_80), .CK(n_3_3), .Q(Data_Size[24]), .QN());
   DFF_X1 \Data_Size_reg[23]  (.D(n_79), .CK(n_3_3), .Q(Data_Size[23]), .QN());
   DFF_X1 \Data_Size_reg[22]  (.D(n_78), .CK(n_3_3), .Q(Data_Size[22]), .QN());
   DFF_X1 \Data_Size_reg[21]  (.D(n_77), .CK(n_3_3), .Q(Data_Size[21]), .QN());
   DFF_X1 \Data_Size_reg[20]  (.D(n_76), .CK(n_3_3), .Q(Data_Size[20]), .QN());
   DFF_X1 \Data_Size_reg[19]  (.D(n_75), .CK(n_3_3), .Q(Data_Size[19]), .QN());
   DFF_X1 \Data_Size_reg[18]  (.D(n_74), .CK(n_3_3), .Q(Data_Size[18]), .QN());
   DFF_X1 \Data_Size_reg[17]  (.D(n_73), .CK(n_3_3), .Q(Data_Size[17]), .QN());
   DFF_X1 \Data_Size_reg[16]  (.D(n_72), .CK(n_3_3), .Q(Data_Size[16]), .QN());
   DFF_X1 \Data_Size_reg[15]  (.D(n_71), .CK(n_3_3), .Q(Data_Size[15]), .QN());
   DFF_X1 \Data_Size_reg[14]  (.D(n_70), .CK(n_3_3), .Q(Data_Size[14]), .QN());
   DFF_X1 \Data_Size_reg[13]  (.D(n_69), .CK(n_3_3), .Q(Data_Size[13]), .QN());
   DFF_X1 \Data_Size_reg[12]  (.D(n_68), .CK(n_3_3), .Q(Data_Size[12]), .QN());
   DFF_X1 \Data_Size_reg[11]  (.D(n_67), .CK(n_3_3), .Q(Data_Size[11]), .QN());
   DFF_X1 \Data_Size_reg[10]  (.D(n_66), .CK(n_3_3), .Q(Data_Size[10]), .QN());
   DFF_X1 \Data_Size_reg[9]  (.D(n_65), .CK(n_3_3), .Q(Data_Size[9]), .QN());
   DFF_X1 \Data_Size_reg[8]  (.D(n_64), .CK(n_3_3), .Q(Data_Size[8]), .QN());
   DFF_X1 \Data_Size_reg[7]  (.D(n_63), .CK(n_3_3), .Q(Data_Size[7]), .QN());
   DFF_X1 \Data_Size_reg[6]  (.D(n_62), .CK(n_3_3), .Q(Data_Size[6]), .QN());
   DFF_X1 \Data_Size_reg[5]  (.D(n_61), .CK(n_3_3), .Q(Data_Size[5]), .QN());
   DFF_X1 \Data_Size_reg[4]  (.D(n_60), .CK(n_3_3), .Q(Data_Size[4]), .QN());
   DFF_X1 \Data_Size_reg[3]  (.D(n_59), .CK(n_3_3), .Q(Data_Size[3]), .QN());
   DFF_X1 \Data_Size_reg[2]  (.D(n_58), .CK(n_3_3), .Q(Data_Size[2]), .QN());
   DFF_X1 \Data_Size_reg[1]  (.D(n_57), .CK(n_3_3), .Q(Data_Size[1]), .QN());
   DFF_X1 \Data_Size_reg[0]  (.D(n_56), .CK(n_3_3), .Q(Data_Size[0]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[31]  (.D(n_125), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[31]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[30]  (.D(n_124), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[30]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[29]  (.D(n_123), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[29]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[28]  (.D(n_122), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[28]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[27]  (.D(n_121), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[27]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[26]  (.D(n_120), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[26]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[25]  (.D(n_119), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[25]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[24]  (.D(n_118), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[24]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[23]  (.D(n_117), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[23]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[22]  (.D(n_116), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[22]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[21]  (.D(n_115), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[21]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[20]  (.D(n_114), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[20]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[19]  (.D(n_113), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[19]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[18]  (.D(n_112), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[18]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[17]  (.D(n_111), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[17]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[16]  (.D(n_110), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[16]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[15]  (.D(n_109), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[15]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[14]  (.D(n_108), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[14]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[13]  (.D(n_107), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[13]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[12]  (.D(n_106), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[12]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[11]  (.D(n_105), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[11]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[10]  (.D(n_104), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[10]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[9]  (.D(n_103), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[9]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[8]  (.D(n_102), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[8]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[7]  (.D(n_101), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[7]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[6]  (.D(n_100), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[6]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[5]  (.D(n_99), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[5]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[4]  (.D(n_98), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[4]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[3]  (.D(n_97), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[3]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[2]  (.D(n_96), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[2]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[1]  (.D(n_95), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[1]), .QN());
   DFF_X1 \Small_Packet_Data_Size_reg[0]  (.D(n_94), .CK(n_3_3), .Q(
      Small_Packet_Data_Size[0]), .QN());
   CLKGATETST_X1 clk_gate_RAM_Data_reg (.CK(CLK), .E(n_189), .SE(1'b0), .GCK(
      n_3_2));
   CLKGATETST_X1 clk_gate_Done_Processing_Current_Packet_reg (.CK(CLK), .E(n_126), 
      .SE(1'b0), .GCK(n_3_3));
   Counter__parameterized0 Rows_Counter (.value(RowsCount), .Enable(n_0_4), 
      .CLK(CLK), .RST(n_0_0));
   DFlipFlop__4_2 Delay (.D(Done_Element), .CLK(CLK), .RST(RST), .Enable(n_0_3), 
      .Q(Done_Element_Delayed));
   Counter Init_Counter (.value(InitCount), .Enable(n_0_2), .CLK(CLK), .RST(RST));
   DFlipFlop Delay2 (.D(Row_Done_Bit), .CLK(CLK), .RST(RST), .Enable(n_0_1), 
      .Q(Row_Done_Bit_Delayed));
   OR2_X1 i_0_0_0 (.A1(RST), .A2(n_323), .ZN(n_0_0));
   NOR4_X1 i_0_0_1 (.A1(n_0_0_15), .A2(n_0_0_10), .A3(n_0_0_5), .A4(n_0_0_0), 
      .ZN(n_323));
   NAND4_X1 i_0_0_2 (.A1(n_0_0_4), .A2(n_0_0_3), .A3(n_0_0_2), .A4(n_0_0_1), 
      .ZN(n_0_0_0));
   XNOR2_X1 i_0_0_3 (.A(RowsNum[3]), .B(RowsCount[3]), .ZN(n_0_0_1));
   XNOR2_X1 i_0_0_4 (.A(RowsNum[11]), .B(RowsCount[11]), .ZN(n_0_0_2));
   XNOR2_X1 i_0_0_5 (.A(RowsNum[0]), .B(RowsCount[0]), .ZN(n_0_0_3));
   XNOR2_X1 i_0_0_6 (.A(RowsNum[12]), .B(RowsCount[12]), .ZN(n_0_0_4));
   NAND4_X1 i_0_0_7 (.A1(n_0_0_9), .A2(n_0_0_8), .A3(n_0_0_7), .A4(n_0_0_6), 
      .ZN(n_0_0_5));
   XNOR2_X1 i_0_0_8 (.A(RowsNum[13]), .B(RowsCount[13]), .ZN(n_0_0_6));
   XNOR2_X1 i_0_0_9 (.A(RowsNum[8]), .B(RowsCount[8]), .ZN(n_0_0_7));
   XNOR2_X1 i_0_0_10 (.A(RowsNum[15]), .B(RowsCount[15]), .ZN(n_0_0_8));
   XNOR2_X1 i_0_0_11 (.A(RowsNum[6]), .B(RowsCount[6]), .ZN(n_0_0_9));
   NAND4_X1 i_0_0_12 (.A1(n_0_0_14), .A2(n_0_0_13), .A3(n_0_0_12), .A4(n_0_0_11), 
      .ZN(n_0_0_10));
   XNOR2_X1 i_0_0_13 (.A(RowsNum[2]), .B(RowsCount[2]), .ZN(n_0_0_11));
   XNOR2_X1 i_0_0_14 (.A(RowsNum[10]), .B(RowsCount[10]), .ZN(n_0_0_12));
   XNOR2_X1 i_0_0_15 (.A(RowsNum[4]), .B(RowsCount[4]), .ZN(n_0_0_13));
   XNOR2_X1 i_0_0_16 (.A(RowsNum[1]), .B(RowsCount[1]), .ZN(n_0_0_14));
   NAND4_X1 i_0_0_17 (.A1(n_0_0_19), .A2(n_0_0_18), .A3(n_0_0_17), .A4(n_0_0_16), 
      .ZN(n_0_0_15));
   XNOR2_X1 i_0_0_18 (.A(RowsNum[5]), .B(RowsCount[5]), .ZN(n_0_0_16));
   XNOR2_X1 i_0_0_19 (.A(RowsNum[7]), .B(RowsCount[7]), .ZN(n_0_0_17));
   XNOR2_X1 i_0_0_20 (.A(RowsNum[14]), .B(RowsCount[14]), .ZN(n_0_0_18));
   XNOR2_X1 i_0_0_21 (.A(RowsNum[9]), .B(RowsCount[9]), .ZN(n_0_0_19));
   INV_X1 i_0_1_0 (.A(n_0_1_0), .ZN(n_0_1));
   AOI21_X1 i_0_1_1 (.A(Row_Done_Bit), .B1(n_324), .B2(Row_Done_Bit_Delayed), 
      .ZN(n_0_1_0));
   NOR2_X1 i_0_1_2 (.A1(Done_Loading), .A2(InitCount[1]), .ZN(n_0_2));
   OR2_X1 i_0_1_3 (.A1(Done_Element), .A2(Done_Element_Delayed), .ZN(n_0_3));
   NOR2_X1 i_0_1_4 (.A1(Done_Loading), .A2(n_0_1_1), .ZN(n_0_4));
   NAND2_X1 i_0_1_5 (.A1(Start_Bit), .A2(Row_Done_Bit), .ZN(n_0_1_1));
   INV_X1 i_0_1_6 (.A(Done_Element), .ZN(n_324));
endmodule

module Results_Sender(RST, CLK, Sending_Enable, CPU_Bus, Done_Sending, 
      RAM_Data_A, RAM_Data_B, RAM_Address_A, RAM_Address_B);
   input RST;
   input CLK;
   input Sending_Enable;
   output [31:0]CPU_Bus;
   output Done_Sending;
   input [63:0]RAM_Data_A;
   input [63:0]RAM_Data_B;
   output [12:0]RAM_Address_A;
   output [12:0]RAM_Address_B;

   wire n_0_0;

   DFF_X1 \CPU_Bus_reg[31]  (.D(n_31), .CK(CLK), .Q(CPU_Bus[31]), .QN());
   DFF_X1 \CPU_Bus_reg[30]  (.D(n_30), .CK(CLK), .Q(CPU_Bus[30]), .QN());
   DFF_X1 \CPU_Bus_reg[29]  (.D(n_29), .CK(CLK), .Q(CPU_Bus[29]), .QN());
   DFF_X1 \CPU_Bus_reg[28]  (.D(n_28), .CK(CLK), .Q(CPU_Bus[28]), .QN());
   DFF_X1 \CPU_Bus_reg[27]  (.D(n_27), .CK(CLK), .Q(CPU_Bus[27]), .QN());
   DFF_X1 \CPU_Bus_reg[26]  (.D(n_26), .CK(CLK), .Q(CPU_Bus[26]), .QN());
   DFF_X1 \CPU_Bus_reg[25]  (.D(n_25), .CK(CLK), .Q(CPU_Bus[25]), .QN());
   DFF_X1 \CPU_Bus_reg[24]  (.D(n_24), .CK(CLK), .Q(CPU_Bus[24]), .QN());
   DFF_X1 \CPU_Bus_reg[23]  (.D(n_23), .CK(CLK), .Q(CPU_Bus[23]), .QN());
   DFF_X1 \CPU_Bus_reg[22]  (.D(n_22), .CK(CLK), .Q(CPU_Bus[22]), .QN());
   DFF_X1 \CPU_Bus_reg[21]  (.D(n_21), .CK(CLK), .Q(CPU_Bus[21]), .QN());
   DFF_X1 \CPU_Bus_reg[20]  (.D(n_20), .CK(CLK), .Q(CPU_Bus[20]), .QN());
   DFF_X1 \CPU_Bus_reg[19]  (.D(n_19), .CK(CLK), .Q(CPU_Bus[19]), .QN());
   DFF_X1 \CPU_Bus_reg[18]  (.D(n_18), .CK(CLK), .Q(CPU_Bus[18]), .QN());
   DFF_X1 \CPU_Bus_reg[17]  (.D(n_17), .CK(CLK), .Q(CPU_Bus[17]), .QN());
   DFF_X1 \CPU_Bus_reg[16]  (.D(n_16), .CK(CLK), .Q(CPU_Bus[16]), .QN());
   DFF_X1 \CPU_Bus_reg[15]  (.D(n_15), .CK(CLK), .Q(CPU_Bus[15]), .QN());
   DFF_X1 \CPU_Bus_reg[14]  (.D(n_14), .CK(CLK), .Q(CPU_Bus[14]), .QN());
   DFF_X1 \CPU_Bus_reg[13]  (.D(n_13), .CK(CLK), .Q(CPU_Bus[13]), .QN());
   DFF_X1 \CPU_Bus_reg[12]  (.D(n_12), .CK(CLK), .Q(CPU_Bus[12]), .QN());
   DFF_X1 \CPU_Bus_reg[11]  (.D(n_11), .CK(CLK), .Q(CPU_Bus[11]), .QN());
   DFF_X1 \CPU_Bus_reg[10]  (.D(n_10), .CK(CLK), .Q(CPU_Bus[10]), .QN());
   DFF_X1 \CPU_Bus_reg[9]  (.D(n_9), .CK(CLK), .Q(CPU_Bus[9]), .QN());
   DFF_X1 \CPU_Bus_reg[8]  (.D(n_8), .CK(CLK), .Q(CPU_Bus[8]), .QN());
   DFF_X1 \CPU_Bus_reg[7]  (.D(n_7), .CK(CLK), .Q(CPU_Bus[7]), .QN());
   DFF_X1 \CPU_Bus_reg[6]  (.D(n_6), .CK(CLK), .Q(CPU_Bus[6]), .QN());
   DFF_X1 \CPU_Bus_reg[5]  (.D(n_5), .CK(CLK), .Q(CPU_Bus[5]), .QN());
   DFF_X1 \CPU_Bus_reg[4]  (.D(n_4), .CK(CLK), .Q(CPU_Bus[4]), .QN());
   DFF_X1 \CPU_Bus_reg[3]  (.D(n_3), .CK(CLK), .Q(CPU_Bus[3]), .QN());
   DFF_X1 \CPU_Bus_reg[2]  (.D(n_2), .CK(CLK), .Q(CPU_Bus[2]), .QN());
   DFF_X1 \CPU_Bus_reg[1]  (.D(n_1), .CK(CLK), .Q(CPU_Bus[1]), .QN());
   DFF_X1 \CPU_Bus_reg[0]  (.D(n_0), .CK(CLK), .Q(CPU_Bus[0]), .QN());
   AND2_X1 i_0_0 (.A1(n_0_0), .A2(RAM_Data_A[0]), .ZN(n_0));
   AND2_X1 i_0_1 (.A1(n_0_0), .A2(RAM_Data_A[1]), .ZN(n_1));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(RAM_Data_A[2]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(RAM_Data_A[3]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(RAM_Data_A[4]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(RAM_Data_A[5]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(RAM_Data_A[6]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(RAM_Data_A[7]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(RAM_Data_A[8]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(RAM_Data_A[9]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(RAM_Data_A[10]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(RAM_Data_A[11]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(RAM_Data_A[12]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(RAM_Data_A[13]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(RAM_Data_A[14]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(RAM_Data_A[15]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(RAM_Data_A[16]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(RAM_Data_A[17]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(RAM_Data_A[18]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(RAM_Data_A[19]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(RAM_Data_A[20]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(RAM_Data_A[21]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(RAM_Data_A[22]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(RAM_Data_A[23]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(RAM_Data_A[24]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(RAM_Data_A[25]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(RAM_Data_A[26]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(RAM_Data_A[27]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(RAM_Data_A[28]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(RAM_Data_A[29]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(RAM_Data_A[30]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(RAM_Data_A[31]), .ZN(n_31));
   INV_X1 i_0_32 (.A(RST), .ZN(n_0_0));
endmodule

module IO_Module(RST, CLK, INT, Load_Process, CPU_Bus, Done_Loading, 
      Done_Processing_Current_Packet, Done_Processing, IO_Memory_WR_Enable, 
      RAM_Data_RD_A, RAM_Data_RD_B, RAM_Data_WR, RAM_Address_RD_A, 
      RAM_Address_RD_B, RAM_Address_WR);
   input RST;
   input CLK;
   input INT;
   input Load_Process;
   inout [31:0]CPU_Bus;
   output Done_Loading;
   output Done_Processing_Current_Packet;
   output Done_Processing;
   output IO_Memory_WR_Enable;
   input [63:0]RAM_Data_RD_A;
   input [63:0]RAM_Data_RD_B;
   output [63:0]RAM_Data_WR;
   output [12:0]RAM_Address_RD_A;
   output [12:0]RAM_Address_RD_B;
   output [12:0]RAM_Address_WR;

   assign RAM_Address_RD_A[12] = 1'b0;
   assign RAM_Address_RD_A[11] = 1'b0;
   assign RAM_Address_RD_A[10] = 1'b0;
   assign RAM_Address_RD_A[9] = 1'b0;
   assign RAM_Address_RD_A[8] = 1'b0;
   assign RAM_Address_RD_A[7] = 1'b0;
   assign RAM_Address_RD_A[6] = 1'b0;
   assign RAM_Address_RD_A[5] = 1'b0;
   assign RAM_Address_RD_A[4] = 1'b0;
   assign RAM_Address_RD_A[3] = 1'b0;
   assign RAM_Address_RD_A[2] = 1'b0;
   assign RAM_Address_RD_A[1] = 1'b0;
   assign RAM_Address_RD_A[0] = 1'b0;
   assign RAM_Address_RD_B[12] = 1'b0;
   assign RAM_Address_RD_B[11] = 1'b0;
   assign RAM_Address_RD_B[10] = 1'b0;
   assign RAM_Address_RD_B[9] = 1'b0;
   assign RAM_Address_RD_B[8] = 1'b0;
   assign RAM_Address_RD_B[7] = 1'b0;
   assign RAM_Address_RD_B[6] = 1'b0;
   assign RAM_Address_RD_B[5] = 1'b0;
   assign RAM_Address_RD_B[4] = 1'b0;
   assign RAM_Address_RD_B[3] = 1'b0;
   assign RAM_Address_RD_B[2] = 1'b0;
   assign RAM_Address_RD_B[1] = 1'b0;
   assign RAM_Address_RD_B[0] = 1'b0;

   Decoder_Receiver DR (.RST(RST), .CLK(CLK), .CPU_Bus(CPU_Bus), .Loading_Enable(), 
      .Done_Loading(Done_Loading), .Done_Processing_Current_Packet(
      Done_Processing_Current_Packet), .Done_Element(IO_Memory_WR_Enable), 
      .RAM_Address(RAM_Address_WR), .RAM_Data(RAM_Data_WR));
   Results_Sender RS (.RST(RST), .CLK(CLK), .Sending_Enable(), .CPU_Bus(CPU_Bus), 
      .Done_Sending(), .RAM_Data_A({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, 
      uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, 
      uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, 
      uc_28, uc_29, uc_30, uc_31, RAM_Data_RD_A[31], RAM_Data_RD_A[30], 
      RAM_Data_RD_A[29], RAM_Data_RD_A[28], RAM_Data_RD_A[27], RAM_Data_RD_A[26], 
      RAM_Data_RD_A[25], RAM_Data_RD_A[24], RAM_Data_RD_A[23], RAM_Data_RD_A[22], 
      RAM_Data_RD_A[21], RAM_Data_RD_A[20], RAM_Data_RD_A[19], RAM_Data_RD_A[18], 
      RAM_Data_RD_A[17], RAM_Data_RD_A[16], RAM_Data_RD_A[15], RAM_Data_RD_A[14], 
      RAM_Data_RD_A[13], RAM_Data_RD_A[12], RAM_Data_RD_A[11], RAM_Data_RD_A[10], 
      RAM_Data_RD_A[9], RAM_Data_RD_A[8], RAM_Data_RD_A[7], RAM_Data_RD_A[6], 
      RAM_Data_RD_A[5], RAM_Data_RD_A[4], RAM_Data_RD_A[3], RAM_Data_RD_A[2], 
      RAM_Data_RD_A[1], RAM_Data_RD_A[0]}), .RAM_Data_B(), .RAM_Address_A(), 
      .RAM_Address_B());
endmodule
