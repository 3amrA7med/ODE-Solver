/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 14:46:43 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 360526778 */

module RAM(CLK, RST, WR_Enable, address_RD1, address_RD2, address_WR, dataOut1, 
      dataOut2, dataIn);
   input CLK;
   input RST;
   input WR_Enable;
   input [12:0]address_RD1;
   input [12:0]address_RD2;
   input [12:0]address_WR;
   output [63:0]dataOut1;
   output [63:0]dataOut2;
   input [63:0]dataIn;

   wire n_0_0;
   wire [63:0]\Memory[16] ;
   wire n_0_1;
   wire [63:0]\Memory[15] ;
   wire n_0_2;
   wire [63:0]\Memory[14] ;
   wire n_0_3;
   wire [63:0]\Memory[13] ;
   wire n_0_4;
   wire [63:0]\Memory[12] ;
   wire n_0_5;
   wire [63:0]\Memory[11] ;
   wire n_0_6;
   wire [63:0]\Memory[10] ;
   wire n_0_7;
   wire [63:0]\Memory[9] ;
   wire n_0_8;
   wire [63:0]\Memory[8] ;
   wire n_0_9;
   wire [63:0]\Memory[7] ;
   wire n_0_10;
   wire [63:0]\Memory[6] ;
   wire n_0_11;
   wire [63:0]\Memory[5] ;
   wire n_0_12;
   wire [63:0]\Memory[4] ;
   wire n_0_13;
   wire [63:0]\Memory[3] ;
   wire n_0_14;
   wire [63:0]\Memory[2] ;
   wire n_0_15;
   wire [63:0]\Memory[1] ;
   wire n_0_16;
   wire [63:0]\Memory[0] ;
   wire n_0_34;
   wire n_0_0_0;
   wire n_0_35;
   wire n_0_0_1;
   wire n_0_36;
   wire n_0_0_2;
   wire n_0_37;
   wire n_0_0_3;
   wire n_0_38;
   wire n_0_0_4;
   wire n_0_39;
   wire n_0_0_5;
   wire n_0_40;
   wire n_0_0_6;
   wire n_0_41;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_42;
   wire n_0_0_10;
   wire n_0_43;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_44;
   wire n_0_0_13;
   wire n_0_45;
   wire n_0_0_14;
   wire n_0_46;
   wire n_0_0_15;
   wire n_0_47;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_48;
   wire n_0_49;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_50;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_2_0;
   wire n_0_2_1;
   wire n_0_2_2;
   wire n_0_2_3;
   wire n_0_2_4;
   wire n_0_2_5;
   wire n_0_2_6;
   wire n_0_2_7;
   wire n_0_2_8;
   wire n_0_2_9;
   wire n_0_2_10;
   wire n_0_2_11;
   wire n_0_2_12;
   wire n_0_2_13;
   wire n_0_2_14;
   wire n_0_2_15;
   wire n_0_2_16;
   wire n_0_2_17;
   wire n_0_2_18;
   wire n_0_2_19;
   wire n_0_2_20;
   wire n_0_2_21;
   wire n_0_2_22;
   wire n_0_2_23;
   wire n_0_2_24;
   wire n_0_2_25;
   wire n_0_2_26;
   wire n_0_2_27;
   wire n_0_2_28;
   wire n_0_2_29;
   wire n_0_2_30;
   wire n_0_2_31;
   wire n_0_2_32;
   wire n_0_2_33;
   wire n_0_2_34;
   wire n_0_2_35;
   wire n_0_2_36;
   wire n_0_2_37;
   wire n_0_2_38;
   wire n_0_2_39;
   wire n_0_2_40;
   wire n_0_2_41;
   wire n_0_2_42;
   wire n_0_2_43;
   wire n_0_2_44;
   wire n_0_2_45;
   wire n_0_2_46;
   wire n_0_2_47;
   wire n_0_2_48;
   wire n_0_2_49;
   wire n_0_2_50;
   wire n_0_2_51;
   wire n_0_2_52;
   wire n_0_2_53;
   wire n_0_2_54;
   wire n_0_2_55;
   wire n_0_2_56;
   wire n_0_2_57;
   wire n_0_2_58;
   wire n_0_2_59;
   wire n_0_2_60;
   wire n_0_2_61;
   wire n_0_2_62;
   wire n_0_2_63;
   wire n_0_2_64;
   wire n_0_2_65;
   wire n_0_2_66;
   wire n_0_2_67;
   wire n_0_2_68;
   wire n_0_2_69;
   wire n_0_2_70;
   wire n_0_2_71;
   wire n_0_2_72;
   wire n_0_2_73;
   wire n_0_2_74;
   wire n_0_2_75;
   wire n_0_2_76;
   wire n_0_2_77;
   wire n_0_2_78;
   wire n_0_2_79;
   wire n_0_2_80;
   wire n_0_2_81;
   wire n_0_2_82;
   wire n_0_2_83;
   wire n_0_2_84;
   wire n_0_2_85;
   wire n_0_2_86;
   wire n_0_2_87;
   wire n_0_2_88;
   wire n_0_2_89;
   wire n_0_2_90;
   wire n_0_2_91;
   wire n_0_2_92;
   wire n_0_2_93;
   wire n_0_2_94;
   wire n_0_2_95;
   wire n_0_2_96;
   wire n_0_2_97;
   wire n_0_2_98;
   wire n_0_2_99;
   wire n_0_2_100;
   wire n_0_2_101;
   wire n_0_2_102;
   wire n_0_2_103;
   wire n_0_2_104;
   wire n_0_2_105;
   wire n_0_2_106;
   wire n_0_2_107;
   wire n_0_2_108;
   wire n_0_2_109;
   wire n_0_2_110;
   wire n_0_2_111;
   wire n_0_2_112;
   wire n_0_2_113;
   wire n_0_2_114;
   wire n_0_2_115;
   wire n_0_2_116;
   wire n_0_2_117;
   wire n_0_2_118;
   wire n_0_2_119;
   wire n_0_2_120;
   wire n_0_2_121;
   wire n_0_2_122;
   wire n_0_2_123;
   wire n_0_2_124;
   wire n_0_2_125;
   wire n_0_2_126;
   wire n_0_2_127;
   wire n_0_2_128;
   wire n_0_2_129;
   wire n_0_2_130;
   wire n_0_2_131;
   wire n_0_2_132;
   wire n_0_2_133;
   wire n_0_2_134;
   wire n_0_2_135;
   wire n_0_2_136;
   wire n_0_2_137;
   wire n_0_2_138;
   wire n_0_2_139;
   wire n_0_2_140;
   wire n_0_2_141;
   wire n_0_2_142;
   wire n_0_2_143;
   wire n_0_2_144;
   wire n_0_2_145;
   wire n_0_2_146;
   wire n_0_2_147;
   wire n_0_2_148;
   wire n_0_2_149;
   wire n_0_2_150;
   wire n_0_2_151;
   wire n_0_2_152;
   wire n_0_2_153;
   wire n_0_2_154;
   wire n_0_2_155;
   wire n_0_2_156;
   wire n_0_2_157;
   wire n_0_2_158;
   wire n_0_2_159;
   wire n_0_2_160;
   wire n_0_2_161;
   wire n_0_2_162;
   wire n_0_2_163;
   wire n_0_2_164;
   wire n_0_2_165;
   wire n_0_2_166;
   wire n_0_2_167;
   wire n_0_2_168;
   wire n_0_2_169;
   wire n_0_2_170;
   wire n_0_2_171;
   wire n_0_2_172;
   wire n_0_2_173;
   wire n_0_2_174;
   wire n_0_2_175;
   wire n_0_2_176;
   wire n_0_2_177;
   wire n_0_2_178;
   wire n_0_2_179;
   wire n_0_2_180;
   wire n_0_2_181;
   wire n_0_2_182;
   wire n_0_2_183;
   wire n_0_2_184;
   wire n_0_2_185;
   wire n_0_2_186;
   wire n_0_2_187;
   wire n_0_2_188;
   wire n_0_2_189;
   wire n_0_2_190;
   wire n_0_2_191;
   wire n_0_2_192;
   wire n_0_2_193;
   wire n_0_2_194;
   wire n_0_2_195;
   wire n_0_2_196;
   wire n_0_2_197;
   wire n_0_2_198;
   wire n_0_2_199;
   wire n_0_2_200;
   wire n_0_2_201;
   wire n_0_2_202;
   wire n_0_2_203;
   wire n_0_2_204;
   wire n_0_2_205;
   wire n_0_2_206;
   wire n_0_2_207;
   wire n_0_2_208;
   wire n_0_2_209;
   wire n_0_2_210;
   wire n_0_2_211;
   wire n_0_2_212;
   wire n_0_2_213;
   wire n_0_2_214;
   wire n_0_2_215;
   wire n_0_2_216;
   wire n_0_2_217;
   wire n_0_2_218;
   wire n_0_2_219;
   wire n_0_2_220;
   wire n_0_2_221;
   wire n_0_2_222;
   wire n_0_2_223;
   wire n_0_2_224;
   wire n_0_2_225;
   wire n_0_2_226;
   wire n_0_2_227;
   wire n_0_2_228;
   wire n_0_2_229;
   wire n_0_2_230;
   wire n_0_2_231;
   wire n_0_2_232;
   wire n_0_2_233;
   wire n_0_2_234;
   wire n_0_2_235;
   wire n_0_2_236;
   wire n_0_2_237;
   wire n_0_2_238;
   wire n_0_2_239;
   wire n_0_2_240;
   wire n_0_2_241;
   wire n_0_2_242;
   wire n_0_2_243;
   wire n_0_2_244;
   wire n_0_2_245;
   wire n_0_2_246;
   wire n_0_2_247;
   wire n_0_2_248;
   wire n_0_2_249;
   wire n_0_2_250;
   wire n_0_2_251;
   wire n_0_2_252;
   wire n_0_2_253;
   wire n_0_2_254;
   wire n_0_2_255;
   wire n_0_2_256;
   wire n_0_2_257;
   wire n_0_2_258;
   wire n_0_2_259;
   wire n_0_2_260;
   wire n_0_2_261;
   wire n_0_2_262;
   wire n_0_2_263;
   wire n_0_2_264;
   wire n_0_2_265;
   wire n_0_2_266;
   wire n_0_2_267;
   wire n_0_2_268;
   wire n_0_2_269;
   wire n_0_2_270;
   wire n_0_2_271;
   wire n_0_2_272;
   wire n_0_2_273;
   wire n_0_2_274;
   wire n_0_2_275;
   wire n_0_2_276;
   wire n_0_2_277;
   wire n_0_2_278;
   wire n_0_2_279;
   wire n_0_2_280;
   wire n_0_2_281;
   wire n_0_2_282;
   wire n_0_2_283;
   wire n_0_2_284;
   wire n_0_2_285;
   wire n_0_2_286;
   wire n_0_2_287;
   wire n_0_2_288;
   wire n_0_2_289;
   wire n_0_2_290;
   wire n_0_2_291;
   wire n_0_2_292;
   wire n_0_2_293;
   wire n_0_2_294;
   wire n_0_2_295;
   wire n_0_2_296;
   wire n_0_2_297;
   wire n_0_2_298;
   wire n_0_2_299;
   wire n_0_2_300;
   wire n_0_2_301;
   wire n_0_2_302;
   wire n_0_2_303;
   wire n_0_2_304;
   wire n_0_2_305;
   wire n_0_2_306;
   wire n_0_2_307;
   wire n_0_2_308;
   wire n_0_2_309;
   wire n_0_2_310;
   wire n_0_2_311;
   wire n_0_2_312;
   wire n_0_2_313;
   wire n_0_2_314;
   wire n_0_2_315;
   wire n_0_2_316;
   wire n_0_2_317;
   wire n_0_2_318;
   wire n_0_2_319;
   wire n_0_2_320;
   wire n_0_2_321;
   wire n_0_2_322;
   wire n_0_2_323;
   wire n_0_2_324;
   wire n_0_2_325;
   wire n_0_2_326;
   wire n_0_2_327;
   wire n_0_2_328;
   wire n_0_2_329;
   wire n_0_2_330;
   wire n_0_2_331;
   wire n_0_2_332;
   wire n_0_2_333;
   wire n_0_2_334;
   wire n_0_2_335;
   wire n_0_2_336;
   wire n_0_2_337;
   wire n_0_2_338;
   wire n_0_2_339;
   wire n_0_2_340;
   wire n_0_2_341;
   wire n_0_2_342;
   wire n_0_2_343;
   wire n_0_2_344;
   wire n_0_2_345;
   wire n_0_2_346;
   wire n_0_2_347;
   wire n_0_2_348;
   wire n_0_2_349;
   wire n_0_2_350;
   wire n_0_2_351;
   wire n_0_2_352;
   wire n_0_2_353;
   wire n_0_2_354;
   wire n_0_2_355;
   wire n_0_2_356;
   wire n_0_2_357;
   wire n_0_2_358;
   wire n_0_2_359;
   wire n_0_2_360;
   wire n_0_2_361;
   wire n_0_2_362;
   wire n_0_2_363;
   wire n_0_2_364;
   wire n_0_2_365;
   wire n_0_2_366;
   wire n_0_2_367;
   wire n_0_2_368;
   wire n_0_2_369;
   wire n_0_2_370;
   wire n_0_2_371;
   wire n_0_2_372;
   wire n_0_2_373;
   wire n_0_2_374;
   wire n_0_2_375;
   wire n_0_2_376;
   wire n_0_2_377;
   wire n_0_2_378;
   wire n_0_2_379;
   wire n_0_2_380;
   wire n_0_2_381;
   wire n_0_2_382;
   wire n_0_2_383;
   wire n_0_2_384;
   wire n_0_2_385;
   wire n_0_2_386;
   wire n_0_2_387;
   wire n_0_2_388;
   wire n_0_2_389;
   wire n_0_2_390;
   wire n_0_2_391;
   wire n_0_2_392;
   wire n_0_2_393;
   wire n_0_2_394;
   wire n_0_2_395;
   wire n_0_2_396;
   wire n_0_2_397;
   wire n_0_2_398;
   wire n_0_2_399;
   wire n_0_2_400;
   wire n_0_2_401;
   wire n_0_2_402;
   wire n_0_2_403;
   wire n_0_2_404;
   wire n_0_2_405;
   wire n_0_2_406;
   wire n_0_2_407;
   wire n_0_2_408;
   wire n_0_2_409;
   wire n_0_2_410;
   wire n_0_2_411;
   wire n_0_2_412;
   wire n_0_2_413;
   wire n_0_2_414;
   wire n_0_2_415;
   wire n_0_2_416;
   wire n_0_2_417;
   wire n_0_2_418;
   wire n_0_2_419;
   wire n_0_2_420;
   wire n_0_2_421;
   wire n_0_2_422;
   wire n_0_2_423;
   wire n_0_2_424;
   wire n_0_2_425;
   wire n_0_2_426;
   wire n_0_2_427;
   wire n_0_2_428;
   wire n_0_2_429;
   wire n_0_2_430;
   wire n_0_2_431;
   wire n_0_2_432;
   wire n_0_2_433;
   wire n_0_2_434;
   wire n_0_2_435;
   wire n_0_2_436;
   wire n_0_2_437;
   wire n_0_2_438;
   wire n_0_2_439;
   wire n_0_2_440;
   wire n_0_2_441;
   wire n_0_2_442;
   wire n_0_2_443;
   wire n_0_2_444;
   wire n_0_2_445;
   wire n_0_2_446;
   wire n_0_2_447;
   wire n_0_2_448;
   wire n_0_2_449;
   wire n_0_2_450;
   wire n_0_2_451;
   wire n_0_2_452;
   wire n_0_2_453;
   wire n_0_2_454;
   wire n_0_2_455;
   wire n_0_2_456;
   wire n_0_2_457;
   wire n_0_2_458;
   wire n_0_2_459;
   wire n_0_2_460;
   wire n_0_2_461;
   wire n_0_2_462;
   wire n_0_2_463;
   wire n_0_2_464;
   wire n_0_2_465;
   wire n_0_2_466;
   wire n_0_2_467;
   wire n_0_2_468;
   wire n_0_2_469;
   wire n_0_2_470;
   wire n_0_2_471;
   wire n_0_2_472;
   wire n_0_2_473;
   wire n_0_2_474;
   wire n_0_2_475;
   wire n_0_2_476;
   wire n_0_2_477;
   wire n_0_2_478;
   wire n_0_2_479;
   wire n_0_2_480;
   wire n_0_2_481;
   wire n_0_2_482;
   wire n_0_2_483;
   wire n_0_2_484;
   wire n_0_2_485;
   wire n_0_2_486;
   wire n_0_2_487;
   wire n_0_2_488;
   wire n_0_2_489;
   wire n_0_2_490;
   wire n_0_2_491;
   wire n_0_2_492;
   wire n_0_2_493;
   wire n_0_2_494;
   wire n_0_2_495;
   wire n_0_2_496;
   wire n_0_2_497;
   wire n_0_2_498;
   wire n_0_2_499;
   wire n_0_2_500;
   wire n_0_2_501;
   wire n_0_2_502;
   wire n_0_2_503;
   wire n_0_2_504;
   wire n_0_2_505;
   wire n_0_2_506;
   wire n_0_2_507;
   wire n_0_2_508;
   wire n_0_2_509;
   wire n_0_2_510;
   wire n_0_2_511;
   wire n_0_2_512;
   wire n_0_2_513;
   wire n_0_2_514;
   wire n_0_2_515;
   wire n_0_2_516;
   wire n_0_2_517;
   wire n_0_2_518;
   wire n_0_2_519;
   wire n_0_2_520;
   wire n_0_2_521;
   wire n_0_2_522;
   wire n_0_2_523;
   wire n_0_2_524;
   wire n_0_2_525;
   wire n_0_2_526;
   wire n_0_2_527;
   wire n_0_2_528;
   wire n_0_2_529;
   wire n_0_2_530;
   wire n_0_2_531;
   wire n_0_2_532;
   wire n_0_2_533;
   wire n_0_2_534;
   wire n_0_2_535;
   wire n_0_2_536;
   wire n_0_2_537;
   wire n_0_2_538;
   wire n_0_2_539;
   wire n_0_2_540;
   wire n_0_2_541;
   wire n_0_2_542;
   wire n_0_2_543;
   wire n_0_2_544;
   wire n_0_2_545;
   wire n_0_2_546;
   wire n_0_2_547;
   wire n_0_2_548;
   wire n_0_2_549;
   wire n_0_2_550;
   wire n_0_2_551;
   wire n_0_2_552;
   wire n_0_2_553;
   wire n_0_2_554;
   wire n_0_2_555;
   wire n_0_2_556;
   wire n_0_2_557;
   wire n_0_2_558;
   wire n_0_2_559;
   wire n_0_2_560;
   wire n_0_2_561;
   wire n_0_2_562;
   wire n_0_2_563;
   wire n_0_2_564;
   wire n_0_2_565;
   wire n_0_2_566;
   wire n_0_2_567;
   wire n_0_2_568;
   wire n_0_2_569;
   wire n_0_2_570;
   wire n_0_2_571;
   wire n_0_2_572;
   wire n_0_2_573;
   wire n_0_2_574;
   wire n_0_2_575;
   wire n_0_2_576;
   wire n_0_2_577;
   wire n_0_2_578;
   wire n_0_2_579;
   wire n_0_2_580;
   wire n_0_2_581;
   wire n_0_2_582;
   wire n_0_2_583;
   wire n_0_2_584;
   wire n_0_2_585;
   wire n_0_2_586;
   wire n_0_2_587;
   wire n_0_2_588;
   wire n_0_2_589;
   wire n_0_2_590;
   wire n_0_2_591;
   wire n_0_2_592;
   wire n_0_2_593;
   wire n_0_2_594;
   wire n_0_2_595;
   wire n_0_2_596;
   wire n_0_2_597;
   wire n_0_2_598;
   wire n_0_2_599;
   wire n_0_2_600;
   wire n_0_2_601;
   wire n_0_2_602;
   wire n_0_2_603;
   wire n_0_2_604;
   wire n_0_2_605;
   wire n_0_2_606;
   wire n_0_2_607;
   wire n_0_2_608;
   wire n_0_2_609;
   wire n_0_2_610;
   wire n_0_2_611;
   wire n_0_2_612;
   wire n_0_2_613;
   wire n_0_2_614;
   wire n_0_2_615;
   wire n_0_2_616;
   wire n_0_2_617;
   wire n_0_2_618;
   wire n_0_2_619;
   wire n_0_2_620;
   wire n_0_2_621;
   wire n_0_2_622;
   wire n_0_2_623;
   wire n_0_2_624;
   wire n_0_2_625;
   wire n_0_2_626;
   wire n_0_2_627;
   wire n_0_2_628;
   wire n_0_2_629;
   wire n_0_2_630;
   wire n_0_2_631;
   wire n_0_2_632;
   wire n_0_2_633;
   wire n_0_2_634;
   wire n_0_2_635;
   wire n_0_2_636;
   wire n_0_2_637;
   wire n_0_2_638;
   wire n_0_2_639;
   wire n_0_2_640;
   wire n_0_2_641;
   wire n_0_2_642;
   wire n_0_2_643;
   wire n_0_2_644;
   wire n_0_2_645;
   wire n_0_2_646;
   wire n_0_2_647;
   wire n_0_2_648;
   wire n_0_2_649;
   wire n_0_2_650;
   wire n_0_2_651;
   wire n_0_2_652;
   wire n_0_2_653;
   wire n_0_2_654;
   wire n_0_2_655;
   wire n_0_2_656;
   wire n_0_2_657;
   wire n_0_2_658;
   wire n_0_2_659;
   wire n_0_2_660;
   wire n_0_2_661;
   wire n_0_2_662;
   wire n_0_2_663;
   wire n_0_2_664;
   wire n_0_2_665;
   wire n_0_2_666;
   wire n_0_2_667;
   wire n_0_2_668;
   wire n_0_2_669;
   wire n_0_2_670;
   wire n_0_2_671;
   wire n_0_2_672;
   wire n_0_2_673;
   wire n_0_2_674;
   wire n_0_2_675;
   wire n_0_2_676;
   wire n_0_2_677;
   wire n_0_2_678;
   wire n_0_2_679;
   wire n_0_2_680;
   wire n_0_2_681;
   wire n_0_2_682;
   wire n_0_2_683;
   wire n_0_2_684;
   wire n_0_2_685;
   wire n_0_2_686;
   wire n_0_2_687;
   wire n_0_2_688;
   wire n_0_2_689;
   wire n_0_2_690;
   wire n_0_2_691;
   wire n_0_2_692;
   wire n_0_2_693;
   wire n_0_2_694;
   wire n_0_2_695;
   wire n_0_2_696;
   wire n_0_2_697;
   wire n_0_2_698;
   wire n_0_2_699;
   wire n_0_2_700;
   wire n_0_2_701;
   wire n_0_2_702;
   wire n_0_2_703;
   wire n_0_2_704;
   wire n_0_2_705;
   wire n_0_2_706;
   wire n_0_2_707;
   wire n_0_2_708;
   wire n_0_2_709;
   wire n_0_2_710;
   wire n_0_2_711;
   wire n_0_2_712;
   wire n_0_2_713;
   wire n_0_2_714;
   wire n_0_2_715;
   wire n_0_2_716;
   wire n_0_2_717;
   wire n_0_2_718;
   wire n_0_2_719;
   wire n_0_2_720;
   wire n_0_2_721;
   wire n_0_2_722;
   wire n_0_2_723;
   wire n_0_2_724;
   wire n_0_2_725;
   wire n_0_2_726;
   wire n_0_2_727;
   wire n_0_2_728;
   wire n_0_2_729;
   wire n_0_2_730;
   wire n_0_2_731;
   wire n_0_2_732;
   wire n_0_2_733;
   wire n_0_2_734;
   wire n_0_2_735;
   wire n_0_2_736;
   wire n_0_2_737;
   wire n_0_2_738;
   wire n_0_2_739;
   wire n_0_2_740;
   wire n_0_2_741;
   wire n_0_2_742;
   wire n_0_2_743;
   wire n_0_2_744;
   wire n_0_2_745;
   wire n_0_2_746;
   wire n_0_2_747;
   wire n_0_2_748;
   wire n_0_2_749;
   wire n_0_2_750;
   wire n_0_2_751;
   wire n_0_2_752;
   wire n_0_2_753;
   wire n_0_2_754;
   wire n_0_2_755;
   wire n_0_2_756;
   wire n_0_2_757;
   wire n_0_2_758;
   wire n_0_2_759;
   wire n_0_2_760;
   wire n_0_2_761;
   wire n_0_2_762;
   wire n_0_2_763;
   wire n_0_2_764;
   wire n_0_2_765;
   wire n_0_2_766;
   wire n_0_2_767;
   wire n_0_2_768;
   wire n_0_2_769;
   wire n_0_2_770;
   wire n_0_2_771;
   wire n_0_2_772;
   wire n_0_2_773;
   wire n_0_2_774;
   wire n_0_2_775;
   wire n_0_2_776;
   wire n_0_2_777;
   wire n_0_2_778;
   wire n_0_2_779;
   wire n_0_2_780;
   wire n_0_2_781;
   wire n_0_2_782;
   wire n_0_2_783;
   wire n_0_2_784;
   wire n_0_2_785;
   wire n_0_2_786;
   wire n_0_2_787;
   wire n_0_2_788;
   wire n_0_2_789;
   wire n_0_2_790;
   wire n_0_2_791;
   wire n_0_2_792;
   wire n_0_2_793;
   wire n_0_2_794;
   wire n_0_2_795;
   wire n_0_2_796;
   wire n_0_2_797;
   wire n_0_2_798;
   wire n_0_2_799;
   wire n_0_2_800;
   wire n_0_2_801;
   wire n_0_2_802;
   wire n_0_2_803;
   wire n_0_2_804;
   wire n_0_2_805;
   wire n_0_2_806;
   wire n_0_2_807;
   wire n_0_2_808;
   wire n_0_2_809;
   wire n_0_2_810;
   wire n_0_2_811;
   wire n_0_2_812;
   wire n_0_2_813;
   wire n_0_2_814;
   wire n_0_2_815;
   wire n_0_2_816;
   wire n_0_2_817;
   wire n_0_2_818;
   wire n_0_2_819;
   wire n_0_2_820;
   wire n_0_2_821;
   wire n_0_2_822;
   wire n_0_2_823;
   wire n_0_2_824;
   wire n_0_2_825;
   wire n_0_2_826;
   wire n_0_2_827;
   wire n_0_2_828;
   wire n_0_2_829;
   wire n_0_2_830;
   wire n_0_2_831;
   wire n_0_2_832;
   wire n_0_2_833;
   wire n_0_2_834;
   wire n_0_2_835;
   wire n_0_2_836;
   wire n_0_2_837;
   wire n_0_2_838;
   wire n_0_2_839;
   wire n_0_2_840;
   wire n_0_2_841;
   wire n_0_2_842;
   wire n_0_2_843;
   wire n_0_2_844;
   wire n_0_2_845;
   wire n_0_2_846;
   wire n_0_2_847;
   wire n_0_2_848;
   wire n_0_2_849;
   wire n_0_2_850;
   wire n_0_2_851;
   wire n_0_2_852;
   wire n_0_2_853;
   wire n_0_2_854;
   wire n_0_2_855;
   wire n_0_2_856;
   wire n_0_2_857;
   wire n_0_2_858;
   wire n_0_2_859;
   wire n_0_2_860;
   wire n_0_2_861;
   wire n_0_2_862;
   wire n_0_2_863;
   wire n_0_2_864;
   wire n_0_2_865;
   wire n_0_2_866;
   wire n_0_2_867;
   wire n_0_2_868;
   wire n_0_2_869;
   wire n_0_2_870;
   wire n_0_2_871;
   wire n_0_2_872;
   wire n_0_2_873;
   wire n_0_2_874;
   wire n_0_2_875;
   wire n_0_2_876;
   wire n_0_2_877;
   wire n_0_2_878;
   wire n_0_2_879;
   wire n_0_2_880;
   wire n_0_2_881;
   wire n_0_2_882;
   wire n_0_2_883;
   wire n_0_2_884;
   wire n_0_2_885;
   wire n_0_2_886;
   wire n_0_2_887;
   wire n_0_2_888;
   wire n_0_2_889;
   wire n_0_2_890;
   wire n_0_2_891;
   wire n_0_2_892;
   wire n_0_2_893;
   wire n_0_2_894;
   wire n_0_2_895;
   wire n_0_2_896;
   wire n_0_2_897;
   wire n_0_2_898;
   wire n_0_2_899;
   wire n_0_2_900;
   wire n_0_2_901;
   wire n_0_2_902;
   wire n_0_2_903;
   wire n_0_2_904;
   wire n_0_2_905;
   wire n_0_2_906;
   wire n_0_2_907;
   wire n_0_2_908;
   wire n_0_2_909;
   wire n_0_2_910;
   wire n_0_2_911;
   wire n_0_2_912;
   wire n_0_2_913;
   wire n_0_2_914;
   wire n_0_2_915;
   wire n_0_2_916;
   wire n_0_2_917;
   wire n_0_2_918;
   wire n_0_2_919;
   wire n_0_2_920;
   wire n_0_2_921;
   wire n_0_2_922;
   wire n_0_2_923;
   wire n_0_2_924;
   wire n_0_2_925;
   wire n_0_2_926;
   wire n_0_2_927;
   wire n_0_2_928;
   wire n_0_2_929;
   wire n_0_2_930;
   wire n_0_2_931;
   wire n_0_2_932;
   wire n_0_2_933;
   wire n_0_2_934;
   wire n_0_2_935;
   wire n_0_2_936;
   wire n_0_2_937;
   wire n_0_2_938;
   wire n_0_2_939;
   wire n_0_2_940;
   wire n_0_2_941;
   wire n_0_2_942;
   wire n_0_2_943;
   wire n_0_2_944;
   wire n_0_2_945;
   wire n_0_2_946;
   wire n_0_2_947;
   wire n_0_2_948;
   wire n_0_2_949;
   wire n_0_2_950;
   wire n_0_2_951;
   wire n_0_2_952;
   wire n_0_2_953;
   wire n_0_2_954;
   wire n_0_2_955;
   wire n_0_2_956;
   wire n_0_2_957;
   wire n_0_2_958;
   wire n_0_2_959;
   wire n_0_2_960;
   wire n_0_2_961;
   wire n_0_2_962;
   wire n_0_2_963;
   wire n_0_2_964;
   wire n_0_2_965;
   wire n_0_2_966;
   wire n_0_2_967;
   wire n_0_2_968;
   wire n_0_2_969;
   wire n_0_2_970;
   wire n_0_2_971;
   wire n_0_2_972;
   wire n_0_2_973;
   wire n_0_2_974;
   wire n_0_2_975;
   wire n_0_2_976;
   wire n_0_2_977;
   wire n_0_2_978;
   wire n_0_2_979;
   wire n_0_2_980;
   wire n_0_2_981;
   wire n_0_2_982;
   wire n_0_2_983;
   wire n_0_2_984;
   wire n_0_2_985;
   wire n_0_2_986;
   wire n_0_2_987;
   wire n_0_2_988;
   wire n_0_2_989;
   wire n_0_2_990;
   wire n_0_2_991;
   wire n_0_2_992;
   wire n_0_2_993;
   wire n_0_2_994;
   wire n_0_2_995;
   wire n_0_2_996;
   wire n_0_2_997;
   wire n_0_2_998;
   wire n_0_2_999;
   wire n_0_2_1000;
   wire n_0_2_1001;
   wire n_0_2_1002;
   wire n_0_2_1003;
   wire n_0_2_1004;
   wire n_0_2_1005;
   wire n_0_2_1006;
   wire n_0_2_1007;
   wire n_0_2_1008;
   wire n_0_2_1009;
   wire n_0_2_1010;
   wire n_0_2_1011;
   wire n_0_2_1012;
   wire n_0_2_1013;
   wire n_0_2_1014;
   wire n_0_2_1015;
   wire n_0_2_1016;
   wire n_0_2_1017;
   wire n_0_2_1018;
   wire n_0_2_1019;
   wire n_0_2_1020;
   wire n_0_2_1021;
   wire n_0_2_1022;
   wire n_0_2_1023;
   wire n_0_2_1024;
   wire n_0_2_1025;
   wire n_0_2_1026;
   wire n_0_2_1027;
   wire n_0_2_1028;
   wire n_0_2_1029;
   wire n_0_2_1030;
   wire n_0_2_1031;
   wire n_0_2_1032;
   wire n_0_2_1033;
   wire n_0_2_1034;
   wire n_0_2_1035;
   wire n_0_2_1036;
   wire n_0_2_1037;
   wire n_0_2_1038;
   wire n_0_2_1039;
   wire n_0_2_1040;
   wire n_0_2_1041;
   wire n_0_2_1042;
   wire n_0_2_1043;
   wire n_0_2_1044;
   wire n_0_2_1045;
   wire n_0_2_1046;
   wire n_0_2_1047;
   wire n_0_2_1048;
   wire n_0_2_1049;
   wire n_0_2_1050;
   wire n_0_2_1051;
   wire n_0_2_1052;
   wire n_0_2_1053;
   wire n_0_2_1054;
   wire n_0_2_1055;
   wire n_0_2_1056;
   wire n_0_2_1057;
   wire n_0_2_1058;
   wire n_0_2_1059;
   wire n_0_2_1060;
   wire n_0_2_1061;
   wire n_0_2_1062;
   wire n_0_2_1063;
   wire n_0_2_1064;
   wire n_0_2_1065;
   wire n_0_2_1066;
   wire n_0_2_1067;
   wire n_0_2_1068;
   wire n_0_2_1069;
   wire n_0_2_1070;
   wire n_0_2_1071;
   wire n_0_2_1072;
   wire n_0_2_1073;
   wire n_0_2_1074;
   wire n_0_2_1075;
   wire n_0_2_1076;
   wire n_0_2_1077;
   wire n_0_2_1078;
   wire n_0_2_1079;
   wire n_0_2_1080;
   wire n_0_2_1081;
   wire n_0_2_1082;
   wire n_0_2_1083;
   wire n_0_2_1084;
   wire n_0_2_1085;
   wire n_0_2_1086;
   wire n_0_2_1087;
   wire n_0_2_1088;
   wire n_0_2_1089;
   wire n_0_2_1090;
   wire n_0_2_1091;
   wire n_0_2_1092;
   wire n_0_2_1093;
   wire n_0_2_1094;
   wire n_0_2_1095;
   wire n_0_2_1096;
   wire n_0_2_1097;
   wire n_0_2_1098;
   wire n_0_2_1099;
   wire n_0_2_1100;
   wire n_0_2_1101;
   wire n_0_2_1102;
   wire n_0_2_1103;
   wire n_0_2_1104;
   wire n_0_2_1105;
   wire n_0_2_1106;
   wire n_0_2_1107;
   wire n_0_2_1108;
   wire n_0_2_1109;
   wire n_0_2_1110;
   wire n_0_2_1111;
   wire n_0_2_1112;
   wire n_0_2_1113;
   wire n_0_2_1114;
   wire n_0_2_1115;
   wire n_0_2_1116;
   wire n_0_2_1117;
   wire n_0_2_1118;
   wire n_0_2_1119;
   wire n_0_2_1120;
   wire n_0_2_1121;
   wire n_0_2_1122;
   wire n_0_2_1123;
   wire n_0_2_1124;
   wire n_0_2_1125;
   wire n_0_2_1126;
   wire n_0_2_1127;
   wire n_0_2_1128;
   wire n_0_2_1129;
   wire n_0_2_1130;
   wire n_0_2_1131;
   wire n_0_2_1132;
   wire n_0_2_1133;
   wire n_0_2_1134;
   wire n_0_2_1135;
   wire n_0_2_1136;
   wire n_0_2_1137;
   wire n_0_2_1138;
   wire n_0_2_1139;
   wire n_0_2_1140;
   wire n_0_2_1141;
   wire n_0_2_1142;
   wire n_0_2_1143;
   wire n_0_2_1144;
   wire n_0_2_1145;
   wire n_0_2_1146;
   wire n_0_2_1147;
   wire n_0_2_1148;
   wire n_0_2_1149;
   wire n_0_2_1150;
   wire n_0_2_1151;
   wire n_0_2_1152;
   wire n_0_2_1153;
   wire n_0_2_1154;
   wire n_0_2_1155;
   wire n_0_2_1156;
   wire n_0_2_1157;
   wire n_0_2_1158;
   wire n_0_2_1159;
   wire n_0_2_1160;
   wire n_0_2_1161;
   wire n_0_2_1162;
   wire n_0_2_1163;
   wire n_0_2_1164;
   wire n_0_2_1165;
   wire n_0_2_1166;
   wire n_0_2_1167;
   wire n_0_2_1168;
   wire n_0_2_1169;
   wire n_0_2_1170;
   wire n_0_2_1171;
   wire n_0_2_1172;
   wire n_0_2_1173;
   wire n_0_2_1174;
   wire n_0_2_1175;
   wire n_0_2_1176;
   wire n_0_2_1177;
   wire n_0_2_1178;
   wire n_0_2_1179;
   wire n_0_2_1180;
   wire n_0_2_1181;
   wire n_0_2_1182;
   wire n_0_2_1183;
   wire n_0_2_1184;
   wire n_0_2_1185;
   wire n_0_2_1186;
   wire n_0_2_1187;
   wire n_0_2_1188;
   wire n_0_2_1189;
   wire n_0_2_1190;
   wire n_0_2_1191;
   wire n_0_2_1192;
   wire n_0_2_1193;
   wire n_0_2_1194;
   wire n_0_2_1195;
   wire n_0_2_1196;
   wire n_0_2_1197;
   wire n_0_2_1198;
   wire n_0_2_1199;
   wire n_0_2_1200;
   wire n_0_2_1201;
   wire n_0_2_1202;
   wire n_0_2_1203;
   wire n_0_2_1204;
   wire n_0_2_1205;
   wire n_0_2_1206;
   wire n_0_2_1207;
   wire n_0_2_1208;
   wire n_0_2_1209;
   wire n_0_2_1210;
   wire n_0_2_1211;
   wire n_0_2_1212;
   wire n_0_2_1213;
   wire n_0_2_1214;
   wire n_0_2_1215;
   wire n_0_2_1216;
   wire n_0_2_1217;
   wire n_0_2_1218;
   wire n_0_2_1219;
   wire n_0_2_1220;
   wire n_0_2_1221;
   wire n_0_2_1222;
   wire n_0_2_1223;
   wire n_0_2_1224;
   wire n_0_2_1225;
   wire n_0_2_1226;
   wire n_0_2_1227;
   wire n_0_2_1228;
   wire n_0_2_1229;
   wire n_0_2_1230;
   wire n_0_2_1231;
   wire n_0_2_1232;
   wire n_0_2_1233;
   wire n_0_2_1234;
   wire n_0_2_1235;
   wire n_0_2_1236;
   wire n_0_2_1237;
   wire n_0_2_1238;
   wire n_0_2_1239;
   wire n_0_2_1240;
   wire n_0_2_1241;
   wire n_0_2_1242;
   wire n_0_2_1243;
   wire n_0_2_1244;
   wire n_0_2_1245;
   wire n_0_2_1246;
   wire n_0_2_1247;
   wire n_0_2_1248;
   wire n_0_2_1249;
   wire n_0_2_1250;
   wire n_0_2_1251;
   wire n_0_2_1252;
   wire n_0_2_1253;
   wire n_0_2_1254;
   wire n_0_2_1255;
   wire n_0_2_1256;
   wire n_0_2_1257;
   wire n_0_2_1258;
   wire n_0_2_1259;
   wire n_0_2_1260;
   wire n_0_2_1261;
   wire n_0_2_1262;
   wire n_0_2_1263;
   wire n_0_2_1264;
   wire n_0_2_1265;
   wire n_0_2_1266;
   wire n_0_2_1267;
   wire n_0_2_1268;
   wire n_0_2_1269;
   wire n_0_2_1270;
   wire n_0_2_1271;
   wire n_0_2_1272;
   wire n_0_2_1273;
   wire n_0_2_1274;
   wire n_0_2_1275;
   wire n_0_2_1276;
   wire n_0_2_1277;
   wire n_0_2_1278;
   wire n_0_2_1279;
   wire n_0_2_1280;
   wire n_0_2_1281;
   wire n_0_2_1282;
   wire n_0_2_1283;
   wire n_0_2_1284;
   wire n_0_2_1285;
   wire n_0_2_1286;
   wire n_0_2_1287;
   wire n_0_2_1288;
   wire n_0_2_1289;
   wire n_0_2_1290;
   wire n_0_2_1291;
   wire n_0_2_1292;
   wire n_0_2_1293;
   wire n_0_2_1294;
   wire n_0_2_1295;
   wire n_0_2_1296;
   wire n_0_2_1297;
   wire n_0_2_1298;
   wire n_0_2_1299;
   wire n_0_2_1300;
   wire n_0_2_1301;
   wire n_0_2_1302;
   wire n_0_2_1303;
   wire n_0_2_1304;
   wire n_0_2_1305;
   wire n_0_2_1306;
   wire n_0_2_1307;
   wire n_0_2_1308;
   wire n_0_2_1309;
   wire n_0_2_1310;
   wire n_0_2_1311;
   wire n_0_2_1312;
   wire n_0_2_1313;
   wire n_0_2_1314;
   wire n_0_2_1315;
   wire n_0_2_1316;
   wire n_0_2_1317;
   wire n_0_2_1318;
   wire n_0_2_1319;
   wire n_0_2_1320;
   wire n_0_2_1321;
   wire n_0_2_1322;
   wire n_0_2_1323;
   wire n_0_2_1324;
   wire n_0_2_1325;
   wire n_0_2_1326;
   wire n_0_2_1327;
   wire n_0_2_1328;
   wire n_0_2_1329;
   wire n_0_2_1330;
   wire n_0_2_1331;
   wire n_0_2_1332;
   wire n_0_2_1333;
   wire n_0_2_1334;
   wire n_0_2_1335;
   wire n_0_2_1336;
   wire n_0_2_1337;
   wire n_0_2_1338;
   wire n_0_2_1339;
   wire n_0_2_1340;
   wire n_0_2_1341;
   wire n_0_2_1342;
   wire n_0_2_1343;
   wire n_0_2_1344;
   wire n_0_2_1345;
   wire n_0_2_1346;
   wire n_0_2_1347;
   wire n_0_2_1348;
   wire n_0_2_1349;
   wire n_0_2_1350;
   wire n_0_2_1351;
   wire n_0_2_1352;
   wire n_0_2_1353;
   wire n_0_2_1354;
   wire n_0_2_1355;
   wire n_0_2_1356;
   wire n_0_2_1357;
   wire n_0_2_1358;
   wire n_0_2_1359;
   wire n_0_2_1360;
   wire n_0_2_1361;
   wire n_0_2_1362;
   wire n_0_2_1363;
   wire n_0_2_1364;
   wire n_0_2_1365;
   wire n_0_2_1366;
   wire n_0_2_1367;
   wire n_0_2_1368;
   wire n_0_2_1369;
   wire n_0_2_1370;
   wire n_0_2_1371;
   wire n_0_2_1372;
   wire n_0_2_1373;
   wire n_0_2_1374;
   wire n_0_2_1375;
   wire n_0_2_1376;
   wire n_0_2_1377;
   wire n_0_2_1378;
   wire n_0_2_1379;
   wire n_0_2_1380;
   wire n_0_2_1381;
   wire n_0_2_1382;
   wire n_0_2_1383;
   wire n_0_2_1384;
   wire n_0_2_1385;
   wire n_0_2_1386;
   wire n_0_2_1387;
   wire n_0_2_1388;
   wire n_0_2_1389;
   wire n_0_2_1390;
   wire n_0_2_1391;
   wire n_0_2_1392;
   wire n_0_2_1393;
   wire n_0_2_1394;
   wire n_0_2_1395;
   wire n_0_2_1396;
   wire n_0_2_1397;
   wire n_0_2_1398;
   wire n_0_2_1399;
   wire n_0_2_1400;
   wire n_0_2_1401;
   wire n_0_2_1402;
   wire n_0_2_1403;
   wire n_0_2_1404;
   wire n_0_2_1405;
   wire n_0_2_1406;
   wire n_0_2_1407;
   wire n_0_2_1408;
   wire n_0_2_1409;
   wire n_0_2_1410;
   wire n_0_2_1411;
   wire n_0_2_1412;
   wire n_0_2_1413;
   wire n_0_2_1414;
   wire n_0_2_1415;
   wire n_0_2_1416;
   wire n_0_2_1417;
   wire n_0_2_1418;
   wire n_0_2_1419;
   wire n_0_2_1420;
   wire n_0_2_1421;
   wire n_0_2_1422;
   wire n_0_2_1423;
   wire n_0_2_1424;
   wire n_0_2_1425;
   wire n_0_2_1426;
   wire n_0_2_1427;
   wire n_0_2_1428;
   wire n_0_2_1429;
   wire n_0_2_1430;
   wire n_0_2_1431;
   wire n_0_2_1432;
   wire n_0_2_1433;
   wire n_0_2_1434;
   wire n_0_2_1435;
   wire n_0_2_1436;
   wire n_0_2_1437;
   wire n_0_2_1438;
   wire n_0_2_1439;
   wire n_0_2_1440;
   wire n_0_2_1441;
   wire n_0_2_1442;
   wire n_0_2_1443;
   wire n_0_2_1444;
   wire n_0_2_1445;
   wire n_0_2_1446;
   wire n_0_2_1447;
   wire n_0_2_1448;
   wire n_0_2_1449;
   wire n_0_2_1450;
   wire n_0_2_1451;
   wire n_0_2_1452;
   wire n_0_2_1453;
   wire n_0_2_1454;
   wire n_0_2_1455;
   wire n_0_2_1456;
   wire n_0_2_1457;
   wire n_0_2_1458;
   wire n_0_2_1459;
   wire n_0_2_1460;
   wire n_0_2_1461;
   wire n_0_2_1462;
   wire n_0_2_1463;
   wire n_0_2_1464;
   wire n_0_2_1465;
   wire n_0_2_1466;
   wire n_0_2_1467;
   wire n_0_2_1468;
   wire n_0_2_1469;
   wire n_0_2_1470;
   wire n_0_2_1471;
   wire n_0_2_1472;
   wire n_0_2_1473;
   wire n_0_2_1474;
   wire n_0_2_1475;
   wire n_0_2_1476;
   wire n_0_2_1477;
   wire n_0_2_1478;
   wire n_0_2_1479;
   wire n_0_2_1480;
   wire n_0_2_1481;
   wire n_0_2_1482;
   wire n_0_2_1483;
   wire n_0_2_1484;
   wire n_0_2_1485;
   wire n_0_2_1486;
   wire n_0_2_1487;
   wire n_0_2_1488;
   wire n_0_2_1489;
   wire n_0_2_1490;
   wire n_0_2_1491;
   wire n_0_2_1492;
   wire n_0_2_1493;
   wire n_0_2_1494;
   wire n_0_2_1495;
   wire n_0_2_1496;
   wire n_0_2_1497;
   wire n_0_2_1498;
   wire n_0_2_1499;
   wire n_0_2_1500;
   wire n_0_2_1501;
   wire n_0_2_1502;
   wire n_0_2_1503;
   wire n_0_2_1504;
   wire n_0_2_1505;
   wire n_0_2_1506;
   wire n_0_2_1507;
   wire n_0_2_1508;
   wire n_0_2_1509;
   wire n_0_2_1510;
   wire n_0_2_1511;
   wire n_0_2_1512;
   wire n_0_2_1513;
   wire n_0_2_1514;
   wire n_0_2_1515;
   wire n_0_2_1516;
   wire n_0_2_1517;
   wire n_0_2_1518;
   wire n_0_2_1519;
   wire n_0_2_1520;
   wire n_0_2_1521;
   wire n_0_2_1522;
   wire n_0_2_1523;
   wire n_0_2_1524;
   wire n_0_2_1525;
   wire n_0_2_1526;
   wire n_0_2_1527;
   wire n_0_2_1528;
   wire n_0_2_1529;
   wire n_0_2_1530;
   wire n_0_2_1531;
   wire n_0_2_1532;
   wire n_0_2_1533;
   wire n_0_2_1534;
   wire n_0_2_1535;
   wire n_0_2_1536;
   wire n_0_2_1537;
   wire n_0_2_1538;
   wire n_0_2_1539;
   wire n_0_2_1540;
   wire n_0_2_1541;
   wire n_0_2_1542;
   wire n_0_2_1543;
   wire n_0_2_1544;
   wire n_0_2_1545;
   wire n_0_2_1546;
   wire n_0_2_1547;
   wire n_0_2_1548;
   wire n_0_2_1549;
   wire n_0_2_1550;
   wire n_0_2_1551;
   wire n_0_2_1552;
   wire n_0_2_1553;
   wire n_0_2_1554;
   wire n_0_2_1555;
   wire n_0_2_1556;
   wire n_0_2_1557;
   wire n_0_2_1558;
   wire n_0_2_1559;
   wire n_0_2_1560;
   wire n_0_2_1561;
   wire n_0_2_1562;
   wire n_0_2_1563;
   wire n_0_2_1564;
   wire n_0_2_1565;
   wire n_0_2_1566;
   wire n_0_2_1567;
   wire n_0_2_1568;
   wire n_0_2_1569;
   wire n_0_2_1570;
   wire n_0_2_1571;
   wire n_0_2_1572;
   wire n_0_2_1573;
   wire n_0_2_1574;
   wire n_0_2_1575;
   wire n_0_2_1576;
   wire n_0_2_1577;
   wire n_0_2_1578;
   wire n_0_2_1579;
   wire n_0_2_1580;
   wire n_0_2_1581;
   wire n_0_2_1582;
   wire n_0_2_1583;
   wire n_0_2_1584;
   wire n_0_2_1585;
   wire n_0_2_1586;
   wire n_0_2_1587;
   wire n_0_2_1588;
   wire n_0_2_1589;
   wire n_0_2_1590;
   wire n_0_2_1591;
   wire n_0_2_1592;
   wire n_0_2_1593;
   wire n_0_2_1594;
   wire n_0_2_1595;
   wire n_0_2_1596;
   wire n_0_2_1597;
   wire n_0_2_1598;
   wire n_0_2_1599;
   wire n_0_51;
   wire n_0_3_0;
   wire n_0_52;
   wire n_0_3_1;
   wire n_0_53;
   wire n_0_3_2;
   wire n_0_54;
   wire n_0_3_3;
   wire n_0_55;
   wire n_0_3_4;
   wire n_0_56;
   wire n_0_3_5;
   wire n_0_57;
   wire n_0_3_6;
   wire n_0_58;
   wire n_0_3_7;
   wire n_0_3_8;
   wire n_0_3_9;
   wire n_0_59;
   wire n_0_3_10;
   wire n_0_60;
   wire n_0_3_11;
   wire n_0_3_12;
   wire n_0_61;
   wire n_0_3_13;
   wire n_0_62;
   wire n_0_3_14;
   wire n_0_63;
   wire n_0_3_15;
   wire n_0_64;
   wire n_0_3_16;
   wire n_0_3_17;
   wire n_0_3_18;
   wire n_0_65;
   wire n_0_66;
   wire n_0_3_19;
   wire n_0_3_20;
   wire n_0_67;
   wire n_0_3_21;
   wire n_0_3_22;
   wire n_0_3_23;
   wire n_0_3_24;
   wire n_0_3_25;
   wire n_0_3_26;
   wire n_0_4_0;
   wire n_0_4_1;
   wire n_0_4_2;
   wire n_0_4_3;
   wire n_0_4_4;
   wire n_0_4_5;
   wire n_0_4_6;
   wire n_0_4_7;
   wire n_0_4_8;
   wire n_0_4_9;
   wire n_0_4_10;
   wire n_0_4_11;
   wire n_0_4_12;
   wire n_0_4_13;
   wire n_0_4_14;
   wire n_0_4_15;
   wire n_0_4_16;
   wire n_0_4_17;
   wire n_0_4_18;
   wire n_0_4_19;
   wire n_0_4_20;
   wire n_0_4_21;
   wire n_0_4_22;
   wire n_0_4_23;
   wire n_0_4_24;
   wire n_0_4_25;
   wire n_0_4_26;
   wire n_0_4_27;
   wire n_0_4_28;
   wire n_0_4_29;
   wire n_0_4_30;
   wire n_0_4_31;
   wire n_0_4_32;
   wire n_0_4_33;
   wire n_0_4_34;
   wire n_0_4_35;
   wire n_0_4_36;
   wire n_0_4_37;
   wire n_0_4_38;
   wire n_0_4_39;
   wire n_0_4_40;
   wire n_0_4_41;
   wire n_0_4_42;
   wire n_0_4_43;
   wire n_0_4_44;
   wire n_0_4_45;
   wire n_0_4_46;
   wire n_0_4_47;
   wire n_0_4_48;
   wire n_0_4_49;
   wire n_0_4_50;
   wire n_0_4_51;
   wire n_0_4_52;
   wire n_0_4_53;
   wire n_0_4_54;
   wire n_0_4_55;
   wire n_0_4_56;
   wire n_0_4_57;
   wire n_0_4_58;
   wire n_0_4_59;
   wire n_0_4_60;
   wire n_0_4_61;
   wire n_0_4_62;
   wire n_0_4_63;
   wire n_0_4_64;
   wire n_0_4_65;
   wire n_0_4_66;
   wire n_0_4_67;
   wire n_0_4_68;
   wire n_0_4_69;
   wire n_0_4_70;
   wire n_0_4_71;
   wire n_0_4_72;
   wire n_0_4_73;
   wire n_0_4_74;
   wire n_0_4_75;
   wire n_0_4_76;
   wire n_0_4_77;
   wire n_0_4_78;
   wire n_0_4_79;
   wire n_0_4_80;
   wire n_0_4_81;
   wire n_0_4_82;
   wire n_0_4_83;
   wire n_0_4_84;
   wire n_0_4_85;
   wire n_0_4_86;
   wire n_0_4_87;
   wire n_0_4_88;
   wire n_0_4_89;
   wire n_0_4_90;
   wire n_0_4_91;
   wire n_0_4_92;
   wire n_0_4_93;
   wire n_0_4_94;
   wire n_0_4_95;
   wire n_0_4_96;
   wire n_0_4_97;
   wire n_0_4_98;
   wire n_0_4_99;
   wire n_0_4_100;
   wire n_0_4_101;
   wire n_0_4_102;
   wire n_0_4_103;
   wire n_0_4_104;
   wire n_0_4_105;
   wire n_0_4_106;
   wire n_0_4_107;
   wire n_0_4_108;
   wire n_0_4_109;
   wire n_0_4_110;
   wire n_0_4_111;
   wire n_0_4_112;
   wire n_0_4_113;
   wire n_0_4_114;
   wire n_0_4_115;
   wire n_0_4_116;
   wire n_0_4_117;
   wire n_0_4_118;
   wire n_0_4_119;
   wire n_0_4_120;
   wire n_0_4_121;
   wire n_0_4_122;
   wire n_0_4_123;
   wire n_0_4_124;
   wire n_0_4_125;
   wire n_0_4_126;
   wire n_0_4_127;
   wire n_0_4_128;
   wire n_0_4_129;
   wire n_0_4_130;
   wire n_0_4_131;
   wire n_0_4_132;
   wire n_0_4_133;
   wire n_0_4_134;
   wire n_0_4_135;
   wire n_0_4_136;
   wire n_0_4_137;
   wire n_0_4_138;
   wire n_0_4_139;
   wire n_0_4_140;
   wire n_0_4_141;
   wire n_0_4_142;
   wire n_0_4_143;
   wire n_0_4_144;
   wire n_0_4_145;
   wire n_0_4_146;
   wire n_0_4_147;
   wire n_0_4_148;
   wire n_0_4_149;
   wire n_0_4_150;
   wire n_0_4_151;
   wire n_0_4_152;
   wire n_0_4_153;
   wire n_0_4_154;
   wire n_0_4_155;
   wire n_0_4_156;
   wire n_0_4_157;
   wire n_0_4_158;
   wire n_0_4_159;
   wire n_0_4_160;
   wire n_0_4_161;
   wire n_0_4_162;
   wire n_0_4_163;
   wire n_0_4_164;
   wire n_0_4_165;
   wire n_0_4_166;
   wire n_0_4_167;
   wire n_0_4_168;
   wire n_0_4_169;
   wire n_0_4_170;
   wire n_0_4_171;
   wire n_0_4_172;
   wire n_0_4_173;
   wire n_0_4_174;
   wire n_0_4_175;
   wire n_0_4_176;
   wire n_0_4_177;
   wire n_0_4_178;
   wire n_0_4_179;
   wire n_0_4_180;
   wire n_0_4_181;
   wire n_0_4_182;
   wire n_0_4_183;
   wire n_0_4_184;
   wire n_0_4_185;
   wire n_0_4_186;
   wire n_0_4_187;
   wire n_0_4_188;
   wire n_0_4_189;
   wire n_0_4_190;
   wire n_0_4_191;
   wire n_0_4_192;
   wire n_0_4_193;
   wire n_0_4_194;
   wire n_0_4_195;
   wire n_0_4_196;
   wire n_0_4_197;
   wire n_0_4_198;
   wire n_0_4_199;
   wire n_0_4_200;
   wire n_0_4_201;
   wire n_0_4_202;
   wire n_0_4_203;
   wire n_0_4_204;
   wire n_0_4_205;
   wire n_0_4_206;
   wire n_0_4_207;
   wire n_0_4_208;
   wire n_0_4_209;
   wire n_0_4_210;
   wire n_0_4_211;
   wire n_0_4_212;
   wire n_0_4_213;
   wire n_0_4_214;
   wire n_0_4_215;
   wire n_0_4_216;
   wire n_0_4_217;
   wire n_0_4_218;
   wire n_0_4_219;
   wire n_0_4_220;
   wire n_0_4_221;
   wire n_0_4_222;
   wire n_0_4_223;
   wire n_0_4_224;
   wire n_0_4_225;
   wire n_0_4_226;
   wire n_0_4_227;
   wire n_0_4_228;
   wire n_0_4_229;
   wire n_0_4_230;
   wire n_0_4_231;
   wire n_0_4_232;
   wire n_0_4_233;
   wire n_0_4_234;
   wire n_0_4_235;
   wire n_0_4_236;
   wire n_0_4_237;
   wire n_0_4_238;
   wire n_0_4_239;
   wire n_0_4_240;
   wire n_0_4_241;
   wire n_0_4_242;
   wire n_0_4_243;
   wire n_0_4_244;
   wire n_0_4_245;
   wire n_0_4_246;
   wire n_0_4_247;
   wire n_0_4_248;
   wire n_0_4_249;
   wire n_0_4_250;
   wire n_0_4_251;
   wire n_0_4_252;
   wire n_0_4_253;
   wire n_0_4_254;
   wire n_0_4_255;
   wire n_0_4_256;
   wire n_0_4_257;
   wire n_0_4_258;
   wire n_0_4_259;
   wire n_0_4_260;
   wire n_0_4_261;
   wire n_0_4_262;
   wire n_0_4_263;
   wire n_0_4_264;
   wire n_0_4_265;
   wire n_0_4_266;
   wire n_0_4_267;
   wire n_0_4_268;
   wire n_0_4_269;
   wire n_0_4_270;
   wire n_0_4_271;
   wire n_0_4_272;
   wire n_0_4_273;
   wire n_0_4_274;
   wire n_0_4_275;
   wire n_0_4_276;
   wire n_0_4_277;
   wire n_0_4_278;
   wire n_0_4_279;
   wire n_0_4_280;
   wire n_0_4_281;
   wire n_0_4_282;
   wire n_0_4_283;
   wire n_0_4_284;
   wire n_0_4_285;
   wire n_0_4_286;
   wire n_0_4_287;
   wire n_0_4_288;
   wire n_0_4_289;
   wire n_0_4_290;
   wire n_0_4_291;
   wire n_0_4_292;
   wire n_0_4_293;
   wire n_0_4_294;
   wire n_0_4_295;
   wire n_0_4_296;
   wire n_0_4_297;
   wire n_0_4_298;
   wire n_0_4_299;
   wire n_0_4_300;
   wire n_0_4_301;
   wire n_0_4_302;
   wire n_0_4_303;
   wire n_0_4_304;
   wire n_0_4_305;
   wire n_0_4_306;
   wire n_0_4_307;
   wire n_0_4_308;
   wire n_0_4_309;
   wire n_0_4_310;
   wire n_0_4_311;
   wire n_0_4_312;
   wire n_0_4_313;
   wire n_0_4_314;
   wire n_0_4_315;
   wire n_0_4_316;
   wire n_0_4_317;
   wire n_0_4_318;
   wire n_0_4_319;
   wire n_0_4_320;
   wire n_0_4_321;
   wire n_0_4_322;
   wire n_0_4_323;
   wire n_0_4_324;
   wire n_0_4_325;
   wire n_0_4_326;
   wire n_0_4_327;
   wire n_0_4_328;
   wire n_0_4_329;
   wire n_0_4_330;
   wire n_0_4_331;
   wire n_0_4_332;
   wire n_0_4_333;
   wire n_0_4_334;
   wire n_0_4_335;
   wire n_0_4_336;
   wire n_0_4_337;
   wire n_0_4_338;
   wire n_0_4_339;
   wire n_0_4_340;
   wire n_0_4_341;
   wire n_0_4_342;
   wire n_0_4_343;
   wire n_0_4_344;
   wire n_0_4_345;
   wire n_0_4_346;
   wire n_0_4_347;
   wire n_0_4_348;
   wire n_0_4_349;
   wire n_0_4_350;
   wire n_0_4_351;
   wire n_0_4_352;
   wire n_0_4_353;
   wire n_0_4_354;
   wire n_0_4_355;
   wire n_0_4_356;
   wire n_0_4_357;
   wire n_0_4_358;
   wire n_0_4_359;
   wire n_0_4_360;
   wire n_0_4_361;
   wire n_0_4_362;
   wire n_0_4_363;
   wire n_0_4_364;
   wire n_0_4_365;
   wire n_0_4_366;
   wire n_0_4_367;
   wire n_0_4_368;
   wire n_0_4_369;
   wire n_0_4_370;
   wire n_0_4_371;
   wire n_0_4_372;
   wire n_0_4_373;
   wire n_0_4_374;
   wire n_0_4_375;
   wire n_0_4_376;
   wire n_0_4_377;
   wire n_0_4_378;
   wire n_0_4_379;
   wire n_0_4_380;
   wire n_0_4_381;
   wire n_0_4_382;
   wire n_0_4_383;
   wire n_0_4_384;
   wire n_0_4_385;
   wire n_0_4_386;
   wire n_0_4_387;
   wire n_0_4_388;
   wire n_0_4_389;
   wire n_0_4_390;
   wire n_0_4_391;
   wire n_0_4_392;
   wire n_0_4_393;
   wire n_0_4_394;
   wire n_0_4_395;
   wire n_0_4_396;
   wire n_0_4_397;
   wire n_0_4_398;
   wire n_0_4_399;
   wire n_0_4_400;
   wire n_0_4_401;
   wire n_0_4_402;
   wire n_0_4_403;
   wire n_0_4_404;
   wire n_0_4_405;
   wire n_0_4_406;
   wire n_0_4_407;
   wire n_0_4_408;
   wire n_0_4_409;
   wire n_0_4_410;
   wire n_0_4_411;
   wire n_0_4_412;
   wire n_0_4_413;
   wire n_0_4_414;
   wire n_0_4_415;
   wire n_0_4_416;
   wire n_0_4_417;
   wire n_0_4_418;
   wire n_0_4_419;
   wire n_0_4_420;
   wire n_0_4_421;
   wire n_0_4_422;
   wire n_0_4_423;
   wire n_0_4_424;
   wire n_0_4_425;
   wire n_0_4_426;
   wire n_0_4_427;
   wire n_0_4_428;
   wire n_0_4_429;
   wire n_0_4_430;
   wire n_0_4_431;
   wire n_0_4_432;
   wire n_0_4_433;
   wire n_0_4_434;
   wire n_0_4_435;
   wire n_0_4_436;
   wire n_0_4_437;
   wire n_0_4_438;
   wire n_0_4_439;
   wire n_0_4_440;
   wire n_0_4_441;
   wire n_0_4_442;
   wire n_0_4_443;
   wire n_0_4_444;
   wire n_0_4_445;
   wire n_0_4_446;
   wire n_0_4_447;
   wire n_0_4_448;
   wire n_0_4_449;
   wire n_0_4_450;
   wire n_0_4_451;
   wire n_0_4_452;
   wire n_0_4_453;
   wire n_0_4_454;
   wire n_0_4_455;
   wire n_0_4_456;
   wire n_0_4_457;
   wire n_0_4_458;
   wire n_0_4_459;
   wire n_0_4_460;
   wire n_0_4_461;
   wire n_0_4_462;
   wire n_0_4_463;
   wire n_0_4_464;
   wire n_0_4_465;
   wire n_0_4_466;
   wire n_0_4_467;
   wire n_0_4_468;
   wire n_0_4_469;
   wire n_0_4_470;
   wire n_0_4_471;
   wire n_0_4_472;
   wire n_0_4_473;
   wire n_0_4_474;
   wire n_0_4_475;
   wire n_0_4_476;
   wire n_0_4_477;
   wire n_0_4_478;
   wire n_0_4_479;
   wire n_0_4_480;
   wire n_0_4_481;
   wire n_0_4_482;
   wire n_0_4_483;
   wire n_0_4_484;
   wire n_0_4_485;
   wire n_0_4_486;
   wire n_0_4_487;
   wire n_0_4_488;
   wire n_0_4_489;
   wire n_0_4_490;
   wire n_0_4_491;
   wire n_0_4_492;
   wire n_0_4_493;
   wire n_0_4_494;
   wire n_0_4_495;
   wire n_0_4_496;
   wire n_0_4_497;
   wire n_0_4_498;
   wire n_0_4_499;
   wire n_0_4_500;
   wire n_0_4_501;
   wire n_0_4_502;
   wire n_0_4_503;
   wire n_0_4_504;
   wire n_0_4_505;
   wire n_0_4_506;
   wire n_0_4_507;
   wire n_0_4_508;
   wire n_0_4_509;
   wire n_0_4_510;
   wire n_0_4_511;
   wire n_0_4_512;
   wire n_0_4_513;
   wire n_0_4_514;
   wire n_0_4_515;
   wire n_0_4_516;
   wire n_0_4_517;
   wire n_0_4_518;
   wire n_0_4_519;
   wire n_0_4_520;
   wire n_0_4_521;
   wire n_0_4_522;
   wire n_0_4_523;
   wire n_0_4_524;
   wire n_0_4_525;
   wire n_0_4_526;
   wire n_0_4_527;
   wire n_0_4_528;
   wire n_0_4_529;
   wire n_0_4_530;
   wire n_0_4_531;
   wire n_0_4_532;
   wire n_0_4_533;
   wire n_0_4_534;
   wire n_0_4_535;
   wire n_0_4_536;
   wire n_0_4_537;
   wire n_0_4_538;
   wire n_0_4_539;
   wire n_0_4_540;
   wire n_0_4_541;
   wire n_0_4_542;
   wire n_0_4_543;
   wire n_0_4_544;
   wire n_0_4_545;
   wire n_0_4_546;
   wire n_0_4_547;
   wire n_0_4_548;
   wire n_0_4_549;
   wire n_0_4_550;
   wire n_0_4_551;
   wire n_0_4_552;
   wire n_0_4_553;
   wire n_0_4_554;
   wire n_0_4_555;
   wire n_0_4_556;
   wire n_0_4_557;
   wire n_0_4_558;
   wire n_0_4_559;
   wire n_0_4_560;
   wire n_0_4_561;
   wire n_0_4_562;
   wire n_0_4_563;
   wire n_0_4_564;
   wire n_0_4_565;
   wire n_0_4_566;
   wire n_0_4_567;
   wire n_0_4_568;
   wire n_0_4_569;
   wire n_0_4_570;
   wire n_0_4_571;
   wire n_0_4_572;
   wire n_0_4_573;
   wire n_0_4_574;
   wire n_0_4_575;
   wire n_0_4_576;
   wire n_0_4_577;
   wire n_0_4_578;
   wire n_0_4_579;
   wire n_0_4_580;
   wire n_0_4_581;
   wire n_0_4_582;
   wire n_0_4_583;
   wire n_0_4_584;
   wire n_0_4_585;
   wire n_0_4_586;
   wire n_0_4_587;
   wire n_0_4_588;
   wire n_0_4_589;
   wire n_0_4_590;
   wire n_0_4_591;
   wire n_0_4_592;
   wire n_0_4_593;
   wire n_0_4_594;
   wire n_0_4_595;
   wire n_0_4_596;
   wire n_0_4_597;
   wire n_0_4_598;
   wire n_0_4_599;
   wire n_0_4_600;
   wire n_0_4_601;
   wire n_0_4_602;
   wire n_0_4_603;
   wire n_0_4_604;
   wire n_0_4_605;
   wire n_0_4_606;
   wire n_0_4_607;
   wire n_0_4_608;
   wire n_0_4_609;
   wire n_0_4_610;
   wire n_0_4_611;
   wire n_0_4_612;
   wire n_0_4_613;
   wire n_0_4_614;
   wire n_0_4_615;
   wire n_0_4_616;
   wire n_0_4_617;
   wire n_0_4_618;
   wire n_0_4_619;
   wire n_0_4_620;
   wire n_0_4_621;
   wire n_0_4_622;
   wire n_0_4_623;
   wire n_0_4_624;
   wire n_0_4_625;
   wire n_0_4_626;
   wire n_0_4_627;
   wire n_0_4_628;
   wire n_0_4_629;
   wire n_0_4_630;
   wire n_0_4_631;
   wire n_0_4_632;
   wire n_0_4_633;
   wire n_0_4_634;
   wire n_0_4_635;
   wire n_0_4_636;
   wire n_0_4_637;
   wire n_0_4_638;
   wire n_0_4_639;
   wire n_0_4_640;
   wire n_0_4_641;
   wire n_0_4_642;
   wire n_0_4_643;
   wire n_0_4_644;
   wire n_0_4_645;
   wire n_0_4_646;
   wire n_0_4_647;
   wire n_0_4_648;
   wire n_0_4_649;
   wire n_0_4_650;
   wire n_0_4_651;
   wire n_0_4_652;
   wire n_0_4_653;
   wire n_0_4_654;
   wire n_0_4_655;
   wire n_0_4_656;
   wire n_0_4_657;
   wire n_0_4_658;
   wire n_0_4_659;
   wire n_0_4_660;
   wire n_0_4_661;
   wire n_0_4_662;
   wire n_0_4_663;
   wire n_0_4_664;
   wire n_0_4_665;
   wire n_0_4_666;
   wire n_0_4_667;
   wire n_0_4_668;
   wire n_0_4_669;
   wire n_0_4_670;
   wire n_0_4_671;
   wire n_0_4_672;
   wire n_0_4_673;
   wire n_0_4_674;
   wire n_0_4_675;
   wire n_0_4_676;
   wire n_0_4_677;
   wire n_0_4_678;
   wire n_0_4_679;
   wire n_0_4_680;
   wire n_0_4_681;
   wire n_0_4_682;
   wire n_0_4_683;
   wire n_0_4_684;
   wire n_0_4_685;
   wire n_0_4_686;
   wire n_0_4_687;
   wire n_0_4_688;
   wire n_0_4_689;
   wire n_0_4_690;
   wire n_0_4_691;
   wire n_0_4_692;
   wire n_0_4_693;
   wire n_0_4_694;
   wire n_0_4_695;
   wire n_0_4_696;
   wire n_0_4_697;
   wire n_0_4_698;
   wire n_0_4_699;
   wire n_0_4_700;
   wire n_0_4_701;
   wire n_0_4_702;
   wire n_0_4_703;
   wire n_0_4_704;
   wire n_0_4_705;
   wire n_0_4_706;
   wire n_0_4_707;
   wire n_0_4_708;
   wire n_0_4_709;
   wire n_0_4_710;
   wire n_0_4_711;
   wire n_0_4_712;
   wire n_0_4_713;
   wire n_0_4_714;
   wire n_0_4_715;
   wire n_0_4_716;
   wire n_0_4_717;
   wire n_0_4_718;
   wire n_0_4_719;
   wire n_0_4_720;
   wire n_0_4_721;
   wire n_0_4_722;
   wire n_0_4_723;
   wire n_0_4_724;
   wire n_0_4_725;
   wire n_0_4_726;
   wire n_0_4_727;
   wire n_0_4_728;
   wire n_0_4_729;
   wire n_0_4_730;
   wire n_0_4_731;
   wire n_0_4_732;
   wire n_0_4_733;
   wire n_0_4_734;
   wire n_0_4_735;
   wire n_0_4_736;
   wire n_0_4_737;
   wire n_0_4_738;
   wire n_0_4_739;
   wire n_0_4_740;
   wire n_0_4_741;
   wire n_0_4_742;
   wire n_0_4_743;
   wire n_0_4_744;
   wire n_0_4_745;
   wire n_0_4_746;
   wire n_0_4_747;
   wire n_0_4_748;
   wire n_0_4_749;
   wire n_0_4_750;
   wire n_0_4_751;
   wire n_0_4_752;
   wire n_0_4_753;
   wire n_0_4_754;
   wire n_0_4_755;
   wire n_0_4_756;
   wire n_0_4_757;
   wire n_0_4_758;
   wire n_0_4_759;
   wire n_0_4_760;
   wire n_0_4_761;
   wire n_0_4_762;
   wire n_0_4_763;
   wire n_0_4_764;
   wire n_0_4_765;
   wire n_0_4_766;
   wire n_0_4_767;
   wire n_0_4_768;
   wire n_0_4_769;
   wire n_0_4_770;
   wire n_0_4_771;
   wire n_0_4_772;
   wire n_0_4_773;
   wire n_0_4_774;
   wire n_0_4_775;
   wire n_0_4_776;
   wire n_0_4_777;
   wire n_0_4_778;
   wire n_0_4_779;
   wire n_0_4_780;
   wire n_0_4_781;
   wire n_0_4_782;
   wire n_0_4_783;
   wire n_0_4_784;
   wire n_0_4_785;
   wire n_0_4_786;
   wire n_0_4_787;
   wire n_0_4_788;
   wire n_0_4_789;
   wire n_0_4_790;
   wire n_0_4_791;
   wire n_0_4_792;
   wire n_0_4_793;
   wire n_0_4_794;
   wire n_0_4_795;
   wire n_0_4_796;
   wire n_0_4_797;
   wire n_0_4_798;
   wire n_0_4_799;
   wire n_0_4_800;
   wire n_0_4_801;
   wire n_0_4_802;
   wire n_0_4_803;
   wire n_0_4_804;
   wire n_0_4_805;
   wire n_0_4_806;
   wire n_0_4_807;
   wire n_0_4_808;
   wire n_0_4_809;
   wire n_0_4_810;
   wire n_0_4_811;
   wire n_0_4_812;
   wire n_0_4_813;
   wire n_0_4_814;
   wire n_0_4_815;
   wire n_0_4_816;
   wire n_0_4_817;
   wire n_0_4_818;
   wire n_0_4_819;
   wire n_0_4_820;
   wire n_0_4_821;
   wire n_0_4_822;
   wire n_0_4_823;
   wire n_0_4_824;
   wire n_0_4_825;
   wire n_0_4_826;
   wire n_0_4_827;
   wire n_0_4_828;
   wire n_0_4_829;
   wire n_0_4_830;
   wire n_0_4_831;
   wire n_0_4_832;
   wire n_0_4_833;
   wire n_0_4_834;
   wire n_0_4_835;
   wire n_0_4_836;
   wire n_0_4_837;
   wire n_0_4_838;
   wire n_0_4_839;
   wire n_0_4_840;
   wire n_0_4_841;
   wire n_0_4_842;
   wire n_0_4_843;
   wire n_0_4_844;
   wire n_0_4_845;
   wire n_0_4_846;
   wire n_0_4_847;
   wire n_0_4_848;
   wire n_0_4_849;
   wire n_0_4_850;
   wire n_0_4_851;
   wire n_0_4_852;
   wire n_0_4_853;
   wire n_0_4_854;
   wire n_0_4_855;
   wire n_0_4_856;
   wire n_0_4_857;
   wire n_0_4_858;
   wire n_0_4_859;
   wire n_0_4_860;
   wire n_0_4_861;
   wire n_0_4_862;
   wire n_0_4_863;
   wire n_0_4_864;
   wire n_0_4_865;
   wire n_0_4_866;
   wire n_0_4_867;
   wire n_0_4_868;
   wire n_0_4_869;
   wire n_0_4_870;
   wire n_0_4_871;
   wire n_0_4_872;
   wire n_0_4_873;
   wire n_0_4_874;
   wire n_0_4_875;
   wire n_0_4_876;
   wire n_0_4_877;
   wire n_0_4_878;
   wire n_0_4_879;
   wire n_0_4_880;
   wire n_0_4_881;
   wire n_0_4_882;
   wire n_0_4_883;
   wire n_0_4_884;
   wire n_0_4_885;
   wire n_0_4_886;
   wire n_0_4_887;
   wire n_0_4_888;
   wire n_0_4_889;
   wire n_0_4_890;
   wire n_0_4_891;
   wire n_0_4_892;
   wire n_0_4_893;
   wire n_0_4_894;
   wire n_0_4_895;
   wire n_0_4_896;
   wire n_0_4_897;
   wire n_0_4_898;
   wire n_0_4_899;
   wire n_0_4_900;
   wire n_0_4_901;
   wire n_0_4_902;
   wire n_0_4_903;
   wire n_0_4_904;
   wire n_0_4_905;
   wire n_0_4_906;
   wire n_0_4_907;
   wire n_0_4_908;
   wire n_0_4_909;
   wire n_0_4_910;
   wire n_0_4_911;
   wire n_0_4_912;
   wire n_0_4_913;
   wire n_0_4_914;
   wire n_0_4_915;
   wire n_0_4_916;
   wire n_0_4_917;
   wire n_0_4_918;
   wire n_0_4_919;
   wire n_0_4_920;
   wire n_0_4_921;
   wire n_0_4_922;
   wire n_0_4_923;
   wire n_0_4_924;
   wire n_0_4_925;
   wire n_0_4_926;
   wire n_0_4_927;
   wire n_0_4_928;
   wire n_0_4_929;
   wire n_0_4_930;
   wire n_0_4_931;
   wire n_0_4_932;
   wire n_0_4_933;
   wire n_0_4_934;
   wire n_0_4_935;
   wire n_0_4_936;
   wire n_0_4_937;
   wire n_0_4_938;
   wire n_0_4_939;
   wire n_0_4_940;
   wire n_0_4_941;
   wire n_0_4_942;
   wire n_0_4_943;
   wire n_0_4_944;
   wire n_0_4_945;
   wire n_0_4_946;
   wire n_0_4_947;
   wire n_0_4_948;
   wire n_0_4_949;
   wire n_0_4_950;
   wire n_0_4_951;
   wire n_0_4_952;
   wire n_0_4_953;
   wire n_0_4_954;
   wire n_0_4_955;
   wire n_0_4_956;
   wire n_0_4_957;
   wire n_0_4_958;
   wire n_0_4_959;
   wire n_0_4_960;
   wire n_0_4_961;
   wire n_0_4_962;
   wire n_0_4_963;
   wire n_0_4_964;
   wire n_0_4_965;
   wire n_0_4_966;
   wire n_0_4_967;
   wire n_0_4_968;
   wire n_0_4_969;
   wire n_0_4_970;
   wire n_0_4_971;
   wire n_0_4_972;
   wire n_0_4_973;
   wire n_0_4_974;
   wire n_0_4_975;
   wire n_0_4_976;
   wire n_0_4_977;
   wire n_0_4_978;
   wire n_0_4_979;
   wire n_0_4_980;
   wire n_0_4_981;
   wire n_0_4_982;
   wire n_0_4_983;
   wire n_0_4_984;
   wire n_0_4_985;
   wire n_0_4_986;
   wire n_0_4_987;
   wire n_0_4_988;
   wire n_0_4_989;
   wire n_0_4_990;
   wire n_0_4_991;
   wire n_0_4_992;
   wire n_0_4_993;
   wire n_0_4_994;
   wire n_0_4_995;
   wire n_0_4_996;
   wire n_0_4_997;
   wire n_0_4_998;
   wire n_0_4_999;
   wire n_0_4_1000;
   wire n_0_4_1001;
   wire n_0_4_1002;
   wire n_0_4_1003;
   wire n_0_4_1004;
   wire n_0_4_1005;
   wire n_0_4_1006;
   wire n_0_4_1007;
   wire n_0_4_1008;
   wire n_0_4_1009;
   wire n_0_4_1010;
   wire n_0_4_1011;
   wire n_0_4_1012;
   wire n_0_4_1013;
   wire n_0_4_1014;
   wire n_0_4_1015;
   wire n_0_4_1016;
   wire n_0_4_1017;
   wire n_0_4_1018;
   wire n_0_4_1019;
   wire n_0_4_1020;
   wire n_0_4_1021;
   wire n_0_4_1022;
   wire n_0_4_1023;
   wire n_0_4_1024;
   wire n_0_4_1025;
   wire n_0_4_1026;
   wire n_0_4_1027;
   wire n_0_4_1028;
   wire n_0_4_1029;
   wire n_0_4_1030;
   wire n_0_4_1031;
   wire n_0_4_1032;
   wire n_0_4_1033;
   wire n_0_4_1034;
   wire n_0_4_1035;
   wire n_0_4_1036;
   wire n_0_4_1037;
   wire n_0_4_1038;
   wire n_0_4_1039;
   wire n_0_4_1040;
   wire n_0_4_1041;
   wire n_0_4_1042;
   wire n_0_4_1043;
   wire n_0_4_1044;
   wire n_0_4_1045;
   wire n_0_4_1046;
   wire n_0_4_1047;
   wire n_0_4_1048;
   wire n_0_4_1049;
   wire n_0_4_1050;
   wire n_0_4_1051;
   wire n_0_4_1052;
   wire n_0_4_1053;
   wire n_0_4_1054;
   wire n_0_4_1055;
   wire n_0_4_1056;
   wire n_0_4_1057;
   wire n_0_4_1058;
   wire n_0_4_1059;
   wire n_0_4_1060;
   wire n_0_4_1061;
   wire n_0_4_1062;
   wire n_0_4_1063;
   wire n_0_4_1064;
   wire n_0_4_1065;
   wire n_0_4_1066;
   wire n_0_4_1067;
   wire n_0_4_1068;
   wire n_0_4_1069;
   wire n_0_4_1070;
   wire n_0_4_1071;
   wire n_0_4_1072;
   wire n_0_4_1073;
   wire n_0_4_1074;
   wire n_0_4_1075;
   wire n_0_4_1076;
   wire n_0_4_1077;
   wire n_0_4_1078;
   wire n_0_4_1079;
   wire n_0_4_1080;
   wire n_0_4_1081;
   wire n_0_4_1082;
   wire n_0_4_1083;
   wire n_0_4_1084;
   wire n_0_4_1085;
   wire n_0_4_1086;
   wire n_0_4_1087;
   wire n_0_4_1088;
   wire n_0_4_1089;
   wire n_0_4_1090;
   wire n_0_4_1091;
   wire n_0_4_1092;
   wire n_0_4_1093;
   wire n_0_4_1094;
   wire n_0_4_1095;
   wire n_0_4_1096;
   wire n_0_4_1097;
   wire n_0_4_1098;
   wire n_0_4_1099;
   wire n_0_4_1100;
   wire n_0_4_1101;
   wire n_0_4_1102;
   wire n_0_4_1103;
   wire n_0_4_1104;
   wire n_0_4_1105;
   wire n_0_4_1106;
   wire n_0_4_1107;
   wire n_0_4_1108;
   wire n_0_4_1109;
   wire n_0_4_1110;
   wire n_0_4_1111;
   wire n_0_4_1112;
   wire n_0_4_1113;
   wire n_0_4_1114;
   wire n_0_4_1115;
   wire n_0_4_1116;
   wire n_0_4_1117;
   wire n_0_4_1118;
   wire n_0_4_1119;
   wire n_0_4_1120;
   wire n_0_4_1121;
   wire n_0_4_1122;
   wire n_0_4_1123;
   wire n_0_4_1124;
   wire n_0_4_1125;
   wire n_0_4_1126;
   wire n_0_4_1127;
   wire n_0_4_1128;
   wire n_0_4_1129;
   wire n_0_4_1130;
   wire n_0_4_1131;
   wire n_0_4_1132;
   wire n_0_4_1133;
   wire n_0_4_1134;
   wire n_0_4_1135;
   wire n_0_4_1136;
   wire n_0_4_1137;
   wire n_0_4_1138;
   wire n_0_4_1139;
   wire n_0_4_1140;
   wire n_0_4_1141;
   wire n_0_4_1142;
   wire n_0_4_1143;
   wire n_0_4_1144;
   wire n_0_4_1145;
   wire n_0_4_1146;
   wire n_0_4_1147;
   wire n_0_4_1148;
   wire n_0_4_1149;
   wire n_0_4_1150;
   wire n_0_4_1151;
   wire n_0_4_1152;
   wire n_0_4_1153;
   wire n_0_4_1154;
   wire n_0_4_1155;
   wire n_0_4_1156;
   wire n_0_4_1157;
   wire n_0_4_1158;
   wire n_0_4_1159;
   wire n_0_4_1160;
   wire n_0_4_1161;
   wire n_0_4_1162;
   wire n_0_4_1163;
   wire n_0_4_1164;
   wire n_0_4_1165;
   wire n_0_4_1166;
   wire n_0_4_1167;
   wire n_0_4_1168;
   wire n_0_4_1169;
   wire n_0_4_1170;
   wire n_0_4_1171;
   wire n_0_4_1172;
   wire n_0_4_1173;
   wire n_0_4_1174;
   wire n_0_4_1175;
   wire n_0_4_1176;
   wire n_0_4_1177;
   wire n_0_4_1178;
   wire n_0_4_1179;
   wire n_0_4_1180;
   wire n_0_4_1181;
   wire n_0_4_1182;
   wire n_0_4_1183;
   wire n_0_4_1184;
   wire n_0_4_1185;
   wire n_0_4_1186;
   wire n_0_4_1187;
   wire n_0_4_1188;
   wire n_0_4_1189;
   wire n_0_4_1190;
   wire n_0_4_1191;
   wire n_0_4_1192;
   wire n_0_4_1193;
   wire n_0_4_1194;
   wire n_0_4_1195;
   wire n_0_4_1196;
   wire n_0_4_1197;
   wire n_0_4_1198;
   wire n_0_4_1199;
   wire n_0_4_1200;
   wire n_0_4_1201;
   wire n_0_4_1202;
   wire n_0_4_1203;
   wire n_0_4_1204;
   wire n_0_4_1205;
   wire n_0_4_1206;
   wire n_0_4_1207;
   wire n_0_4_1208;
   wire n_0_4_1209;
   wire n_0_4_1210;
   wire n_0_4_1211;
   wire n_0_4_1212;
   wire n_0_4_1213;
   wire n_0_4_1214;
   wire n_0_4_1215;
   wire n_0_4_1216;
   wire n_0_4_1217;
   wire n_0_4_1218;
   wire n_0_4_1219;
   wire n_0_4_1220;
   wire n_0_4_1221;
   wire n_0_4_1222;
   wire n_0_4_1223;
   wire n_0_4_1224;
   wire n_0_4_1225;
   wire n_0_4_1226;
   wire n_0_4_1227;
   wire n_0_4_1228;
   wire n_0_4_1229;
   wire n_0_4_1230;
   wire n_0_4_1231;
   wire n_0_4_1232;
   wire n_0_4_1233;
   wire n_0_4_1234;
   wire n_0_4_1235;
   wire n_0_4_1236;
   wire n_0_4_1237;
   wire n_0_4_1238;
   wire n_0_4_1239;
   wire n_0_4_1240;
   wire n_0_4_1241;
   wire n_0_4_1242;
   wire n_0_4_1243;
   wire n_0_4_1244;
   wire n_0_4_1245;
   wire n_0_4_1246;
   wire n_0_4_1247;
   wire n_0_4_1248;
   wire n_0_4_1249;
   wire n_0_4_1250;
   wire n_0_4_1251;
   wire n_0_4_1252;
   wire n_0_4_1253;
   wire n_0_4_1254;
   wire n_0_4_1255;
   wire n_0_4_1256;
   wire n_0_4_1257;
   wire n_0_4_1258;
   wire n_0_4_1259;
   wire n_0_4_1260;
   wire n_0_4_1261;
   wire n_0_4_1262;
   wire n_0_4_1263;
   wire n_0_4_1264;
   wire n_0_4_1265;
   wire n_0_4_1266;
   wire n_0_4_1267;
   wire n_0_4_1268;
   wire n_0_4_1269;
   wire n_0_4_1270;
   wire n_0_4_1271;
   wire n_0_4_1272;
   wire n_0_4_1273;
   wire n_0_4_1274;
   wire n_0_4_1275;
   wire n_0_4_1276;
   wire n_0_4_1277;
   wire n_0_4_1278;
   wire n_0_4_1279;
   wire n_0_4_1280;
   wire n_0_4_1281;
   wire n_0_4_1282;
   wire n_0_4_1283;
   wire n_0_4_1284;
   wire n_0_4_1285;
   wire n_0_4_1286;
   wire n_0_4_1287;
   wire n_0_4_1288;
   wire n_0_4_1289;
   wire n_0_4_1290;
   wire n_0_4_1291;
   wire n_0_4_1292;
   wire n_0_4_1293;
   wire n_0_4_1294;
   wire n_0_4_1295;
   wire n_0_4_1296;
   wire n_0_4_1297;
   wire n_0_4_1298;
   wire n_0_4_1299;
   wire n_0_4_1300;
   wire n_0_4_1301;
   wire n_0_4_1302;
   wire n_0_4_1303;
   wire n_0_4_1304;
   wire n_0_4_1305;
   wire n_0_4_1306;
   wire n_0_4_1307;
   wire n_0_4_1308;
   wire n_0_4_1309;
   wire n_0_4_1310;
   wire n_0_4_1311;
   wire n_0_4_1312;
   wire n_0_4_1313;
   wire n_0_4_1314;
   wire n_0_4_1315;
   wire n_0_4_1316;
   wire n_0_4_1317;
   wire n_0_4_1318;
   wire n_0_4_1319;
   wire n_0_4_1320;
   wire n_0_4_1321;
   wire n_0_4_1322;
   wire n_0_4_1323;
   wire n_0_4_1324;
   wire n_0_4_1325;
   wire n_0_4_1326;
   wire n_0_4_1327;
   wire n_0_4_1328;
   wire n_0_4_1329;
   wire n_0_4_1330;
   wire n_0_4_1331;
   wire n_0_4_1332;
   wire n_0_4_1333;
   wire n_0_4_1334;
   wire n_0_4_1335;
   wire n_0_4_1336;
   wire n_0_4_1337;
   wire n_0_4_1338;
   wire n_0_4_1339;
   wire n_0_4_1340;
   wire n_0_4_1341;
   wire n_0_4_1342;
   wire n_0_4_1343;
   wire n_0_4_1344;
   wire n_0_4_1345;
   wire n_0_4_1346;
   wire n_0_4_1347;
   wire n_0_4_1348;
   wire n_0_4_1349;
   wire n_0_4_1350;
   wire n_0_4_1351;
   wire n_0_4_1352;
   wire n_0_4_1353;
   wire n_0_4_1354;
   wire n_0_4_1355;
   wire n_0_4_1356;
   wire n_0_4_1357;
   wire n_0_4_1358;
   wire n_0_4_1359;
   wire n_0_4_1360;
   wire n_0_4_1361;
   wire n_0_4_1362;
   wire n_0_4_1363;
   wire n_0_4_1364;
   wire n_0_4_1365;
   wire n_0_4_1366;
   wire n_0_4_1367;
   wire n_0_4_1368;
   wire n_0_4_1369;
   wire n_0_4_1370;
   wire n_0_4_1371;
   wire n_0_4_1372;
   wire n_0_4_1373;
   wire n_0_4_1374;
   wire n_0_4_1375;
   wire n_0_4_1376;
   wire n_0_4_1377;
   wire n_0_4_1378;
   wire n_0_4_1379;
   wire n_0_4_1380;
   wire n_0_4_1381;
   wire n_0_4_1382;
   wire n_0_4_1383;
   wire n_0_4_1384;
   wire n_0_4_1385;
   wire n_0_4_1386;
   wire n_0_4_1387;
   wire n_0_4_1388;
   wire n_0_4_1389;
   wire n_0_4_1390;
   wire n_0_4_1391;
   wire n_0_4_1392;
   wire n_0_4_1393;
   wire n_0_4_1394;
   wire n_0_4_1395;
   wire n_0_4_1396;
   wire n_0_4_1397;
   wire n_0_4_1398;
   wire n_0_4_1399;
   wire n_0_4_1400;
   wire n_0_4_1401;
   wire n_0_4_1402;
   wire n_0_4_1403;
   wire n_0_4_1404;
   wire n_0_4_1405;
   wire n_0_4_1406;
   wire n_0_4_1407;
   wire n_0_4_1408;
   wire n_0_4_1409;
   wire n_0_4_1410;
   wire n_0_4_1411;
   wire n_0_4_1412;
   wire n_0_4_1413;
   wire n_0_4_1414;
   wire n_0_4_1415;
   wire n_0_4_1416;
   wire n_0_4_1417;
   wire n_0_4_1418;
   wire n_0_4_1419;
   wire n_0_4_1420;
   wire n_0_4_1421;
   wire n_0_4_1422;
   wire n_0_4_1423;
   wire n_0_4_1424;
   wire n_0_4_1425;
   wire n_0_4_1426;
   wire n_0_4_1427;
   wire n_0_4_1428;
   wire n_0_4_1429;
   wire n_0_4_1430;
   wire n_0_4_1431;
   wire n_0_4_1432;
   wire n_0_4_1433;
   wire n_0_4_1434;
   wire n_0_4_1435;
   wire n_0_4_1436;
   wire n_0_4_1437;
   wire n_0_4_1438;
   wire n_0_4_1439;
   wire n_0_4_1440;
   wire n_0_4_1441;
   wire n_0_4_1442;
   wire n_0_4_1443;
   wire n_0_4_1444;
   wire n_0_4_1445;
   wire n_0_4_1446;
   wire n_0_4_1447;
   wire n_0_4_1448;
   wire n_0_4_1449;
   wire n_0_4_1450;
   wire n_0_4_1451;
   wire n_0_4_1452;
   wire n_0_4_1453;
   wire n_0_4_1454;
   wire n_0_4_1455;
   wire n_0_4_1456;
   wire n_0_4_1457;
   wire n_0_4_1458;
   wire n_0_4_1459;
   wire n_0_4_1460;
   wire n_0_4_1461;
   wire n_0_4_1462;
   wire n_0_4_1463;
   wire n_0_4_1464;
   wire n_0_4_1465;
   wire n_0_4_1466;
   wire n_0_4_1467;
   wire n_0_4_1468;
   wire n_0_4_1469;
   wire n_0_4_1470;
   wire n_0_4_1471;
   wire n_0_4_1472;
   wire n_0_4_1473;
   wire n_0_4_1474;
   wire n_0_4_1475;
   wire n_0_4_1476;
   wire n_0_4_1477;
   wire n_0_4_1478;
   wire n_0_4_1479;
   wire n_0_4_1480;
   wire n_0_4_1481;
   wire n_0_4_1482;
   wire n_0_4_1483;
   wire n_0_4_1484;
   wire n_0_4_1485;
   wire n_0_4_1486;
   wire n_0_4_1487;
   wire n_0_4_1488;
   wire n_0_4_1489;
   wire n_0_4_1490;
   wire n_0_4_1491;
   wire n_0_4_1492;
   wire n_0_4_1493;
   wire n_0_4_1494;
   wire n_0_4_1495;
   wire n_0_4_1496;
   wire n_0_4_1497;
   wire n_0_4_1498;
   wire n_0_4_1499;
   wire n_0_4_1500;
   wire n_0_4_1501;
   wire n_0_4_1502;
   wire n_0_4_1503;
   wire n_0_4_1504;
   wire n_0_4_1505;
   wire n_0_4_1506;
   wire n_0_4_1507;
   wire n_0_4_1508;
   wire n_0_4_1509;
   wire n_0_4_1510;
   wire n_0_4_1511;
   wire n_0_4_1512;
   wire n_0_4_1513;
   wire n_0_4_1514;
   wire n_0_4_1515;
   wire n_0_4_1516;
   wire n_0_4_1517;
   wire n_0_4_1518;
   wire n_0_4_1519;
   wire n_0_4_1520;
   wire n_0_4_1521;
   wire n_0_4_1522;
   wire n_0_4_1523;
   wire n_0_4_1524;
   wire n_0_4_1525;
   wire n_0_4_1526;
   wire n_0_4_1527;
   wire n_0_4_1528;
   wire n_0_4_1529;
   wire n_0_4_1530;
   wire n_0_4_1531;
   wire n_0_4_1532;
   wire n_0_4_1533;
   wire n_0_4_1534;
   wire n_0_4_1535;
   wire n_0_4_1536;
   wire n_0_4_1537;
   wire n_0_4_1538;
   wire n_0_4_1539;
   wire n_0_4_1540;
   wire n_0_4_1541;
   wire n_0_4_1542;
   wire n_0_4_1543;
   wire n_0_4_1544;
   wire n_0_4_1545;
   wire n_0_4_1546;
   wire n_0_4_1547;
   wire n_0_4_1548;
   wire n_0_4_1549;
   wire n_0_4_1550;
   wire n_0_4_1551;
   wire n_0_4_1552;
   wire n_0_4_1553;
   wire n_0_4_1554;
   wire n_0_4_1555;
   wire n_0_4_1556;
   wire n_0_4_1557;
   wire n_0_4_1558;
   wire n_0_4_1559;
   wire n_0_4_1560;
   wire n_0_4_1561;
   wire n_0_4_1562;
   wire n_0_4_1563;
   wire n_0_4_1564;
   wire n_0_4_1565;
   wire n_0_4_1566;
   wire n_0_4_1567;
   wire n_0_4_1568;
   wire n_0_4_1569;
   wire n_0_4_1570;
   wire n_0_4_1571;
   wire n_0_4_1572;
   wire n_0_4_1573;
   wire n_0_4_1574;
   wire n_0_4_1575;
   wire n_0_4_1576;
   wire n_0_4_1577;
   wire n_0_4_1578;
   wire n_0_4_1579;
   wire n_0_4_1580;
   wire n_0_4_1581;
   wire n_0_4_1582;
   wire n_0_4_1583;
   wire n_0_4_1584;
   wire n_0_4_1585;
   wire n_0_4_1586;
   wire n_0_4_1587;
   wire n_0_4_1588;
   wire n_0_4_1589;
   wire n_0_4_1590;
   wire n_0_4_1591;
   wire n_0_4_1592;
   wire n_0_4_1593;
   wire n_0_4_1594;
   wire n_0_4_1595;
   wire n_0_4_1596;
   wire n_0_4_1597;
   wire n_0_4_1598;
   wire n_0_4_1599;
   wire [63:0]Memory;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_1_0;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_1_1;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_1_2;
   wire n_0_1_3;
   wire n_0_29;
   wire n_0_30;
   wire n_0_1_4;
   wire n_0_31;
   wire n_0_1_5;
   wire n_0_32;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_1_8;
   wire n_0_1_9;
   wire n_0_33;
   wire n_0_1_10;
   wire n_0_1_11;
   wire n_0_1_12;
   wire n_0_1_13;
   wire n_0_1_14;
   wire n_0_1_15;
   wire n_0_1_16;
   wire n_0_1_17;
   wire n_0_1_18;
   wire n_0_1_19;
   wire n_0_1_20;
   wire n_0_1_21;

   CLKGATETST_X1 \clk_gate_Memory_reg[16]_reg  (.CK(CLK), .E(n_0_33), .SE(1'b0), 
      .GCK(n_0_0));
   DFF_X1 \Memory_reg[16][63]  (.D(dataIn[63]), .CK(n_0_0), .Q(\Memory[16] [63]), 
      .QN());
   DFF_X1 \Memory_reg[16][62]  (.D(dataIn[62]), .CK(n_0_0), .Q(\Memory[16] [62]), 
      .QN());
   DFF_X1 \Memory_reg[16][61]  (.D(dataIn[61]), .CK(n_0_0), .Q(\Memory[16] [61]), 
      .QN());
   DFF_X1 \Memory_reg[16][60]  (.D(dataIn[60]), .CK(n_0_0), .Q(\Memory[16] [60]), 
      .QN());
   DFF_X1 \Memory_reg[16][59]  (.D(dataIn[59]), .CK(n_0_0), .Q(\Memory[16] [59]), 
      .QN());
   DFF_X1 \Memory_reg[16][58]  (.D(dataIn[58]), .CK(n_0_0), .Q(\Memory[16] [58]), 
      .QN());
   DFF_X1 \Memory_reg[16][57]  (.D(dataIn[57]), .CK(n_0_0), .Q(\Memory[16] [57]), 
      .QN());
   DFF_X1 \Memory_reg[16][56]  (.D(dataIn[56]), .CK(n_0_0), .Q(\Memory[16] [56]), 
      .QN());
   DFF_X1 \Memory_reg[16][55]  (.D(dataIn[55]), .CK(n_0_0), .Q(\Memory[16] [55]), 
      .QN());
   DFF_X1 \Memory_reg[16][54]  (.D(dataIn[54]), .CK(n_0_0), .Q(\Memory[16] [54]), 
      .QN());
   DFF_X1 \Memory_reg[16][53]  (.D(dataIn[53]), .CK(n_0_0), .Q(\Memory[16] [53]), 
      .QN());
   DFF_X1 \Memory_reg[16][52]  (.D(dataIn[52]), .CK(n_0_0), .Q(\Memory[16] [52]), 
      .QN());
   DFF_X1 \Memory_reg[16][51]  (.D(dataIn[51]), .CK(n_0_0), .Q(\Memory[16] [51]), 
      .QN());
   DFF_X1 \Memory_reg[16][50]  (.D(dataIn[50]), .CK(n_0_0), .Q(\Memory[16] [50]), 
      .QN());
   DFF_X1 \Memory_reg[16][49]  (.D(dataIn[49]), .CK(n_0_0), .Q(\Memory[16] [49]), 
      .QN());
   DFF_X1 \Memory_reg[16][48]  (.D(dataIn[48]), .CK(n_0_0), .Q(\Memory[16] [48]), 
      .QN());
   DFF_X1 \Memory_reg[16][47]  (.D(dataIn[47]), .CK(n_0_0), .Q(\Memory[16] [47]), 
      .QN());
   DFF_X1 \Memory_reg[16][46]  (.D(dataIn[46]), .CK(n_0_0), .Q(\Memory[16] [46]), 
      .QN());
   DFF_X1 \Memory_reg[16][45]  (.D(dataIn[45]), .CK(n_0_0), .Q(\Memory[16] [45]), 
      .QN());
   DFF_X1 \Memory_reg[16][44]  (.D(dataIn[44]), .CK(n_0_0), .Q(\Memory[16] [44]), 
      .QN());
   DFF_X1 \Memory_reg[16][43]  (.D(dataIn[43]), .CK(n_0_0), .Q(\Memory[16] [43]), 
      .QN());
   DFF_X1 \Memory_reg[16][42]  (.D(dataIn[42]), .CK(n_0_0), .Q(\Memory[16] [42]), 
      .QN());
   DFF_X1 \Memory_reg[16][41]  (.D(dataIn[41]), .CK(n_0_0), .Q(\Memory[16] [41]), 
      .QN());
   DFF_X1 \Memory_reg[16][40]  (.D(dataIn[40]), .CK(n_0_0), .Q(\Memory[16] [40]), 
      .QN());
   DFF_X1 \Memory_reg[16][39]  (.D(dataIn[39]), .CK(n_0_0), .Q(\Memory[16] [39]), 
      .QN());
   DFF_X1 \Memory_reg[16][38]  (.D(dataIn[38]), .CK(n_0_0), .Q(\Memory[16] [38]), 
      .QN());
   DFF_X1 \Memory_reg[16][37]  (.D(dataIn[37]), .CK(n_0_0), .Q(\Memory[16] [37]), 
      .QN());
   DFF_X1 \Memory_reg[16][36]  (.D(dataIn[36]), .CK(n_0_0), .Q(\Memory[16] [36]), 
      .QN());
   DFF_X1 \Memory_reg[16][35]  (.D(dataIn[35]), .CK(n_0_0), .Q(\Memory[16] [35]), 
      .QN());
   DFF_X1 \Memory_reg[16][34]  (.D(dataIn[34]), .CK(n_0_0), .Q(\Memory[16] [34]), 
      .QN());
   DFF_X1 \Memory_reg[16][33]  (.D(dataIn[33]), .CK(n_0_0), .Q(\Memory[16] [33]), 
      .QN());
   DFF_X1 \Memory_reg[16][32]  (.D(dataIn[32]), .CK(n_0_0), .Q(\Memory[16] [32]), 
      .QN());
   DFF_X1 \Memory_reg[16][31]  (.D(dataIn[31]), .CK(n_0_0), .Q(\Memory[16] [31]), 
      .QN());
   DFF_X1 \Memory_reg[16][30]  (.D(dataIn[30]), .CK(n_0_0), .Q(\Memory[16] [30]), 
      .QN());
   DFF_X1 \Memory_reg[16][29]  (.D(dataIn[29]), .CK(n_0_0), .Q(\Memory[16] [29]), 
      .QN());
   DFF_X1 \Memory_reg[16][28]  (.D(dataIn[28]), .CK(n_0_0), .Q(\Memory[16] [28]), 
      .QN());
   DFF_X1 \Memory_reg[16][27]  (.D(dataIn[27]), .CK(n_0_0), .Q(\Memory[16] [27]), 
      .QN());
   DFF_X1 \Memory_reg[16][26]  (.D(dataIn[26]), .CK(n_0_0), .Q(\Memory[16] [26]), 
      .QN());
   DFF_X1 \Memory_reg[16][25]  (.D(dataIn[25]), .CK(n_0_0), .Q(\Memory[16] [25]), 
      .QN());
   DFF_X1 \Memory_reg[16][24]  (.D(dataIn[24]), .CK(n_0_0), .Q(\Memory[16] [24]), 
      .QN());
   DFF_X1 \Memory_reg[16][23]  (.D(dataIn[23]), .CK(n_0_0), .Q(\Memory[16] [23]), 
      .QN());
   DFF_X1 \Memory_reg[16][22]  (.D(dataIn[22]), .CK(n_0_0), .Q(\Memory[16] [22]), 
      .QN());
   DFF_X1 \Memory_reg[16][21]  (.D(dataIn[21]), .CK(n_0_0), .Q(\Memory[16] [21]), 
      .QN());
   DFF_X1 \Memory_reg[16][20]  (.D(dataIn[20]), .CK(n_0_0), .Q(\Memory[16] [20]), 
      .QN());
   DFF_X1 \Memory_reg[16][19]  (.D(dataIn[19]), .CK(n_0_0), .Q(\Memory[16] [19]), 
      .QN());
   DFF_X1 \Memory_reg[16][18]  (.D(dataIn[18]), .CK(n_0_0), .Q(\Memory[16] [18]), 
      .QN());
   DFF_X1 \Memory_reg[16][17]  (.D(dataIn[17]), .CK(n_0_0), .Q(\Memory[16] [17]), 
      .QN());
   DFF_X1 \Memory_reg[16][16]  (.D(dataIn[16]), .CK(n_0_0), .Q(\Memory[16] [16]), 
      .QN());
   DFF_X1 \Memory_reg[16][15]  (.D(dataIn[15]), .CK(n_0_0), .Q(\Memory[16] [15]), 
      .QN());
   DFF_X1 \Memory_reg[16][14]  (.D(dataIn[14]), .CK(n_0_0), .Q(\Memory[16] [14]), 
      .QN());
   DFF_X1 \Memory_reg[16][13]  (.D(dataIn[13]), .CK(n_0_0), .Q(\Memory[16] [13]), 
      .QN());
   DFF_X1 \Memory_reg[16][12]  (.D(dataIn[12]), .CK(n_0_0), .Q(\Memory[16] [12]), 
      .QN());
   DFF_X1 \Memory_reg[16][11]  (.D(dataIn[11]), .CK(n_0_0), .Q(\Memory[16] [11]), 
      .QN());
   DFF_X1 \Memory_reg[16][10]  (.D(dataIn[10]), .CK(n_0_0), .Q(\Memory[16] [10]), 
      .QN());
   DFF_X1 \Memory_reg[16][9]  (.D(dataIn[9]), .CK(n_0_0), .Q(\Memory[16] [9]), 
      .QN());
   DFF_X1 \Memory_reg[16][8]  (.D(dataIn[8]), .CK(n_0_0), .Q(\Memory[16] [8]), 
      .QN());
   DFF_X1 \Memory_reg[16][7]  (.D(dataIn[7]), .CK(n_0_0), .Q(\Memory[16] [7]), 
      .QN());
   DFF_X1 \Memory_reg[16][6]  (.D(dataIn[6]), .CK(n_0_0), .Q(\Memory[16] [6]), 
      .QN());
   DFF_X1 \Memory_reg[16][5]  (.D(dataIn[5]), .CK(n_0_0), .Q(\Memory[16] [5]), 
      .QN());
   DFF_X1 \Memory_reg[16][4]  (.D(dataIn[4]), .CK(n_0_0), .Q(\Memory[16] [4]), 
      .QN());
   DFF_X1 \Memory_reg[16][3]  (.D(dataIn[3]), .CK(n_0_0), .Q(\Memory[16] [3]), 
      .QN());
   DFF_X1 \Memory_reg[16][2]  (.D(dataIn[2]), .CK(n_0_0), .Q(\Memory[16] [2]), 
      .QN());
   DFF_X1 \Memory_reg[16][1]  (.D(dataIn[1]), .CK(n_0_0), .Q(\Memory[16] [1]), 
      .QN());
   DFF_X1 \Memory_reg[16][0]  (.D(dataIn[0]), .CK(n_0_0), .Q(\Memory[16] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[15]_reg  (.CK(CLK), .E(n_0_32), .SE(1'b0), 
      .GCK(n_0_1));
   DFF_X1 \Memory_reg[15][63]  (.D(Memory[63]), .CK(n_0_1), .Q(\Memory[15] [63]), 
      .QN());
   DFF_X1 \Memory_reg[15][62]  (.D(Memory[62]), .CK(n_0_1), .Q(\Memory[15] [62]), 
      .QN());
   DFF_X1 \Memory_reg[15][61]  (.D(Memory[61]), .CK(n_0_1), .Q(\Memory[15] [61]), 
      .QN());
   DFF_X1 \Memory_reg[15][60]  (.D(Memory[60]), .CK(n_0_1), .Q(\Memory[15] [60]), 
      .QN());
   DFF_X1 \Memory_reg[15][59]  (.D(Memory[59]), .CK(n_0_1), .Q(\Memory[15] [59]), 
      .QN());
   DFF_X1 \Memory_reg[15][58]  (.D(Memory[58]), .CK(n_0_1), .Q(\Memory[15] [58]), 
      .QN());
   DFF_X1 \Memory_reg[15][57]  (.D(Memory[57]), .CK(n_0_1), .Q(\Memory[15] [57]), 
      .QN());
   DFF_X1 \Memory_reg[15][56]  (.D(Memory[56]), .CK(n_0_1), .Q(\Memory[15] [56]), 
      .QN());
   DFF_X1 \Memory_reg[15][55]  (.D(Memory[55]), .CK(n_0_1), .Q(\Memory[15] [55]), 
      .QN());
   DFF_X1 \Memory_reg[15][54]  (.D(Memory[54]), .CK(n_0_1), .Q(\Memory[15] [54]), 
      .QN());
   DFF_X1 \Memory_reg[15][53]  (.D(Memory[53]), .CK(n_0_1), .Q(\Memory[15] [53]), 
      .QN());
   DFF_X1 \Memory_reg[15][52]  (.D(Memory[52]), .CK(n_0_1), .Q(\Memory[15] [52]), 
      .QN());
   DFF_X1 \Memory_reg[15][51]  (.D(Memory[51]), .CK(n_0_1), .Q(\Memory[15] [51]), 
      .QN());
   DFF_X1 \Memory_reg[15][50]  (.D(Memory[50]), .CK(n_0_1), .Q(\Memory[15] [50]), 
      .QN());
   DFF_X1 \Memory_reg[15][49]  (.D(Memory[49]), .CK(n_0_1), .Q(\Memory[15] [49]), 
      .QN());
   DFF_X1 \Memory_reg[15][48]  (.D(Memory[48]), .CK(n_0_1), .Q(\Memory[15] [48]), 
      .QN());
   DFF_X1 \Memory_reg[15][47]  (.D(Memory[47]), .CK(n_0_1), .Q(\Memory[15] [47]), 
      .QN());
   DFF_X1 \Memory_reg[15][46]  (.D(Memory[46]), .CK(n_0_1), .Q(\Memory[15] [46]), 
      .QN());
   DFF_X1 \Memory_reg[15][45]  (.D(Memory[45]), .CK(n_0_1), .Q(\Memory[15] [45]), 
      .QN());
   DFF_X1 \Memory_reg[15][44]  (.D(Memory[44]), .CK(n_0_1), .Q(\Memory[15] [44]), 
      .QN());
   DFF_X1 \Memory_reg[15][43]  (.D(Memory[43]), .CK(n_0_1), .Q(\Memory[15] [43]), 
      .QN());
   DFF_X1 \Memory_reg[15][42]  (.D(Memory[42]), .CK(n_0_1), .Q(\Memory[15] [42]), 
      .QN());
   DFF_X1 \Memory_reg[15][41]  (.D(Memory[41]), .CK(n_0_1), .Q(\Memory[15] [41]), 
      .QN());
   DFF_X1 \Memory_reg[15][40]  (.D(Memory[40]), .CK(n_0_1), .Q(\Memory[15] [40]), 
      .QN());
   DFF_X1 \Memory_reg[15][39]  (.D(Memory[39]), .CK(n_0_1), .Q(\Memory[15] [39]), 
      .QN());
   DFF_X1 \Memory_reg[15][38]  (.D(Memory[38]), .CK(n_0_1), .Q(\Memory[15] [38]), 
      .QN());
   DFF_X1 \Memory_reg[15][37]  (.D(Memory[37]), .CK(n_0_1), .Q(\Memory[15] [37]), 
      .QN());
   DFF_X1 \Memory_reg[15][36]  (.D(Memory[36]), .CK(n_0_1), .Q(\Memory[15] [36]), 
      .QN());
   DFF_X1 \Memory_reg[15][35]  (.D(Memory[35]), .CK(n_0_1), .Q(\Memory[15] [35]), 
      .QN());
   DFF_X1 \Memory_reg[15][34]  (.D(Memory[34]), .CK(n_0_1), .Q(\Memory[15] [34]), 
      .QN());
   DFF_X1 \Memory_reg[15][33]  (.D(Memory[33]), .CK(n_0_1), .Q(\Memory[15] [33]), 
      .QN());
   DFF_X1 \Memory_reg[15][32]  (.D(Memory[32]), .CK(n_0_1), .Q(\Memory[15] [32]), 
      .QN());
   DFF_X1 \Memory_reg[15][31]  (.D(Memory[31]), .CK(n_0_1), .Q(\Memory[15] [31]), 
      .QN());
   DFF_X1 \Memory_reg[15][30]  (.D(Memory[30]), .CK(n_0_1), .Q(\Memory[15] [30]), 
      .QN());
   DFF_X1 \Memory_reg[15][29]  (.D(Memory[29]), .CK(n_0_1), .Q(\Memory[15] [29]), 
      .QN());
   DFF_X1 \Memory_reg[15][28]  (.D(Memory[28]), .CK(n_0_1), .Q(\Memory[15] [28]), 
      .QN());
   DFF_X1 \Memory_reg[15][27]  (.D(Memory[27]), .CK(n_0_1), .Q(\Memory[15] [27]), 
      .QN());
   DFF_X1 \Memory_reg[15][26]  (.D(Memory[26]), .CK(n_0_1), .Q(\Memory[15] [26]), 
      .QN());
   DFF_X1 \Memory_reg[15][25]  (.D(Memory[25]), .CK(n_0_1), .Q(\Memory[15] [25]), 
      .QN());
   DFF_X1 \Memory_reg[15][24]  (.D(Memory[24]), .CK(n_0_1), .Q(\Memory[15] [24]), 
      .QN());
   DFF_X1 \Memory_reg[15][23]  (.D(Memory[23]), .CK(n_0_1), .Q(\Memory[15] [23]), 
      .QN());
   DFF_X1 \Memory_reg[15][22]  (.D(Memory[22]), .CK(n_0_1), .Q(\Memory[15] [22]), 
      .QN());
   DFF_X1 \Memory_reg[15][21]  (.D(Memory[21]), .CK(n_0_1), .Q(\Memory[15] [21]), 
      .QN());
   DFF_X1 \Memory_reg[15][20]  (.D(Memory[20]), .CK(n_0_1), .Q(\Memory[15] [20]), 
      .QN());
   DFF_X1 \Memory_reg[15][19]  (.D(Memory[19]), .CK(n_0_1), .Q(\Memory[15] [19]), 
      .QN());
   DFF_X1 \Memory_reg[15][18]  (.D(Memory[18]), .CK(n_0_1), .Q(\Memory[15] [18]), 
      .QN());
   DFF_X1 \Memory_reg[15][17]  (.D(Memory[17]), .CK(n_0_1), .Q(\Memory[15] [17]), 
      .QN());
   DFF_X1 \Memory_reg[15][16]  (.D(Memory[16]), .CK(n_0_1), .Q(\Memory[15] [16]), 
      .QN());
   DFF_X1 \Memory_reg[15][15]  (.D(Memory[15]), .CK(n_0_1), .Q(\Memory[15] [15]), 
      .QN());
   DFF_X1 \Memory_reg[15][14]  (.D(Memory[14]), .CK(n_0_1), .Q(\Memory[15] [14]), 
      .QN());
   DFF_X1 \Memory_reg[15][13]  (.D(Memory[13]), .CK(n_0_1), .Q(\Memory[15] [13]), 
      .QN());
   DFF_X1 \Memory_reg[15][12]  (.D(Memory[12]), .CK(n_0_1), .Q(\Memory[15] [12]), 
      .QN());
   DFF_X1 \Memory_reg[15][11]  (.D(Memory[11]), .CK(n_0_1), .Q(\Memory[15] [11]), 
      .QN());
   DFF_X1 \Memory_reg[15][10]  (.D(Memory[10]), .CK(n_0_1), .Q(\Memory[15] [10]), 
      .QN());
   DFF_X1 \Memory_reg[15][9]  (.D(Memory[9]), .CK(n_0_1), .Q(\Memory[15] [9]), 
      .QN());
   DFF_X1 \Memory_reg[15][8]  (.D(Memory[8]), .CK(n_0_1), .Q(\Memory[15] [8]), 
      .QN());
   DFF_X1 \Memory_reg[15][7]  (.D(Memory[7]), .CK(n_0_1), .Q(\Memory[15] [7]), 
      .QN());
   DFF_X1 \Memory_reg[15][6]  (.D(Memory[6]), .CK(n_0_1), .Q(\Memory[15] [6]), 
      .QN());
   DFF_X1 \Memory_reg[15][5]  (.D(Memory[5]), .CK(n_0_1), .Q(\Memory[15] [5]), 
      .QN());
   DFF_X1 \Memory_reg[15][4]  (.D(Memory[4]), .CK(n_0_1), .Q(\Memory[15] [4]), 
      .QN());
   DFF_X1 \Memory_reg[15][3]  (.D(Memory[3]), .CK(n_0_1), .Q(\Memory[15] [3]), 
      .QN());
   DFF_X1 \Memory_reg[15][2]  (.D(Memory[2]), .CK(n_0_1), .Q(\Memory[15] [2]), 
      .QN());
   DFF_X1 \Memory_reg[15][1]  (.D(Memory[1]), .CK(n_0_1), .Q(\Memory[15] [1]), 
      .QN());
   DFF_X1 \Memory_reg[15][0]  (.D(Memory[0]), .CK(n_0_1), .Q(\Memory[15] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[14]_reg  (.CK(CLK), .E(n_0_31), .SE(1'b0), 
      .GCK(n_0_2));
   DFF_X1 \Memory_reg[14][63]  (.D(Memory[63]), .CK(n_0_2), .Q(\Memory[14] [63]), 
      .QN());
   DFF_X1 \Memory_reg[14][62]  (.D(Memory[62]), .CK(n_0_2), .Q(\Memory[14] [62]), 
      .QN());
   DFF_X1 \Memory_reg[14][61]  (.D(Memory[61]), .CK(n_0_2), .Q(\Memory[14] [61]), 
      .QN());
   DFF_X1 \Memory_reg[14][60]  (.D(Memory[60]), .CK(n_0_2), .Q(\Memory[14] [60]), 
      .QN());
   DFF_X1 \Memory_reg[14][59]  (.D(Memory[59]), .CK(n_0_2), .Q(\Memory[14] [59]), 
      .QN());
   DFF_X1 \Memory_reg[14][58]  (.D(Memory[58]), .CK(n_0_2), .Q(\Memory[14] [58]), 
      .QN());
   DFF_X1 \Memory_reg[14][57]  (.D(Memory[57]), .CK(n_0_2), .Q(\Memory[14] [57]), 
      .QN());
   DFF_X1 \Memory_reg[14][56]  (.D(Memory[56]), .CK(n_0_2), .Q(\Memory[14] [56]), 
      .QN());
   DFF_X1 \Memory_reg[14][55]  (.D(Memory[55]), .CK(n_0_2), .Q(\Memory[14] [55]), 
      .QN());
   DFF_X1 \Memory_reg[14][54]  (.D(Memory[54]), .CK(n_0_2), .Q(\Memory[14] [54]), 
      .QN());
   DFF_X1 \Memory_reg[14][53]  (.D(Memory[53]), .CK(n_0_2), .Q(\Memory[14] [53]), 
      .QN());
   DFF_X1 \Memory_reg[14][52]  (.D(Memory[52]), .CK(n_0_2), .Q(\Memory[14] [52]), 
      .QN());
   DFF_X1 \Memory_reg[14][51]  (.D(Memory[51]), .CK(n_0_2), .Q(\Memory[14] [51]), 
      .QN());
   DFF_X1 \Memory_reg[14][50]  (.D(Memory[50]), .CK(n_0_2), .Q(\Memory[14] [50]), 
      .QN());
   DFF_X1 \Memory_reg[14][49]  (.D(Memory[49]), .CK(n_0_2), .Q(\Memory[14] [49]), 
      .QN());
   DFF_X1 \Memory_reg[14][48]  (.D(Memory[48]), .CK(n_0_2), .Q(\Memory[14] [48]), 
      .QN());
   DFF_X1 \Memory_reg[14][47]  (.D(Memory[47]), .CK(n_0_2), .Q(\Memory[14] [47]), 
      .QN());
   DFF_X1 \Memory_reg[14][46]  (.D(Memory[46]), .CK(n_0_2), .Q(\Memory[14] [46]), 
      .QN());
   DFF_X1 \Memory_reg[14][45]  (.D(Memory[45]), .CK(n_0_2), .Q(\Memory[14] [45]), 
      .QN());
   DFF_X1 \Memory_reg[14][44]  (.D(Memory[44]), .CK(n_0_2), .Q(\Memory[14] [44]), 
      .QN());
   DFF_X1 \Memory_reg[14][43]  (.D(Memory[43]), .CK(n_0_2), .Q(\Memory[14] [43]), 
      .QN());
   DFF_X1 \Memory_reg[14][42]  (.D(Memory[42]), .CK(n_0_2), .Q(\Memory[14] [42]), 
      .QN());
   DFF_X1 \Memory_reg[14][41]  (.D(Memory[41]), .CK(n_0_2), .Q(\Memory[14] [41]), 
      .QN());
   DFF_X1 \Memory_reg[14][40]  (.D(Memory[40]), .CK(n_0_2), .Q(\Memory[14] [40]), 
      .QN());
   DFF_X1 \Memory_reg[14][39]  (.D(Memory[39]), .CK(n_0_2), .Q(\Memory[14] [39]), 
      .QN());
   DFF_X1 \Memory_reg[14][38]  (.D(Memory[38]), .CK(n_0_2), .Q(\Memory[14] [38]), 
      .QN());
   DFF_X1 \Memory_reg[14][37]  (.D(Memory[37]), .CK(n_0_2), .Q(\Memory[14] [37]), 
      .QN());
   DFF_X1 \Memory_reg[14][36]  (.D(Memory[36]), .CK(n_0_2), .Q(\Memory[14] [36]), 
      .QN());
   DFF_X1 \Memory_reg[14][35]  (.D(Memory[35]), .CK(n_0_2), .Q(\Memory[14] [35]), 
      .QN());
   DFF_X1 \Memory_reg[14][34]  (.D(Memory[34]), .CK(n_0_2), .Q(\Memory[14] [34]), 
      .QN());
   DFF_X1 \Memory_reg[14][33]  (.D(Memory[33]), .CK(n_0_2), .Q(\Memory[14] [33]), 
      .QN());
   DFF_X1 \Memory_reg[14][32]  (.D(Memory[32]), .CK(n_0_2), .Q(\Memory[14] [32]), 
      .QN());
   DFF_X1 \Memory_reg[14][31]  (.D(Memory[31]), .CK(n_0_2), .Q(\Memory[14] [31]), 
      .QN());
   DFF_X1 \Memory_reg[14][30]  (.D(Memory[30]), .CK(n_0_2), .Q(\Memory[14] [30]), 
      .QN());
   DFF_X1 \Memory_reg[14][29]  (.D(Memory[29]), .CK(n_0_2), .Q(\Memory[14] [29]), 
      .QN());
   DFF_X1 \Memory_reg[14][28]  (.D(Memory[28]), .CK(n_0_2), .Q(\Memory[14] [28]), 
      .QN());
   DFF_X1 \Memory_reg[14][27]  (.D(Memory[27]), .CK(n_0_2), .Q(\Memory[14] [27]), 
      .QN());
   DFF_X1 \Memory_reg[14][26]  (.D(Memory[26]), .CK(n_0_2), .Q(\Memory[14] [26]), 
      .QN());
   DFF_X1 \Memory_reg[14][25]  (.D(Memory[25]), .CK(n_0_2), .Q(\Memory[14] [25]), 
      .QN());
   DFF_X1 \Memory_reg[14][24]  (.D(Memory[24]), .CK(n_0_2), .Q(\Memory[14] [24]), 
      .QN());
   DFF_X1 \Memory_reg[14][23]  (.D(Memory[23]), .CK(n_0_2), .Q(\Memory[14] [23]), 
      .QN());
   DFF_X1 \Memory_reg[14][22]  (.D(Memory[22]), .CK(n_0_2), .Q(\Memory[14] [22]), 
      .QN());
   DFF_X1 \Memory_reg[14][21]  (.D(Memory[21]), .CK(n_0_2), .Q(\Memory[14] [21]), 
      .QN());
   DFF_X1 \Memory_reg[14][20]  (.D(Memory[20]), .CK(n_0_2), .Q(\Memory[14] [20]), 
      .QN());
   DFF_X1 \Memory_reg[14][19]  (.D(Memory[19]), .CK(n_0_2), .Q(\Memory[14] [19]), 
      .QN());
   DFF_X1 \Memory_reg[14][18]  (.D(Memory[18]), .CK(n_0_2), .Q(\Memory[14] [18]), 
      .QN());
   DFF_X1 \Memory_reg[14][17]  (.D(Memory[17]), .CK(n_0_2), .Q(\Memory[14] [17]), 
      .QN());
   DFF_X1 \Memory_reg[14][16]  (.D(Memory[16]), .CK(n_0_2), .Q(\Memory[14] [16]), 
      .QN());
   DFF_X1 \Memory_reg[14][15]  (.D(Memory[15]), .CK(n_0_2), .Q(\Memory[14] [15]), 
      .QN());
   DFF_X1 \Memory_reg[14][14]  (.D(Memory[14]), .CK(n_0_2), .Q(\Memory[14] [14]), 
      .QN());
   DFF_X1 \Memory_reg[14][13]  (.D(Memory[13]), .CK(n_0_2), .Q(\Memory[14] [13]), 
      .QN());
   DFF_X1 \Memory_reg[14][12]  (.D(Memory[12]), .CK(n_0_2), .Q(\Memory[14] [12]), 
      .QN());
   DFF_X1 \Memory_reg[14][11]  (.D(Memory[11]), .CK(n_0_2), .Q(\Memory[14] [11]), 
      .QN());
   DFF_X1 \Memory_reg[14][10]  (.D(Memory[10]), .CK(n_0_2), .Q(\Memory[14] [10]), 
      .QN());
   DFF_X1 \Memory_reg[14][9]  (.D(Memory[9]), .CK(n_0_2), .Q(\Memory[14] [9]), 
      .QN());
   DFF_X1 \Memory_reg[14][8]  (.D(Memory[8]), .CK(n_0_2), .Q(\Memory[14] [8]), 
      .QN());
   DFF_X1 \Memory_reg[14][7]  (.D(Memory[7]), .CK(n_0_2), .Q(\Memory[14] [7]), 
      .QN());
   DFF_X1 \Memory_reg[14][6]  (.D(Memory[6]), .CK(n_0_2), .Q(\Memory[14] [6]), 
      .QN());
   DFF_X1 \Memory_reg[14][5]  (.D(Memory[5]), .CK(n_0_2), .Q(\Memory[14] [5]), 
      .QN());
   DFF_X1 \Memory_reg[14][4]  (.D(Memory[4]), .CK(n_0_2), .Q(\Memory[14] [4]), 
      .QN());
   DFF_X1 \Memory_reg[14][3]  (.D(Memory[3]), .CK(n_0_2), .Q(\Memory[14] [3]), 
      .QN());
   DFF_X1 \Memory_reg[14][2]  (.D(Memory[2]), .CK(n_0_2), .Q(\Memory[14] [2]), 
      .QN());
   DFF_X1 \Memory_reg[14][1]  (.D(Memory[1]), .CK(n_0_2), .Q(\Memory[14] [1]), 
      .QN());
   DFF_X1 \Memory_reg[14][0]  (.D(Memory[0]), .CK(n_0_2), .Q(\Memory[14] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[13]_reg  (.CK(CLK), .E(n_0_30), .SE(1'b0), 
      .GCK(n_0_3));
   DFF_X1 \Memory_reg[13][63]  (.D(Memory[63]), .CK(n_0_3), .Q(\Memory[13] [63]), 
      .QN());
   DFF_X1 \Memory_reg[13][62]  (.D(Memory[62]), .CK(n_0_3), .Q(\Memory[13] [62]), 
      .QN());
   DFF_X1 \Memory_reg[13][61]  (.D(Memory[61]), .CK(n_0_3), .Q(\Memory[13] [61]), 
      .QN());
   DFF_X1 \Memory_reg[13][60]  (.D(Memory[60]), .CK(n_0_3), .Q(\Memory[13] [60]), 
      .QN());
   DFF_X1 \Memory_reg[13][59]  (.D(Memory[59]), .CK(n_0_3), .Q(\Memory[13] [59]), 
      .QN());
   DFF_X1 \Memory_reg[13][58]  (.D(Memory[58]), .CK(n_0_3), .Q(\Memory[13] [58]), 
      .QN());
   DFF_X1 \Memory_reg[13][57]  (.D(Memory[57]), .CK(n_0_3), .Q(\Memory[13] [57]), 
      .QN());
   DFF_X1 \Memory_reg[13][56]  (.D(Memory[56]), .CK(n_0_3), .Q(\Memory[13] [56]), 
      .QN());
   DFF_X1 \Memory_reg[13][55]  (.D(Memory[55]), .CK(n_0_3), .Q(\Memory[13] [55]), 
      .QN());
   DFF_X1 \Memory_reg[13][54]  (.D(Memory[54]), .CK(n_0_3), .Q(\Memory[13] [54]), 
      .QN());
   DFF_X1 \Memory_reg[13][53]  (.D(Memory[53]), .CK(n_0_3), .Q(\Memory[13] [53]), 
      .QN());
   DFF_X1 \Memory_reg[13][52]  (.D(Memory[52]), .CK(n_0_3), .Q(\Memory[13] [52]), 
      .QN());
   DFF_X1 \Memory_reg[13][51]  (.D(Memory[51]), .CK(n_0_3), .Q(\Memory[13] [51]), 
      .QN());
   DFF_X1 \Memory_reg[13][50]  (.D(Memory[50]), .CK(n_0_3), .Q(\Memory[13] [50]), 
      .QN());
   DFF_X1 \Memory_reg[13][49]  (.D(Memory[49]), .CK(n_0_3), .Q(\Memory[13] [49]), 
      .QN());
   DFF_X1 \Memory_reg[13][48]  (.D(Memory[48]), .CK(n_0_3), .Q(\Memory[13] [48]), 
      .QN());
   DFF_X1 \Memory_reg[13][47]  (.D(Memory[47]), .CK(n_0_3), .Q(\Memory[13] [47]), 
      .QN());
   DFF_X1 \Memory_reg[13][46]  (.D(Memory[46]), .CK(n_0_3), .Q(\Memory[13] [46]), 
      .QN());
   DFF_X1 \Memory_reg[13][45]  (.D(Memory[45]), .CK(n_0_3), .Q(\Memory[13] [45]), 
      .QN());
   DFF_X1 \Memory_reg[13][44]  (.D(Memory[44]), .CK(n_0_3), .Q(\Memory[13] [44]), 
      .QN());
   DFF_X1 \Memory_reg[13][43]  (.D(Memory[43]), .CK(n_0_3), .Q(\Memory[13] [43]), 
      .QN());
   DFF_X1 \Memory_reg[13][42]  (.D(Memory[42]), .CK(n_0_3), .Q(\Memory[13] [42]), 
      .QN());
   DFF_X1 \Memory_reg[13][41]  (.D(Memory[41]), .CK(n_0_3), .Q(\Memory[13] [41]), 
      .QN());
   DFF_X1 \Memory_reg[13][40]  (.D(Memory[40]), .CK(n_0_3), .Q(\Memory[13] [40]), 
      .QN());
   DFF_X1 \Memory_reg[13][39]  (.D(Memory[39]), .CK(n_0_3), .Q(\Memory[13] [39]), 
      .QN());
   DFF_X1 \Memory_reg[13][38]  (.D(Memory[38]), .CK(n_0_3), .Q(\Memory[13] [38]), 
      .QN());
   DFF_X1 \Memory_reg[13][37]  (.D(Memory[37]), .CK(n_0_3), .Q(\Memory[13] [37]), 
      .QN());
   DFF_X1 \Memory_reg[13][36]  (.D(Memory[36]), .CK(n_0_3), .Q(\Memory[13] [36]), 
      .QN());
   DFF_X1 \Memory_reg[13][35]  (.D(Memory[35]), .CK(n_0_3), .Q(\Memory[13] [35]), 
      .QN());
   DFF_X1 \Memory_reg[13][34]  (.D(Memory[34]), .CK(n_0_3), .Q(\Memory[13] [34]), 
      .QN());
   DFF_X1 \Memory_reg[13][33]  (.D(Memory[33]), .CK(n_0_3), .Q(\Memory[13] [33]), 
      .QN());
   DFF_X1 \Memory_reg[13][32]  (.D(Memory[32]), .CK(n_0_3), .Q(\Memory[13] [32]), 
      .QN());
   DFF_X1 \Memory_reg[13][31]  (.D(Memory[31]), .CK(n_0_3), .Q(\Memory[13] [31]), 
      .QN());
   DFF_X1 \Memory_reg[13][30]  (.D(Memory[30]), .CK(n_0_3), .Q(\Memory[13] [30]), 
      .QN());
   DFF_X1 \Memory_reg[13][29]  (.D(Memory[29]), .CK(n_0_3), .Q(\Memory[13] [29]), 
      .QN());
   DFF_X1 \Memory_reg[13][28]  (.D(Memory[28]), .CK(n_0_3), .Q(\Memory[13] [28]), 
      .QN());
   DFF_X1 \Memory_reg[13][27]  (.D(Memory[27]), .CK(n_0_3), .Q(\Memory[13] [27]), 
      .QN());
   DFF_X1 \Memory_reg[13][26]  (.D(Memory[26]), .CK(n_0_3), .Q(\Memory[13] [26]), 
      .QN());
   DFF_X1 \Memory_reg[13][25]  (.D(Memory[25]), .CK(n_0_3), .Q(\Memory[13] [25]), 
      .QN());
   DFF_X1 \Memory_reg[13][24]  (.D(Memory[24]), .CK(n_0_3), .Q(\Memory[13] [24]), 
      .QN());
   DFF_X1 \Memory_reg[13][23]  (.D(Memory[23]), .CK(n_0_3), .Q(\Memory[13] [23]), 
      .QN());
   DFF_X1 \Memory_reg[13][22]  (.D(Memory[22]), .CK(n_0_3), .Q(\Memory[13] [22]), 
      .QN());
   DFF_X1 \Memory_reg[13][21]  (.D(Memory[21]), .CK(n_0_3), .Q(\Memory[13] [21]), 
      .QN());
   DFF_X1 \Memory_reg[13][20]  (.D(Memory[20]), .CK(n_0_3), .Q(\Memory[13] [20]), 
      .QN());
   DFF_X1 \Memory_reg[13][19]  (.D(Memory[19]), .CK(n_0_3), .Q(\Memory[13] [19]), 
      .QN());
   DFF_X1 \Memory_reg[13][18]  (.D(Memory[18]), .CK(n_0_3), .Q(\Memory[13] [18]), 
      .QN());
   DFF_X1 \Memory_reg[13][17]  (.D(Memory[17]), .CK(n_0_3), .Q(\Memory[13] [17]), 
      .QN());
   DFF_X1 \Memory_reg[13][16]  (.D(Memory[16]), .CK(n_0_3), .Q(\Memory[13] [16]), 
      .QN());
   DFF_X1 \Memory_reg[13][15]  (.D(Memory[15]), .CK(n_0_3), .Q(\Memory[13] [15]), 
      .QN());
   DFF_X1 \Memory_reg[13][14]  (.D(Memory[14]), .CK(n_0_3), .Q(\Memory[13] [14]), 
      .QN());
   DFF_X1 \Memory_reg[13][13]  (.D(Memory[13]), .CK(n_0_3), .Q(\Memory[13] [13]), 
      .QN());
   DFF_X1 \Memory_reg[13][12]  (.D(Memory[12]), .CK(n_0_3), .Q(\Memory[13] [12]), 
      .QN());
   DFF_X1 \Memory_reg[13][11]  (.D(Memory[11]), .CK(n_0_3), .Q(\Memory[13] [11]), 
      .QN());
   DFF_X1 \Memory_reg[13][10]  (.D(Memory[10]), .CK(n_0_3), .Q(\Memory[13] [10]), 
      .QN());
   DFF_X1 \Memory_reg[13][9]  (.D(Memory[9]), .CK(n_0_3), .Q(\Memory[13] [9]), 
      .QN());
   DFF_X1 \Memory_reg[13][8]  (.D(Memory[8]), .CK(n_0_3), .Q(\Memory[13] [8]), 
      .QN());
   DFF_X1 \Memory_reg[13][7]  (.D(Memory[7]), .CK(n_0_3), .Q(\Memory[13] [7]), 
      .QN());
   DFF_X1 \Memory_reg[13][6]  (.D(Memory[6]), .CK(n_0_3), .Q(\Memory[13] [6]), 
      .QN());
   DFF_X1 \Memory_reg[13][5]  (.D(Memory[5]), .CK(n_0_3), .Q(\Memory[13] [5]), 
      .QN());
   DFF_X1 \Memory_reg[13][4]  (.D(Memory[4]), .CK(n_0_3), .Q(\Memory[13] [4]), 
      .QN());
   DFF_X1 \Memory_reg[13][3]  (.D(Memory[3]), .CK(n_0_3), .Q(\Memory[13] [3]), 
      .QN());
   DFF_X1 \Memory_reg[13][2]  (.D(Memory[2]), .CK(n_0_3), .Q(\Memory[13] [2]), 
      .QN());
   DFF_X1 \Memory_reg[13][1]  (.D(Memory[1]), .CK(n_0_3), .Q(\Memory[13] [1]), 
      .QN());
   DFF_X1 \Memory_reg[13][0]  (.D(Memory[0]), .CK(n_0_3), .Q(\Memory[13] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[12]_reg  (.CK(CLK), .E(n_0_29), .SE(1'b0), 
      .GCK(n_0_4));
   DFF_X1 \Memory_reg[12][63]  (.D(Memory[63]), .CK(n_0_4), .Q(\Memory[12] [63]), 
      .QN());
   DFF_X1 \Memory_reg[12][62]  (.D(Memory[62]), .CK(n_0_4), .Q(\Memory[12] [62]), 
      .QN());
   DFF_X1 \Memory_reg[12][61]  (.D(Memory[61]), .CK(n_0_4), .Q(\Memory[12] [61]), 
      .QN());
   DFF_X1 \Memory_reg[12][60]  (.D(Memory[60]), .CK(n_0_4), .Q(\Memory[12] [60]), 
      .QN());
   DFF_X1 \Memory_reg[12][59]  (.D(Memory[59]), .CK(n_0_4), .Q(\Memory[12] [59]), 
      .QN());
   DFF_X1 \Memory_reg[12][58]  (.D(Memory[58]), .CK(n_0_4), .Q(\Memory[12] [58]), 
      .QN());
   DFF_X1 \Memory_reg[12][57]  (.D(Memory[57]), .CK(n_0_4), .Q(\Memory[12] [57]), 
      .QN());
   DFF_X1 \Memory_reg[12][56]  (.D(Memory[56]), .CK(n_0_4), .Q(\Memory[12] [56]), 
      .QN());
   DFF_X1 \Memory_reg[12][55]  (.D(Memory[55]), .CK(n_0_4), .Q(\Memory[12] [55]), 
      .QN());
   DFF_X1 \Memory_reg[12][54]  (.D(Memory[54]), .CK(n_0_4), .Q(\Memory[12] [54]), 
      .QN());
   DFF_X1 \Memory_reg[12][53]  (.D(Memory[53]), .CK(n_0_4), .Q(\Memory[12] [53]), 
      .QN());
   DFF_X1 \Memory_reg[12][52]  (.D(Memory[52]), .CK(n_0_4), .Q(\Memory[12] [52]), 
      .QN());
   DFF_X1 \Memory_reg[12][51]  (.D(Memory[51]), .CK(n_0_4), .Q(\Memory[12] [51]), 
      .QN());
   DFF_X1 \Memory_reg[12][50]  (.D(Memory[50]), .CK(n_0_4), .Q(\Memory[12] [50]), 
      .QN());
   DFF_X1 \Memory_reg[12][49]  (.D(Memory[49]), .CK(n_0_4), .Q(\Memory[12] [49]), 
      .QN());
   DFF_X1 \Memory_reg[12][48]  (.D(Memory[48]), .CK(n_0_4), .Q(\Memory[12] [48]), 
      .QN());
   DFF_X1 \Memory_reg[12][47]  (.D(Memory[47]), .CK(n_0_4), .Q(\Memory[12] [47]), 
      .QN());
   DFF_X1 \Memory_reg[12][46]  (.D(Memory[46]), .CK(n_0_4), .Q(\Memory[12] [46]), 
      .QN());
   DFF_X1 \Memory_reg[12][45]  (.D(Memory[45]), .CK(n_0_4), .Q(\Memory[12] [45]), 
      .QN());
   DFF_X1 \Memory_reg[12][44]  (.D(Memory[44]), .CK(n_0_4), .Q(\Memory[12] [44]), 
      .QN());
   DFF_X1 \Memory_reg[12][43]  (.D(Memory[43]), .CK(n_0_4), .Q(\Memory[12] [43]), 
      .QN());
   DFF_X1 \Memory_reg[12][42]  (.D(Memory[42]), .CK(n_0_4), .Q(\Memory[12] [42]), 
      .QN());
   DFF_X1 \Memory_reg[12][41]  (.D(Memory[41]), .CK(n_0_4), .Q(\Memory[12] [41]), 
      .QN());
   DFF_X1 \Memory_reg[12][40]  (.D(Memory[40]), .CK(n_0_4), .Q(\Memory[12] [40]), 
      .QN());
   DFF_X1 \Memory_reg[12][39]  (.D(Memory[39]), .CK(n_0_4), .Q(\Memory[12] [39]), 
      .QN());
   DFF_X1 \Memory_reg[12][38]  (.D(Memory[38]), .CK(n_0_4), .Q(\Memory[12] [38]), 
      .QN());
   DFF_X1 \Memory_reg[12][37]  (.D(Memory[37]), .CK(n_0_4), .Q(\Memory[12] [37]), 
      .QN());
   DFF_X1 \Memory_reg[12][36]  (.D(Memory[36]), .CK(n_0_4), .Q(\Memory[12] [36]), 
      .QN());
   DFF_X1 \Memory_reg[12][35]  (.D(Memory[35]), .CK(n_0_4), .Q(\Memory[12] [35]), 
      .QN());
   DFF_X1 \Memory_reg[12][34]  (.D(Memory[34]), .CK(n_0_4), .Q(\Memory[12] [34]), 
      .QN());
   DFF_X1 \Memory_reg[12][33]  (.D(Memory[33]), .CK(n_0_4), .Q(\Memory[12] [33]), 
      .QN());
   DFF_X1 \Memory_reg[12][32]  (.D(Memory[32]), .CK(n_0_4), .Q(\Memory[12] [32]), 
      .QN());
   DFF_X1 \Memory_reg[12][31]  (.D(Memory[31]), .CK(n_0_4), .Q(\Memory[12] [31]), 
      .QN());
   DFF_X1 \Memory_reg[12][30]  (.D(Memory[30]), .CK(n_0_4), .Q(\Memory[12] [30]), 
      .QN());
   DFF_X1 \Memory_reg[12][29]  (.D(Memory[29]), .CK(n_0_4), .Q(\Memory[12] [29]), 
      .QN());
   DFF_X1 \Memory_reg[12][28]  (.D(Memory[28]), .CK(n_0_4), .Q(\Memory[12] [28]), 
      .QN());
   DFF_X1 \Memory_reg[12][27]  (.D(Memory[27]), .CK(n_0_4), .Q(\Memory[12] [27]), 
      .QN());
   DFF_X1 \Memory_reg[12][26]  (.D(Memory[26]), .CK(n_0_4), .Q(\Memory[12] [26]), 
      .QN());
   DFF_X1 \Memory_reg[12][25]  (.D(Memory[25]), .CK(n_0_4), .Q(\Memory[12] [25]), 
      .QN());
   DFF_X1 \Memory_reg[12][24]  (.D(Memory[24]), .CK(n_0_4), .Q(\Memory[12] [24]), 
      .QN());
   DFF_X1 \Memory_reg[12][23]  (.D(Memory[23]), .CK(n_0_4), .Q(\Memory[12] [23]), 
      .QN());
   DFF_X1 \Memory_reg[12][22]  (.D(Memory[22]), .CK(n_0_4), .Q(\Memory[12] [22]), 
      .QN());
   DFF_X1 \Memory_reg[12][21]  (.D(Memory[21]), .CK(n_0_4), .Q(\Memory[12] [21]), 
      .QN());
   DFF_X1 \Memory_reg[12][20]  (.D(Memory[20]), .CK(n_0_4), .Q(\Memory[12] [20]), 
      .QN());
   DFF_X1 \Memory_reg[12][19]  (.D(Memory[19]), .CK(n_0_4), .Q(\Memory[12] [19]), 
      .QN());
   DFF_X1 \Memory_reg[12][18]  (.D(Memory[18]), .CK(n_0_4), .Q(\Memory[12] [18]), 
      .QN());
   DFF_X1 \Memory_reg[12][17]  (.D(Memory[17]), .CK(n_0_4), .Q(\Memory[12] [17]), 
      .QN());
   DFF_X1 \Memory_reg[12][16]  (.D(Memory[16]), .CK(n_0_4), .Q(\Memory[12] [16]), 
      .QN());
   DFF_X1 \Memory_reg[12][15]  (.D(Memory[15]), .CK(n_0_4), .Q(\Memory[12] [15]), 
      .QN());
   DFF_X1 \Memory_reg[12][14]  (.D(Memory[14]), .CK(n_0_4), .Q(\Memory[12] [14]), 
      .QN());
   DFF_X1 \Memory_reg[12][13]  (.D(Memory[13]), .CK(n_0_4), .Q(\Memory[12] [13]), 
      .QN());
   DFF_X1 \Memory_reg[12][12]  (.D(Memory[12]), .CK(n_0_4), .Q(\Memory[12] [12]), 
      .QN());
   DFF_X1 \Memory_reg[12][11]  (.D(Memory[11]), .CK(n_0_4), .Q(\Memory[12] [11]), 
      .QN());
   DFF_X1 \Memory_reg[12][10]  (.D(Memory[10]), .CK(n_0_4), .Q(\Memory[12] [10]), 
      .QN());
   DFF_X1 \Memory_reg[12][9]  (.D(Memory[9]), .CK(n_0_4), .Q(\Memory[12] [9]), 
      .QN());
   DFF_X1 \Memory_reg[12][8]  (.D(Memory[8]), .CK(n_0_4), .Q(\Memory[12] [8]), 
      .QN());
   DFF_X1 \Memory_reg[12][7]  (.D(Memory[7]), .CK(n_0_4), .Q(\Memory[12] [7]), 
      .QN());
   DFF_X1 \Memory_reg[12][6]  (.D(Memory[6]), .CK(n_0_4), .Q(\Memory[12] [6]), 
      .QN());
   DFF_X1 \Memory_reg[12][5]  (.D(Memory[5]), .CK(n_0_4), .Q(\Memory[12] [5]), 
      .QN());
   DFF_X1 \Memory_reg[12][4]  (.D(Memory[4]), .CK(n_0_4), .Q(\Memory[12] [4]), 
      .QN());
   DFF_X1 \Memory_reg[12][3]  (.D(Memory[3]), .CK(n_0_4), .Q(\Memory[12] [3]), 
      .QN());
   DFF_X1 \Memory_reg[12][2]  (.D(Memory[2]), .CK(n_0_4), .Q(\Memory[12] [2]), 
      .QN());
   DFF_X1 \Memory_reg[12][1]  (.D(Memory[1]), .CK(n_0_4), .Q(\Memory[12] [1]), 
      .QN());
   DFF_X1 \Memory_reg[12][0]  (.D(Memory[0]), .CK(n_0_4), .Q(\Memory[12] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[11]_reg  (.CK(CLK), .E(n_0_28), .SE(1'b0), 
      .GCK(n_0_5));
   DFF_X1 \Memory_reg[11][63]  (.D(Memory[63]), .CK(n_0_5), .Q(\Memory[11] [63]), 
      .QN());
   DFF_X1 \Memory_reg[11][62]  (.D(Memory[62]), .CK(n_0_5), .Q(\Memory[11] [62]), 
      .QN());
   DFF_X1 \Memory_reg[11][61]  (.D(Memory[61]), .CK(n_0_5), .Q(\Memory[11] [61]), 
      .QN());
   DFF_X1 \Memory_reg[11][60]  (.D(Memory[60]), .CK(n_0_5), .Q(\Memory[11] [60]), 
      .QN());
   DFF_X1 \Memory_reg[11][59]  (.D(Memory[59]), .CK(n_0_5), .Q(\Memory[11] [59]), 
      .QN());
   DFF_X1 \Memory_reg[11][58]  (.D(Memory[58]), .CK(n_0_5), .Q(\Memory[11] [58]), 
      .QN());
   DFF_X1 \Memory_reg[11][57]  (.D(Memory[57]), .CK(n_0_5), .Q(\Memory[11] [57]), 
      .QN());
   DFF_X1 \Memory_reg[11][56]  (.D(Memory[56]), .CK(n_0_5), .Q(\Memory[11] [56]), 
      .QN());
   DFF_X1 \Memory_reg[11][55]  (.D(Memory[55]), .CK(n_0_5), .Q(\Memory[11] [55]), 
      .QN());
   DFF_X1 \Memory_reg[11][54]  (.D(Memory[54]), .CK(n_0_5), .Q(\Memory[11] [54]), 
      .QN());
   DFF_X1 \Memory_reg[11][53]  (.D(Memory[53]), .CK(n_0_5), .Q(\Memory[11] [53]), 
      .QN());
   DFF_X1 \Memory_reg[11][52]  (.D(Memory[52]), .CK(n_0_5), .Q(\Memory[11] [52]), 
      .QN());
   DFF_X1 \Memory_reg[11][51]  (.D(Memory[51]), .CK(n_0_5), .Q(\Memory[11] [51]), 
      .QN());
   DFF_X1 \Memory_reg[11][50]  (.D(Memory[50]), .CK(n_0_5), .Q(\Memory[11] [50]), 
      .QN());
   DFF_X1 \Memory_reg[11][49]  (.D(Memory[49]), .CK(n_0_5), .Q(\Memory[11] [49]), 
      .QN());
   DFF_X1 \Memory_reg[11][48]  (.D(Memory[48]), .CK(n_0_5), .Q(\Memory[11] [48]), 
      .QN());
   DFF_X1 \Memory_reg[11][47]  (.D(Memory[47]), .CK(n_0_5), .Q(\Memory[11] [47]), 
      .QN());
   DFF_X1 \Memory_reg[11][46]  (.D(Memory[46]), .CK(n_0_5), .Q(\Memory[11] [46]), 
      .QN());
   DFF_X1 \Memory_reg[11][45]  (.D(Memory[45]), .CK(n_0_5), .Q(\Memory[11] [45]), 
      .QN());
   DFF_X1 \Memory_reg[11][44]  (.D(Memory[44]), .CK(n_0_5), .Q(\Memory[11] [44]), 
      .QN());
   DFF_X1 \Memory_reg[11][43]  (.D(Memory[43]), .CK(n_0_5), .Q(\Memory[11] [43]), 
      .QN());
   DFF_X1 \Memory_reg[11][42]  (.D(Memory[42]), .CK(n_0_5), .Q(\Memory[11] [42]), 
      .QN());
   DFF_X1 \Memory_reg[11][41]  (.D(Memory[41]), .CK(n_0_5), .Q(\Memory[11] [41]), 
      .QN());
   DFF_X1 \Memory_reg[11][40]  (.D(Memory[40]), .CK(n_0_5), .Q(\Memory[11] [40]), 
      .QN());
   DFF_X1 \Memory_reg[11][39]  (.D(Memory[39]), .CK(n_0_5), .Q(\Memory[11] [39]), 
      .QN());
   DFF_X1 \Memory_reg[11][38]  (.D(Memory[38]), .CK(n_0_5), .Q(\Memory[11] [38]), 
      .QN());
   DFF_X1 \Memory_reg[11][37]  (.D(Memory[37]), .CK(n_0_5), .Q(\Memory[11] [37]), 
      .QN());
   DFF_X1 \Memory_reg[11][36]  (.D(Memory[36]), .CK(n_0_5), .Q(\Memory[11] [36]), 
      .QN());
   DFF_X1 \Memory_reg[11][35]  (.D(Memory[35]), .CK(n_0_5), .Q(\Memory[11] [35]), 
      .QN());
   DFF_X1 \Memory_reg[11][34]  (.D(Memory[34]), .CK(n_0_5), .Q(\Memory[11] [34]), 
      .QN());
   DFF_X1 \Memory_reg[11][33]  (.D(Memory[33]), .CK(n_0_5), .Q(\Memory[11] [33]), 
      .QN());
   DFF_X1 \Memory_reg[11][32]  (.D(Memory[32]), .CK(n_0_5), .Q(\Memory[11] [32]), 
      .QN());
   DFF_X1 \Memory_reg[11][31]  (.D(Memory[31]), .CK(n_0_5), .Q(\Memory[11] [31]), 
      .QN());
   DFF_X1 \Memory_reg[11][30]  (.D(Memory[30]), .CK(n_0_5), .Q(\Memory[11] [30]), 
      .QN());
   DFF_X1 \Memory_reg[11][29]  (.D(Memory[29]), .CK(n_0_5), .Q(\Memory[11] [29]), 
      .QN());
   DFF_X1 \Memory_reg[11][28]  (.D(Memory[28]), .CK(n_0_5), .Q(\Memory[11] [28]), 
      .QN());
   DFF_X1 \Memory_reg[11][27]  (.D(Memory[27]), .CK(n_0_5), .Q(\Memory[11] [27]), 
      .QN());
   DFF_X1 \Memory_reg[11][26]  (.D(Memory[26]), .CK(n_0_5), .Q(\Memory[11] [26]), 
      .QN());
   DFF_X1 \Memory_reg[11][25]  (.D(Memory[25]), .CK(n_0_5), .Q(\Memory[11] [25]), 
      .QN());
   DFF_X1 \Memory_reg[11][24]  (.D(Memory[24]), .CK(n_0_5), .Q(\Memory[11] [24]), 
      .QN());
   DFF_X1 \Memory_reg[11][23]  (.D(Memory[23]), .CK(n_0_5), .Q(\Memory[11] [23]), 
      .QN());
   DFF_X1 \Memory_reg[11][22]  (.D(Memory[22]), .CK(n_0_5), .Q(\Memory[11] [22]), 
      .QN());
   DFF_X1 \Memory_reg[11][21]  (.D(Memory[21]), .CK(n_0_5), .Q(\Memory[11] [21]), 
      .QN());
   DFF_X1 \Memory_reg[11][20]  (.D(Memory[20]), .CK(n_0_5), .Q(\Memory[11] [20]), 
      .QN());
   DFF_X1 \Memory_reg[11][19]  (.D(Memory[19]), .CK(n_0_5), .Q(\Memory[11] [19]), 
      .QN());
   DFF_X1 \Memory_reg[11][18]  (.D(Memory[18]), .CK(n_0_5), .Q(\Memory[11] [18]), 
      .QN());
   DFF_X1 \Memory_reg[11][17]  (.D(Memory[17]), .CK(n_0_5), .Q(\Memory[11] [17]), 
      .QN());
   DFF_X1 \Memory_reg[11][16]  (.D(Memory[16]), .CK(n_0_5), .Q(\Memory[11] [16]), 
      .QN());
   DFF_X1 \Memory_reg[11][15]  (.D(Memory[15]), .CK(n_0_5), .Q(\Memory[11] [15]), 
      .QN());
   DFF_X1 \Memory_reg[11][14]  (.D(Memory[14]), .CK(n_0_5), .Q(\Memory[11] [14]), 
      .QN());
   DFF_X1 \Memory_reg[11][13]  (.D(Memory[13]), .CK(n_0_5), .Q(\Memory[11] [13]), 
      .QN());
   DFF_X1 \Memory_reg[11][12]  (.D(Memory[12]), .CK(n_0_5), .Q(\Memory[11] [12]), 
      .QN());
   DFF_X1 \Memory_reg[11][11]  (.D(Memory[11]), .CK(n_0_5), .Q(\Memory[11] [11]), 
      .QN());
   DFF_X1 \Memory_reg[11][10]  (.D(Memory[10]), .CK(n_0_5), .Q(\Memory[11] [10]), 
      .QN());
   DFF_X1 \Memory_reg[11][9]  (.D(Memory[9]), .CK(n_0_5), .Q(\Memory[11] [9]), 
      .QN());
   DFF_X1 \Memory_reg[11][8]  (.D(Memory[8]), .CK(n_0_5), .Q(\Memory[11] [8]), 
      .QN());
   DFF_X1 \Memory_reg[11][7]  (.D(Memory[7]), .CK(n_0_5), .Q(\Memory[11] [7]), 
      .QN());
   DFF_X1 \Memory_reg[11][6]  (.D(Memory[6]), .CK(n_0_5), .Q(\Memory[11] [6]), 
      .QN());
   DFF_X1 \Memory_reg[11][5]  (.D(Memory[5]), .CK(n_0_5), .Q(\Memory[11] [5]), 
      .QN());
   DFF_X1 \Memory_reg[11][4]  (.D(Memory[4]), .CK(n_0_5), .Q(\Memory[11] [4]), 
      .QN());
   DFF_X1 \Memory_reg[11][3]  (.D(Memory[3]), .CK(n_0_5), .Q(\Memory[11] [3]), 
      .QN());
   DFF_X1 \Memory_reg[11][2]  (.D(Memory[2]), .CK(n_0_5), .Q(\Memory[11] [2]), 
      .QN());
   DFF_X1 \Memory_reg[11][1]  (.D(Memory[1]), .CK(n_0_5), .Q(\Memory[11] [1]), 
      .QN());
   DFF_X1 \Memory_reg[11][0]  (.D(Memory[0]), .CK(n_0_5), .Q(\Memory[11] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[10]_reg  (.CK(CLK), .E(n_0_27), .SE(1'b0), 
      .GCK(n_0_6));
   DFF_X1 \Memory_reg[10][63]  (.D(Memory[63]), .CK(n_0_6), .Q(\Memory[10] [63]), 
      .QN());
   DFF_X1 \Memory_reg[10][62]  (.D(Memory[62]), .CK(n_0_6), .Q(\Memory[10] [62]), 
      .QN());
   DFF_X1 \Memory_reg[10][61]  (.D(Memory[61]), .CK(n_0_6), .Q(\Memory[10] [61]), 
      .QN());
   DFF_X1 \Memory_reg[10][60]  (.D(Memory[60]), .CK(n_0_6), .Q(\Memory[10] [60]), 
      .QN());
   DFF_X1 \Memory_reg[10][59]  (.D(Memory[59]), .CK(n_0_6), .Q(\Memory[10] [59]), 
      .QN());
   DFF_X1 \Memory_reg[10][58]  (.D(Memory[58]), .CK(n_0_6), .Q(\Memory[10] [58]), 
      .QN());
   DFF_X1 \Memory_reg[10][57]  (.D(Memory[57]), .CK(n_0_6), .Q(\Memory[10] [57]), 
      .QN());
   DFF_X1 \Memory_reg[10][56]  (.D(Memory[56]), .CK(n_0_6), .Q(\Memory[10] [56]), 
      .QN());
   DFF_X1 \Memory_reg[10][55]  (.D(Memory[55]), .CK(n_0_6), .Q(\Memory[10] [55]), 
      .QN());
   DFF_X1 \Memory_reg[10][54]  (.D(Memory[54]), .CK(n_0_6), .Q(\Memory[10] [54]), 
      .QN());
   DFF_X1 \Memory_reg[10][53]  (.D(Memory[53]), .CK(n_0_6), .Q(\Memory[10] [53]), 
      .QN());
   DFF_X1 \Memory_reg[10][52]  (.D(Memory[52]), .CK(n_0_6), .Q(\Memory[10] [52]), 
      .QN());
   DFF_X1 \Memory_reg[10][51]  (.D(Memory[51]), .CK(n_0_6), .Q(\Memory[10] [51]), 
      .QN());
   DFF_X1 \Memory_reg[10][50]  (.D(Memory[50]), .CK(n_0_6), .Q(\Memory[10] [50]), 
      .QN());
   DFF_X1 \Memory_reg[10][49]  (.D(Memory[49]), .CK(n_0_6), .Q(\Memory[10] [49]), 
      .QN());
   DFF_X1 \Memory_reg[10][48]  (.D(Memory[48]), .CK(n_0_6), .Q(\Memory[10] [48]), 
      .QN());
   DFF_X1 \Memory_reg[10][47]  (.D(Memory[47]), .CK(n_0_6), .Q(\Memory[10] [47]), 
      .QN());
   DFF_X1 \Memory_reg[10][46]  (.D(Memory[46]), .CK(n_0_6), .Q(\Memory[10] [46]), 
      .QN());
   DFF_X1 \Memory_reg[10][45]  (.D(Memory[45]), .CK(n_0_6), .Q(\Memory[10] [45]), 
      .QN());
   DFF_X1 \Memory_reg[10][44]  (.D(Memory[44]), .CK(n_0_6), .Q(\Memory[10] [44]), 
      .QN());
   DFF_X1 \Memory_reg[10][43]  (.D(Memory[43]), .CK(n_0_6), .Q(\Memory[10] [43]), 
      .QN());
   DFF_X1 \Memory_reg[10][42]  (.D(Memory[42]), .CK(n_0_6), .Q(\Memory[10] [42]), 
      .QN());
   DFF_X1 \Memory_reg[10][41]  (.D(Memory[41]), .CK(n_0_6), .Q(\Memory[10] [41]), 
      .QN());
   DFF_X1 \Memory_reg[10][40]  (.D(Memory[40]), .CK(n_0_6), .Q(\Memory[10] [40]), 
      .QN());
   DFF_X1 \Memory_reg[10][39]  (.D(Memory[39]), .CK(n_0_6), .Q(\Memory[10] [39]), 
      .QN());
   DFF_X1 \Memory_reg[10][38]  (.D(Memory[38]), .CK(n_0_6), .Q(\Memory[10] [38]), 
      .QN());
   DFF_X1 \Memory_reg[10][37]  (.D(Memory[37]), .CK(n_0_6), .Q(\Memory[10] [37]), 
      .QN());
   DFF_X1 \Memory_reg[10][36]  (.D(Memory[36]), .CK(n_0_6), .Q(\Memory[10] [36]), 
      .QN());
   DFF_X1 \Memory_reg[10][35]  (.D(Memory[35]), .CK(n_0_6), .Q(\Memory[10] [35]), 
      .QN());
   DFF_X1 \Memory_reg[10][34]  (.D(Memory[34]), .CK(n_0_6), .Q(\Memory[10] [34]), 
      .QN());
   DFF_X1 \Memory_reg[10][33]  (.D(Memory[33]), .CK(n_0_6), .Q(\Memory[10] [33]), 
      .QN());
   DFF_X1 \Memory_reg[10][32]  (.D(Memory[32]), .CK(n_0_6), .Q(\Memory[10] [32]), 
      .QN());
   DFF_X1 \Memory_reg[10][31]  (.D(Memory[31]), .CK(n_0_6), .Q(\Memory[10] [31]), 
      .QN());
   DFF_X1 \Memory_reg[10][30]  (.D(Memory[30]), .CK(n_0_6), .Q(\Memory[10] [30]), 
      .QN());
   DFF_X1 \Memory_reg[10][29]  (.D(Memory[29]), .CK(n_0_6), .Q(\Memory[10] [29]), 
      .QN());
   DFF_X1 \Memory_reg[10][28]  (.D(Memory[28]), .CK(n_0_6), .Q(\Memory[10] [28]), 
      .QN());
   DFF_X1 \Memory_reg[10][27]  (.D(Memory[27]), .CK(n_0_6), .Q(\Memory[10] [27]), 
      .QN());
   DFF_X1 \Memory_reg[10][26]  (.D(Memory[26]), .CK(n_0_6), .Q(\Memory[10] [26]), 
      .QN());
   DFF_X1 \Memory_reg[10][25]  (.D(Memory[25]), .CK(n_0_6), .Q(\Memory[10] [25]), 
      .QN());
   DFF_X1 \Memory_reg[10][24]  (.D(Memory[24]), .CK(n_0_6), .Q(\Memory[10] [24]), 
      .QN());
   DFF_X1 \Memory_reg[10][23]  (.D(Memory[23]), .CK(n_0_6), .Q(\Memory[10] [23]), 
      .QN());
   DFF_X1 \Memory_reg[10][22]  (.D(Memory[22]), .CK(n_0_6), .Q(\Memory[10] [22]), 
      .QN());
   DFF_X1 \Memory_reg[10][21]  (.D(Memory[21]), .CK(n_0_6), .Q(\Memory[10] [21]), 
      .QN());
   DFF_X1 \Memory_reg[10][20]  (.D(Memory[20]), .CK(n_0_6), .Q(\Memory[10] [20]), 
      .QN());
   DFF_X1 \Memory_reg[10][19]  (.D(Memory[19]), .CK(n_0_6), .Q(\Memory[10] [19]), 
      .QN());
   DFF_X1 \Memory_reg[10][18]  (.D(Memory[18]), .CK(n_0_6), .Q(\Memory[10] [18]), 
      .QN());
   DFF_X1 \Memory_reg[10][17]  (.D(Memory[17]), .CK(n_0_6), .Q(\Memory[10] [17]), 
      .QN());
   DFF_X1 \Memory_reg[10][16]  (.D(Memory[16]), .CK(n_0_6), .Q(\Memory[10] [16]), 
      .QN());
   DFF_X1 \Memory_reg[10][15]  (.D(Memory[15]), .CK(n_0_6), .Q(\Memory[10] [15]), 
      .QN());
   DFF_X1 \Memory_reg[10][14]  (.D(Memory[14]), .CK(n_0_6), .Q(\Memory[10] [14]), 
      .QN());
   DFF_X1 \Memory_reg[10][13]  (.D(Memory[13]), .CK(n_0_6), .Q(\Memory[10] [13]), 
      .QN());
   DFF_X1 \Memory_reg[10][12]  (.D(Memory[12]), .CK(n_0_6), .Q(\Memory[10] [12]), 
      .QN());
   DFF_X1 \Memory_reg[10][11]  (.D(Memory[11]), .CK(n_0_6), .Q(\Memory[10] [11]), 
      .QN());
   DFF_X1 \Memory_reg[10][10]  (.D(Memory[10]), .CK(n_0_6), .Q(\Memory[10] [10]), 
      .QN());
   DFF_X1 \Memory_reg[10][9]  (.D(Memory[9]), .CK(n_0_6), .Q(\Memory[10] [9]), 
      .QN());
   DFF_X1 \Memory_reg[10][8]  (.D(Memory[8]), .CK(n_0_6), .Q(\Memory[10] [8]), 
      .QN());
   DFF_X1 \Memory_reg[10][7]  (.D(Memory[7]), .CK(n_0_6), .Q(\Memory[10] [7]), 
      .QN());
   DFF_X1 \Memory_reg[10][6]  (.D(Memory[6]), .CK(n_0_6), .Q(\Memory[10] [6]), 
      .QN());
   DFF_X1 \Memory_reg[10][5]  (.D(Memory[5]), .CK(n_0_6), .Q(\Memory[10] [5]), 
      .QN());
   DFF_X1 \Memory_reg[10][4]  (.D(Memory[4]), .CK(n_0_6), .Q(\Memory[10] [4]), 
      .QN());
   DFF_X1 \Memory_reg[10][3]  (.D(Memory[3]), .CK(n_0_6), .Q(\Memory[10] [3]), 
      .QN());
   DFF_X1 \Memory_reg[10][2]  (.D(Memory[2]), .CK(n_0_6), .Q(\Memory[10] [2]), 
      .QN());
   DFF_X1 \Memory_reg[10][1]  (.D(Memory[1]), .CK(n_0_6), .Q(\Memory[10] [1]), 
      .QN());
   DFF_X1 \Memory_reg[10][0]  (.D(Memory[0]), .CK(n_0_6), .Q(\Memory[10] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[9]_reg  (.CK(CLK), .E(n_0_26), .SE(1'b0), 
      .GCK(n_0_7));
   DFF_X1 \Memory_reg[9][63]  (.D(Memory[63]), .CK(n_0_7), .Q(\Memory[9] [63]), 
      .QN());
   DFF_X1 \Memory_reg[9][62]  (.D(Memory[62]), .CK(n_0_7), .Q(\Memory[9] [62]), 
      .QN());
   DFF_X1 \Memory_reg[9][61]  (.D(Memory[61]), .CK(n_0_7), .Q(\Memory[9] [61]), 
      .QN());
   DFF_X1 \Memory_reg[9][60]  (.D(Memory[60]), .CK(n_0_7), .Q(\Memory[9] [60]), 
      .QN());
   DFF_X1 \Memory_reg[9][59]  (.D(Memory[59]), .CK(n_0_7), .Q(\Memory[9] [59]), 
      .QN());
   DFF_X1 \Memory_reg[9][58]  (.D(Memory[58]), .CK(n_0_7), .Q(\Memory[9] [58]), 
      .QN());
   DFF_X1 \Memory_reg[9][57]  (.D(Memory[57]), .CK(n_0_7), .Q(\Memory[9] [57]), 
      .QN());
   DFF_X1 \Memory_reg[9][56]  (.D(Memory[56]), .CK(n_0_7), .Q(\Memory[9] [56]), 
      .QN());
   DFF_X1 \Memory_reg[9][55]  (.D(Memory[55]), .CK(n_0_7), .Q(\Memory[9] [55]), 
      .QN());
   DFF_X1 \Memory_reg[9][54]  (.D(Memory[54]), .CK(n_0_7), .Q(\Memory[9] [54]), 
      .QN());
   DFF_X1 \Memory_reg[9][53]  (.D(Memory[53]), .CK(n_0_7), .Q(\Memory[9] [53]), 
      .QN());
   DFF_X1 \Memory_reg[9][52]  (.D(Memory[52]), .CK(n_0_7), .Q(\Memory[9] [52]), 
      .QN());
   DFF_X1 \Memory_reg[9][51]  (.D(Memory[51]), .CK(n_0_7), .Q(\Memory[9] [51]), 
      .QN());
   DFF_X1 \Memory_reg[9][50]  (.D(Memory[50]), .CK(n_0_7), .Q(\Memory[9] [50]), 
      .QN());
   DFF_X1 \Memory_reg[9][49]  (.D(Memory[49]), .CK(n_0_7), .Q(\Memory[9] [49]), 
      .QN());
   DFF_X1 \Memory_reg[9][48]  (.D(Memory[48]), .CK(n_0_7), .Q(\Memory[9] [48]), 
      .QN());
   DFF_X1 \Memory_reg[9][47]  (.D(Memory[47]), .CK(n_0_7), .Q(\Memory[9] [47]), 
      .QN());
   DFF_X1 \Memory_reg[9][46]  (.D(Memory[46]), .CK(n_0_7), .Q(\Memory[9] [46]), 
      .QN());
   DFF_X1 \Memory_reg[9][45]  (.D(Memory[45]), .CK(n_0_7), .Q(\Memory[9] [45]), 
      .QN());
   DFF_X1 \Memory_reg[9][44]  (.D(Memory[44]), .CK(n_0_7), .Q(\Memory[9] [44]), 
      .QN());
   DFF_X1 \Memory_reg[9][43]  (.D(Memory[43]), .CK(n_0_7), .Q(\Memory[9] [43]), 
      .QN());
   DFF_X1 \Memory_reg[9][42]  (.D(Memory[42]), .CK(n_0_7), .Q(\Memory[9] [42]), 
      .QN());
   DFF_X1 \Memory_reg[9][41]  (.D(Memory[41]), .CK(n_0_7), .Q(\Memory[9] [41]), 
      .QN());
   DFF_X1 \Memory_reg[9][40]  (.D(Memory[40]), .CK(n_0_7), .Q(\Memory[9] [40]), 
      .QN());
   DFF_X1 \Memory_reg[9][39]  (.D(Memory[39]), .CK(n_0_7), .Q(\Memory[9] [39]), 
      .QN());
   DFF_X1 \Memory_reg[9][38]  (.D(Memory[38]), .CK(n_0_7), .Q(\Memory[9] [38]), 
      .QN());
   DFF_X1 \Memory_reg[9][37]  (.D(Memory[37]), .CK(n_0_7), .Q(\Memory[9] [37]), 
      .QN());
   DFF_X1 \Memory_reg[9][36]  (.D(Memory[36]), .CK(n_0_7), .Q(\Memory[9] [36]), 
      .QN());
   DFF_X1 \Memory_reg[9][35]  (.D(Memory[35]), .CK(n_0_7), .Q(\Memory[9] [35]), 
      .QN());
   DFF_X1 \Memory_reg[9][34]  (.D(Memory[34]), .CK(n_0_7), .Q(\Memory[9] [34]), 
      .QN());
   DFF_X1 \Memory_reg[9][33]  (.D(Memory[33]), .CK(n_0_7), .Q(\Memory[9] [33]), 
      .QN());
   DFF_X1 \Memory_reg[9][32]  (.D(Memory[32]), .CK(n_0_7), .Q(\Memory[9] [32]), 
      .QN());
   DFF_X1 \Memory_reg[9][31]  (.D(Memory[31]), .CK(n_0_7), .Q(\Memory[9] [31]), 
      .QN());
   DFF_X1 \Memory_reg[9][30]  (.D(Memory[30]), .CK(n_0_7), .Q(\Memory[9] [30]), 
      .QN());
   DFF_X1 \Memory_reg[9][29]  (.D(Memory[29]), .CK(n_0_7), .Q(\Memory[9] [29]), 
      .QN());
   DFF_X1 \Memory_reg[9][28]  (.D(Memory[28]), .CK(n_0_7), .Q(\Memory[9] [28]), 
      .QN());
   DFF_X1 \Memory_reg[9][27]  (.D(Memory[27]), .CK(n_0_7), .Q(\Memory[9] [27]), 
      .QN());
   DFF_X1 \Memory_reg[9][26]  (.D(Memory[26]), .CK(n_0_7), .Q(\Memory[9] [26]), 
      .QN());
   DFF_X1 \Memory_reg[9][25]  (.D(Memory[25]), .CK(n_0_7), .Q(\Memory[9] [25]), 
      .QN());
   DFF_X1 \Memory_reg[9][24]  (.D(Memory[24]), .CK(n_0_7), .Q(\Memory[9] [24]), 
      .QN());
   DFF_X1 \Memory_reg[9][23]  (.D(Memory[23]), .CK(n_0_7), .Q(\Memory[9] [23]), 
      .QN());
   DFF_X1 \Memory_reg[9][22]  (.D(Memory[22]), .CK(n_0_7), .Q(\Memory[9] [22]), 
      .QN());
   DFF_X1 \Memory_reg[9][21]  (.D(Memory[21]), .CK(n_0_7), .Q(\Memory[9] [21]), 
      .QN());
   DFF_X1 \Memory_reg[9][20]  (.D(Memory[20]), .CK(n_0_7), .Q(\Memory[9] [20]), 
      .QN());
   DFF_X1 \Memory_reg[9][19]  (.D(Memory[19]), .CK(n_0_7), .Q(\Memory[9] [19]), 
      .QN());
   DFF_X1 \Memory_reg[9][18]  (.D(Memory[18]), .CK(n_0_7), .Q(\Memory[9] [18]), 
      .QN());
   DFF_X1 \Memory_reg[9][17]  (.D(Memory[17]), .CK(n_0_7), .Q(\Memory[9] [17]), 
      .QN());
   DFF_X1 \Memory_reg[9][16]  (.D(Memory[16]), .CK(n_0_7), .Q(\Memory[9] [16]), 
      .QN());
   DFF_X1 \Memory_reg[9][15]  (.D(Memory[15]), .CK(n_0_7), .Q(\Memory[9] [15]), 
      .QN());
   DFF_X1 \Memory_reg[9][14]  (.D(Memory[14]), .CK(n_0_7), .Q(\Memory[9] [14]), 
      .QN());
   DFF_X1 \Memory_reg[9][13]  (.D(Memory[13]), .CK(n_0_7), .Q(\Memory[9] [13]), 
      .QN());
   DFF_X1 \Memory_reg[9][12]  (.D(Memory[12]), .CK(n_0_7), .Q(\Memory[9] [12]), 
      .QN());
   DFF_X1 \Memory_reg[9][11]  (.D(Memory[11]), .CK(n_0_7), .Q(\Memory[9] [11]), 
      .QN());
   DFF_X1 \Memory_reg[9][10]  (.D(Memory[10]), .CK(n_0_7), .Q(\Memory[9] [10]), 
      .QN());
   DFF_X1 \Memory_reg[9][9]  (.D(Memory[9]), .CK(n_0_7), .Q(\Memory[9] [9]), 
      .QN());
   DFF_X1 \Memory_reg[9][8]  (.D(Memory[8]), .CK(n_0_7), .Q(\Memory[9] [8]), 
      .QN());
   DFF_X1 \Memory_reg[9][7]  (.D(Memory[7]), .CK(n_0_7), .Q(\Memory[9] [7]), 
      .QN());
   DFF_X1 \Memory_reg[9][6]  (.D(Memory[6]), .CK(n_0_7), .Q(\Memory[9] [6]), 
      .QN());
   DFF_X1 \Memory_reg[9][5]  (.D(Memory[5]), .CK(n_0_7), .Q(\Memory[9] [5]), 
      .QN());
   DFF_X1 \Memory_reg[9][4]  (.D(Memory[4]), .CK(n_0_7), .Q(\Memory[9] [4]), 
      .QN());
   DFF_X1 \Memory_reg[9][3]  (.D(Memory[3]), .CK(n_0_7), .Q(\Memory[9] [3]), 
      .QN());
   DFF_X1 \Memory_reg[9][2]  (.D(Memory[2]), .CK(n_0_7), .Q(\Memory[9] [2]), 
      .QN());
   DFF_X1 \Memory_reg[9][1]  (.D(Memory[1]), .CK(n_0_7), .Q(\Memory[9] [1]), 
      .QN());
   DFF_X1 \Memory_reg[9][0]  (.D(Memory[0]), .CK(n_0_7), .Q(\Memory[9] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[8]_reg  (.CK(CLK), .E(n_0_25), .SE(1'b0), 
      .GCK(n_0_8));
   DFF_X1 \Memory_reg[8][63]  (.D(Memory[63]), .CK(n_0_8), .Q(\Memory[8] [63]), 
      .QN());
   DFF_X1 \Memory_reg[8][62]  (.D(Memory[62]), .CK(n_0_8), .Q(\Memory[8] [62]), 
      .QN());
   DFF_X1 \Memory_reg[8][61]  (.D(Memory[61]), .CK(n_0_8), .Q(\Memory[8] [61]), 
      .QN());
   DFF_X1 \Memory_reg[8][60]  (.D(Memory[60]), .CK(n_0_8), .Q(\Memory[8] [60]), 
      .QN());
   DFF_X1 \Memory_reg[8][59]  (.D(Memory[59]), .CK(n_0_8), .Q(\Memory[8] [59]), 
      .QN());
   DFF_X1 \Memory_reg[8][58]  (.D(Memory[58]), .CK(n_0_8), .Q(\Memory[8] [58]), 
      .QN());
   DFF_X1 \Memory_reg[8][57]  (.D(Memory[57]), .CK(n_0_8), .Q(\Memory[8] [57]), 
      .QN());
   DFF_X1 \Memory_reg[8][56]  (.D(Memory[56]), .CK(n_0_8), .Q(\Memory[8] [56]), 
      .QN());
   DFF_X1 \Memory_reg[8][55]  (.D(Memory[55]), .CK(n_0_8), .Q(\Memory[8] [55]), 
      .QN());
   DFF_X1 \Memory_reg[8][54]  (.D(Memory[54]), .CK(n_0_8), .Q(\Memory[8] [54]), 
      .QN());
   DFF_X1 \Memory_reg[8][53]  (.D(Memory[53]), .CK(n_0_8), .Q(\Memory[8] [53]), 
      .QN());
   DFF_X1 \Memory_reg[8][52]  (.D(Memory[52]), .CK(n_0_8), .Q(\Memory[8] [52]), 
      .QN());
   DFF_X1 \Memory_reg[8][51]  (.D(Memory[51]), .CK(n_0_8), .Q(\Memory[8] [51]), 
      .QN());
   DFF_X1 \Memory_reg[8][50]  (.D(Memory[50]), .CK(n_0_8), .Q(\Memory[8] [50]), 
      .QN());
   DFF_X1 \Memory_reg[8][49]  (.D(Memory[49]), .CK(n_0_8), .Q(\Memory[8] [49]), 
      .QN());
   DFF_X1 \Memory_reg[8][48]  (.D(Memory[48]), .CK(n_0_8), .Q(\Memory[8] [48]), 
      .QN());
   DFF_X1 \Memory_reg[8][47]  (.D(Memory[47]), .CK(n_0_8), .Q(\Memory[8] [47]), 
      .QN());
   DFF_X1 \Memory_reg[8][46]  (.D(Memory[46]), .CK(n_0_8), .Q(\Memory[8] [46]), 
      .QN());
   DFF_X1 \Memory_reg[8][45]  (.D(Memory[45]), .CK(n_0_8), .Q(\Memory[8] [45]), 
      .QN());
   DFF_X1 \Memory_reg[8][44]  (.D(Memory[44]), .CK(n_0_8), .Q(\Memory[8] [44]), 
      .QN());
   DFF_X1 \Memory_reg[8][43]  (.D(Memory[43]), .CK(n_0_8), .Q(\Memory[8] [43]), 
      .QN());
   DFF_X1 \Memory_reg[8][42]  (.D(Memory[42]), .CK(n_0_8), .Q(\Memory[8] [42]), 
      .QN());
   DFF_X1 \Memory_reg[8][41]  (.D(Memory[41]), .CK(n_0_8), .Q(\Memory[8] [41]), 
      .QN());
   DFF_X1 \Memory_reg[8][40]  (.D(Memory[40]), .CK(n_0_8), .Q(\Memory[8] [40]), 
      .QN());
   DFF_X1 \Memory_reg[8][39]  (.D(Memory[39]), .CK(n_0_8), .Q(\Memory[8] [39]), 
      .QN());
   DFF_X1 \Memory_reg[8][38]  (.D(Memory[38]), .CK(n_0_8), .Q(\Memory[8] [38]), 
      .QN());
   DFF_X1 \Memory_reg[8][37]  (.D(Memory[37]), .CK(n_0_8), .Q(\Memory[8] [37]), 
      .QN());
   DFF_X1 \Memory_reg[8][36]  (.D(Memory[36]), .CK(n_0_8), .Q(\Memory[8] [36]), 
      .QN());
   DFF_X1 \Memory_reg[8][35]  (.D(Memory[35]), .CK(n_0_8), .Q(\Memory[8] [35]), 
      .QN());
   DFF_X1 \Memory_reg[8][34]  (.D(Memory[34]), .CK(n_0_8), .Q(\Memory[8] [34]), 
      .QN());
   DFF_X1 \Memory_reg[8][33]  (.D(Memory[33]), .CK(n_0_8), .Q(\Memory[8] [33]), 
      .QN());
   DFF_X1 \Memory_reg[8][32]  (.D(Memory[32]), .CK(n_0_8), .Q(\Memory[8] [32]), 
      .QN());
   DFF_X1 \Memory_reg[8][31]  (.D(Memory[31]), .CK(n_0_8), .Q(\Memory[8] [31]), 
      .QN());
   DFF_X1 \Memory_reg[8][30]  (.D(Memory[30]), .CK(n_0_8), .Q(\Memory[8] [30]), 
      .QN());
   DFF_X1 \Memory_reg[8][29]  (.D(Memory[29]), .CK(n_0_8), .Q(\Memory[8] [29]), 
      .QN());
   DFF_X1 \Memory_reg[8][28]  (.D(Memory[28]), .CK(n_0_8), .Q(\Memory[8] [28]), 
      .QN());
   DFF_X1 \Memory_reg[8][27]  (.D(Memory[27]), .CK(n_0_8), .Q(\Memory[8] [27]), 
      .QN());
   DFF_X1 \Memory_reg[8][26]  (.D(Memory[26]), .CK(n_0_8), .Q(\Memory[8] [26]), 
      .QN());
   DFF_X1 \Memory_reg[8][25]  (.D(Memory[25]), .CK(n_0_8), .Q(\Memory[8] [25]), 
      .QN());
   DFF_X1 \Memory_reg[8][24]  (.D(Memory[24]), .CK(n_0_8), .Q(\Memory[8] [24]), 
      .QN());
   DFF_X1 \Memory_reg[8][23]  (.D(Memory[23]), .CK(n_0_8), .Q(\Memory[8] [23]), 
      .QN());
   DFF_X1 \Memory_reg[8][22]  (.D(Memory[22]), .CK(n_0_8), .Q(\Memory[8] [22]), 
      .QN());
   DFF_X1 \Memory_reg[8][21]  (.D(Memory[21]), .CK(n_0_8), .Q(\Memory[8] [21]), 
      .QN());
   DFF_X1 \Memory_reg[8][20]  (.D(Memory[20]), .CK(n_0_8), .Q(\Memory[8] [20]), 
      .QN());
   DFF_X1 \Memory_reg[8][19]  (.D(Memory[19]), .CK(n_0_8), .Q(\Memory[8] [19]), 
      .QN());
   DFF_X1 \Memory_reg[8][18]  (.D(Memory[18]), .CK(n_0_8), .Q(\Memory[8] [18]), 
      .QN());
   DFF_X1 \Memory_reg[8][17]  (.D(Memory[17]), .CK(n_0_8), .Q(\Memory[8] [17]), 
      .QN());
   DFF_X1 \Memory_reg[8][16]  (.D(Memory[16]), .CK(n_0_8), .Q(\Memory[8] [16]), 
      .QN());
   DFF_X1 \Memory_reg[8][15]  (.D(Memory[15]), .CK(n_0_8), .Q(\Memory[8] [15]), 
      .QN());
   DFF_X1 \Memory_reg[8][14]  (.D(Memory[14]), .CK(n_0_8), .Q(\Memory[8] [14]), 
      .QN());
   DFF_X1 \Memory_reg[8][13]  (.D(Memory[13]), .CK(n_0_8), .Q(\Memory[8] [13]), 
      .QN());
   DFF_X1 \Memory_reg[8][12]  (.D(Memory[12]), .CK(n_0_8), .Q(\Memory[8] [12]), 
      .QN());
   DFF_X1 \Memory_reg[8][11]  (.D(Memory[11]), .CK(n_0_8), .Q(\Memory[8] [11]), 
      .QN());
   DFF_X1 \Memory_reg[8][10]  (.D(Memory[10]), .CK(n_0_8), .Q(\Memory[8] [10]), 
      .QN());
   DFF_X1 \Memory_reg[8][9]  (.D(Memory[9]), .CK(n_0_8), .Q(\Memory[8] [9]), 
      .QN());
   DFF_X1 \Memory_reg[8][8]  (.D(Memory[8]), .CK(n_0_8), .Q(\Memory[8] [8]), 
      .QN());
   DFF_X1 \Memory_reg[8][7]  (.D(Memory[7]), .CK(n_0_8), .Q(\Memory[8] [7]), 
      .QN());
   DFF_X1 \Memory_reg[8][6]  (.D(Memory[6]), .CK(n_0_8), .Q(\Memory[8] [6]), 
      .QN());
   DFF_X1 \Memory_reg[8][5]  (.D(Memory[5]), .CK(n_0_8), .Q(\Memory[8] [5]), 
      .QN());
   DFF_X1 \Memory_reg[8][4]  (.D(Memory[4]), .CK(n_0_8), .Q(\Memory[8] [4]), 
      .QN());
   DFF_X1 \Memory_reg[8][3]  (.D(Memory[3]), .CK(n_0_8), .Q(\Memory[8] [3]), 
      .QN());
   DFF_X1 \Memory_reg[8][2]  (.D(Memory[2]), .CK(n_0_8), .Q(\Memory[8] [2]), 
      .QN());
   DFF_X1 \Memory_reg[8][1]  (.D(Memory[1]), .CK(n_0_8), .Q(\Memory[8] [1]), 
      .QN());
   DFF_X1 \Memory_reg[8][0]  (.D(Memory[0]), .CK(n_0_8), .Q(\Memory[8] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[7]_reg  (.CK(CLK), .E(n_0_24), .SE(1'b0), 
      .GCK(n_0_9));
   DFF_X1 \Memory_reg[7][63]  (.D(Memory[63]), .CK(n_0_9), .Q(\Memory[7] [63]), 
      .QN());
   DFF_X1 \Memory_reg[7][62]  (.D(Memory[62]), .CK(n_0_9), .Q(\Memory[7] [62]), 
      .QN());
   DFF_X1 \Memory_reg[7][61]  (.D(Memory[61]), .CK(n_0_9), .Q(\Memory[7] [61]), 
      .QN());
   DFF_X1 \Memory_reg[7][60]  (.D(Memory[60]), .CK(n_0_9), .Q(\Memory[7] [60]), 
      .QN());
   DFF_X1 \Memory_reg[7][59]  (.D(Memory[59]), .CK(n_0_9), .Q(\Memory[7] [59]), 
      .QN());
   DFF_X1 \Memory_reg[7][58]  (.D(Memory[58]), .CK(n_0_9), .Q(\Memory[7] [58]), 
      .QN());
   DFF_X1 \Memory_reg[7][57]  (.D(Memory[57]), .CK(n_0_9), .Q(\Memory[7] [57]), 
      .QN());
   DFF_X1 \Memory_reg[7][56]  (.D(Memory[56]), .CK(n_0_9), .Q(\Memory[7] [56]), 
      .QN());
   DFF_X1 \Memory_reg[7][55]  (.D(Memory[55]), .CK(n_0_9), .Q(\Memory[7] [55]), 
      .QN());
   DFF_X1 \Memory_reg[7][54]  (.D(Memory[54]), .CK(n_0_9), .Q(\Memory[7] [54]), 
      .QN());
   DFF_X1 \Memory_reg[7][53]  (.D(Memory[53]), .CK(n_0_9), .Q(\Memory[7] [53]), 
      .QN());
   DFF_X1 \Memory_reg[7][52]  (.D(Memory[52]), .CK(n_0_9), .Q(\Memory[7] [52]), 
      .QN());
   DFF_X1 \Memory_reg[7][51]  (.D(Memory[51]), .CK(n_0_9), .Q(\Memory[7] [51]), 
      .QN());
   DFF_X1 \Memory_reg[7][50]  (.D(Memory[50]), .CK(n_0_9), .Q(\Memory[7] [50]), 
      .QN());
   DFF_X1 \Memory_reg[7][49]  (.D(Memory[49]), .CK(n_0_9), .Q(\Memory[7] [49]), 
      .QN());
   DFF_X1 \Memory_reg[7][48]  (.D(Memory[48]), .CK(n_0_9), .Q(\Memory[7] [48]), 
      .QN());
   DFF_X1 \Memory_reg[7][47]  (.D(Memory[47]), .CK(n_0_9), .Q(\Memory[7] [47]), 
      .QN());
   DFF_X1 \Memory_reg[7][46]  (.D(Memory[46]), .CK(n_0_9), .Q(\Memory[7] [46]), 
      .QN());
   DFF_X1 \Memory_reg[7][45]  (.D(Memory[45]), .CK(n_0_9), .Q(\Memory[7] [45]), 
      .QN());
   DFF_X1 \Memory_reg[7][44]  (.D(Memory[44]), .CK(n_0_9), .Q(\Memory[7] [44]), 
      .QN());
   DFF_X1 \Memory_reg[7][43]  (.D(Memory[43]), .CK(n_0_9), .Q(\Memory[7] [43]), 
      .QN());
   DFF_X1 \Memory_reg[7][42]  (.D(Memory[42]), .CK(n_0_9), .Q(\Memory[7] [42]), 
      .QN());
   DFF_X1 \Memory_reg[7][41]  (.D(Memory[41]), .CK(n_0_9), .Q(\Memory[7] [41]), 
      .QN());
   DFF_X1 \Memory_reg[7][40]  (.D(Memory[40]), .CK(n_0_9), .Q(\Memory[7] [40]), 
      .QN());
   DFF_X1 \Memory_reg[7][39]  (.D(Memory[39]), .CK(n_0_9), .Q(\Memory[7] [39]), 
      .QN());
   DFF_X1 \Memory_reg[7][38]  (.D(Memory[38]), .CK(n_0_9), .Q(\Memory[7] [38]), 
      .QN());
   DFF_X1 \Memory_reg[7][37]  (.D(Memory[37]), .CK(n_0_9), .Q(\Memory[7] [37]), 
      .QN());
   DFF_X1 \Memory_reg[7][36]  (.D(Memory[36]), .CK(n_0_9), .Q(\Memory[7] [36]), 
      .QN());
   DFF_X1 \Memory_reg[7][35]  (.D(Memory[35]), .CK(n_0_9), .Q(\Memory[7] [35]), 
      .QN());
   DFF_X1 \Memory_reg[7][34]  (.D(Memory[34]), .CK(n_0_9), .Q(\Memory[7] [34]), 
      .QN());
   DFF_X1 \Memory_reg[7][33]  (.D(Memory[33]), .CK(n_0_9), .Q(\Memory[7] [33]), 
      .QN());
   DFF_X1 \Memory_reg[7][32]  (.D(Memory[32]), .CK(n_0_9), .Q(\Memory[7] [32]), 
      .QN());
   DFF_X1 \Memory_reg[7][31]  (.D(Memory[31]), .CK(n_0_9), .Q(\Memory[7] [31]), 
      .QN());
   DFF_X1 \Memory_reg[7][30]  (.D(Memory[30]), .CK(n_0_9), .Q(\Memory[7] [30]), 
      .QN());
   DFF_X1 \Memory_reg[7][29]  (.D(Memory[29]), .CK(n_0_9), .Q(\Memory[7] [29]), 
      .QN());
   DFF_X1 \Memory_reg[7][28]  (.D(Memory[28]), .CK(n_0_9), .Q(\Memory[7] [28]), 
      .QN());
   DFF_X1 \Memory_reg[7][27]  (.D(Memory[27]), .CK(n_0_9), .Q(\Memory[7] [27]), 
      .QN());
   DFF_X1 \Memory_reg[7][26]  (.D(Memory[26]), .CK(n_0_9), .Q(\Memory[7] [26]), 
      .QN());
   DFF_X1 \Memory_reg[7][25]  (.D(Memory[25]), .CK(n_0_9), .Q(\Memory[7] [25]), 
      .QN());
   DFF_X1 \Memory_reg[7][24]  (.D(Memory[24]), .CK(n_0_9), .Q(\Memory[7] [24]), 
      .QN());
   DFF_X1 \Memory_reg[7][23]  (.D(Memory[23]), .CK(n_0_9), .Q(\Memory[7] [23]), 
      .QN());
   DFF_X1 \Memory_reg[7][22]  (.D(Memory[22]), .CK(n_0_9), .Q(\Memory[7] [22]), 
      .QN());
   DFF_X1 \Memory_reg[7][21]  (.D(Memory[21]), .CK(n_0_9), .Q(\Memory[7] [21]), 
      .QN());
   DFF_X1 \Memory_reg[7][20]  (.D(Memory[20]), .CK(n_0_9), .Q(\Memory[7] [20]), 
      .QN());
   DFF_X1 \Memory_reg[7][19]  (.D(Memory[19]), .CK(n_0_9), .Q(\Memory[7] [19]), 
      .QN());
   DFF_X1 \Memory_reg[7][18]  (.D(Memory[18]), .CK(n_0_9), .Q(\Memory[7] [18]), 
      .QN());
   DFF_X1 \Memory_reg[7][17]  (.D(Memory[17]), .CK(n_0_9), .Q(\Memory[7] [17]), 
      .QN());
   DFF_X1 \Memory_reg[7][16]  (.D(Memory[16]), .CK(n_0_9), .Q(\Memory[7] [16]), 
      .QN());
   DFF_X1 \Memory_reg[7][15]  (.D(Memory[15]), .CK(n_0_9), .Q(\Memory[7] [15]), 
      .QN());
   DFF_X1 \Memory_reg[7][14]  (.D(Memory[14]), .CK(n_0_9), .Q(\Memory[7] [14]), 
      .QN());
   DFF_X1 \Memory_reg[7][13]  (.D(Memory[13]), .CK(n_0_9), .Q(\Memory[7] [13]), 
      .QN());
   DFF_X1 \Memory_reg[7][12]  (.D(Memory[12]), .CK(n_0_9), .Q(\Memory[7] [12]), 
      .QN());
   DFF_X1 \Memory_reg[7][11]  (.D(Memory[11]), .CK(n_0_9), .Q(\Memory[7] [11]), 
      .QN());
   DFF_X1 \Memory_reg[7][10]  (.D(Memory[10]), .CK(n_0_9), .Q(\Memory[7] [10]), 
      .QN());
   DFF_X1 \Memory_reg[7][9]  (.D(Memory[9]), .CK(n_0_9), .Q(\Memory[7] [9]), 
      .QN());
   DFF_X1 \Memory_reg[7][8]  (.D(Memory[8]), .CK(n_0_9), .Q(\Memory[7] [8]), 
      .QN());
   DFF_X1 \Memory_reg[7][7]  (.D(Memory[7]), .CK(n_0_9), .Q(\Memory[7] [7]), 
      .QN());
   DFF_X1 \Memory_reg[7][6]  (.D(Memory[6]), .CK(n_0_9), .Q(\Memory[7] [6]), 
      .QN());
   DFF_X1 \Memory_reg[7][5]  (.D(Memory[5]), .CK(n_0_9), .Q(\Memory[7] [5]), 
      .QN());
   DFF_X1 \Memory_reg[7][4]  (.D(Memory[4]), .CK(n_0_9), .Q(\Memory[7] [4]), 
      .QN());
   DFF_X1 \Memory_reg[7][3]  (.D(Memory[3]), .CK(n_0_9), .Q(\Memory[7] [3]), 
      .QN());
   DFF_X1 \Memory_reg[7][2]  (.D(Memory[2]), .CK(n_0_9), .Q(\Memory[7] [2]), 
      .QN());
   DFF_X1 \Memory_reg[7][1]  (.D(Memory[1]), .CK(n_0_9), .Q(\Memory[7] [1]), 
      .QN());
   DFF_X1 \Memory_reg[7][0]  (.D(Memory[0]), .CK(n_0_9), .Q(\Memory[7] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[6]_reg  (.CK(CLK), .E(n_0_23), .SE(1'b0), 
      .GCK(n_0_10));
   DFF_X1 \Memory_reg[6][63]  (.D(Memory[63]), .CK(n_0_10), .Q(\Memory[6] [63]), 
      .QN());
   DFF_X1 \Memory_reg[6][62]  (.D(Memory[62]), .CK(n_0_10), .Q(\Memory[6] [62]), 
      .QN());
   DFF_X1 \Memory_reg[6][61]  (.D(Memory[61]), .CK(n_0_10), .Q(\Memory[6] [61]), 
      .QN());
   DFF_X1 \Memory_reg[6][60]  (.D(Memory[60]), .CK(n_0_10), .Q(\Memory[6] [60]), 
      .QN());
   DFF_X1 \Memory_reg[6][59]  (.D(Memory[59]), .CK(n_0_10), .Q(\Memory[6] [59]), 
      .QN());
   DFF_X1 \Memory_reg[6][58]  (.D(Memory[58]), .CK(n_0_10), .Q(\Memory[6] [58]), 
      .QN());
   DFF_X1 \Memory_reg[6][57]  (.D(Memory[57]), .CK(n_0_10), .Q(\Memory[6] [57]), 
      .QN());
   DFF_X1 \Memory_reg[6][56]  (.D(Memory[56]), .CK(n_0_10), .Q(\Memory[6] [56]), 
      .QN());
   DFF_X1 \Memory_reg[6][55]  (.D(Memory[55]), .CK(n_0_10), .Q(\Memory[6] [55]), 
      .QN());
   DFF_X1 \Memory_reg[6][54]  (.D(Memory[54]), .CK(n_0_10), .Q(\Memory[6] [54]), 
      .QN());
   DFF_X1 \Memory_reg[6][53]  (.D(Memory[53]), .CK(n_0_10), .Q(\Memory[6] [53]), 
      .QN());
   DFF_X1 \Memory_reg[6][52]  (.D(Memory[52]), .CK(n_0_10), .Q(\Memory[6] [52]), 
      .QN());
   DFF_X1 \Memory_reg[6][51]  (.D(Memory[51]), .CK(n_0_10), .Q(\Memory[6] [51]), 
      .QN());
   DFF_X1 \Memory_reg[6][50]  (.D(Memory[50]), .CK(n_0_10), .Q(\Memory[6] [50]), 
      .QN());
   DFF_X1 \Memory_reg[6][49]  (.D(Memory[49]), .CK(n_0_10), .Q(\Memory[6] [49]), 
      .QN());
   DFF_X1 \Memory_reg[6][48]  (.D(Memory[48]), .CK(n_0_10), .Q(\Memory[6] [48]), 
      .QN());
   DFF_X1 \Memory_reg[6][47]  (.D(Memory[47]), .CK(n_0_10), .Q(\Memory[6] [47]), 
      .QN());
   DFF_X1 \Memory_reg[6][46]  (.D(Memory[46]), .CK(n_0_10), .Q(\Memory[6] [46]), 
      .QN());
   DFF_X1 \Memory_reg[6][45]  (.D(Memory[45]), .CK(n_0_10), .Q(\Memory[6] [45]), 
      .QN());
   DFF_X1 \Memory_reg[6][44]  (.D(Memory[44]), .CK(n_0_10), .Q(\Memory[6] [44]), 
      .QN());
   DFF_X1 \Memory_reg[6][43]  (.D(Memory[43]), .CK(n_0_10), .Q(\Memory[6] [43]), 
      .QN());
   DFF_X1 \Memory_reg[6][42]  (.D(Memory[42]), .CK(n_0_10), .Q(\Memory[6] [42]), 
      .QN());
   DFF_X1 \Memory_reg[6][41]  (.D(Memory[41]), .CK(n_0_10), .Q(\Memory[6] [41]), 
      .QN());
   DFF_X1 \Memory_reg[6][40]  (.D(Memory[40]), .CK(n_0_10), .Q(\Memory[6] [40]), 
      .QN());
   DFF_X1 \Memory_reg[6][39]  (.D(Memory[39]), .CK(n_0_10), .Q(\Memory[6] [39]), 
      .QN());
   DFF_X1 \Memory_reg[6][38]  (.D(Memory[38]), .CK(n_0_10), .Q(\Memory[6] [38]), 
      .QN());
   DFF_X1 \Memory_reg[6][37]  (.D(Memory[37]), .CK(n_0_10), .Q(\Memory[6] [37]), 
      .QN());
   DFF_X1 \Memory_reg[6][36]  (.D(Memory[36]), .CK(n_0_10), .Q(\Memory[6] [36]), 
      .QN());
   DFF_X1 \Memory_reg[6][35]  (.D(Memory[35]), .CK(n_0_10), .Q(\Memory[6] [35]), 
      .QN());
   DFF_X1 \Memory_reg[6][34]  (.D(Memory[34]), .CK(n_0_10), .Q(\Memory[6] [34]), 
      .QN());
   DFF_X1 \Memory_reg[6][33]  (.D(Memory[33]), .CK(n_0_10), .Q(\Memory[6] [33]), 
      .QN());
   DFF_X1 \Memory_reg[6][32]  (.D(Memory[32]), .CK(n_0_10), .Q(\Memory[6] [32]), 
      .QN());
   DFF_X1 \Memory_reg[6][31]  (.D(Memory[31]), .CK(n_0_10), .Q(\Memory[6] [31]), 
      .QN());
   DFF_X1 \Memory_reg[6][30]  (.D(Memory[30]), .CK(n_0_10), .Q(\Memory[6] [30]), 
      .QN());
   DFF_X1 \Memory_reg[6][29]  (.D(Memory[29]), .CK(n_0_10), .Q(\Memory[6] [29]), 
      .QN());
   DFF_X1 \Memory_reg[6][28]  (.D(Memory[28]), .CK(n_0_10), .Q(\Memory[6] [28]), 
      .QN());
   DFF_X1 \Memory_reg[6][27]  (.D(Memory[27]), .CK(n_0_10), .Q(\Memory[6] [27]), 
      .QN());
   DFF_X1 \Memory_reg[6][26]  (.D(Memory[26]), .CK(n_0_10), .Q(\Memory[6] [26]), 
      .QN());
   DFF_X1 \Memory_reg[6][25]  (.D(Memory[25]), .CK(n_0_10), .Q(\Memory[6] [25]), 
      .QN());
   DFF_X1 \Memory_reg[6][24]  (.D(Memory[24]), .CK(n_0_10), .Q(\Memory[6] [24]), 
      .QN());
   DFF_X1 \Memory_reg[6][23]  (.D(Memory[23]), .CK(n_0_10), .Q(\Memory[6] [23]), 
      .QN());
   DFF_X1 \Memory_reg[6][22]  (.D(Memory[22]), .CK(n_0_10), .Q(\Memory[6] [22]), 
      .QN());
   DFF_X1 \Memory_reg[6][21]  (.D(Memory[21]), .CK(n_0_10), .Q(\Memory[6] [21]), 
      .QN());
   DFF_X1 \Memory_reg[6][20]  (.D(Memory[20]), .CK(n_0_10), .Q(\Memory[6] [20]), 
      .QN());
   DFF_X1 \Memory_reg[6][19]  (.D(Memory[19]), .CK(n_0_10), .Q(\Memory[6] [19]), 
      .QN());
   DFF_X1 \Memory_reg[6][18]  (.D(Memory[18]), .CK(n_0_10), .Q(\Memory[6] [18]), 
      .QN());
   DFF_X1 \Memory_reg[6][17]  (.D(Memory[17]), .CK(n_0_10), .Q(\Memory[6] [17]), 
      .QN());
   DFF_X1 \Memory_reg[6][16]  (.D(Memory[16]), .CK(n_0_10), .Q(\Memory[6] [16]), 
      .QN());
   DFF_X1 \Memory_reg[6][15]  (.D(Memory[15]), .CK(n_0_10), .Q(\Memory[6] [15]), 
      .QN());
   DFF_X1 \Memory_reg[6][14]  (.D(Memory[14]), .CK(n_0_10), .Q(\Memory[6] [14]), 
      .QN());
   DFF_X1 \Memory_reg[6][13]  (.D(Memory[13]), .CK(n_0_10), .Q(\Memory[6] [13]), 
      .QN());
   DFF_X1 \Memory_reg[6][12]  (.D(Memory[12]), .CK(n_0_10), .Q(\Memory[6] [12]), 
      .QN());
   DFF_X1 \Memory_reg[6][11]  (.D(Memory[11]), .CK(n_0_10), .Q(\Memory[6] [11]), 
      .QN());
   DFF_X1 \Memory_reg[6][10]  (.D(Memory[10]), .CK(n_0_10), .Q(\Memory[6] [10]), 
      .QN());
   DFF_X1 \Memory_reg[6][9]  (.D(Memory[9]), .CK(n_0_10), .Q(\Memory[6] [9]), 
      .QN());
   DFF_X1 \Memory_reg[6][8]  (.D(Memory[8]), .CK(n_0_10), .Q(\Memory[6] [8]), 
      .QN());
   DFF_X1 \Memory_reg[6][7]  (.D(Memory[7]), .CK(n_0_10), .Q(\Memory[6] [7]), 
      .QN());
   DFF_X1 \Memory_reg[6][6]  (.D(Memory[6]), .CK(n_0_10), .Q(\Memory[6] [6]), 
      .QN());
   DFF_X1 \Memory_reg[6][5]  (.D(Memory[5]), .CK(n_0_10), .Q(\Memory[6] [5]), 
      .QN());
   DFF_X1 \Memory_reg[6][4]  (.D(Memory[4]), .CK(n_0_10), .Q(\Memory[6] [4]), 
      .QN());
   DFF_X1 \Memory_reg[6][3]  (.D(Memory[3]), .CK(n_0_10), .Q(\Memory[6] [3]), 
      .QN());
   DFF_X1 \Memory_reg[6][2]  (.D(Memory[2]), .CK(n_0_10), .Q(\Memory[6] [2]), 
      .QN());
   DFF_X1 \Memory_reg[6][1]  (.D(Memory[1]), .CK(n_0_10), .Q(\Memory[6] [1]), 
      .QN());
   DFF_X1 \Memory_reg[6][0]  (.D(Memory[0]), .CK(n_0_10), .Q(\Memory[6] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[5]_reg  (.CK(CLK), .E(n_0_22), .SE(1'b0), 
      .GCK(n_0_11));
   DFF_X1 \Memory_reg[5][63]  (.D(Memory[63]), .CK(n_0_11), .Q(\Memory[5] [63]), 
      .QN());
   DFF_X1 \Memory_reg[5][62]  (.D(Memory[62]), .CK(n_0_11), .Q(\Memory[5] [62]), 
      .QN());
   DFF_X1 \Memory_reg[5][61]  (.D(Memory[61]), .CK(n_0_11), .Q(\Memory[5] [61]), 
      .QN());
   DFF_X1 \Memory_reg[5][60]  (.D(Memory[60]), .CK(n_0_11), .Q(\Memory[5] [60]), 
      .QN());
   DFF_X1 \Memory_reg[5][59]  (.D(Memory[59]), .CK(n_0_11), .Q(\Memory[5] [59]), 
      .QN());
   DFF_X1 \Memory_reg[5][58]  (.D(Memory[58]), .CK(n_0_11), .Q(\Memory[5] [58]), 
      .QN());
   DFF_X1 \Memory_reg[5][57]  (.D(Memory[57]), .CK(n_0_11), .Q(\Memory[5] [57]), 
      .QN());
   DFF_X1 \Memory_reg[5][56]  (.D(Memory[56]), .CK(n_0_11), .Q(\Memory[5] [56]), 
      .QN());
   DFF_X1 \Memory_reg[5][55]  (.D(Memory[55]), .CK(n_0_11), .Q(\Memory[5] [55]), 
      .QN());
   DFF_X1 \Memory_reg[5][54]  (.D(Memory[54]), .CK(n_0_11), .Q(\Memory[5] [54]), 
      .QN());
   DFF_X1 \Memory_reg[5][53]  (.D(Memory[53]), .CK(n_0_11), .Q(\Memory[5] [53]), 
      .QN());
   DFF_X1 \Memory_reg[5][52]  (.D(Memory[52]), .CK(n_0_11), .Q(\Memory[5] [52]), 
      .QN());
   DFF_X1 \Memory_reg[5][51]  (.D(Memory[51]), .CK(n_0_11), .Q(\Memory[5] [51]), 
      .QN());
   DFF_X1 \Memory_reg[5][50]  (.D(Memory[50]), .CK(n_0_11), .Q(\Memory[5] [50]), 
      .QN());
   DFF_X1 \Memory_reg[5][49]  (.D(Memory[49]), .CK(n_0_11), .Q(\Memory[5] [49]), 
      .QN());
   DFF_X1 \Memory_reg[5][48]  (.D(Memory[48]), .CK(n_0_11), .Q(\Memory[5] [48]), 
      .QN());
   DFF_X1 \Memory_reg[5][47]  (.D(Memory[47]), .CK(n_0_11), .Q(\Memory[5] [47]), 
      .QN());
   DFF_X1 \Memory_reg[5][46]  (.D(Memory[46]), .CK(n_0_11), .Q(\Memory[5] [46]), 
      .QN());
   DFF_X1 \Memory_reg[5][45]  (.D(Memory[45]), .CK(n_0_11), .Q(\Memory[5] [45]), 
      .QN());
   DFF_X1 \Memory_reg[5][44]  (.D(Memory[44]), .CK(n_0_11), .Q(\Memory[5] [44]), 
      .QN());
   DFF_X1 \Memory_reg[5][43]  (.D(Memory[43]), .CK(n_0_11), .Q(\Memory[5] [43]), 
      .QN());
   DFF_X1 \Memory_reg[5][42]  (.D(Memory[42]), .CK(n_0_11), .Q(\Memory[5] [42]), 
      .QN());
   DFF_X1 \Memory_reg[5][41]  (.D(Memory[41]), .CK(n_0_11), .Q(\Memory[5] [41]), 
      .QN());
   DFF_X1 \Memory_reg[5][40]  (.D(Memory[40]), .CK(n_0_11), .Q(\Memory[5] [40]), 
      .QN());
   DFF_X1 \Memory_reg[5][39]  (.D(Memory[39]), .CK(n_0_11), .Q(\Memory[5] [39]), 
      .QN());
   DFF_X1 \Memory_reg[5][38]  (.D(Memory[38]), .CK(n_0_11), .Q(\Memory[5] [38]), 
      .QN());
   DFF_X1 \Memory_reg[5][37]  (.D(Memory[37]), .CK(n_0_11), .Q(\Memory[5] [37]), 
      .QN());
   DFF_X1 \Memory_reg[5][36]  (.D(Memory[36]), .CK(n_0_11), .Q(\Memory[5] [36]), 
      .QN());
   DFF_X1 \Memory_reg[5][35]  (.D(Memory[35]), .CK(n_0_11), .Q(\Memory[5] [35]), 
      .QN());
   DFF_X1 \Memory_reg[5][34]  (.D(Memory[34]), .CK(n_0_11), .Q(\Memory[5] [34]), 
      .QN());
   DFF_X1 \Memory_reg[5][33]  (.D(Memory[33]), .CK(n_0_11), .Q(\Memory[5] [33]), 
      .QN());
   DFF_X1 \Memory_reg[5][32]  (.D(Memory[32]), .CK(n_0_11), .Q(\Memory[5] [32]), 
      .QN());
   DFF_X1 \Memory_reg[5][31]  (.D(Memory[31]), .CK(n_0_11), .Q(\Memory[5] [31]), 
      .QN());
   DFF_X1 \Memory_reg[5][30]  (.D(Memory[30]), .CK(n_0_11), .Q(\Memory[5] [30]), 
      .QN());
   DFF_X1 \Memory_reg[5][29]  (.D(Memory[29]), .CK(n_0_11), .Q(\Memory[5] [29]), 
      .QN());
   DFF_X1 \Memory_reg[5][28]  (.D(Memory[28]), .CK(n_0_11), .Q(\Memory[5] [28]), 
      .QN());
   DFF_X1 \Memory_reg[5][27]  (.D(Memory[27]), .CK(n_0_11), .Q(\Memory[5] [27]), 
      .QN());
   DFF_X1 \Memory_reg[5][26]  (.D(Memory[26]), .CK(n_0_11), .Q(\Memory[5] [26]), 
      .QN());
   DFF_X1 \Memory_reg[5][25]  (.D(Memory[25]), .CK(n_0_11), .Q(\Memory[5] [25]), 
      .QN());
   DFF_X1 \Memory_reg[5][24]  (.D(Memory[24]), .CK(n_0_11), .Q(\Memory[5] [24]), 
      .QN());
   DFF_X1 \Memory_reg[5][23]  (.D(Memory[23]), .CK(n_0_11), .Q(\Memory[5] [23]), 
      .QN());
   DFF_X1 \Memory_reg[5][22]  (.D(Memory[22]), .CK(n_0_11), .Q(\Memory[5] [22]), 
      .QN());
   DFF_X1 \Memory_reg[5][21]  (.D(Memory[21]), .CK(n_0_11), .Q(\Memory[5] [21]), 
      .QN());
   DFF_X1 \Memory_reg[5][20]  (.D(Memory[20]), .CK(n_0_11), .Q(\Memory[5] [20]), 
      .QN());
   DFF_X1 \Memory_reg[5][19]  (.D(Memory[19]), .CK(n_0_11), .Q(\Memory[5] [19]), 
      .QN());
   DFF_X1 \Memory_reg[5][18]  (.D(Memory[18]), .CK(n_0_11), .Q(\Memory[5] [18]), 
      .QN());
   DFF_X1 \Memory_reg[5][17]  (.D(Memory[17]), .CK(n_0_11), .Q(\Memory[5] [17]), 
      .QN());
   DFF_X1 \Memory_reg[5][16]  (.D(Memory[16]), .CK(n_0_11), .Q(\Memory[5] [16]), 
      .QN());
   DFF_X1 \Memory_reg[5][15]  (.D(Memory[15]), .CK(n_0_11), .Q(\Memory[5] [15]), 
      .QN());
   DFF_X1 \Memory_reg[5][14]  (.D(Memory[14]), .CK(n_0_11), .Q(\Memory[5] [14]), 
      .QN());
   DFF_X1 \Memory_reg[5][13]  (.D(Memory[13]), .CK(n_0_11), .Q(\Memory[5] [13]), 
      .QN());
   DFF_X1 \Memory_reg[5][12]  (.D(Memory[12]), .CK(n_0_11), .Q(\Memory[5] [12]), 
      .QN());
   DFF_X1 \Memory_reg[5][11]  (.D(Memory[11]), .CK(n_0_11), .Q(\Memory[5] [11]), 
      .QN());
   DFF_X1 \Memory_reg[5][10]  (.D(Memory[10]), .CK(n_0_11), .Q(\Memory[5] [10]), 
      .QN());
   DFF_X1 \Memory_reg[5][9]  (.D(Memory[9]), .CK(n_0_11), .Q(\Memory[5] [9]), 
      .QN());
   DFF_X1 \Memory_reg[5][8]  (.D(Memory[8]), .CK(n_0_11), .Q(\Memory[5] [8]), 
      .QN());
   DFF_X1 \Memory_reg[5][7]  (.D(Memory[7]), .CK(n_0_11), .Q(\Memory[5] [7]), 
      .QN());
   DFF_X1 \Memory_reg[5][6]  (.D(Memory[6]), .CK(n_0_11), .Q(\Memory[5] [6]), 
      .QN());
   DFF_X1 \Memory_reg[5][5]  (.D(Memory[5]), .CK(n_0_11), .Q(\Memory[5] [5]), 
      .QN());
   DFF_X1 \Memory_reg[5][4]  (.D(Memory[4]), .CK(n_0_11), .Q(\Memory[5] [4]), 
      .QN());
   DFF_X1 \Memory_reg[5][3]  (.D(Memory[3]), .CK(n_0_11), .Q(\Memory[5] [3]), 
      .QN());
   DFF_X1 \Memory_reg[5][2]  (.D(Memory[2]), .CK(n_0_11), .Q(\Memory[5] [2]), 
      .QN());
   DFF_X1 \Memory_reg[5][1]  (.D(Memory[1]), .CK(n_0_11), .Q(\Memory[5] [1]), 
      .QN());
   DFF_X1 \Memory_reg[5][0]  (.D(Memory[0]), .CK(n_0_11), .Q(\Memory[5] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[4]_reg  (.CK(CLK), .E(n_0_21), .SE(1'b0), 
      .GCK(n_0_12));
   DFF_X1 \Memory_reg[4][63]  (.D(Memory[63]), .CK(n_0_12), .Q(\Memory[4] [63]), 
      .QN());
   DFF_X1 \Memory_reg[4][62]  (.D(Memory[62]), .CK(n_0_12), .Q(\Memory[4] [62]), 
      .QN());
   DFF_X1 \Memory_reg[4][61]  (.D(Memory[61]), .CK(n_0_12), .Q(\Memory[4] [61]), 
      .QN());
   DFF_X1 \Memory_reg[4][60]  (.D(Memory[60]), .CK(n_0_12), .Q(\Memory[4] [60]), 
      .QN());
   DFF_X1 \Memory_reg[4][59]  (.D(Memory[59]), .CK(n_0_12), .Q(\Memory[4] [59]), 
      .QN());
   DFF_X1 \Memory_reg[4][58]  (.D(Memory[58]), .CK(n_0_12), .Q(\Memory[4] [58]), 
      .QN());
   DFF_X1 \Memory_reg[4][57]  (.D(Memory[57]), .CK(n_0_12), .Q(\Memory[4] [57]), 
      .QN());
   DFF_X1 \Memory_reg[4][56]  (.D(Memory[56]), .CK(n_0_12), .Q(\Memory[4] [56]), 
      .QN());
   DFF_X1 \Memory_reg[4][55]  (.D(Memory[55]), .CK(n_0_12), .Q(\Memory[4] [55]), 
      .QN());
   DFF_X1 \Memory_reg[4][54]  (.D(Memory[54]), .CK(n_0_12), .Q(\Memory[4] [54]), 
      .QN());
   DFF_X1 \Memory_reg[4][53]  (.D(Memory[53]), .CK(n_0_12), .Q(\Memory[4] [53]), 
      .QN());
   DFF_X1 \Memory_reg[4][52]  (.D(Memory[52]), .CK(n_0_12), .Q(\Memory[4] [52]), 
      .QN());
   DFF_X1 \Memory_reg[4][51]  (.D(Memory[51]), .CK(n_0_12), .Q(\Memory[4] [51]), 
      .QN());
   DFF_X1 \Memory_reg[4][50]  (.D(Memory[50]), .CK(n_0_12), .Q(\Memory[4] [50]), 
      .QN());
   DFF_X1 \Memory_reg[4][49]  (.D(Memory[49]), .CK(n_0_12), .Q(\Memory[4] [49]), 
      .QN());
   DFF_X1 \Memory_reg[4][48]  (.D(Memory[48]), .CK(n_0_12), .Q(\Memory[4] [48]), 
      .QN());
   DFF_X1 \Memory_reg[4][47]  (.D(Memory[47]), .CK(n_0_12), .Q(\Memory[4] [47]), 
      .QN());
   DFF_X1 \Memory_reg[4][46]  (.D(Memory[46]), .CK(n_0_12), .Q(\Memory[4] [46]), 
      .QN());
   DFF_X1 \Memory_reg[4][45]  (.D(Memory[45]), .CK(n_0_12), .Q(\Memory[4] [45]), 
      .QN());
   DFF_X1 \Memory_reg[4][44]  (.D(Memory[44]), .CK(n_0_12), .Q(\Memory[4] [44]), 
      .QN());
   DFF_X1 \Memory_reg[4][43]  (.D(Memory[43]), .CK(n_0_12), .Q(\Memory[4] [43]), 
      .QN());
   DFF_X1 \Memory_reg[4][42]  (.D(Memory[42]), .CK(n_0_12), .Q(\Memory[4] [42]), 
      .QN());
   DFF_X1 \Memory_reg[4][41]  (.D(Memory[41]), .CK(n_0_12), .Q(\Memory[4] [41]), 
      .QN());
   DFF_X1 \Memory_reg[4][40]  (.D(Memory[40]), .CK(n_0_12), .Q(\Memory[4] [40]), 
      .QN());
   DFF_X1 \Memory_reg[4][39]  (.D(Memory[39]), .CK(n_0_12), .Q(\Memory[4] [39]), 
      .QN());
   DFF_X1 \Memory_reg[4][38]  (.D(Memory[38]), .CK(n_0_12), .Q(\Memory[4] [38]), 
      .QN());
   DFF_X1 \Memory_reg[4][37]  (.D(Memory[37]), .CK(n_0_12), .Q(\Memory[4] [37]), 
      .QN());
   DFF_X1 \Memory_reg[4][36]  (.D(Memory[36]), .CK(n_0_12), .Q(\Memory[4] [36]), 
      .QN());
   DFF_X1 \Memory_reg[4][35]  (.D(Memory[35]), .CK(n_0_12), .Q(\Memory[4] [35]), 
      .QN());
   DFF_X1 \Memory_reg[4][34]  (.D(Memory[34]), .CK(n_0_12), .Q(\Memory[4] [34]), 
      .QN());
   DFF_X1 \Memory_reg[4][33]  (.D(Memory[33]), .CK(n_0_12), .Q(\Memory[4] [33]), 
      .QN());
   DFF_X1 \Memory_reg[4][32]  (.D(Memory[32]), .CK(n_0_12), .Q(\Memory[4] [32]), 
      .QN());
   DFF_X1 \Memory_reg[4][31]  (.D(Memory[31]), .CK(n_0_12), .Q(\Memory[4] [31]), 
      .QN());
   DFF_X1 \Memory_reg[4][30]  (.D(Memory[30]), .CK(n_0_12), .Q(\Memory[4] [30]), 
      .QN());
   DFF_X1 \Memory_reg[4][29]  (.D(Memory[29]), .CK(n_0_12), .Q(\Memory[4] [29]), 
      .QN());
   DFF_X1 \Memory_reg[4][28]  (.D(Memory[28]), .CK(n_0_12), .Q(\Memory[4] [28]), 
      .QN());
   DFF_X1 \Memory_reg[4][27]  (.D(Memory[27]), .CK(n_0_12), .Q(\Memory[4] [27]), 
      .QN());
   DFF_X1 \Memory_reg[4][26]  (.D(Memory[26]), .CK(n_0_12), .Q(\Memory[4] [26]), 
      .QN());
   DFF_X1 \Memory_reg[4][25]  (.D(Memory[25]), .CK(n_0_12), .Q(\Memory[4] [25]), 
      .QN());
   DFF_X1 \Memory_reg[4][24]  (.D(Memory[24]), .CK(n_0_12), .Q(\Memory[4] [24]), 
      .QN());
   DFF_X1 \Memory_reg[4][23]  (.D(Memory[23]), .CK(n_0_12), .Q(\Memory[4] [23]), 
      .QN());
   DFF_X1 \Memory_reg[4][22]  (.D(Memory[22]), .CK(n_0_12), .Q(\Memory[4] [22]), 
      .QN());
   DFF_X1 \Memory_reg[4][21]  (.D(Memory[21]), .CK(n_0_12), .Q(\Memory[4] [21]), 
      .QN());
   DFF_X1 \Memory_reg[4][20]  (.D(Memory[20]), .CK(n_0_12), .Q(\Memory[4] [20]), 
      .QN());
   DFF_X1 \Memory_reg[4][19]  (.D(Memory[19]), .CK(n_0_12), .Q(\Memory[4] [19]), 
      .QN());
   DFF_X1 \Memory_reg[4][18]  (.D(Memory[18]), .CK(n_0_12), .Q(\Memory[4] [18]), 
      .QN());
   DFF_X1 \Memory_reg[4][17]  (.D(Memory[17]), .CK(n_0_12), .Q(\Memory[4] [17]), 
      .QN());
   DFF_X1 \Memory_reg[4][16]  (.D(Memory[16]), .CK(n_0_12), .Q(\Memory[4] [16]), 
      .QN());
   DFF_X1 \Memory_reg[4][15]  (.D(Memory[15]), .CK(n_0_12), .Q(\Memory[4] [15]), 
      .QN());
   DFF_X1 \Memory_reg[4][14]  (.D(Memory[14]), .CK(n_0_12), .Q(\Memory[4] [14]), 
      .QN());
   DFF_X1 \Memory_reg[4][13]  (.D(Memory[13]), .CK(n_0_12), .Q(\Memory[4] [13]), 
      .QN());
   DFF_X1 \Memory_reg[4][12]  (.D(Memory[12]), .CK(n_0_12), .Q(\Memory[4] [12]), 
      .QN());
   DFF_X1 \Memory_reg[4][11]  (.D(Memory[11]), .CK(n_0_12), .Q(\Memory[4] [11]), 
      .QN());
   DFF_X1 \Memory_reg[4][10]  (.D(Memory[10]), .CK(n_0_12), .Q(\Memory[4] [10]), 
      .QN());
   DFF_X1 \Memory_reg[4][9]  (.D(Memory[9]), .CK(n_0_12), .Q(\Memory[4] [9]), 
      .QN());
   DFF_X1 \Memory_reg[4][8]  (.D(Memory[8]), .CK(n_0_12), .Q(\Memory[4] [8]), 
      .QN());
   DFF_X1 \Memory_reg[4][7]  (.D(Memory[7]), .CK(n_0_12), .Q(\Memory[4] [7]), 
      .QN());
   DFF_X1 \Memory_reg[4][6]  (.D(Memory[6]), .CK(n_0_12), .Q(\Memory[4] [6]), 
      .QN());
   DFF_X1 \Memory_reg[4][5]  (.D(Memory[5]), .CK(n_0_12), .Q(\Memory[4] [5]), 
      .QN());
   DFF_X1 \Memory_reg[4][4]  (.D(Memory[4]), .CK(n_0_12), .Q(\Memory[4] [4]), 
      .QN());
   DFF_X1 \Memory_reg[4][3]  (.D(Memory[3]), .CK(n_0_12), .Q(\Memory[4] [3]), 
      .QN());
   DFF_X1 \Memory_reg[4][2]  (.D(Memory[2]), .CK(n_0_12), .Q(\Memory[4] [2]), 
      .QN());
   DFF_X1 \Memory_reg[4][1]  (.D(Memory[1]), .CK(n_0_12), .Q(\Memory[4] [1]), 
      .QN());
   DFF_X1 \Memory_reg[4][0]  (.D(Memory[0]), .CK(n_0_12), .Q(\Memory[4] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[3]_reg  (.CK(CLK), .E(n_0_20), .SE(1'b0), 
      .GCK(n_0_13));
   DFF_X1 \Memory_reg[3][63]  (.D(Memory[63]), .CK(n_0_13), .Q(\Memory[3] [63]), 
      .QN());
   DFF_X1 \Memory_reg[3][62]  (.D(Memory[62]), .CK(n_0_13), .Q(\Memory[3] [62]), 
      .QN());
   DFF_X1 \Memory_reg[3][61]  (.D(Memory[61]), .CK(n_0_13), .Q(\Memory[3] [61]), 
      .QN());
   DFF_X1 \Memory_reg[3][60]  (.D(Memory[60]), .CK(n_0_13), .Q(\Memory[3] [60]), 
      .QN());
   DFF_X1 \Memory_reg[3][59]  (.D(Memory[59]), .CK(n_0_13), .Q(\Memory[3] [59]), 
      .QN());
   DFF_X1 \Memory_reg[3][58]  (.D(Memory[58]), .CK(n_0_13), .Q(\Memory[3] [58]), 
      .QN());
   DFF_X1 \Memory_reg[3][57]  (.D(Memory[57]), .CK(n_0_13), .Q(\Memory[3] [57]), 
      .QN());
   DFF_X1 \Memory_reg[3][56]  (.D(Memory[56]), .CK(n_0_13), .Q(\Memory[3] [56]), 
      .QN());
   DFF_X1 \Memory_reg[3][55]  (.D(Memory[55]), .CK(n_0_13), .Q(\Memory[3] [55]), 
      .QN());
   DFF_X1 \Memory_reg[3][54]  (.D(Memory[54]), .CK(n_0_13), .Q(\Memory[3] [54]), 
      .QN());
   DFF_X1 \Memory_reg[3][53]  (.D(Memory[53]), .CK(n_0_13), .Q(\Memory[3] [53]), 
      .QN());
   DFF_X1 \Memory_reg[3][52]  (.D(Memory[52]), .CK(n_0_13), .Q(\Memory[3] [52]), 
      .QN());
   DFF_X1 \Memory_reg[3][51]  (.D(Memory[51]), .CK(n_0_13), .Q(\Memory[3] [51]), 
      .QN());
   DFF_X1 \Memory_reg[3][50]  (.D(Memory[50]), .CK(n_0_13), .Q(\Memory[3] [50]), 
      .QN());
   DFF_X1 \Memory_reg[3][49]  (.D(Memory[49]), .CK(n_0_13), .Q(\Memory[3] [49]), 
      .QN());
   DFF_X1 \Memory_reg[3][48]  (.D(Memory[48]), .CK(n_0_13), .Q(\Memory[3] [48]), 
      .QN());
   DFF_X1 \Memory_reg[3][47]  (.D(Memory[47]), .CK(n_0_13), .Q(\Memory[3] [47]), 
      .QN());
   DFF_X1 \Memory_reg[3][46]  (.D(Memory[46]), .CK(n_0_13), .Q(\Memory[3] [46]), 
      .QN());
   DFF_X1 \Memory_reg[3][45]  (.D(Memory[45]), .CK(n_0_13), .Q(\Memory[3] [45]), 
      .QN());
   DFF_X1 \Memory_reg[3][44]  (.D(Memory[44]), .CK(n_0_13), .Q(\Memory[3] [44]), 
      .QN());
   DFF_X1 \Memory_reg[3][43]  (.D(Memory[43]), .CK(n_0_13), .Q(\Memory[3] [43]), 
      .QN());
   DFF_X1 \Memory_reg[3][42]  (.D(Memory[42]), .CK(n_0_13), .Q(\Memory[3] [42]), 
      .QN());
   DFF_X1 \Memory_reg[3][41]  (.D(Memory[41]), .CK(n_0_13), .Q(\Memory[3] [41]), 
      .QN());
   DFF_X1 \Memory_reg[3][40]  (.D(Memory[40]), .CK(n_0_13), .Q(\Memory[3] [40]), 
      .QN());
   DFF_X1 \Memory_reg[3][39]  (.D(Memory[39]), .CK(n_0_13), .Q(\Memory[3] [39]), 
      .QN());
   DFF_X1 \Memory_reg[3][38]  (.D(Memory[38]), .CK(n_0_13), .Q(\Memory[3] [38]), 
      .QN());
   DFF_X1 \Memory_reg[3][37]  (.D(Memory[37]), .CK(n_0_13), .Q(\Memory[3] [37]), 
      .QN());
   DFF_X1 \Memory_reg[3][36]  (.D(Memory[36]), .CK(n_0_13), .Q(\Memory[3] [36]), 
      .QN());
   DFF_X1 \Memory_reg[3][35]  (.D(Memory[35]), .CK(n_0_13), .Q(\Memory[3] [35]), 
      .QN());
   DFF_X1 \Memory_reg[3][34]  (.D(Memory[34]), .CK(n_0_13), .Q(\Memory[3] [34]), 
      .QN());
   DFF_X1 \Memory_reg[3][33]  (.D(Memory[33]), .CK(n_0_13), .Q(\Memory[3] [33]), 
      .QN());
   DFF_X1 \Memory_reg[3][32]  (.D(Memory[32]), .CK(n_0_13), .Q(\Memory[3] [32]), 
      .QN());
   DFF_X1 \Memory_reg[3][31]  (.D(Memory[31]), .CK(n_0_13), .Q(\Memory[3] [31]), 
      .QN());
   DFF_X1 \Memory_reg[3][30]  (.D(Memory[30]), .CK(n_0_13), .Q(\Memory[3] [30]), 
      .QN());
   DFF_X1 \Memory_reg[3][29]  (.D(Memory[29]), .CK(n_0_13), .Q(\Memory[3] [29]), 
      .QN());
   DFF_X1 \Memory_reg[3][28]  (.D(Memory[28]), .CK(n_0_13), .Q(\Memory[3] [28]), 
      .QN());
   DFF_X1 \Memory_reg[3][27]  (.D(Memory[27]), .CK(n_0_13), .Q(\Memory[3] [27]), 
      .QN());
   DFF_X1 \Memory_reg[3][26]  (.D(Memory[26]), .CK(n_0_13), .Q(\Memory[3] [26]), 
      .QN());
   DFF_X1 \Memory_reg[3][25]  (.D(Memory[25]), .CK(n_0_13), .Q(\Memory[3] [25]), 
      .QN());
   DFF_X1 \Memory_reg[3][24]  (.D(Memory[24]), .CK(n_0_13), .Q(\Memory[3] [24]), 
      .QN());
   DFF_X1 \Memory_reg[3][23]  (.D(Memory[23]), .CK(n_0_13), .Q(\Memory[3] [23]), 
      .QN());
   DFF_X1 \Memory_reg[3][22]  (.D(Memory[22]), .CK(n_0_13), .Q(\Memory[3] [22]), 
      .QN());
   DFF_X1 \Memory_reg[3][21]  (.D(Memory[21]), .CK(n_0_13), .Q(\Memory[3] [21]), 
      .QN());
   DFF_X1 \Memory_reg[3][20]  (.D(Memory[20]), .CK(n_0_13), .Q(\Memory[3] [20]), 
      .QN());
   DFF_X1 \Memory_reg[3][19]  (.D(Memory[19]), .CK(n_0_13), .Q(\Memory[3] [19]), 
      .QN());
   DFF_X1 \Memory_reg[3][18]  (.D(Memory[18]), .CK(n_0_13), .Q(\Memory[3] [18]), 
      .QN());
   DFF_X1 \Memory_reg[3][17]  (.D(Memory[17]), .CK(n_0_13), .Q(\Memory[3] [17]), 
      .QN());
   DFF_X1 \Memory_reg[3][16]  (.D(Memory[16]), .CK(n_0_13), .Q(\Memory[3] [16]), 
      .QN());
   DFF_X1 \Memory_reg[3][15]  (.D(Memory[15]), .CK(n_0_13), .Q(\Memory[3] [15]), 
      .QN());
   DFF_X1 \Memory_reg[3][14]  (.D(Memory[14]), .CK(n_0_13), .Q(\Memory[3] [14]), 
      .QN());
   DFF_X1 \Memory_reg[3][13]  (.D(Memory[13]), .CK(n_0_13), .Q(\Memory[3] [13]), 
      .QN());
   DFF_X1 \Memory_reg[3][12]  (.D(Memory[12]), .CK(n_0_13), .Q(\Memory[3] [12]), 
      .QN());
   DFF_X1 \Memory_reg[3][11]  (.D(Memory[11]), .CK(n_0_13), .Q(\Memory[3] [11]), 
      .QN());
   DFF_X1 \Memory_reg[3][10]  (.D(Memory[10]), .CK(n_0_13), .Q(\Memory[3] [10]), 
      .QN());
   DFF_X1 \Memory_reg[3][9]  (.D(Memory[9]), .CK(n_0_13), .Q(\Memory[3] [9]), 
      .QN());
   DFF_X1 \Memory_reg[3][8]  (.D(Memory[8]), .CK(n_0_13), .Q(\Memory[3] [8]), 
      .QN());
   DFF_X1 \Memory_reg[3][7]  (.D(Memory[7]), .CK(n_0_13), .Q(\Memory[3] [7]), 
      .QN());
   DFF_X1 \Memory_reg[3][6]  (.D(Memory[6]), .CK(n_0_13), .Q(\Memory[3] [6]), 
      .QN());
   DFF_X1 \Memory_reg[3][5]  (.D(Memory[5]), .CK(n_0_13), .Q(\Memory[3] [5]), 
      .QN());
   DFF_X1 \Memory_reg[3][4]  (.D(Memory[4]), .CK(n_0_13), .Q(\Memory[3] [4]), 
      .QN());
   DFF_X1 \Memory_reg[3][3]  (.D(Memory[3]), .CK(n_0_13), .Q(\Memory[3] [3]), 
      .QN());
   DFF_X1 \Memory_reg[3][2]  (.D(Memory[2]), .CK(n_0_13), .Q(\Memory[3] [2]), 
      .QN());
   DFF_X1 \Memory_reg[3][1]  (.D(Memory[1]), .CK(n_0_13), .Q(\Memory[3] [1]), 
      .QN());
   DFF_X1 \Memory_reg[3][0]  (.D(Memory[0]), .CK(n_0_13), .Q(\Memory[3] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[2]_reg  (.CK(CLK), .E(n_0_19), .SE(1'b0), 
      .GCK(n_0_14));
   DFF_X1 \Memory_reg[2][63]  (.D(Memory[63]), .CK(n_0_14), .Q(\Memory[2] [63]), 
      .QN());
   DFF_X1 \Memory_reg[2][62]  (.D(Memory[62]), .CK(n_0_14), .Q(\Memory[2] [62]), 
      .QN());
   DFF_X1 \Memory_reg[2][61]  (.D(Memory[61]), .CK(n_0_14), .Q(\Memory[2] [61]), 
      .QN());
   DFF_X1 \Memory_reg[2][60]  (.D(Memory[60]), .CK(n_0_14), .Q(\Memory[2] [60]), 
      .QN());
   DFF_X1 \Memory_reg[2][59]  (.D(Memory[59]), .CK(n_0_14), .Q(\Memory[2] [59]), 
      .QN());
   DFF_X1 \Memory_reg[2][58]  (.D(Memory[58]), .CK(n_0_14), .Q(\Memory[2] [58]), 
      .QN());
   DFF_X1 \Memory_reg[2][57]  (.D(Memory[57]), .CK(n_0_14), .Q(\Memory[2] [57]), 
      .QN());
   DFF_X1 \Memory_reg[2][56]  (.D(Memory[56]), .CK(n_0_14), .Q(\Memory[2] [56]), 
      .QN());
   DFF_X1 \Memory_reg[2][55]  (.D(Memory[55]), .CK(n_0_14), .Q(\Memory[2] [55]), 
      .QN());
   DFF_X1 \Memory_reg[2][54]  (.D(Memory[54]), .CK(n_0_14), .Q(\Memory[2] [54]), 
      .QN());
   DFF_X1 \Memory_reg[2][53]  (.D(Memory[53]), .CK(n_0_14), .Q(\Memory[2] [53]), 
      .QN());
   DFF_X1 \Memory_reg[2][52]  (.D(Memory[52]), .CK(n_0_14), .Q(\Memory[2] [52]), 
      .QN());
   DFF_X1 \Memory_reg[2][51]  (.D(Memory[51]), .CK(n_0_14), .Q(\Memory[2] [51]), 
      .QN());
   DFF_X1 \Memory_reg[2][50]  (.D(Memory[50]), .CK(n_0_14), .Q(\Memory[2] [50]), 
      .QN());
   DFF_X1 \Memory_reg[2][49]  (.D(Memory[49]), .CK(n_0_14), .Q(\Memory[2] [49]), 
      .QN());
   DFF_X1 \Memory_reg[2][48]  (.D(Memory[48]), .CK(n_0_14), .Q(\Memory[2] [48]), 
      .QN());
   DFF_X1 \Memory_reg[2][47]  (.D(Memory[47]), .CK(n_0_14), .Q(\Memory[2] [47]), 
      .QN());
   DFF_X1 \Memory_reg[2][46]  (.D(Memory[46]), .CK(n_0_14), .Q(\Memory[2] [46]), 
      .QN());
   DFF_X1 \Memory_reg[2][45]  (.D(Memory[45]), .CK(n_0_14), .Q(\Memory[2] [45]), 
      .QN());
   DFF_X1 \Memory_reg[2][44]  (.D(Memory[44]), .CK(n_0_14), .Q(\Memory[2] [44]), 
      .QN());
   DFF_X1 \Memory_reg[2][43]  (.D(Memory[43]), .CK(n_0_14), .Q(\Memory[2] [43]), 
      .QN());
   DFF_X1 \Memory_reg[2][42]  (.D(Memory[42]), .CK(n_0_14), .Q(\Memory[2] [42]), 
      .QN());
   DFF_X1 \Memory_reg[2][41]  (.D(Memory[41]), .CK(n_0_14), .Q(\Memory[2] [41]), 
      .QN());
   DFF_X1 \Memory_reg[2][40]  (.D(Memory[40]), .CK(n_0_14), .Q(\Memory[2] [40]), 
      .QN());
   DFF_X1 \Memory_reg[2][39]  (.D(Memory[39]), .CK(n_0_14), .Q(\Memory[2] [39]), 
      .QN());
   DFF_X1 \Memory_reg[2][38]  (.D(Memory[38]), .CK(n_0_14), .Q(\Memory[2] [38]), 
      .QN());
   DFF_X1 \Memory_reg[2][37]  (.D(Memory[37]), .CK(n_0_14), .Q(\Memory[2] [37]), 
      .QN());
   DFF_X1 \Memory_reg[2][36]  (.D(Memory[36]), .CK(n_0_14), .Q(\Memory[2] [36]), 
      .QN());
   DFF_X1 \Memory_reg[2][35]  (.D(Memory[35]), .CK(n_0_14), .Q(\Memory[2] [35]), 
      .QN());
   DFF_X1 \Memory_reg[2][34]  (.D(Memory[34]), .CK(n_0_14), .Q(\Memory[2] [34]), 
      .QN());
   DFF_X1 \Memory_reg[2][33]  (.D(Memory[33]), .CK(n_0_14), .Q(\Memory[2] [33]), 
      .QN());
   DFF_X1 \Memory_reg[2][32]  (.D(Memory[32]), .CK(n_0_14), .Q(\Memory[2] [32]), 
      .QN());
   DFF_X1 \Memory_reg[2][31]  (.D(Memory[31]), .CK(n_0_14), .Q(\Memory[2] [31]), 
      .QN());
   DFF_X1 \Memory_reg[2][30]  (.D(Memory[30]), .CK(n_0_14), .Q(\Memory[2] [30]), 
      .QN());
   DFF_X1 \Memory_reg[2][29]  (.D(Memory[29]), .CK(n_0_14), .Q(\Memory[2] [29]), 
      .QN());
   DFF_X1 \Memory_reg[2][28]  (.D(Memory[28]), .CK(n_0_14), .Q(\Memory[2] [28]), 
      .QN());
   DFF_X1 \Memory_reg[2][27]  (.D(Memory[27]), .CK(n_0_14), .Q(\Memory[2] [27]), 
      .QN());
   DFF_X1 \Memory_reg[2][26]  (.D(Memory[26]), .CK(n_0_14), .Q(\Memory[2] [26]), 
      .QN());
   DFF_X1 \Memory_reg[2][25]  (.D(Memory[25]), .CK(n_0_14), .Q(\Memory[2] [25]), 
      .QN());
   DFF_X1 \Memory_reg[2][24]  (.D(Memory[24]), .CK(n_0_14), .Q(\Memory[2] [24]), 
      .QN());
   DFF_X1 \Memory_reg[2][23]  (.D(Memory[23]), .CK(n_0_14), .Q(\Memory[2] [23]), 
      .QN());
   DFF_X1 \Memory_reg[2][22]  (.D(Memory[22]), .CK(n_0_14), .Q(\Memory[2] [22]), 
      .QN());
   DFF_X1 \Memory_reg[2][21]  (.D(Memory[21]), .CK(n_0_14), .Q(\Memory[2] [21]), 
      .QN());
   DFF_X1 \Memory_reg[2][20]  (.D(Memory[20]), .CK(n_0_14), .Q(\Memory[2] [20]), 
      .QN());
   DFF_X1 \Memory_reg[2][19]  (.D(Memory[19]), .CK(n_0_14), .Q(\Memory[2] [19]), 
      .QN());
   DFF_X1 \Memory_reg[2][18]  (.D(Memory[18]), .CK(n_0_14), .Q(\Memory[2] [18]), 
      .QN());
   DFF_X1 \Memory_reg[2][17]  (.D(Memory[17]), .CK(n_0_14), .Q(\Memory[2] [17]), 
      .QN());
   DFF_X1 \Memory_reg[2][16]  (.D(Memory[16]), .CK(n_0_14), .Q(\Memory[2] [16]), 
      .QN());
   DFF_X1 \Memory_reg[2][15]  (.D(Memory[15]), .CK(n_0_14), .Q(\Memory[2] [15]), 
      .QN());
   DFF_X1 \Memory_reg[2][14]  (.D(Memory[14]), .CK(n_0_14), .Q(\Memory[2] [14]), 
      .QN());
   DFF_X1 \Memory_reg[2][13]  (.D(Memory[13]), .CK(n_0_14), .Q(\Memory[2] [13]), 
      .QN());
   DFF_X1 \Memory_reg[2][12]  (.D(Memory[12]), .CK(n_0_14), .Q(\Memory[2] [12]), 
      .QN());
   DFF_X1 \Memory_reg[2][11]  (.D(Memory[11]), .CK(n_0_14), .Q(\Memory[2] [11]), 
      .QN());
   DFF_X1 \Memory_reg[2][10]  (.D(Memory[10]), .CK(n_0_14), .Q(\Memory[2] [10]), 
      .QN());
   DFF_X1 \Memory_reg[2][9]  (.D(Memory[9]), .CK(n_0_14), .Q(\Memory[2] [9]), 
      .QN());
   DFF_X1 \Memory_reg[2][8]  (.D(Memory[8]), .CK(n_0_14), .Q(\Memory[2] [8]), 
      .QN());
   DFF_X1 \Memory_reg[2][7]  (.D(Memory[7]), .CK(n_0_14), .Q(\Memory[2] [7]), 
      .QN());
   DFF_X1 \Memory_reg[2][6]  (.D(Memory[6]), .CK(n_0_14), .Q(\Memory[2] [6]), 
      .QN());
   DFF_X1 \Memory_reg[2][5]  (.D(Memory[5]), .CK(n_0_14), .Q(\Memory[2] [5]), 
      .QN());
   DFF_X1 \Memory_reg[2][4]  (.D(Memory[4]), .CK(n_0_14), .Q(\Memory[2] [4]), 
      .QN());
   DFF_X1 \Memory_reg[2][3]  (.D(Memory[3]), .CK(n_0_14), .Q(\Memory[2] [3]), 
      .QN());
   DFF_X1 \Memory_reg[2][2]  (.D(Memory[2]), .CK(n_0_14), .Q(\Memory[2] [2]), 
      .QN());
   DFF_X1 \Memory_reg[2][1]  (.D(Memory[1]), .CK(n_0_14), .Q(\Memory[2] [1]), 
      .QN());
   DFF_X1 \Memory_reg[2][0]  (.D(Memory[0]), .CK(n_0_14), .Q(\Memory[2] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[1]_reg  (.CK(CLK), .E(n_0_18), .SE(1'b0), 
      .GCK(n_0_15));
   DFF_X1 \Memory_reg[1][63]  (.D(Memory[63]), .CK(n_0_15), .Q(\Memory[1] [63]), 
      .QN());
   DFF_X1 \Memory_reg[1][62]  (.D(Memory[62]), .CK(n_0_15), .Q(\Memory[1] [62]), 
      .QN());
   DFF_X1 \Memory_reg[1][61]  (.D(Memory[61]), .CK(n_0_15), .Q(\Memory[1] [61]), 
      .QN());
   DFF_X1 \Memory_reg[1][60]  (.D(Memory[60]), .CK(n_0_15), .Q(\Memory[1] [60]), 
      .QN());
   DFF_X1 \Memory_reg[1][59]  (.D(Memory[59]), .CK(n_0_15), .Q(\Memory[1] [59]), 
      .QN());
   DFF_X1 \Memory_reg[1][58]  (.D(Memory[58]), .CK(n_0_15), .Q(\Memory[1] [58]), 
      .QN());
   DFF_X1 \Memory_reg[1][57]  (.D(Memory[57]), .CK(n_0_15), .Q(\Memory[1] [57]), 
      .QN());
   DFF_X1 \Memory_reg[1][56]  (.D(Memory[56]), .CK(n_0_15), .Q(\Memory[1] [56]), 
      .QN());
   DFF_X1 \Memory_reg[1][55]  (.D(Memory[55]), .CK(n_0_15), .Q(\Memory[1] [55]), 
      .QN());
   DFF_X1 \Memory_reg[1][54]  (.D(Memory[54]), .CK(n_0_15), .Q(\Memory[1] [54]), 
      .QN());
   DFF_X1 \Memory_reg[1][53]  (.D(Memory[53]), .CK(n_0_15), .Q(\Memory[1] [53]), 
      .QN());
   DFF_X1 \Memory_reg[1][52]  (.D(Memory[52]), .CK(n_0_15), .Q(\Memory[1] [52]), 
      .QN());
   DFF_X1 \Memory_reg[1][51]  (.D(Memory[51]), .CK(n_0_15), .Q(\Memory[1] [51]), 
      .QN());
   DFF_X1 \Memory_reg[1][50]  (.D(Memory[50]), .CK(n_0_15), .Q(\Memory[1] [50]), 
      .QN());
   DFF_X1 \Memory_reg[1][49]  (.D(Memory[49]), .CK(n_0_15), .Q(\Memory[1] [49]), 
      .QN());
   DFF_X1 \Memory_reg[1][48]  (.D(Memory[48]), .CK(n_0_15), .Q(\Memory[1] [48]), 
      .QN());
   DFF_X1 \Memory_reg[1][47]  (.D(Memory[47]), .CK(n_0_15), .Q(\Memory[1] [47]), 
      .QN());
   DFF_X1 \Memory_reg[1][46]  (.D(Memory[46]), .CK(n_0_15), .Q(\Memory[1] [46]), 
      .QN());
   DFF_X1 \Memory_reg[1][45]  (.D(Memory[45]), .CK(n_0_15), .Q(\Memory[1] [45]), 
      .QN());
   DFF_X1 \Memory_reg[1][44]  (.D(Memory[44]), .CK(n_0_15), .Q(\Memory[1] [44]), 
      .QN());
   DFF_X1 \Memory_reg[1][43]  (.D(Memory[43]), .CK(n_0_15), .Q(\Memory[1] [43]), 
      .QN());
   DFF_X1 \Memory_reg[1][42]  (.D(Memory[42]), .CK(n_0_15), .Q(\Memory[1] [42]), 
      .QN());
   DFF_X1 \Memory_reg[1][41]  (.D(Memory[41]), .CK(n_0_15), .Q(\Memory[1] [41]), 
      .QN());
   DFF_X1 \Memory_reg[1][40]  (.D(Memory[40]), .CK(n_0_15), .Q(\Memory[1] [40]), 
      .QN());
   DFF_X1 \Memory_reg[1][39]  (.D(Memory[39]), .CK(n_0_15), .Q(\Memory[1] [39]), 
      .QN());
   DFF_X1 \Memory_reg[1][38]  (.D(Memory[38]), .CK(n_0_15), .Q(\Memory[1] [38]), 
      .QN());
   DFF_X1 \Memory_reg[1][37]  (.D(Memory[37]), .CK(n_0_15), .Q(\Memory[1] [37]), 
      .QN());
   DFF_X1 \Memory_reg[1][36]  (.D(Memory[36]), .CK(n_0_15), .Q(\Memory[1] [36]), 
      .QN());
   DFF_X1 \Memory_reg[1][35]  (.D(Memory[35]), .CK(n_0_15), .Q(\Memory[1] [35]), 
      .QN());
   DFF_X1 \Memory_reg[1][34]  (.D(Memory[34]), .CK(n_0_15), .Q(\Memory[1] [34]), 
      .QN());
   DFF_X1 \Memory_reg[1][33]  (.D(Memory[33]), .CK(n_0_15), .Q(\Memory[1] [33]), 
      .QN());
   DFF_X1 \Memory_reg[1][32]  (.D(Memory[32]), .CK(n_0_15), .Q(\Memory[1] [32]), 
      .QN());
   DFF_X1 \Memory_reg[1][31]  (.D(Memory[31]), .CK(n_0_15), .Q(\Memory[1] [31]), 
      .QN());
   DFF_X1 \Memory_reg[1][30]  (.D(Memory[30]), .CK(n_0_15), .Q(\Memory[1] [30]), 
      .QN());
   DFF_X1 \Memory_reg[1][29]  (.D(Memory[29]), .CK(n_0_15), .Q(\Memory[1] [29]), 
      .QN());
   DFF_X1 \Memory_reg[1][28]  (.D(Memory[28]), .CK(n_0_15), .Q(\Memory[1] [28]), 
      .QN());
   DFF_X1 \Memory_reg[1][27]  (.D(Memory[27]), .CK(n_0_15), .Q(\Memory[1] [27]), 
      .QN());
   DFF_X1 \Memory_reg[1][26]  (.D(Memory[26]), .CK(n_0_15), .Q(\Memory[1] [26]), 
      .QN());
   DFF_X1 \Memory_reg[1][25]  (.D(Memory[25]), .CK(n_0_15), .Q(\Memory[1] [25]), 
      .QN());
   DFF_X1 \Memory_reg[1][24]  (.D(Memory[24]), .CK(n_0_15), .Q(\Memory[1] [24]), 
      .QN());
   DFF_X1 \Memory_reg[1][23]  (.D(Memory[23]), .CK(n_0_15), .Q(\Memory[1] [23]), 
      .QN());
   DFF_X1 \Memory_reg[1][22]  (.D(Memory[22]), .CK(n_0_15), .Q(\Memory[1] [22]), 
      .QN());
   DFF_X1 \Memory_reg[1][21]  (.D(Memory[21]), .CK(n_0_15), .Q(\Memory[1] [21]), 
      .QN());
   DFF_X1 \Memory_reg[1][20]  (.D(Memory[20]), .CK(n_0_15), .Q(\Memory[1] [20]), 
      .QN());
   DFF_X1 \Memory_reg[1][19]  (.D(Memory[19]), .CK(n_0_15), .Q(\Memory[1] [19]), 
      .QN());
   DFF_X1 \Memory_reg[1][18]  (.D(Memory[18]), .CK(n_0_15), .Q(\Memory[1] [18]), 
      .QN());
   DFF_X1 \Memory_reg[1][17]  (.D(Memory[17]), .CK(n_0_15), .Q(\Memory[1] [17]), 
      .QN());
   DFF_X1 \Memory_reg[1][16]  (.D(Memory[16]), .CK(n_0_15), .Q(\Memory[1] [16]), 
      .QN());
   DFF_X1 \Memory_reg[1][15]  (.D(Memory[15]), .CK(n_0_15), .Q(\Memory[1] [15]), 
      .QN());
   DFF_X1 \Memory_reg[1][14]  (.D(Memory[14]), .CK(n_0_15), .Q(\Memory[1] [14]), 
      .QN());
   DFF_X1 \Memory_reg[1][13]  (.D(Memory[13]), .CK(n_0_15), .Q(\Memory[1] [13]), 
      .QN());
   DFF_X1 \Memory_reg[1][12]  (.D(Memory[12]), .CK(n_0_15), .Q(\Memory[1] [12]), 
      .QN());
   DFF_X1 \Memory_reg[1][11]  (.D(Memory[11]), .CK(n_0_15), .Q(\Memory[1] [11]), 
      .QN());
   DFF_X1 \Memory_reg[1][10]  (.D(Memory[10]), .CK(n_0_15), .Q(\Memory[1] [10]), 
      .QN());
   DFF_X1 \Memory_reg[1][9]  (.D(Memory[9]), .CK(n_0_15), .Q(\Memory[1] [9]), 
      .QN());
   DFF_X1 \Memory_reg[1][8]  (.D(Memory[8]), .CK(n_0_15), .Q(\Memory[1] [8]), 
      .QN());
   DFF_X1 \Memory_reg[1][7]  (.D(Memory[7]), .CK(n_0_15), .Q(\Memory[1] [7]), 
      .QN());
   DFF_X1 \Memory_reg[1][6]  (.D(Memory[6]), .CK(n_0_15), .Q(\Memory[1] [6]), 
      .QN());
   DFF_X1 \Memory_reg[1][5]  (.D(Memory[5]), .CK(n_0_15), .Q(\Memory[1] [5]), 
      .QN());
   DFF_X1 \Memory_reg[1][4]  (.D(Memory[4]), .CK(n_0_15), .Q(\Memory[1] [4]), 
      .QN());
   DFF_X1 \Memory_reg[1][3]  (.D(Memory[3]), .CK(n_0_15), .Q(\Memory[1] [3]), 
      .QN());
   DFF_X1 \Memory_reg[1][2]  (.D(Memory[2]), .CK(n_0_15), .Q(\Memory[1] [2]), 
      .QN());
   DFF_X1 \Memory_reg[1][1]  (.D(Memory[1]), .CK(n_0_15), .Q(\Memory[1] [1]), 
      .QN());
   DFF_X1 \Memory_reg[1][0]  (.D(Memory[0]), .CK(n_0_15), .Q(\Memory[1] [0]), 
      .QN());
   CLKGATETST_X1 \clk_gate_Memory_reg[0]_reg  (.CK(CLK), .E(n_0_17), .SE(1'b0), 
      .GCK(n_0_16));
   DFF_X1 \Memory_reg[0][63]  (.D(Memory[63]), .CK(n_0_16), .Q(\Memory[0] [63]), 
      .QN());
   DFF_X1 \Memory_reg[0][62]  (.D(Memory[62]), .CK(n_0_16), .Q(\Memory[0] [62]), 
      .QN());
   DFF_X1 \Memory_reg[0][61]  (.D(Memory[61]), .CK(n_0_16), .Q(\Memory[0] [61]), 
      .QN());
   DFF_X1 \Memory_reg[0][60]  (.D(Memory[60]), .CK(n_0_16), .Q(\Memory[0] [60]), 
      .QN());
   DFF_X1 \Memory_reg[0][59]  (.D(Memory[59]), .CK(n_0_16), .Q(\Memory[0] [59]), 
      .QN());
   DFF_X1 \Memory_reg[0][58]  (.D(Memory[58]), .CK(n_0_16), .Q(\Memory[0] [58]), 
      .QN());
   DFF_X1 \Memory_reg[0][57]  (.D(Memory[57]), .CK(n_0_16), .Q(\Memory[0] [57]), 
      .QN());
   DFF_X1 \Memory_reg[0][56]  (.D(Memory[56]), .CK(n_0_16), .Q(\Memory[0] [56]), 
      .QN());
   DFF_X1 \Memory_reg[0][55]  (.D(Memory[55]), .CK(n_0_16), .Q(\Memory[0] [55]), 
      .QN());
   DFF_X1 \Memory_reg[0][54]  (.D(Memory[54]), .CK(n_0_16), .Q(\Memory[0] [54]), 
      .QN());
   DFF_X1 \Memory_reg[0][53]  (.D(Memory[53]), .CK(n_0_16), .Q(\Memory[0] [53]), 
      .QN());
   DFF_X1 \Memory_reg[0][52]  (.D(Memory[52]), .CK(n_0_16), .Q(\Memory[0] [52]), 
      .QN());
   DFF_X1 \Memory_reg[0][51]  (.D(Memory[51]), .CK(n_0_16), .Q(\Memory[0] [51]), 
      .QN());
   DFF_X1 \Memory_reg[0][50]  (.D(Memory[50]), .CK(n_0_16), .Q(\Memory[0] [50]), 
      .QN());
   DFF_X1 \Memory_reg[0][49]  (.D(Memory[49]), .CK(n_0_16), .Q(\Memory[0] [49]), 
      .QN());
   DFF_X1 \Memory_reg[0][48]  (.D(Memory[48]), .CK(n_0_16), .Q(\Memory[0] [48]), 
      .QN());
   DFF_X1 \Memory_reg[0][47]  (.D(Memory[47]), .CK(n_0_16), .Q(\Memory[0] [47]), 
      .QN());
   DFF_X1 \Memory_reg[0][46]  (.D(Memory[46]), .CK(n_0_16), .Q(\Memory[0] [46]), 
      .QN());
   DFF_X1 \Memory_reg[0][45]  (.D(Memory[45]), .CK(n_0_16), .Q(\Memory[0] [45]), 
      .QN());
   DFF_X1 \Memory_reg[0][44]  (.D(Memory[44]), .CK(n_0_16), .Q(\Memory[0] [44]), 
      .QN());
   DFF_X1 \Memory_reg[0][43]  (.D(Memory[43]), .CK(n_0_16), .Q(\Memory[0] [43]), 
      .QN());
   DFF_X1 \Memory_reg[0][42]  (.D(Memory[42]), .CK(n_0_16), .Q(\Memory[0] [42]), 
      .QN());
   DFF_X1 \Memory_reg[0][41]  (.D(Memory[41]), .CK(n_0_16), .Q(\Memory[0] [41]), 
      .QN());
   DFF_X1 \Memory_reg[0][40]  (.D(Memory[40]), .CK(n_0_16), .Q(\Memory[0] [40]), 
      .QN());
   DFF_X1 \Memory_reg[0][39]  (.D(Memory[39]), .CK(n_0_16), .Q(\Memory[0] [39]), 
      .QN());
   DFF_X1 \Memory_reg[0][38]  (.D(Memory[38]), .CK(n_0_16), .Q(\Memory[0] [38]), 
      .QN());
   DFF_X1 \Memory_reg[0][37]  (.D(Memory[37]), .CK(n_0_16), .Q(\Memory[0] [37]), 
      .QN());
   DFF_X1 \Memory_reg[0][36]  (.D(Memory[36]), .CK(n_0_16), .Q(\Memory[0] [36]), 
      .QN());
   DFF_X1 \Memory_reg[0][35]  (.D(Memory[35]), .CK(n_0_16), .Q(\Memory[0] [35]), 
      .QN());
   DFF_X1 \Memory_reg[0][34]  (.D(Memory[34]), .CK(n_0_16), .Q(\Memory[0] [34]), 
      .QN());
   DFF_X1 \Memory_reg[0][33]  (.D(Memory[33]), .CK(n_0_16), .Q(\Memory[0] [33]), 
      .QN());
   DFF_X1 \Memory_reg[0][32]  (.D(Memory[32]), .CK(n_0_16), .Q(\Memory[0] [32]), 
      .QN());
   DFF_X1 \Memory_reg[0][31]  (.D(Memory[31]), .CK(n_0_16), .Q(\Memory[0] [31]), 
      .QN());
   DFF_X1 \Memory_reg[0][30]  (.D(Memory[30]), .CK(n_0_16), .Q(\Memory[0] [30]), 
      .QN());
   DFF_X1 \Memory_reg[0][29]  (.D(Memory[29]), .CK(n_0_16), .Q(\Memory[0] [29]), 
      .QN());
   DFF_X1 \Memory_reg[0][28]  (.D(Memory[28]), .CK(n_0_16), .Q(\Memory[0] [28]), 
      .QN());
   DFF_X1 \Memory_reg[0][27]  (.D(Memory[27]), .CK(n_0_16), .Q(\Memory[0] [27]), 
      .QN());
   DFF_X1 \Memory_reg[0][26]  (.D(Memory[26]), .CK(n_0_16), .Q(\Memory[0] [26]), 
      .QN());
   DFF_X1 \Memory_reg[0][25]  (.D(Memory[25]), .CK(n_0_16), .Q(\Memory[0] [25]), 
      .QN());
   DFF_X1 \Memory_reg[0][24]  (.D(Memory[24]), .CK(n_0_16), .Q(\Memory[0] [24]), 
      .QN());
   DFF_X1 \Memory_reg[0][23]  (.D(Memory[23]), .CK(n_0_16), .Q(\Memory[0] [23]), 
      .QN());
   DFF_X1 \Memory_reg[0][22]  (.D(Memory[22]), .CK(n_0_16), .Q(\Memory[0] [22]), 
      .QN());
   DFF_X1 \Memory_reg[0][21]  (.D(Memory[21]), .CK(n_0_16), .Q(\Memory[0] [21]), 
      .QN());
   DFF_X1 \Memory_reg[0][20]  (.D(Memory[20]), .CK(n_0_16), .Q(\Memory[0] [20]), 
      .QN());
   DFF_X1 \Memory_reg[0][19]  (.D(Memory[19]), .CK(n_0_16), .Q(\Memory[0] [19]), 
      .QN());
   DFF_X1 \Memory_reg[0][18]  (.D(Memory[18]), .CK(n_0_16), .Q(\Memory[0] [18]), 
      .QN());
   DFF_X1 \Memory_reg[0][17]  (.D(Memory[17]), .CK(n_0_16), .Q(\Memory[0] [17]), 
      .QN());
   DFF_X1 \Memory_reg[0][16]  (.D(Memory[16]), .CK(n_0_16), .Q(\Memory[0] [16]), 
      .QN());
   DFF_X1 \Memory_reg[0][15]  (.D(Memory[15]), .CK(n_0_16), .Q(\Memory[0] [15]), 
      .QN());
   DFF_X1 \Memory_reg[0][14]  (.D(Memory[14]), .CK(n_0_16), .Q(\Memory[0] [14]), 
      .QN());
   DFF_X1 \Memory_reg[0][13]  (.D(Memory[13]), .CK(n_0_16), .Q(\Memory[0] [13]), 
      .QN());
   DFF_X1 \Memory_reg[0][12]  (.D(Memory[12]), .CK(n_0_16), .Q(\Memory[0] [12]), 
      .QN());
   DFF_X1 \Memory_reg[0][11]  (.D(Memory[11]), .CK(n_0_16), .Q(\Memory[0] [11]), 
      .QN());
   DFF_X1 \Memory_reg[0][10]  (.D(Memory[10]), .CK(n_0_16), .Q(\Memory[0] [10]), 
      .QN());
   DFF_X1 \Memory_reg[0][9]  (.D(Memory[9]), .CK(n_0_16), .Q(\Memory[0] [9]), 
      .QN());
   DFF_X1 \Memory_reg[0][8]  (.D(Memory[8]), .CK(n_0_16), .Q(\Memory[0] [8]), 
      .QN());
   DFF_X1 \Memory_reg[0][7]  (.D(Memory[7]), .CK(n_0_16), .Q(\Memory[0] [7]), 
      .QN());
   DFF_X1 \Memory_reg[0][6]  (.D(Memory[6]), .CK(n_0_16), .Q(\Memory[0] [6]), 
      .QN());
   DFF_X1 \Memory_reg[0][5]  (.D(Memory[5]), .CK(n_0_16), .Q(\Memory[0] [5]), 
      .QN());
   DFF_X1 \Memory_reg[0][4]  (.D(Memory[4]), .CK(n_0_16), .Q(\Memory[0] [4]), 
      .QN());
   DFF_X1 \Memory_reg[0][3]  (.D(Memory[3]), .CK(n_0_16), .Q(\Memory[0] [3]), 
      .QN());
   DFF_X1 \Memory_reg[0][2]  (.D(Memory[2]), .CK(n_0_16), .Q(\Memory[0] [2]), 
      .QN());
   DFF_X1 \Memory_reg[0][1]  (.D(Memory[1]), .CK(n_0_16), .Q(\Memory[0] [1]), 
      .QN());
   DFF_X1 \Memory_reg[0][0]  (.D(Memory[0]), .CK(n_0_16), .Q(\Memory[0] [0]), 
      .QN());
   INV_X1 i_0_0_0 (.A(n_0_0_0), .ZN(n_0_34));
   NAND3_X1 i_0_0_1 (.A1(n_0_0_12), .A2(n_0_0_8), .A3(n_0_0_22), .ZN(n_0_0_0));
   INV_X1 i_0_0_2 (.A(n_0_0_1), .ZN(n_0_35));
   NAND3_X1 i_0_0_3 (.A1(n_0_0_12), .A2(n_0_0_8), .A3(address_RD1[0]), .ZN(
      n_0_0_1));
   INV_X1 i_0_0_4 (.A(n_0_0_2), .ZN(n_0_36));
   NAND4_X1 i_0_0_5 (.A1(n_0_0_8), .A2(n_0_0_26), .A3(address_RD1[1]), .A4(
      n_0_0_22), .ZN(n_0_0_2));
   INV_X1 i_0_0_6 (.A(n_0_0_3), .ZN(n_0_37));
   NAND4_X1 i_0_0_7 (.A1(n_0_0_8), .A2(n_0_0_26), .A3(address_RD1[1]), .A4(
      address_RD1[0]), .ZN(n_0_0_3));
   INV_X1 i_0_0_8 (.A(n_0_0_4), .ZN(n_0_38));
   NAND4_X1 i_0_0_9 (.A1(n_0_0_8), .A2(address_RD1[2]), .A3(n_0_0_25), .A4(
      n_0_0_22), .ZN(n_0_0_4));
   INV_X1 i_0_0_10 (.A(n_0_0_5), .ZN(n_0_39));
   NAND4_X1 i_0_0_11 (.A1(n_0_0_8), .A2(address_RD1[2]), .A3(n_0_0_25), .A4(
      address_RD1[0]), .ZN(n_0_0_5));
   INV_X1 i_0_0_12 (.A(n_0_0_6), .ZN(n_0_40));
   NAND4_X1 i_0_0_13 (.A1(n_0_0_8), .A2(address_RD1[2]), .A3(address_RD1[1]), 
      .A4(n_0_0_22), .ZN(n_0_0_6));
   INV_X1 i_0_0_14 (.A(n_0_0_7), .ZN(n_0_41));
   NAND4_X1 i_0_0_15 (.A1(n_0_0_8), .A2(address_RD1[2]), .A3(address_RD1[1]), 
      .A4(address_RD1[0]), .ZN(n_0_0_7));
   INV_X1 i_0_0_16 (.A(n_0_0_9), .ZN(n_0_0_8));
   NAND2_X1 i_0_0_17 (.A1(n_0_0_20), .A2(n_0_0_23), .ZN(n_0_0_9));
   INV_X1 i_0_0_18 (.A(n_0_0_10), .ZN(n_0_42));
   NAND3_X1 i_0_0_19 (.A1(n_0_0_12), .A2(n_0_0_17), .A3(n_0_0_22), .ZN(n_0_0_10));
   INV_X1 i_0_0_20 (.A(n_0_0_11), .ZN(n_0_43));
   NAND3_X1 i_0_0_21 (.A1(n_0_0_12), .A2(n_0_0_17), .A3(address_RD1[0]), 
      .ZN(n_0_0_11));
   INV_X1 i_0_0_22 (.A(n_0_0_24), .ZN(n_0_0_12));
   INV_X1 i_0_0_23 (.A(n_0_0_13), .ZN(n_0_44));
   NAND4_X1 i_0_0_24 (.A1(n_0_0_17), .A2(n_0_0_26), .A3(address_RD1[1]), 
      .A4(n_0_0_22), .ZN(n_0_0_13));
   INV_X1 i_0_0_25 (.A(n_0_0_14), .ZN(n_0_45));
   NAND4_X1 i_0_0_26 (.A1(n_0_0_17), .A2(n_0_0_26), .A3(address_RD1[1]), 
      .A4(address_RD1[0]), .ZN(n_0_0_14));
   INV_X1 i_0_0_27 (.A(n_0_0_15), .ZN(n_0_46));
   NAND4_X1 i_0_0_28 (.A1(n_0_0_17), .A2(address_RD1[2]), .A3(n_0_0_25), 
      .A4(n_0_0_22), .ZN(n_0_0_15));
   INV_X1 i_0_0_29 (.A(n_0_0_16), .ZN(n_0_47));
   NAND4_X1 i_0_0_30 (.A1(n_0_0_17), .A2(address_RD1[2]), .A3(n_0_0_25), 
      .A4(address_RD1[0]), .ZN(n_0_0_16));
   INV_X1 i_0_0_31 (.A(n_0_0_18), .ZN(n_0_0_17));
   NAND2_X1 i_0_0_32 (.A1(n_0_0_20), .A2(address_RD1[3]), .ZN(n_0_0_18));
   NOR2_X1 i_0_0_33 (.A1(n_0_0_19), .A2(address_RD1[0]), .ZN(n_0_48));
   NOR2_X1 i_0_0_34 (.A1(n_0_0_19), .A2(n_0_0_22), .ZN(n_0_49));
   NAND4_X1 i_0_0_35 (.A1(n_0_0_20), .A2(address_RD1[3]), .A3(address_RD1[2]), 
      .A4(address_RD1[1]), .ZN(n_0_0_19));
   INV_X1 i_0_0_36 (.A(address_RD1[4]), .ZN(n_0_0_20));
   NOR2_X1 i_0_0_37 (.A1(n_0_0_21), .A2(n_0_0_24), .ZN(n_0_50));
   NAND3_X1 i_0_0_38 (.A1(n_0_0_23), .A2(n_0_0_22), .A3(address_RD1[4]), 
      .ZN(n_0_0_21));
   INV_X1 i_0_0_39 (.A(address_RD1[0]), .ZN(n_0_0_22));
   INV_X1 i_0_0_40 (.A(address_RD1[3]), .ZN(n_0_0_23));
   NAND2_X1 i_0_0_41 (.A1(n_0_0_26), .A2(n_0_0_25), .ZN(n_0_0_24));
   INV_X1 i_0_0_42 (.A(address_RD1[1]), .ZN(n_0_0_25));
   INV_X1 i_0_0_43 (.A(address_RD1[2]), .ZN(n_0_0_26));
   NAND2_X1 i_0_2_0 (.A1(n_0_38), .A2(\Memory[4] [0]), .ZN(n_0_2_0));
   NAND2_X1 i_0_2_1 (.A1(n_0_41), .A2(\Memory[7] [0]), .ZN(n_0_2_1));
   NAND2_X1 i_0_2_2 (.A1(n_0_37), .A2(\Memory[3] [0]), .ZN(n_0_2_2));
   NAND2_X1 i_0_2_3 (.A1(n_0_36), .A2(\Memory[2] [0]), .ZN(n_0_2_3));
   NAND4_X1 i_0_2_4 (.A1(n_0_2_0), .A2(n_0_2_1), .A3(n_0_2_2), .A4(n_0_2_3), 
      .ZN(n_0_2_4));
   INV_X1 i_0_2_5 (.A(n_0_2_4), .ZN(n_0_2_5));
   NAND2_X1 i_0_2_6 (.A1(n_0_50), .A2(\Memory[16] [0]), .ZN(n_0_2_6));
   NAND2_X1 i_0_2_7 (.A1(n_0_40), .A2(\Memory[6] [0]), .ZN(n_0_2_7));
   NAND2_X1 i_0_2_8 (.A1(n_0_39), .A2(\Memory[5] [0]), .ZN(n_0_2_8));
   NAND3_X1 i_0_2_9 (.A1(n_0_2_6), .A2(n_0_2_7), .A3(n_0_2_8), .ZN(n_0_2_9));
   NAND2_X1 i_0_2_10 (.A1(n_0_42), .A2(\Memory[8] [0]), .ZN(n_0_2_10));
   NAND2_X1 i_0_2_11 (.A1(n_0_35), .A2(\Memory[1] [0]), .ZN(n_0_2_11));
   NAND2_X1 i_0_2_12 (.A1(n_0_44), .A2(\Memory[10] [0]), .ZN(n_0_2_12));
   NAND3_X1 i_0_2_13 (.A1(n_0_2_10), .A2(n_0_2_11), .A3(n_0_2_12), .ZN(n_0_2_13));
   NOR2_X1 i_0_2_14 (.A1(n_0_2_9), .A2(n_0_2_13), .ZN(n_0_2_14));
   NAND2_X1 i_0_2_15 (.A1(n_0_48), .A2(\Memory[14] [0]), .ZN(n_0_2_15));
   NAND2_X1 i_0_2_16 (.A1(n_0_49), .A2(\Memory[15] [0]), .ZN(n_0_2_16));
   NAND2_X1 i_0_2_17 (.A1(n_0_34), .A2(\Memory[0] [0]), .ZN(n_0_2_17));
   NAND2_X1 i_0_2_18 (.A1(n_0_43), .A2(\Memory[9] [0]), .ZN(n_0_2_18));
   NAND4_X1 i_0_2_19 (.A1(n_0_2_15), .A2(n_0_2_16), .A3(n_0_2_17), .A4(n_0_2_18), 
      .ZN(n_0_2_19));
   NAND2_X1 i_0_2_20 (.A1(n_0_47), .A2(\Memory[13] [0]), .ZN(n_0_2_20));
   NAND2_X1 i_0_2_21 (.A1(n_0_46), .A2(\Memory[12] [0]), .ZN(n_0_2_21));
   NAND2_X1 i_0_2_22 (.A1(n_0_45), .A2(\Memory[11] [0]), .ZN(n_0_2_22));
   NAND3_X1 i_0_2_23 (.A1(n_0_2_20), .A2(n_0_2_21), .A3(n_0_2_22), .ZN(n_0_2_23));
   NOR2_X1 i_0_2_24 (.A1(n_0_2_19), .A2(n_0_2_23), .ZN(n_0_2_24));
   NAND3_X1 i_0_2_25 (.A1(n_0_2_5), .A2(n_0_2_14), .A3(n_0_2_24), .ZN(
      dataOut1[0]));
   NAND2_X1 i_0_2_26 (.A1(n_0_38), .A2(\Memory[4] [1]), .ZN(n_0_2_25));
   NAND2_X1 i_0_2_27 (.A1(n_0_41), .A2(\Memory[7] [1]), .ZN(n_0_2_26));
   NAND2_X1 i_0_2_28 (.A1(n_0_37), .A2(\Memory[3] [1]), .ZN(n_0_2_27));
   NAND2_X1 i_0_2_29 (.A1(n_0_36), .A2(\Memory[2] [1]), .ZN(n_0_2_28));
   NAND4_X1 i_0_2_30 (.A1(n_0_2_25), .A2(n_0_2_26), .A3(n_0_2_27), .A4(n_0_2_28), 
      .ZN(n_0_2_29));
   INV_X1 i_0_2_31 (.A(n_0_2_29), .ZN(n_0_2_30));
   NAND2_X1 i_0_2_32 (.A1(n_0_50), .A2(\Memory[16] [1]), .ZN(n_0_2_31));
   NAND2_X1 i_0_2_33 (.A1(n_0_40), .A2(\Memory[6] [1]), .ZN(n_0_2_32));
   NAND2_X1 i_0_2_34 (.A1(n_0_39), .A2(\Memory[5] [1]), .ZN(n_0_2_33));
   NAND3_X1 i_0_2_35 (.A1(n_0_2_31), .A2(n_0_2_32), .A3(n_0_2_33), .ZN(n_0_2_34));
   NAND2_X1 i_0_2_36 (.A1(n_0_42), .A2(\Memory[8] [1]), .ZN(n_0_2_35));
   NAND2_X1 i_0_2_37 (.A1(n_0_35), .A2(\Memory[1] [1]), .ZN(n_0_2_36));
   NAND2_X1 i_0_2_38 (.A1(n_0_44), .A2(\Memory[10] [1]), .ZN(n_0_2_37));
   NAND3_X1 i_0_2_39 (.A1(n_0_2_35), .A2(n_0_2_36), .A3(n_0_2_37), .ZN(n_0_2_38));
   NOR2_X1 i_0_2_40 (.A1(n_0_2_34), .A2(n_0_2_38), .ZN(n_0_2_39));
   NAND2_X1 i_0_2_41 (.A1(n_0_48), .A2(\Memory[14] [1]), .ZN(n_0_2_40));
   NAND2_X1 i_0_2_42 (.A1(n_0_49), .A2(\Memory[15] [1]), .ZN(n_0_2_41));
   NAND2_X1 i_0_2_43 (.A1(n_0_34), .A2(\Memory[0] [1]), .ZN(n_0_2_42));
   NAND2_X1 i_0_2_44 (.A1(n_0_43), .A2(\Memory[9] [1]), .ZN(n_0_2_43));
   NAND4_X1 i_0_2_45 (.A1(n_0_2_40), .A2(n_0_2_41), .A3(n_0_2_42), .A4(n_0_2_43), 
      .ZN(n_0_2_44));
   NAND2_X1 i_0_2_46 (.A1(n_0_47), .A2(\Memory[13] [1]), .ZN(n_0_2_45));
   NAND2_X1 i_0_2_47 (.A1(n_0_46), .A2(\Memory[12] [1]), .ZN(n_0_2_46));
   NAND2_X1 i_0_2_48 (.A1(n_0_45), .A2(\Memory[11] [1]), .ZN(n_0_2_47));
   NAND3_X1 i_0_2_49 (.A1(n_0_2_45), .A2(n_0_2_46), .A3(n_0_2_47), .ZN(n_0_2_48));
   NOR2_X1 i_0_2_50 (.A1(n_0_2_44), .A2(n_0_2_48), .ZN(n_0_2_49));
   NAND3_X1 i_0_2_51 (.A1(n_0_2_30), .A2(n_0_2_39), .A3(n_0_2_49), .ZN(
      dataOut1[1]));
   NAND2_X1 i_0_2_52 (.A1(n_0_38), .A2(\Memory[4] [2]), .ZN(n_0_2_50));
   NAND2_X1 i_0_2_53 (.A1(n_0_41), .A2(\Memory[7] [2]), .ZN(n_0_2_51));
   NAND2_X1 i_0_2_54 (.A1(n_0_37), .A2(\Memory[3] [2]), .ZN(n_0_2_52));
   NAND2_X1 i_0_2_55 (.A1(n_0_36), .A2(\Memory[2] [2]), .ZN(n_0_2_53));
   NAND4_X1 i_0_2_56 (.A1(n_0_2_50), .A2(n_0_2_51), .A3(n_0_2_52), .A4(n_0_2_53), 
      .ZN(n_0_2_54));
   INV_X1 i_0_2_57 (.A(n_0_2_54), .ZN(n_0_2_55));
   NAND2_X1 i_0_2_58 (.A1(n_0_50), .A2(\Memory[16] [2]), .ZN(n_0_2_56));
   NAND2_X1 i_0_2_59 (.A1(n_0_40), .A2(\Memory[6] [2]), .ZN(n_0_2_57));
   NAND2_X1 i_0_2_60 (.A1(n_0_39), .A2(\Memory[5] [2]), .ZN(n_0_2_58));
   NAND3_X1 i_0_2_61 (.A1(n_0_2_56), .A2(n_0_2_57), .A3(n_0_2_58), .ZN(n_0_2_59));
   NAND2_X1 i_0_2_62 (.A1(n_0_42), .A2(\Memory[8] [2]), .ZN(n_0_2_60));
   NAND2_X1 i_0_2_63 (.A1(n_0_35), .A2(\Memory[1] [2]), .ZN(n_0_2_61));
   NAND2_X1 i_0_2_64 (.A1(n_0_44), .A2(\Memory[10] [2]), .ZN(n_0_2_62));
   NAND3_X1 i_0_2_65 (.A1(n_0_2_60), .A2(n_0_2_61), .A3(n_0_2_62), .ZN(n_0_2_63));
   NOR2_X1 i_0_2_66 (.A1(n_0_2_59), .A2(n_0_2_63), .ZN(n_0_2_64));
   NAND2_X1 i_0_2_67 (.A1(n_0_48), .A2(\Memory[14] [2]), .ZN(n_0_2_65));
   NAND2_X1 i_0_2_68 (.A1(n_0_49), .A2(\Memory[15] [2]), .ZN(n_0_2_66));
   NAND2_X1 i_0_2_69 (.A1(n_0_34), .A2(\Memory[0] [2]), .ZN(n_0_2_67));
   NAND2_X1 i_0_2_70 (.A1(n_0_43), .A2(\Memory[9] [2]), .ZN(n_0_2_68));
   NAND4_X1 i_0_2_71 (.A1(n_0_2_65), .A2(n_0_2_66), .A3(n_0_2_67), .A4(n_0_2_68), 
      .ZN(n_0_2_69));
   NAND2_X1 i_0_2_72 (.A1(n_0_47), .A2(\Memory[13] [2]), .ZN(n_0_2_70));
   NAND2_X1 i_0_2_73 (.A1(n_0_46), .A2(\Memory[12] [2]), .ZN(n_0_2_71));
   NAND2_X1 i_0_2_74 (.A1(n_0_45), .A2(\Memory[11] [2]), .ZN(n_0_2_72));
   NAND3_X1 i_0_2_75 (.A1(n_0_2_70), .A2(n_0_2_71), .A3(n_0_2_72), .ZN(n_0_2_73));
   NOR2_X1 i_0_2_76 (.A1(n_0_2_69), .A2(n_0_2_73), .ZN(n_0_2_74));
   NAND3_X1 i_0_2_77 (.A1(n_0_2_55), .A2(n_0_2_64), .A3(n_0_2_74), .ZN(
      dataOut1[2]));
   NAND2_X1 i_0_2_78 (.A1(n_0_38), .A2(\Memory[4] [3]), .ZN(n_0_2_75));
   NAND2_X1 i_0_2_79 (.A1(n_0_41), .A2(\Memory[7] [3]), .ZN(n_0_2_76));
   NAND2_X1 i_0_2_80 (.A1(n_0_37), .A2(\Memory[3] [3]), .ZN(n_0_2_77));
   NAND2_X1 i_0_2_81 (.A1(n_0_36), .A2(\Memory[2] [3]), .ZN(n_0_2_78));
   NAND4_X1 i_0_2_82 (.A1(n_0_2_75), .A2(n_0_2_76), .A3(n_0_2_77), .A4(n_0_2_78), 
      .ZN(n_0_2_79));
   INV_X1 i_0_2_83 (.A(n_0_2_79), .ZN(n_0_2_80));
   NAND2_X1 i_0_2_84 (.A1(n_0_50), .A2(\Memory[16] [3]), .ZN(n_0_2_81));
   NAND2_X1 i_0_2_85 (.A1(n_0_40), .A2(\Memory[6] [3]), .ZN(n_0_2_82));
   NAND2_X1 i_0_2_86 (.A1(n_0_39), .A2(\Memory[5] [3]), .ZN(n_0_2_83));
   NAND3_X1 i_0_2_87 (.A1(n_0_2_81), .A2(n_0_2_82), .A3(n_0_2_83), .ZN(n_0_2_84));
   NAND2_X1 i_0_2_88 (.A1(n_0_42), .A2(\Memory[8] [3]), .ZN(n_0_2_85));
   NAND2_X1 i_0_2_89 (.A1(n_0_35), .A2(\Memory[1] [3]), .ZN(n_0_2_86));
   NAND2_X1 i_0_2_90 (.A1(n_0_44), .A2(\Memory[10] [3]), .ZN(n_0_2_87));
   NAND3_X1 i_0_2_91 (.A1(n_0_2_85), .A2(n_0_2_86), .A3(n_0_2_87), .ZN(n_0_2_88));
   NOR2_X1 i_0_2_92 (.A1(n_0_2_84), .A2(n_0_2_88), .ZN(n_0_2_89));
   NAND2_X1 i_0_2_93 (.A1(n_0_48), .A2(\Memory[14] [3]), .ZN(n_0_2_90));
   NAND2_X1 i_0_2_94 (.A1(n_0_49), .A2(\Memory[15] [3]), .ZN(n_0_2_91));
   NAND2_X1 i_0_2_95 (.A1(n_0_34), .A2(\Memory[0] [3]), .ZN(n_0_2_92));
   NAND2_X1 i_0_2_96 (.A1(n_0_43), .A2(\Memory[9] [3]), .ZN(n_0_2_93));
   NAND4_X1 i_0_2_97 (.A1(n_0_2_90), .A2(n_0_2_91), .A3(n_0_2_92), .A4(n_0_2_93), 
      .ZN(n_0_2_94));
   NAND2_X1 i_0_2_98 (.A1(n_0_47), .A2(\Memory[13] [3]), .ZN(n_0_2_95));
   NAND2_X1 i_0_2_99 (.A1(n_0_46), .A2(\Memory[12] [3]), .ZN(n_0_2_96));
   NAND2_X1 i_0_2_100 (.A1(n_0_45), .A2(\Memory[11] [3]), .ZN(n_0_2_97));
   NAND3_X1 i_0_2_101 (.A1(n_0_2_95), .A2(n_0_2_96), .A3(n_0_2_97), .ZN(n_0_2_98));
   NOR2_X1 i_0_2_102 (.A1(n_0_2_94), .A2(n_0_2_98), .ZN(n_0_2_99));
   NAND3_X1 i_0_2_103 (.A1(n_0_2_80), .A2(n_0_2_89), .A3(n_0_2_99), .ZN(
      dataOut1[3]));
   NAND2_X1 i_0_2_104 (.A1(n_0_38), .A2(\Memory[4] [4]), .ZN(n_0_2_100));
   NAND2_X1 i_0_2_105 (.A1(n_0_41), .A2(\Memory[7] [4]), .ZN(n_0_2_101));
   NAND2_X1 i_0_2_106 (.A1(n_0_37), .A2(\Memory[3] [4]), .ZN(n_0_2_102));
   NAND2_X1 i_0_2_107 (.A1(n_0_36), .A2(\Memory[2] [4]), .ZN(n_0_2_103));
   NAND4_X1 i_0_2_108 (.A1(n_0_2_100), .A2(n_0_2_101), .A3(n_0_2_102), .A4(
      n_0_2_103), .ZN(n_0_2_104));
   INV_X1 i_0_2_109 (.A(n_0_2_104), .ZN(n_0_2_105));
   NAND2_X1 i_0_2_110 (.A1(n_0_50), .A2(\Memory[16] [4]), .ZN(n_0_2_106));
   NAND2_X1 i_0_2_111 (.A1(n_0_40), .A2(\Memory[6] [4]), .ZN(n_0_2_107));
   NAND2_X1 i_0_2_112 (.A1(n_0_39), .A2(\Memory[5] [4]), .ZN(n_0_2_108));
   NAND3_X1 i_0_2_113 (.A1(n_0_2_106), .A2(n_0_2_107), .A3(n_0_2_108), .ZN(
      n_0_2_109));
   NAND2_X1 i_0_2_114 (.A1(n_0_42), .A2(\Memory[8] [4]), .ZN(n_0_2_110));
   NAND2_X1 i_0_2_115 (.A1(n_0_35), .A2(\Memory[1] [4]), .ZN(n_0_2_111));
   NAND2_X1 i_0_2_116 (.A1(n_0_44), .A2(\Memory[10] [4]), .ZN(n_0_2_112));
   NAND3_X1 i_0_2_117 (.A1(n_0_2_110), .A2(n_0_2_111), .A3(n_0_2_112), .ZN(
      n_0_2_113));
   NOR2_X1 i_0_2_118 (.A1(n_0_2_109), .A2(n_0_2_113), .ZN(n_0_2_114));
   NAND2_X1 i_0_2_119 (.A1(n_0_48), .A2(\Memory[14] [4]), .ZN(n_0_2_115));
   NAND2_X1 i_0_2_120 (.A1(n_0_49), .A2(\Memory[15] [4]), .ZN(n_0_2_116));
   NAND2_X1 i_0_2_121 (.A1(n_0_34), .A2(\Memory[0] [4]), .ZN(n_0_2_117));
   NAND2_X1 i_0_2_122 (.A1(n_0_43), .A2(\Memory[9] [4]), .ZN(n_0_2_118));
   NAND4_X1 i_0_2_123 (.A1(n_0_2_115), .A2(n_0_2_116), .A3(n_0_2_117), .A4(
      n_0_2_118), .ZN(n_0_2_119));
   NAND2_X1 i_0_2_124 (.A1(n_0_47), .A2(\Memory[13] [4]), .ZN(n_0_2_120));
   NAND2_X1 i_0_2_125 (.A1(n_0_46), .A2(\Memory[12] [4]), .ZN(n_0_2_121));
   NAND2_X1 i_0_2_126 (.A1(n_0_45), .A2(\Memory[11] [4]), .ZN(n_0_2_122));
   NAND3_X1 i_0_2_127 (.A1(n_0_2_120), .A2(n_0_2_121), .A3(n_0_2_122), .ZN(
      n_0_2_123));
   NOR2_X1 i_0_2_128 (.A1(n_0_2_119), .A2(n_0_2_123), .ZN(n_0_2_124));
   NAND3_X1 i_0_2_129 (.A1(n_0_2_105), .A2(n_0_2_114), .A3(n_0_2_124), .ZN(
      dataOut1[4]));
   NAND2_X1 i_0_2_130 (.A1(n_0_38), .A2(\Memory[4] [5]), .ZN(n_0_2_125));
   NAND2_X1 i_0_2_131 (.A1(n_0_41), .A2(\Memory[7] [5]), .ZN(n_0_2_126));
   NAND2_X1 i_0_2_132 (.A1(n_0_37), .A2(\Memory[3] [5]), .ZN(n_0_2_127));
   NAND2_X1 i_0_2_133 (.A1(n_0_36), .A2(\Memory[2] [5]), .ZN(n_0_2_128));
   NAND4_X1 i_0_2_134 (.A1(n_0_2_125), .A2(n_0_2_126), .A3(n_0_2_127), .A4(
      n_0_2_128), .ZN(n_0_2_129));
   INV_X1 i_0_2_135 (.A(n_0_2_129), .ZN(n_0_2_130));
   NAND2_X1 i_0_2_136 (.A1(n_0_50), .A2(\Memory[16] [5]), .ZN(n_0_2_131));
   NAND2_X1 i_0_2_137 (.A1(n_0_40), .A2(\Memory[6] [5]), .ZN(n_0_2_132));
   NAND2_X1 i_0_2_138 (.A1(n_0_39), .A2(\Memory[5] [5]), .ZN(n_0_2_133));
   NAND3_X1 i_0_2_139 (.A1(n_0_2_131), .A2(n_0_2_132), .A3(n_0_2_133), .ZN(
      n_0_2_134));
   NAND2_X1 i_0_2_140 (.A1(n_0_42), .A2(\Memory[8] [5]), .ZN(n_0_2_135));
   NAND2_X1 i_0_2_141 (.A1(n_0_35), .A2(\Memory[1] [5]), .ZN(n_0_2_136));
   NAND2_X1 i_0_2_142 (.A1(n_0_44), .A2(\Memory[10] [5]), .ZN(n_0_2_137));
   NAND3_X1 i_0_2_143 (.A1(n_0_2_135), .A2(n_0_2_136), .A3(n_0_2_137), .ZN(
      n_0_2_138));
   NOR2_X1 i_0_2_144 (.A1(n_0_2_134), .A2(n_0_2_138), .ZN(n_0_2_139));
   NAND2_X1 i_0_2_145 (.A1(n_0_48), .A2(\Memory[14] [5]), .ZN(n_0_2_140));
   NAND2_X1 i_0_2_146 (.A1(n_0_49), .A2(\Memory[15] [5]), .ZN(n_0_2_141));
   NAND2_X1 i_0_2_147 (.A1(n_0_34), .A2(\Memory[0] [5]), .ZN(n_0_2_142));
   NAND2_X1 i_0_2_148 (.A1(n_0_43), .A2(\Memory[9] [5]), .ZN(n_0_2_143));
   NAND4_X1 i_0_2_149 (.A1(n_0_2_140), .A2(n_0_2_141), .A3(n_0_2_142), .A4(
      n_0_2_143), .ZN(n_0_2_144));
   NAND2_X1 i_0_2_150 (.A1(n_0_47), .A2(\Memory[13] [5]), .ZN(n_0_2_145));
   NAND2_X1 i_0_2_151 (.A1(n_0_46), .A2(\Memory[12] [5]), .ZN(n_0_2_146));
   NAND2_X1 i_0_2_152 (.A1(n_0_45), .A2(\Memory[11] [5]), .ZN(n_0_2_147));
   NAND3_X1 i_0_2_153 (.A1(n_0_2_145), .A2(n_0_2_146), .A3(n_0_2_147), .ZN(
      n_0_2_148));
   NOR2_X1 i_0_2_154 (.A1(n_0_2_144), .A2(n_0_2_148), .ZN(n_0_2_149));
   NAND3_X1 i_0_2_155 (.A1(n_0_2_130), .A2(n_0_2_139), .A3(n_0_2_149), .ZN(
      dataOut1[5]));
   NAND2_X1 i_0_2_156 (.A1(n_0_38), .A2(\Memory[4] [6]), .ZN(n_0_2_150));
   NAND2_X1 i_0_2_157 (.A1(n_0_41), .A2(\Memory[7] [6]), .ZN(n_0_2_151));
   NAND2_X1 i_0_2_158 (.A1(n_0_37), .A2(\Memory[3] [6]), .ZN(n_0_2_152));
   NAND2_X1 i_0_2_159 (.A1(n_0_36), .A2(\Memory[2] [6]), .ZN(n_0_2_153));
   NAND4_X1 i_0_2_160 (.A1(n_0_2_150), .A2(n_0_2_151), .A3(n_0_2_152), .A4(
      n_0_2_153), .ZN(n_0_2_154));
   INV_X1 i_0_2_161 (.A(n_0_2_154), .ZN(n_0_2_155));
   NAND2_X1 i_0_2_162 (.A1(n_0_50), .A2(\Memory[16] [6]), .ZN(n_0_2_156));
   NAND2_X1 i_0_2_163 (.A1(n_0_40), .A2(\Memory[6] [6]), .ZN(n_0_2_157));
   NAND2_X1 i_0_2_164 (.A1(n_0_39), .A2(\Memory[5] [6]), .ZN(n_0_2_158));
   NAND3_X1 i_0_2_165 (.A1(n_0_2_156), .A2(n_0_2_157), .A3(n_0_2_158), .ZN(
      n_0_2_159));
   NAND2_X1 i_0_2_166 (.A1(n_0_42), .A2(\Memory[8] [6]), .ZN(n_0_2_160));
   NAND2_X1 i_0_2_167 (.A1(n_0_35), .A2(\Memory[1] [6]), .ZN(n_0_2_161));
   NAND2_X1 i_0_2_168 (.A1(n_0_44), .A2(\Memory[10] [6]), .ZN(n_0_2_162));
   NAND3_X1 i_0_2_169 (.A1(n_0_2_160), .A2(n_0_2_161), .A3(n_0_2_162), .ZN(
      n_0_2_163));
   NOR2_X1 i_0_2_170 (.A1(n_0_2_159), .A2(n_0_2_163), .ZN(n_0_2_164));
   NAND2_X1 i_0_2_171 (.A1(n_0_48), .A2(\Memory[14] [6]), .ZN(n_0_2_165));
   NAND2_X1 i_0_2_172 (.A1(n_0_49), .A2(\Memory[15] [6]), .ZN(n_0_2_166));
   NAND2_X1 i_0_2_173 (.A1(n_0_34), .A2(\Memory[0] [6]), .ZN(n_0_2_167));
   NAND2_X1 i_0_2_174 (.A1(n_0_43), .A2(\Memory[9] [6]), .ZN(n_0_2_168));
   NAND4_X1 i_0_2_175 (.A1(n_0_2_165), .A2(n_0_2_166), .A3(n_0_2_167), .A4(
      n_0_2_168), .ZN(n_0_2_169));
   NAND2_X1 i_0_2_176 (.A1(n_0_47), .A2(\Memory[13] [6]), .ZN(n_0_2_170));
   NAND2_X1 i_0_2_177 (.A1(n_0_46), .A2(\Memory[12] [6]), .ZN(n_0_2_171));
   NAND2_X1 i_0_2_178 (.A1(n_0_45), .A2(\Memory[11] [6]), .ZN(n_0_2_172));
   NAND3_X1 i_0_2_179 (.A1(n_0_2_170), .A2(n_0_2_171), .A3(n_0_2_172), .ZN(
      n_0_2_173));
   NOR2_X1 i_0_2_180 (.A1(n_0_2_169), .A2(n_0_2_173), .ZN(n_0_2_174));
   NAND3_X1 i_0_2_181 (.A1(n_0_2_155), .A2(n_0_2_164), .A3(n_0_2_174), .ZN(
      dataOut1[6]));
   NAND2_X1 i_0_2_182 (.A1(n_0_38), .A2(\Memory[4] [7]), .ZN(n_0_2_175));
   NAND2_X1 i_0_2_183 (.A1(n_0_41), .A2(\Memory[7] [7]), .ZN(n_0_2_176));
   NAND2_X1 i_0_2_184 (.A1(n_0_37), .A2(\Memory[3] [7]), .ZN(n_0_2_177));
   NAND2_X1 i_0_2_185 (.A1(n_0_36), .A2(\Memory[2] [7]), .ZN(n_0_2_178));
   NAND4_X1 i_0_2_186 (.A1(n_0_2_175), .A2(n_0_2_176), .A3(n_0_2_177), .A4(
      n_0_2_178), .ZN(n_0_2_179));
   INV_X1 i_0_2_187 (.A(n_0_2_179), .ZN(n_0_2_180));
   NAND2_X1 i_0_2_188 (.A1(n_0_50), .A2(\Memory[16] [7]), .ZN(n_0_2_181));
   NAND2_X1 i_0_2_189 (.A1(n_0_40), .A2(\Memory[6] [7]), .ZN(n_0_2_182));
   NAND2_X1 i_0_2_190 (.A1(n_0_39), .A2(\Memory[5] [7]), .ZN(n_0_2_183));
   NAND3_X1 i_0_2_191 (.A1(n_0_2_181), .A2(n_0_2_182), .A3(n_0_2_183), .ZN(
      n_0_2_184));
   NAND2_X1 i_0_2_192 (.A1(n_0_42), .A2(\Memory[8] [7]), .ZN(n_0_2_185));
   NAND2_X1 i_0_2_193 (.A1(n_0_35), .A2(\Memory[1] [7]), .ZN(n_0_2_186));
   NAND2_X1 i_0_2_194 (.A1(n_0_44), .A2(\Memory[10] [7]), .ZN(n_0_2_187));
   NAND3_X1 i_0_2_195 (.A1(n_0_2_185), .A2(n_0_2_186), .A3(n_0_2_187), .ZN(
      n_0_2_188));
   NOR2_X1 i_0_2_196 (.A1(n_0_2_184), .A2(n_0_2_188), .ZN(n_0_2_189));
   NAND2_X1 i_0_2_197 (.A1(n_0_48), .A2(\Memory[14] [7]), .ZN(n_0_2_190));
   NAND2_X1 i_0_2_198 (.A1(n_0_49), .A2(\Memory[15] [7]), .ZN(n_0_2_191));
   NAND2_X1 i_0_2_199 (.A1(n_0_34), .A2(\Memory[0] [7]), .ZN(n_0_2_192));
   NAND2_X1 i_0_2_200 (.A1(n_0_43), .A2(\Memory[9] [7]), .ZN(n_0_2_193));
   NAND4_X1 i_0_2_201 (.A1(n_0_2_190), .A2(n_0_2_191), .A3(n_0_2_192), .A4(
      n_0_2_193), .ZN(n_0_2_194));
   NAND2_X1 i_0_2_202 (.A1(n_0_47), .A2(\Memory[13] [7]), .ZN(n_0_2_195));
   NAND2_X1 i_0_2_203 (.A1(n_0_46), .A2(\Memory[12] [7]), .ZN(n_0_2_196));
   NAND2_X1 i_0_2_204 (.A1(n_0_45), .A2(\Memory[11] [7]), .ZN(n_0_2_197));
   NAND3_X1 i_0_2_205 (.A1(n_0_2_195), .A2(n_0_2_196), .A3(n_0_2_197), .ZN(
      n_0_2_198));
   NOR2_X1 i_0_2_206 (.A1(n_0_2_194), .A2(n_0_2_198), .ZN(n_0_2_199));
   NAND3_X1 i_0_2_207 (.A1(n_0_2_180), .A2(n_0_2_189), .A3(n_0_2_199), .ZN(
      dataOut1[7]));
   NAND2_X1 i_0_2_208 (.A1(n_0_38), .A2(\Memory[4] [8]), .ZN(n_0_2_200));
   NAND2_X1 i_0_2_209 (.A1(n_0_41), .A2(\Memory[7] [8]), .ZN(n_0_2_201));
   NAND2_X1 i_0_2_210 (.A1(n_0_37), .A2(\Memory[3] [8]), .ZN(n_0_2_202));
   NAND2_X1 i_0_2_211 (.A1(n_0_36), .A2(\Memory[2] [8]), .ZN(n_0_2_203));
   NAND4_X1 i_0_2_212 (.A1(n_0_2_200), .A2(n_0_2_201), .A3(n_0_2_202), .A4(
      n_0_2_203), .ZN(n_0_2_204));
   INV_X1 i_0_2_213 (.A(n_0_2_204), .ZN(n_0_2_205));
   NAND2_X1 i_0_2_214 (.A1(n_0_50), .A2(\Memory[16] [8]), .ZN(n_0_2_206));
   NAND2_X1 i_0_2_215 (.A1(n_0_40), .A2(\Memory[6] [8]), .ZN(n_0_2_207));
   NAND2_X1 i_0_2_216 (.A1(n_0_39), .A2(\Memory[5] [8]), .ZN(n_0_2_208));
   NAND3_X1 i_0_2_217 (.A1(n_0_2_206), .A2(n_0_2_207), .A3(n_0_2_208), .ZN(
      n_0_2_209));
   NAND2_X1 i_0_2_218 (.A1(n_0_42), .A2(\Memory[8] [8]), .ZN(n_0_2_210));
   NAND2_X1 i_0_2_219 (.A1(n_0_35), .A2(\Memory[1] [8]), .ZN(n_0_2_211));
   NAND2_X1 i_0_2_220 (.A1(n_0_44), .A2(\Memory[10] [8]), .ZN(n_0_2_212));
   NAND3_X1 i_0_2_221 (.A1(n_0_2_210), .A2(n_0_2_211), .A3(n_0_2_212), .ZN(
      n_0_2_213));
   NOR2_X1 i_0_2_222 (.A1(n_0_2_209), .A2(n_0_2_213), .ZN(n_0_2_214));
   NAND2_X1 i_0_2_223 (.A1(n_0_48), .A2(\Memory[14] [8]), .ZN(n_0_2_215));
   NAND2_X1 i_0_2_224 (.A1(n_0_49), .A2(\Memory[15] [8]), .ZN(n_0_2_216));
   NAND2_X1 i_0_2_225 (.A1(n_0_34), .A2(\Memory[0] [8]), .ZN(n_0_2_217));
   NAND2_X1 i_0_2_226 (.A1(n_0_43), .A2(\Memory[9] [8]), .ZN(n_0_2_218));
   NAND4_X1 i_0_2_227 (.A1(n_0_2_215), .A2(n_0_2_216), .A3(n_0_2_217), .A4(
      n_0_2_218), .ZN(n_0_2_219));
   NAND2_X1 i_0_2_228 (.A1(n_0_47), .A2(\Memory[13] [8]), .ZN(n_0_2_220));
   NAND2_X1 i_0_2_229 (.A1(n_0_46), .A2(\Memory[12] [8]), .ZN(n_0_2_221));
   NAND2_X1 i_0_2_230 (.A1(n_0_45), .A2(\Memory[11] [8]), .ZN(n_0_2_222));
   NAND3_X1 i_0_2_231 (.A1(n_0_2_220), .A2(n_0_2_221), .A3(n_0_2_222), .ZN(
      n_0_2_223));
   NOR2_X1 i_0_2_232 (.A1(n_0_2_219), .A2(n_0_2_223), .ZN(n_0_2_224));
   NAND3_X1 i_0_2_233 (.A1(n_0_2_205), .A2(n_0_2_214), .A3(n_0_2_224), .ZN(
      dataOut1[8]));
   NAND2_X1 i_0_2_234 (.A1(n_0_38), .A2(\Memory[4] [9]), .ZN(n_0_2_225));
   NAND2_X1 i_0_2_235 (.A1(n_0_41), .A2(\Memory[7] [9]), .ZN(n_0_2_226));
   NAND2_X1 i_0_2_236 (.A1(n_0_37), .A2(\Memory[3] [9]), .ZN(n_0_2_227));
   NAND2_X1 i_0_2_237 (.A1(n_0_36), .A2(\Memory[2] [9]), .ZN(n_0_2_228));
   NAND4_X1 i_0_2_238 (.A1(n_0_2_225), .A2(n_0_2_226), .A3(n_0_2_227), .A4(
      n_0_2_228), .ZN(n_0_2_229));
   INV_X1 i_0_2_239 (.A(n_0_2_229), .ZN(n_0_2_230));
   NAND2_X1 i_0_2_240 (.A1(n_0_50), .A2(\Memory[16] [9]), .ZN(n_0_2_231));
   NAND2_X1 i_0_2_241 (.A1(n_0_40), .A2(\Memory[6] [9]), .ZN(n_0_2_232));
   NAND2_X1 i_0_2_242 (.A1(n_0_39), .A2(\Memory[5] [9]), .ZN(n_0_2_233));
   NAND3_X1 i_0_2_243 (.A1(n_0_2_231), .A2(n_0_2_232), .A3(n_0_2_233), .ZN(
      n_0_2_234));
   NAND2_X1 i_0_2_244 (.A1(n_0_42), .A2(\Memory[8] [9]), .ZN(n_0_2_235));
   NAND2_X1 i_0_2_245 (.A1(n_0_35), .A2(\Memory[1] [9]), .ZN(n_0_2_236));
   NAND2_X1 i_0_2_246 (.A1(n_0_44), .A2(\Memory[10] [9]), .ZN(n_0_2_237));
   NAND3_X1 i_0_2_247 (.A1(n_0_2_235), .A2(n_0_2_236), .A3(n_0_2_237), .ZN(
      n_0_2_238));
   NOR2_X1 i_0_2_248 (.A1(n_0_2_234), .A2(n_0_2_238), .ZN(n_0_2_239));
   NAND2_X1 i_0_2_249 (.A1(n_0_48), .A2(\Memory[14] [9]), .ZN(n_0_2_240));
   NAND2_X1 i_0_2_250 (.A1(n_0_49), .A2(\Memory[15] [9]), .ZN(n_0_2_241));
   NAND2_X1 i_0_2_251 (.A1(n_0_34), .A2(\Memory[0] [9]), .ZN(n_0_2_242));
   NAND2_X1 i_0_2_252 (.A1(n_0_43), .A2(\Memory[9] [9]), .ZN(n_0_2_243));
   NAND4_X1 i_0_2_253 (.A1(n_0_2_240), .A2(n_0_2_241), .A3(n_0_2_242), .A4(
      n_0_2_243), .ZN(n_0_2_244));
   NAND2_X1 i_0_2_254 (.A1(n_0_47), .A2(\Memory[13] [9]), .ZN(n_0_2_245));
   NAND2_X1 i_0_2_255 (.A1(n_0_46), .A2(\Memory[12] [9]), .ZN(n_0_2_246));
   NAND2_X1 i_0_2_256 (.A1(n_0_45), .A2(\Memory[11] [9]), .ZN(n_0_2_247));
   NAND3_X1 i_0_2_257 (.A1(n_0_2_245), .A2(n_0_2_246), .A3(n_0_2_247), .ZN(
      n_0_2_248));
   NOR2_X1 i_0_2_258 (.A1(n_0_2_244), .A2(n_0_2_248), .ZN(n_0_2_249));
   NAND3_X1 i_0_2_259 (.A1(n_0_2_230), .A2(n_0_2_239), .A3(n_0_2_249), .ZN(
      dataOut1[9]));
   NAND2_X1 i_0_2_260 (.A1(n_0_38), .A2(\Memory[4] [10]), .ZN(n_0_2_250));
   NAND2_X1 i_0_2_261 (.A1(n_0_41), .A2(\Memory[7] [10]), .ZN(n_0_2_251));
   NAND2_X1 i_0_2_262 (.A1(n_0_37), .A2(\Memory[3] [10]), .ZN(n_0_2_252));
   NAND2_X1 i_0_2_263 (.A1(n_0_36), .A2(\Memory[2] [10]), .ZN(n_0_2_253));
   NAND4_X1 i_0_2_264 (.A1(n_0_2_250), .A2(n_0_2_251), .A3(n_0_2_252), .A4(
      n_0_2_253), .ZN(n_0_2_254));
   INV_X1 i_0_2_265 (.A(n_0_2_254), .ZN(n_0_2_255));
   NAND2_X1 i_0_2_266 (.A1(n_0_50), .A2(\Memory[16] [10]), .ZN(n_0_2_256));
   NAND2_X1 i_0_2_267 (.A1(n_0_40), .A2(\Memory[6] [10]), .ZN(n_0_2_257));
   NAND2_X1 i_0_2_268 (.A1(n_0_39), .A2(\Memory[5] [10]), .ZN(n_0_2_258));
   NAND3_X1 i_0_2_269 (.A1(n_0_2_256), .A2(n_0_2_257), .A3(n_0_2_258), .ZN(
      n_0_2_259));
   NAND2_X1 i_0_2_270 (.A1(n_0_42), .A2(\Memory[8] [10]), .ZN(n_0_2_260));
   NAND2_X1 i_0_2_271 (.A1(n_0_35), .A2(\Memory[1] [10]), .ZN(n_0_2_261));
   NAND2_X1 i_0_2_272 (.A1(n_0_44), .A2(\Memory[10] [10]), .ZN(n_0_2_262));
   NAND3_X1 i_0_2_273 (.A1(n_0_2_260), .A2(n_0_2_261), .A3(n_0_2_262), .ZN(
      n_0_2_263));
   NOR2_X1 i_0_2_274 (.A1(n_0_2_259), .A2(n_0_2_263), .ZN(n_0_2_264));
   NAND2_X1 i_0_2_275 (.A1(n_0_48), .A2(\Memory[14] [10]), .ZN(n_0_2_265));
   NAND2_X1 i_0_2_276 (.A1(n_0_49), .A2(\Memory[15] [10]), .ZN(n_0_2_266));
   NAND2_X1 i_0_2_277 (.A1(n_0_34), .A2(\Memory[0] [10]), .ZN(n_0_2_267));
   NAND2_X1 i_0_2_278 (.A1(n_0_43), .A2(\Memory[9] [10]), .ZN(n_0_2_268));
   NAND4_X1 i_0_2_279 (.A1(n_0_2_265), .A2(n_0_2_266), .A3(n_0_2_267), .A4(
      n_0_2_268), .ZN(n_0_2_269));
   NAND2_X1 i_0_2_280 (.A1(n_0_47), .A2(\Memory[13] [10]), .ZN(n_0_2_270));
   NAND2_X1 i_0_2_281 (.A1(n_0_46), .A2(\Memory[12] [10]), .ZN(n_0_2_271));
   NAND2_X1 i_0_2_282 (.A1(n_0_45), .A2(\Memory[11] [10]), .ZN(n_0_2_272));
   NAND3_X1 i_0_2_283 (.A1(n_0_2_270), .A2(n_0_2_271), .A3(n_0_2_272), .ZN(
      n_0_2_273));
   NOR2_X1 i_0_2_284 (.A1(n_0_2_269), .A2(n_0_2_273), .ZN(n_0_2_274));
   NAND3_X1 i_0_2_285 (.A1(n_0_2_255), .A2(n_0_2_264), .A3(n_0_2_274), .ZN(
      dataOut1[10]));
   NAND2_X1 i_0_2_286 (.A1(n_0_38), .A2(\Memory[4] [11]), .ZN(n_0_2_275));
   NAND2_X1 i_0_2_287 (.A1(n_0_41), .A2(\Memory[7] [11]), .ZN(n_0_2_276));
   NAND2_X1 i_0_2_288 (.A1(n_0_37), .A2(\Memory[3] [11]), .ZN(n_0_2_277));
   NAND2_X1 i_0_2_289 (.A1(n_0_36), .A2(\Memory[2] [11]), .ZN(n_0_2_278));
   NAND4_X1 i_0_2_290 (.A1(n_0_2_275), .A2(n_0_2_276), .A3(n_0_2_277), .A4(
      n_0_2_278), .ZN(n_0_2_279));
   INV_X1 i_0_2_291 (.A(n_0_2_279), .ZN(n_0_2_280));
   NAND2_X1 i_0_2_292 (.A1(n_0_50), .A2(\Memory[16] [11]), .ZN(n_0_2_281));
   NAND2_X1 i_0_2_293 (.A1(n_0_40), .A2(\Memory[6] [11]), .ZN(n_0_2_282));
   NAND2_X1 i_0_2_294 (.A1(n_0_39), .A2(\Memory[5] [11]), .ZN(n_0_2_283));
   NAND3_X1 i_0_2_295 (.A1(n_0_2_281), .A2(n_0_2_282), .A3(n_0_2_283), .ZN(
      n_0_2_284));
   NAND2_X1 i_0_2_296 (.A1(n_0_42), .A2(\Memory[8] [11]), .ZN(n_0_2_285));
   NAND2_X1 i_0_2_297 (.A1(n_0_35), .A2(\Memory[1] [11]), .ZN(n_0_2_286));
   NAND2_X1 i_0_2_298 (.A1(n_0_44), .A2(\Memory[10] [11]), .ZN(n_0_2_287));
   NAND3_X1 i_0_2_299 (.A1(n_0_2_285), .A2(n_0_2_286), .A3(n_0_2_287), .ZN(
      n_0_2_288));
   NOR2_X1 i_0_2_300 (.A1(n_0_2_284), .A2(n_0_2_288), .ZN(n_0_2_289));
   NAND2_X1 i_0_2_301 (.A1(n_0_48), .A2(\Memory[14] [11]), .ZN(n_0_2_290));
   NAND2_X1 i_0_2_302 (.A1(n_0_49), .A2(\Memory[15] [11]), .ZN(n_0_2_291));
   NAND2_X1 i_0_2_303 (.A1(n_0_34), .A2(\Memory[0] [11]), .ZN(n_0_2_292));
   NAND2_X1 i_0_2_304 (.A1(n_0_43), .A2(\Memory[9] [11]), .ZN(n_0_2_293));
   NAND4_X1 i_0_2_305 (.A1(n_0_2_290), .A2(n_0_2_291), .A3(n_0_2_292), .A4(
      n_0_2_293), .ZN(n_0_2_294));
   NAND2_X1 i_0_2_306 (.A1(n_0_47), .A2(\Memory[13] [11]), .ZN(n_0_2_295));
   NAND2_X1 i_0_2_307 (.A1(n_0_46), .A2(\Memory[12] [11]), .ZN(n_0_2_296));
   NAND2_X1 i_0_2_308 (.A1(n_0_45), .A2(\Memory[11] [11]), .ZN(n_0_2_297));
   NAND3_X1 i_0_2_309 (.A1(n_0_2_295), .A2(n_0_2_296), .A3(n_0_2_297), .ZN(
      n_0_2_298));
   NOR2_X1 i_0_2_310 (.A1(n_0_2_294), .A2(n_0_2_298), .ZN(n_0_2_299));
   NAND3_X1 i_0_2_311 (.A1(n_0_2_280), .A2(n_0_2_289), .A3(n_0_2_299), .ZN(
      dataOut1[11]));
   NAND2_X1 i_0_2_312 (.A1(n_0_38), .A2(\Memory[4] [12]), .ZN(n_0_2_300));
   NAND2_X1 i_0_2_313 (.A1(n_0_41), .A2(\Memory[7] [12]), .ZN(n_0_2_301));
   NAND2_X1 i_0_2_314 (.A1(n_0_37), .A2(\Memory[3] [12]), .ZN(n_0_2_302));
   NAND2_X1 i_0_2_315 (.A1(n_0_36), .A2(\Memory[2] [12]), .ZN(n_0_2_303));
   NAND4_X1 i_0_2_316 (.A1(n_0_2_300), .A2(n_0_2_301), .A3(n_0_2_302), .A4(
      n_0_2_303), .ZN(n_0_2_304));
   INV_X1 i_0_2_317 (.A(n_0_2_304), .ZN(n_0_2_305));
   NAND2_X1 i_0_2_318 (.A1(n_0_50), .A2(\Memory[16] [12]), .ZN(n_0_2_306));
   NAND2_X1 i_0_2_319 (.A1(n_0_40), .A2(\Memory[6] [12]), .ZN(n_0_2_307));
   NAND2_X1 i_0_2_320 (.A1(n_0_39), .A2(\Memory[5] [12]), .ZN(n_0_2_308));
   NAND3_X1 i_0_2_321 (.A1(n_0_2_306), .A2(n_0_2_307), .A3(n_0_2_308), .ZN(
      n_0_2_309));
   NAND2_X1 i_0_2_322 (.A1(n_0_42), .A2(\Memory[8] [12]), .ZN(n_0_2_310));
   NAND2_X1 i_0_2_323 (.A1(n_0_35), .A2(\Memory[1] [12]), .ZN(n_0_2_311));
   NAND2_X1 i_0_2_324 (.A1(n_0_44), .A2(\Memory[10] [12]), .ZN(n_0_2_312));
   NAND3_X1 i_0_2_325 (.A1(n_0_2_310), .A2(n_0_2_311), .A3(n_0_2_312), .ZN(
      n_0_2_313));
   NOR2_X1 i_0_2_326 (.A1(n_0_2_309), .A2(n_0_2_313), .ZN(n_0_2_314));
   NAND2_X1 i_0_2_327 (.A1(n_0_48), .A2(\Memory[14] [12]), .ZN(n_0_2_315));
   NAND2_X1 i_0_2_328 (.A1(n_0_49), .A2(\Memory[15] [12]), .ZN(n_0_2_316));
   NAND2_X1 i_0_2_329 (.A1(n_0_34), .A2(\Memory[0] [12]), .ZN(n_0_2_317));
   NAND2_X1 i_0_2_330 (.A1(n_0_43), .A2(\Memory[9] [12]), .ZN(n_0_2_318));
   NAND4_X1 i_0_2_331 (.A1(n_0_2_315), .A2(n_0_2_316), .A3(n_0_2_317), .A4(
      n_0_2_318), .ZN(n_0_2_319));
   NAND2_X1 i_0_2_332 (.A1(n_0_47), .A2(\Memory[13] [12]), .ZN(n_0_2_320));
   NAND2_X1 i_0_2_333 (.A1(n_0_46), .A2(\Memory[12] [12]), .ZN(n_0_2_321));
   NAND2_X1 i_0_2_334 (.A1(n_0_45), .A2(\Memory[11] [12]), .ZN(n_0_2_322));
   NAND3_X1 i_0_2_335 (.A1(n_0_2_320), .A2(n_0_2_321), .A3(n_0_2_322), .ZN(
      n_0_2_323));
   NOR2_X1 i_0_2_336 (.A1(n_0_2_319), .A2(n_0_2_323), .ZN(n_0_2_324));
   NAND3_X1 i_0_2_337 (.A1(n_0_2_305), .A2(n_0_2_314), .A3(n_0_2_324), .ZN(
      dataOut1[12]));
   NAND2_X1 i_0_2_338 (.A1(n_0_38), .A2(\Memory[4] [13]), .ZN(n_0_2_325));
   NAND2_X1 i_0_2_339 (.A1(n_0_41), .A2(\Memory[7] [13]), .ZN(n_0_2_326));
   NAND2_X1 i_0_2_340 (.A1(n_0_37), .A2(\Memory[3] [13]), .ZN(n_0_2_327));
   NAND2_X1 i_0_2_341 (.A1(n_0_36), .A2(\Memory[2] [13]), .ZN(n_0_2_328));
   NAND4_X1 i_0_2_342 (.A1(n_0_2_325), .A2(n_0_2_326), .A3(n_0_2_327), .A4(
      n_0_2_328), .ZN(n_0_2_329));
   INV_X1 i_0_2_343 (.A(n_0_2_329), .ZN(n_0_2_330));
   NAND2_X1 i_0_2_344 (.A1(n_0_50), .A2(\Memory[16] [13]), .ZN(n_0_2_331));
   NAND2_X1 i_0_2_345 (.A1(n_0_40), .A2(\Memory[6] [13]), .ZN(n_0_2_332));
   NAND2_X1 i_0_2_346 (.A1(n_0_39), .A2(\Memory[5] [13]), .ZN(n_0_2_333));
   NAND3_X1 i_0_2_347 (.A1(n_0_2_331), .A2(n_0_2_332), .A3(n_0_2_333), .ZN(
      n_0_2_334));
   NAND2_X1 i_0_2_348 (.A1(n_0_42), .A2(\Memory[8] [13]), .ZN(n_0_2_335));
   NAND2_X1 i_0_2_349 (.A1(n_0_35), .A2(\Memory[1] [13]), .ZN(n_0_2_336));
   NAND2_X1 i_0_2_350 (.A1(n_0_44), .A2(\Memory[10] [13]), .ZN(n_0_2_337));
   NAND3_X1 i_0_2_351 (.A1(n_0_2_335), .A2(n_0_2_336), .A3(n_0_2_337), .ZN(
      n_0_2_338));
   NOR2_X1 i_0_2_352 (.A1(n_0_2_334), .A2(n_0_2_338), .ZN(n_0_2_339));
   NAND2_X1 i_0_2_353 (.A1(n_0_48), .A2(\Memory[14] [13]), .ZN(n_0_2_340));
   NAND2_X1 i_0_2_354 (.A1(n_0_49), .A2(\Memory[15] [13]), .ZN(n_0_2_341));
   NAND2_X1 i_0_2_355 (.A1(n_0_34), .A2(\Memory[0] [13]), .ZN(n_0_2_342));
   NAND2_X1 i_0_2_356 (.A1(n_0_43), .A2(\Memory[9] [13]), .ZN(n_0_2_343));
   NAND4_X1 i_0_2_357 (.A1(n_0_2_340), .A2(n_0_2_341), .A3(n_0_2_342), .A4(
      n_0_2_343), .ZN(n_0_2_344));
   NAND2_X1 i_0_2_358 (.A1(n_0_47), .A2(\Memory[13] [13]), .ZN(n_0_2_345));
   NAND2_X1 i_0_2_359 (.A1(n_0_46), .A2(\Memory[12] [13]), .ZN(n_0_2_346));
   NAND2_X1 i_0_2_360 (.A1(n_0_45), .A2(\Memory[11] [13]), .ZN(n_0_2_347));
   NAND3_X1 i_0_2_361 (.A1(n_0_2_345), .A2(n_0_2_346), .A3(n_0_2_347), .ZN(
      n_0_2_348));
   NOR2_X1 i_0_2_362 (.A1(n_0_2_344), .A2(n_0_2_348), .ZN(n_0_2_349));
   NAND3_X1 i_0_2_363 (.A1(n_0_2_330), .A2(n_0_2_339), .A3(n_0_2_349), .ZN(
      dataOut1[13]));
   NAND2_X1 i_0_2_364 (.A1(n_0_38), .A2(\Memory[4] [14]), .ZN(n_0_2_350));
   NAND2_X1 i_0_2_365 (.A1(n_0_41), .A2(\Memory[7] [14]), .ZN(n_0_2_351));
   NAND2_X1 i_0_2_366 (.A1(n_0_37), .A2(\Memory[3] [14]), .ZN(n_0_2_352));
   NAND2_X1 i_0_2_367 (.A1(n_0_36), .A2(\Memory[2] [14]), .ZN(n_0_2_353));
   NAND4_X1 i_0_2_368 (.A1(n_0_2_350), .A2(n_0_2_351), .A3(n_0_2_352), .A4(
      n_0_2_353), .ZN(n_0_2_354));
   INV_X1 i_0_2_369 (.A(n_0_2_354), .ZN(n_0_2_355));
   NAND2_X1 i_0_2_370 (.A1(n_0_50), .A2(\Memory[16] [14]), .ZN(n_0_2_356));
   NAND2_X1 i_0_2_371 (.A1(n_0_40), .A2(\Memory[6] [14]), .ZN(n_0_2_357));
   NAND2_X1 i_0_2_372 (.A1(n_0_39), .A2(\Memory[5] [14]), .ZN(n_0_2_358));
   NAND3_X1 i_0_2_373 (.A1(n_0_2_356), .A2(n_0_2_357), .A3(n_0_2_358), .ZN(
      n_0_2_359));
   NAND2_X1 i_0_2_374 (.A1(n_0_42), .A2(\Memory[8] [14]), .ZN(n_0_2_360));
   NAND2_X1 i_0_2_375 (.A1(n_0_35), .A2(\Memory[1] [14]), .ZN(n_0_2_361));
   NAND2_X1 i_0_2_376 (.A1(n_0_44), .A2(\Memory[10] [14]), .ZN(n_0_2_362));
   NAND3_X1 i_0_2_377 (.A1(n_0_2_360), .A2(n_0_2_361), .A3(n_0_2_362), .ZN(
      n_0_2_363));
   NOR2_X1 i_0_2_378 (.A1(n_0_2_359), .A2(n_0_2_363), .ZN(n_0_2_364));
   NAND2_X1 i_0_2_379 (.A1(n_0_48), .A2(\Memory[14] [14]), .ZN(n_0_2_365));
   NAND2_X1 i_0_2_380 (.A1(n_0_49), .A2(\Memory[15] [14]), .ZN(n_0_2_366));
   NAND2_X1 i_0_2_381 (.A1(n_0_34), .A2(\Memory[0] [14]), .ZN(n_0_2_367));
   NAND2_X1 i_0_2_382 (.A1(n_0_43), .A2(\Memory[9] [14]), .ZN(n_0_2_368));
   NAND4_X1 i_0_2_383 (.A1(n_0_2_365), .A2(n_0_2_366), .A3(n_0_2_367), .A4(
      n_0_2_368), .ZN(n_0_2_369));
   NAND2_X1 i_0_2_384 (.A1(n_0_47), .A2(\Memory[13] [14]), .ZN(n_0_2_370));
   NAND2_X1 i_0_2_385 (.A1(n_0_46), .A2(\Memory[12] [14]), .ZN(n_0_2_371));
   NAND2_X1 i_0_2_386 (.A1(n_0_45), .A2(\Memory[11] [14]), .ZN(n_0_2_372));
   NAND3_X1 i_0_2_387 (.A1(n_0_2_370), .A2(n_0_2_371), .A3(n_0_2_372), .ZN(
      n_0_2_373));
   NOR2_X1 i_0_2_388 (.A1(n_0_2_369), .A2(n_0_2_373), .ZN(n_0_2_374));
   NAND3_X1 i_0_2_389 (.A1(n_0_2_355), .A2(n_0_2_364), .A3(n_0_2_374), .ZN(
      dataOut1[14]));
   NAND2_X1 i_0_2_390 (.A1(n_0_38), .A2(\Memory[4] [15]), .ZN(n_0_2_375));
   NAND2_X1 i_0_2_391 (.A1(n_0_41), .A2(\Memory[7] [15]), .ZN(n_0_2_376));
   NAND2_X1 i_0_2_392 (.A1(n_0_37), .A2(\Memory[3] [15]), .ZN(n_0_2_377));
   NAND2_X1 i_0_2_393 (.A1(n_0_36), .A2(\Memory[2] [15]), .ZN(n_0_2_378));
   NAND4_X1 i_0_2_394 (.A1(n_0_2_375), .A2(n_0_2_376), .A3(n_0_2_377), .A4(
      n_0_2_378), .ZN(n_0_2_379));
   INV_X1 i_0_2_395 (.A(n_0_2_379), .ZN(n_0_2_380));
   NAND2_X1 i_0_2_396 (.A1(n_0_50), .A2(\Memory[16] [15]), .ZN(n_0_2_381));
   NAND2_X1 i_0_2_397 (.A1(n_0_40), .A2(\Memory[6] [15]), .ZN(n_0_2_382));
   NAND2_X1 i_0_2_398 (.A1(n_0_39), .A2(\Memory[5] [15]), .ZN(n_0_2_383));
   NAND3_X1 i_0_2_399 (.A1(n_0_2_381), .A2(n_0_2_382), .A3(n_0_2_383), .ZN(
      n_0_2_384));
   NAND2_X1 i_0_2_400 (.A1(n_0_42), .A2(\Memory[8] [15]), .ZN(n_0_2_385));
   NAND2_X1 i_0_2_401 (.A1(n_0_35), .A2(\Memory[1] [15]), .ZN(n_0_2_386));
   NAND2_X1 i_0_2_402 (.A1(n_0_44), .A2(\Memory[10] [15]), .ZN(n_0_2_387));
   NAND3_X1 i_0_2_403 (.A1(n_0_2_385), .A2(n_0_2_386), .A3(n_0_2_387), .ZN(
      n_0_2_388));
   NOR2_X1 i_0_2_404 (.A1(n_0_2_384), .A2(n_0_2_388), .ZN(n_0_2_389));
   NAND2_X1 i_0_2_405 (.A1(n_0_48), .A2(\Memory[14] [15]), .ZN(n_0_2_390));
   NAND2_X1 i_0_2_406 (.A1(n_0_49), .A2(\Memory[15] [15]), .ZN(n_0_2_391));
   NAND2_X1 i_0_2_407 (.A1(n_0_34), .A2(\Memory[0] [15]), .ZN(n_0_2_392));
   NAND2_X1 i_0_2_408 (.A1(n_0_43), .A2(\Memory[9] [15]), .ZN(n_0_2_393));
   NAND4_X1 i_0_2_409 (.A1(n_0_2_390), .A2(n_0_2_391), .A3(n_0_2_392), .A4(
      n_0_2_393), .ZN(n_0_2_394));
   NAND2_X1 i_0_2_410 (.A1(n_0_47), .A2(\Memory[13] [15]), .ZN(n_0_2_395));
   NAND2_X1 i_0_2_411 (.A1(n_0_46), .A2(\Memory[12] [15]), .ZN(n_0_2_396));
   NAND2_X1 i_0_2_412 (.A1(n_0_45), .A2(\Memory[11] [15]), .ZN(n_0_2_397));
   NAND3_X1 i_0_2_413 (.A1(n_0_2_395), .A2(n_0_2_396), .A3(n_0_2_397), .ZN(
      n_0_2_398));
   NOR2_X1 i_0_2_414 (.A1(n_0_2_394), .A2(n_0_2_398), .ZN(n_0_2_399));
   NAND3_X1 i_0_2_415 (.A1(n_0_2_380), .A2(n_0_2_389), .A3(n_0_2_399), .ZN(
      dataOut1[15]));
   NAND2_X1 i_0_2_416 (.A1(n_0_38), .A2(\Memory[4] [16]), .ZN(n_0_2_400));
   NAND2_X1 i_0_2_417 (.A1(n_0_41), .A2(\Memory[7] [16]), .ZN(n_0_2_401));
   NAND2_X1 i_0_2_418 (.A1(n_0_37), .A2(\Memory[3] [16]), .ZN(n_0_2_402));
   NAND2_X1 i_0_2_419 (.A1(n_0_36), .A2(\Memory[2] [16]), .ZN(n_0_2_403));
   NAND4_X1 i_0_2_420 (.A1(n_0_2_400), .A2(n_0_2_401), .A3(n_0_2_402), .A4(
      n_0_2_403), .ZN(n_0_2_404));
   INV_X1 i_0_2_421 (.A(n_0_2_404), .ZN(n_0_2_405));
   NAND2_X1 i_0_2_422 (.A1(n_0_50), .A2(\Memory[16] [16]), .ZN(n_0_2_406));
   NAND2_X1 i_0_2_423 (.A1(n_0_40), .A2(\Memory[6] [16]), .ZN(n_0_2_407));
   NAND2_X1 i_0_2_424 (.A1(n_0_39), .A2(\Memory[5] [16]), .ZN(n_0_2_408));
   NAND3_X1 i_0_2_425 (.A1(n_0_2_406), .A2(n_0_2_407), .A3(n_0_2_408), .ZN(
      n_0_2_409));
   NAND2_X1 i_0_2_426 (.A1(n_0_42), .A2(\Memory[8] [16]), .ZN(n_0_2_410));
   NAND2_X1 i_0_2_427 (.A1(n_0_35), .A2(\Memory[1] [16]), .ZN(n_0_2_411));
   NAND2_X1 i_0_2_428 (.A1(n_0_44), .A2(\Memory[10] [16]), .ZN(n_0_2_412));
   NAND3_X1 i_0_2_429 (.A1(n_0_2_410), .A2(n_0_2_411), .A3(n_0_2_412), .ZN(
      n_0_2_413));
   NOR2_X1 i_0_2_430 (.A1(n_0_2_409), .A2(n_0_2_413), .ZN(n_0_2_414));
   NAND2_X1 i_0_2_431 (.A1(n_0_48), .A2(\Memory[14] [16]), .ZN(n_0_2_415));
   NAND2_X1 i_0_2_432 (.A1(n_0_49), .A2(\Memory[15] [16]), .ZN(n_0_2_416));
   NAND2_X1 i_0_2_433 (.A1(n_0_34), .A2(\Memory[0] [16]), .ZN(n_0_2_417));
   NAND2_X1 i_0_2_434 (.A1(n_0_43), .A2(\Memory[9] [16]), .ZN(n_0_2_418));
   NAND4_X1 i_0_2_435 (.A1(n_0_2_415), .A2(n_0_2_416), .A3(n_0_2_417), .A4(
      n_0_2_418), .ZN(n_0_2_419));
   NAND2_X1 i_0_2_436 (.A1(n_0_47), .A2(\Memory[13] [16]), .ZN(n_0_2_420));
   NAND2_X1 i_0_2_437 (.A1(n_0_46), .A2(\Memory[12] [16]), .ZN(n_0_2_421));
   NAND2_X1 i_0_2_438 (.A1(n_0_45), .A2(\Memory[11] [16]), .ZN(n_0_2_422));
   NAND3_X1 i_0_2_439 (.A1(n_0_2_420), .A2(n_0_2_421), .A3(n_0_2_422), .ZN(
      n_0_2_423));
   NOR2_X1 i_0_2_440 (.A1(n_0_2_419), .A2(n_0_2_423), .ZN(n_0_2_424));
   NAND3_X1 i_0_2_441 (.A1(n_0_2_405), .A2(n_0_2_414), .A3(n_0_2_424), .ZN(
      dataOut1[16]));
   NAND2_X1 i_0_2_442 (.A1(n_0_38), .A2(\Memory[4] [17]), .ZN(n_0_2_425));
   NAND2_X1 i_0_2_443 (.A1(n_0_41), .A2(\Memory[7] [17]), .ZN(n_0_2_426));
   NAND2_X1 i_0_2_444 (.A1(n_0_37), .A2(\Memory[3] [17]), .ZN(n_0_2_427));
   NAND2_X1 i_0_2_445 (.A1(n_0_36), .A2(\Memory[2] [17]), .ZN(n_0_2_428));
   NAND4_X1 i_0_2_446 (.A1(n_0_2_425), .A2(n_0_2_426), .A3(n_0_2_427), .A4(
      n_0_2_428), .ZN(n_0_2_429));
   INV_X1 i_0_2_447 (.A(n_0_2_429), .ZN(n_0_2_430));
   NAND2_X1 i_0_2_448 (.A1(n_0_50), .A2(\Memory[16] [17]), .ZN(n_0_2_431));
   NAND2_X1 i_0_2_449 (.A1(n_0_40), .A2(\Memory[6] [17]), .ZN(n_0_2_432));
   NAND2_X1 i_0_2_450 (.A1(n_0_39), .A2(\Memory[5] [17]), .ZN(n_0_2_433));
   NAND3_X1 i_0_2_451 (.A1(n_0_2_431), .A2(n_0_2_432), .A3(n_0_2_433), .ZN(
      n_0_2_434));
   NAND2_X1 i_0_2_452 (.A1(n_0_42), .A2(\Memory[8] [17]), .ZN(n_0_2_435));
   NAND2_X1 i_0_2_453 (.A1(n_0_35), .A2(\Memory[1] [17]), .ZN(n_0_2_436));
   NAND2_X1 i_0_2_454 (.A1(n_0_44), .A2(\Memory[10] [17]), .ZN(n_0_2_437));
   NAND3_X1 i_0_2_455 (.A1(n_0_2_435), .A2(n_0_2_436), .A3(n_0_2_437), .ZN(
      n_0_2_438));
   NOR2_X1 i_0_2_456 (.A1(n_0_2_434), .A2(n_0_2_438), .ZN(n_0_2_439));
   NAND2_X1 i_0_2_457 (.A1(n_0_48), .A2(\Memory[14] [17]), .ZN(n_0_2_440));
   NAND2_X1 i_0_2_458 (.A1(n_0_49), .A2(\Memory[15] [17]), .ZN(n_0_2_441));
   NAND2_X1 i_0_2_459 (.A1(n_0_34), .A2(\Memory[0] [17]), .ZN(n_0_2_442));
   NAND2_X1 i_0_2_460 (.A1(n_0_43), .A2(\Memory[9] [17]), .ZN(n_0_2_443));
   NAND4_X1 i_0_2_461 (.A1(n_0_2_440), .A2(n_0_2_441), .A3(n_0_2_442), .A4(
      n_0_2_443), .ZN(n_0_2_444));
   NAND2_X1 i_0_2_462 (.A1(n_0_47), .A2(\Memory[13] [17]), .ZN(n_0_2_445));
   NAND2_X1 i_0_2_463 (.A1(n_0_46), .A2(\Memory[12] [17]), .ZN(n_0_2_446));
   NAND2_X1 i_0_2_464 (.A1(n_0_45), .A2(\Memory[11] [17]), .ZN(n_0_2_447));
   NAND3_X1 i_0_2_465 (.A1(n_0_2_445), .A2(n_0_2_446), .A3(n_0_2_447), .ZN(
      n_0_2_448));
   NOR2_X1 i_0_2_466 (.A1(n_0_2_444), .A2(n_0_2_448), .ZN(n_0_2_449));
   NAND3_X1 i_0_2_467 (.A1(n_0_2_430), .A2(n_0_2_439), .A3(n_0_2_449), .ZN(
      dataOut1[17]));
   NAND2_X1 i_0_2_468 (.A1(n_0_38), .A2(\Memory[4] [18]), .ZN(n_0_2_450));
   NAND2_X1 i_0_2_469 (.A1(n_0_41), .A2(\Memory[7] [18]), .ZN(n_0_2_451));
   NAND2_X1 i_0_2_470 (.A1(n_0_37), .A2(\Memory[3] [18]), .ZN(n_0_2_452));
   NAND2_X1 i_0_2_471 (.A1(n_0_36), .A2(\Memory[2] [18]), .ZN(n_0_2_453));
   NAND4_X1 i_0_2_472 (.A1(n_0_2_450), .A2(n_0_2_451), .A3(n_0_2_452), .A4(
      n_0_2_453), .ZN(n_0_2_454));
   INV_X1 i_0_2_473 (.A(n_0_2_454), .ZN(n_0_2_455));
   NAND2_X1 i_0_2_474 (.A1(n_0_50), .A2(\Memory[16] [18]), .ZN(n_0_2_456));
   NAND2_X1 i_0_2_475 (.A1(n_0_40), .A2(\Memory[6] [18]), .ZN(n_0_2_457));
   NAND2_X1 i_0_2_476 (.A1(n_0_39), .A2(\Memory[5] [18]), .ZN(n_0_2_458));
   NAND3_X1 i_0_2_477 (.A1(n_0_2_456), .A2(n_0_2_457), .A3(n_0_2_458), .ZN(
      n_0_2_459));
   NAND2_X1 i_0_2_478 (.A1(n_0_42), .A2(\Memory[8] [18]), .ZN(n_0_2_460));
   NAND2_X1 i_0_2_479 (.A1(n_0_35), .A2(\Memory[1] [18]), .ZN(n_0_2_461));
   NAND2_X1 i_0_2_480 (.A1(n_0_44), .A2(\Memory[10] [18]), .ZN(n_0_2_462));
   NAND3_X1 i_0_2_481 (.A1(n_0_2_460), .A2(n_0_2_461), .A3(n_0_2_462), .ZN(
      n_0_2_463));
   NOR2_X1 i_0_2_482 (.A1(n_0_2_459), .A2(n_0_2_463), .ZN(n_0_2_464));
   NAND2_X1 i_0_2_483 (.A1(n_0_48), .A2(\Memory[14] [18]), .ZN(n_0_2_465));
   NAND2_X1 i_0_2_484 (.A1(n_0_49), .A2(\Memory[15] [18]), .ZN(n_0_2_466));
   NAND2_X1 i_0_2_485 (.A1(n_0_34), .A2(\Memory[0] [18]), .ZN(n_0_2_467));
   NAND2_X1 i_0_2_486 (.A1(n_0_43), .A2(\Memory[9] [18]), .ZN(n_0_2_468));
   NAND4_X1 i_0_2_487 (.A1(n_0_2_465), .A2(n_0_2_466), .A3(n_0_2_467), .A4(
      n_0_2_468), .ZN(n_0_2_469));
   NAND2_X1 i_0_2_488 (.A1(n_0_47), .A2(\Memory[13] [18]), .ZN(n_0_2_470));
   NAND2_X1 i_0_2_489 (.A1(n_0_46), .A2(\Memory[12] [18]), .ZN(n_0_2_471));
   NAND2_X1 i_0_2_490 (.A1(n_0_45), .A2(\Memory[11] [18]), .ZN(n_0_2_472));
   NAND3_X1 i_0_2_491 (.A1(n_0_2_470), .A2(n_0_2_471), .A3(n_0_2_472), .ZN(
      n_0_2_473));
   NOR2_X1 i_0_2_492 (.A1(n_0_2_469), .A2(n_0_2_473), .ZN(n_0_2_474));
   NAND3_X1 i_0_2_493 (.A1(n_0_2_455), .A2(n_0_2_464), .A3(n_0_2_474), .ZN(
      dataOut1[18]));
   NAND2_X1 i_0_2_494 (.A1(n_0_38), .A2(\Memory[4] [19]), .ZN(n_0_2_475));
   NAND2_X1 i_0_2_495 (.A1(n_0_41), .A2(\Memory[7] [19]), .ZN(n_0_2_476));
   NAND2_X1 i_0_2_496 (.A1(n_0_37), .A2(\Memory[3] [19]), .ZN(n_0_2_477));
   NAND2_X1 i_0_2_497 (.A1(n_0_36), .A2(\Memory[2] [19]), .ZN(n_0_2_478));
   NAND4_X1 i_0_2_498 (.A1(n_0_2_475), .A2(n_0_2_476), .A3(n_0_2_477), .A4(
      n_0_2_478), .ZN(n_0_2_479));
   INV_X1 i_0_2_499 (.A(n_0_2_479), .ZN(n_0_2_480));
   NAND2_X1 i_0_2_500 (.A1(n_0_50), .A2(\Memory[16] [19]), .ZN(n_0_2_481));
   NAND2_X1 i_0_2_501 (.A1(n_0_40), .A2(\Memory[6] [19]), .ZN(n_0_2_482));
   NAND2_X1 i_0_2_502 (.A1(n_0_39), .A2(\Memory[5] [19]), .ZN(n_0_2_483));
   NAND3_X1 i_0_2_503 (.A1(n_0_2_481), .A2(n_0_2_482), .A3(n_0_2_483), .ZN(
      n_0_2_484));
   NAND2_X1 i_0_2_504 (.A1(n_0_42), .A2(\Memory[8] [19]), .ZN(n_0_2_485));
   NAND2_X1 i_0_2_505 (.A1(n_0_35), .A2(\Memory[1] [19]), .ZN(n_0_2_486));
   NAND2_X1 i_0_2_506 (.A1(n_0_44), .A2(\Memory[10] [19]), .ZN(n_0_2_487));
   NAND3_X1 i_0_2_507 (.A1(n_0_2_485), .A2(n_0_2_486), .A3(n_0_2_487), .ZN(
      n_0_2_488));
   NOR2_X1 i_0_2_508 (.A1(n_0_2_484), .A2(n_0_2_488), .ZN(n_0_2_489));
   NAND2_X1 i_0_2_509 (.A1(n_0_48), .A2(\Memory[14] [19]), .ZN(n_0_2_490));
   NAND2_X1 i_0_2_510 (.A1(n_0_49), .A2(\Memory[15] [19]), .ZN(n_0_2_491));
   NAND2_X1 i_0_2_511 (.A1(n_0_34), .A2(\Memory[0] [19]), .ZN(n_0_2_492));
   NAND2_X1 i_0_2_512 (.A1(n_0_43), .A2(\Memory[9] [19]), .ZN(n_0_2_493));
   NAND4_X1 i_0_2_513 (.A1(n_0_2_490), .A2(n_0_2_491), .A3(n_0_2_492), .A4(
      n_0_2_493), .ZN(n_0_2_494));
   NAND2_X1 i_0_2_514 (.A1(n_0_47), .A2(\Memory[13] [19]), .ZN(n_0_2_495));
   NAND2_X1 i_0_2_515 (.A1(n_0_46), .A2(\Memory[12] [19]), .ZN(n_0_2_496));
   NAND2_X1 i_0_2_516 (.A1(n_0_45), .A2(\Memory[11] [19]), .ZN(n_0_2_497));
   NAND3_X1 i_0_2_517 (.A1(n_0_2_495), .A2(n_0_2_496), .A3(n_0_2_497), .ZN(
      n_0_2_498));
   NOR2_X1 i_0_2_518 (.A1(n_0_2_494), .A2(n_0_2_498), .ZN(n_0_2_499));
   NAND3_X1 i_0_2_519 (.A1(n_0_2_480), .A2(n_0_2_489), .A3(n_0_2_499), .ZN(
      dataOut1[19]));
   NAND2_X1 i_0_2_520 (.A1(n_0_38), .A2(\Memory[4] [20]), .ZN(n_0_2_500));
   NAND2_X1 i_0_2_521 (.A1(n_0_41), .A2(\Memory[7] [20]), .ZN(n_0_2_501));
   NAND2_X1 i_0_2_522 (.A1(n_0_37), .A2(\Memory[3] [20]), .ZN(n_0_2_502));
   NAND2_X1 i_0_2_523 (.A1(n_0_36), .A2(\Memory[2] [20]), .ZN(n_0_2_503));
   NAND4_X1 i_0_2_524 (.A1(n_0_2_500), .A2(n_0_2_501), .A3(n_0_2_502), .A4(
      n_0_2_503), .ZN(n_0_2_504));
   INV_X1 i_0_2_525 (.A(n_0_2_504), .ZN(n_0_2_505));
   NAND2_X1 i_0_2_526 (.A1(n_0_50), .A2(\Memory[16] [20]), .ZN(n_0_2_506));
   NAND2_X1 i_0_2_527 (.A1(n_0_40), .A2(\Memory[6] [20]), .ZN(n_0_2_507));
   NAND2_X1 i_0_2_528 (.A1(n_0_39), .A2(\Memory[5] [20]), .ZN(n_0_2_508));
   NAND3_X1 i_0_2_529 (.A1(n_0_2_506), .A2(n_0_2_507), .A3(n_0_2_508), .ZN(
      n_0_2_509));
   NAND2_X1 i_0_2_530 (.A1(n_0_42), .A2(\Memory[8] [20]), .ZN(n_0_2_510));
   NAND2_X1 i_0_2_531 (.A1(n_0_35), .A2(\Memory[1] [20]), .ZN(n_0_2_511));
   NAND2_X1 i_0_2_532 (.A1(n_0_44), .A2(\Memory[10] [20]), .ZN(n_0_2_512));
   NAND3_X1 i_0_2_533 (.A1(n_0_2_510), .A2(n_0_2_511), .A3(n_0_2_512), .ZN(
      n_0_2_513));
   NOR2_X1 i_0_2_534 (.A1(n_0_2_509), .A2(n_0_2_513), .ZN(n_0_2_514));
   NAND2_X1 i_0_2_535 (.A1(n_0_48), .A2(\Memory[14] [20]), .ZN(n_0_2_515));
   NAND2_X1 i_0_2_536 (.A1(n_0_49), .A2(\Memory[15] [20]), .ZN(n_0_2_516));
   NAND2_X1 i_0_2_537 (.A1(n_0_34), .A2(\Memory[0] [20]), .ZN(n_0_2_517));
   NAND2_X1 i_0_2_538 (.A1(n_0_43), .A2(\Memory[9] [20]), .ZN(n_0_2_518));
   NAND4_X1 i_0_2_539 (.A1(n_0_2_515), .A2(n_0_2_516), .A3(n_0_2_517), .A4(
      n_0_2_518), .ZN(n_0_2_519));
   NAND2_X1 i_0_2_540 (.A1(n_0_47), .A2(\Memory[13] [20]), .ZN(n_0_2_520));
   NAND2_X1 i_0_2_541 (.A1(n_0_46), .A2(\Memory[12] [20]), .ZN(n_0_2_521));
   NAND2_X1 i_0_2_542 (.A1(n_0_45), .A2(\Memory[11] [20]), .ZN(n_0_2_522));
   NAND3_X1 i_0_2_543 (.A1(n_0_2_520), .A2(n_0_2_521), .A3(n_0_2_522), .ZN(
      n_0_2_523));
   NOR2_X1 i_0_2_544 (.A1(n_0_2_519), .A2(n_0_2_523), .ZN(n_0_2_524));
   NAND3_X1 i_0_2_545 (.A1(n_0_2_505), .A2(n_0_2_514), .A3(n_0_2_524), .ZN(
      dataOut1[20]));
   NAND2_X1 i_0_2_546 (.A1(n_0_38), .A2(\Memory[4] [21]), .ZN(n_0_2_525));
   NAND2_X1 i_0_2_547 (.A1(n_0_41), .A2(\Memory[7] [21]), .ZN(n_0_2_526));
   NAND2_X1 i_0_2_548 (.A1(n_0_37), .A2(\Memory[3] [21]), .ZN(n_0_2_527));
   NAND2_X1 i_0_2_549 (.A1(n_0_36), .A2(\Memory[2] [21]), .ZN(n_0_2_528));
   NAND4_X1 i_0_2_550 (.A1(n_0_2_525), .A2(n_0_2_526), .A3(n_0_2_527), .A4(
      n_0_2_528), .ZN(n_0_2_529));
   INV_X1 i_0_2_551 (.A(n_0_2_529), .ZN(n_0_2_530));
   NAND2_X1 i_0_2_552 (.A1(n_0_50), .A2(\Memory[16] [21]), .ZN(n_0_2_531));
   NAND2_X1 i_0_2_553 (.A1(n_0_40), .A2(\Memory[6] [21]), .ZN(n_0_2_532));
   NAND2_X1 i_0_2_554 (.A1(n_0_39), .A2(\Memory[5] [21]), .ZN(n_0_2_533));
   NAND3_X1 i_0_2_555 (.A1(n_0_2_531), .A2(n_0_2_532), .A3(n_0_2_533), .ZN(
      n_0_2_534));
   NAND2_X1 i_0_2_556 (.A1(n_0_42), .A2(\Memory[8] [21]), .ZN(n_0_2_535));
   NAND2_X1 i_0_2_557 (.A1(n_0_35), .A2(\Memory[1] [21]), .ZN(n_0_2_536));
   NAND2_X1 i_0_2_558 (.A1(n_0_44), .A2(\Memory[10] [21]), .ZN(n_0_2_537));
   NAND3_X1 i_0_2_559 (.A1(n_0_2_535), .A2(n_0_2_536), .A3(n_0_2_537), .ZN(
      n_0_2_538));
   NOR2_X1 i_0_2_560 (.A1(n_0_2_534), .A2(n_0_2_538), .ZN(n_0_2_539));
   NAND2_X1 i_0_2_561 (.A1(n_0_48), .A2(\Memory[14] [21]), .ZN(n_0_2_540));
   NAND2_X1 i_0_2_562 (.A1(n_0_49), .A2(\Memory[15] [21]), .ZN(n_0_2_541));
   NAND2_X1 i_0_2_563 (.A1(n_0_34), .A2(\Memory[0] [21]), .ZN(n_0_2_542));
   NAND2_X1 i_0_2_564 (.A1(n_0_43), .A2(\Memory[9] [21]), .ZN(n_0_2_543));
   NAND4_X1 i_0_2_565 (.A1(n_0_2_540), .A2(n_0_2_541), .A3(n_0_2_542), .A4(
      n_0_2_543), .ZN(n_0_2_544));
   NAND2_X1 i_0_2_566 (.A1(n_0_47), .A2(\Memory[13] [21]), .ZN(n_0_2_545));
   NAND2_X1 i_0_2_567 (.A1(n_0_46), .A2(\Memory[12] [21]), .ZN(n_0_2_546));
   NAND2_X1 i_0_2_568 (.A1(n_0_45), .A2(\Memory[11] [21]), .ZN(n_0_2_547));
   NAND3_X1 i_0_2_569 (.A1(n_0_2_545), .A2(n_0_2_546), .A3(n_0_2_547), .ZN(
      n_0_2_548));
   NOR2_X1 i_0_2_570 (.A1(n_0_2_544), .A2(n_0_2_548), .ZN(n_0_2_549));
   NAND3_X1 i_0_2_571 (.A1(n_0_2_530), .A2(n_0_2_539), .A3(n_0_2_549), .ZN(
      dataOut1[21]));
   NAND2_X1 i_0_2_572 (.A1(n_0_38), .A2(\Memory[4] [22]), .ZN(n_0_2_550));
   NAND2_X1 i_0_2_573 (.A1(n_0_41), .A2(\Memory[7] [22]), .ZN(n_0_2_551));
   NAND2_X1 i_0_2_574 (.A1(n_0_37), .A2(\Memory[3] [22]), .ZN(n_0_2_552));
   NAND2_X1 i_0_2_575 (.A1(n_0_36), .A2(\Memory[2] [22]), .ZN(n_0_2_553));
   NAND4_X1 i_0_2_576 (.A1(n_0_2_550), .A2(n_0_2_551), .A3(n_0_2_552), .A4(
      n_0_2_553), .ZN(n_0_2_554));
   INV_X1 i_0_2_577 (.A(n_0_2_554), .ZN(n_0_2_555));
   NAND2_X1 i_0_2_578 (.A1(n_0_50), .A2(\Memory[16] [22]), .ZN(n_0_2_556));
   NAND2_X1 i_0_2_579 (.A1(n_0_40), .A2(\Memory[6] [22]), .ZN(n_0_2_557));
   NAND2_X1 i_0_2_580 (.A1(n_0_39), .A2(\Memory[5] [22]), .ZN(n_0_2_558));
   NAND3_X1 i_0_2_581 (.A1(n_0_2_556), .A2(n_0_2_557), .A3(n_0_2_558), .ZN(
      n_0_2_559));
   NAND2_X1 i_0_2_582 (.A1(n_0_42), .A2(\Memory[8] [22]), .ZN(n_0_2_560));
   NAND2_X1 i_0_2_583 (.A1(n_0_35), .A2(\Memory[1] [22]), .ZN(n_0_2_561));
   NAND2_X1 i_0_2_584 (.A1(n_0_44), .A2(\Memory[10] [22]), .ZN(n_0_2_562));
   NAND3_X1 i_0_2_585 (.A1(n_0_2_560), .A2(n_0_2_561), .A3(n_0_2_562), .ZN(
      n_0_2_563));
   NOR2_X1 i_0_2_586 (.A1(n_0_2_559), .A2(n_0_2_563), .ZN(n_0_2_564));
   NAND2_X1 i_0_2_587 (.A1(n_0_48), .A2(\Memory[14] [22]), .ZN(n_0_2_565));
   NAND2_X1 i_0_2_588 (.A1(n_0_49), .A2(\Memory[15] [22]), .ZN(n_0_2_566));
   NAND2_X1 i_0_2_589 (.A1(n_0_34), .A2(\Memory[0] [22]), .ZN(n_0_2_567));
   NAND2_X1 i_0_2_590 (.A1(n_0_43), .A2(\Memory[9] [22]), .ZN(n_0_2_568));
   NAND4_X1 i_0_2_591 (.A1(n_0_2_565), .A2(n_0_2_566), .A3(n_0_2_567), .A4(
      n_0_2_568), .ZN(n_0_2_569));
   NAND2_X1 i_0_2_592 (.A1(n_0_47), .A2(\Memory[13] [22]), .ZN(n_0_2_570));
   NAND2_X1 i_0_2_593 (.A1(n_0_46), .A2(\Memory[12] [22]), .ZN(n_0_2_571));
   NAND2_X1 i_0_2_594 (.A1(n_0_45), .A2(\Memory[11] [22]), .ZN(n_0_2_572));
   NAND3_X1 i_0_2_595 (.A1(n_0_2_570), .A2(n_0_2_571), .A3(n_0_2_572), .ZN(
      n_0_2_573));
   NOR2_X1 i_0_2_596 (.A1(n_0_2_569), .A2(n_0_2_573), .ZN(n_0_2_574));
   NAND3_X1 i_0_2_597 (.A1(n_0_2_555), .A2(n_0_2_564), .A3(n_0_2_574), .ZN(
      dataOut1[22]));
   NAND2_X1 i_0_2_598 (.A1(n_0_38), .A2(\Memory[4] [23]), .ZN(n_0_2_575));
   NAND2_X1 i_0_2_599 (.A1(n_0_41), .A2(\Memory[7] [23]), .ZN(n_0_2_576));
   NAND2_X1 i_0_2_600 (.A1(n_0_37), .A2(\Memory[3] [23]), .ZN(n_0_2_577));
   NAND2_X1 i_0_2_601 (.A1(n_0_36), .A2(\Memory[2] [23]), .ZN(n_0_2_578));
   NAND4_X1 i_0_2_602 (.A1(n_0_2_575), .A2(n_0_2_576), .A3(n_0_2_577), .A4(
      n_0_2_578), .ZN(n_0_2_579));
   INV_X1 i_0_2_603 (.A(n_0_2_579), .ZN(n_0_2_580));
   NAND2_X1 i_0_2_604 (.A1(n_0_50), .A2(\Memory[16] [23]), .ZN(n_0_2_581));
   NAND2_X1 i_0_2_605 (.A1(n_0_40), .A2(\Memory[6] [23]), .ZN(n_0_2_582));
   NAND2_X1 i_0_2_606 (.A1(n_0_39), .A2(\Memory[5] [23]), .ZN(n_0_2_583));
   NAND3_X1 i_0_2_607 (.A1(n_0_2_581), .A2(n_0_2_582), .A3(n_0_2_583), .ZN(
      n_0_2_584));
   NAND2_X1 i_0_2_608 (.A1(n_0_42), .A2(\Memory[8] [23]), .ZN(n_0_2_585));
   NAND2_X1 i_0_2_609 (.A1(n_0_35), .A2(\Memory[1] [23]), .ZN(n_0_2_586));
   NAND2_X1 i_0_2_610 (.A1(n_0_44), .A2(\Memory[10] [23]), .ZN(n_0_2_587));
   NAND3_X1 i_0_2_611 (.A1(n_0_2_585), .A2(n_0_2_586), .A3(n_0_2_587), .ZN(
      n_0_2_588));
   NOR2_X1 i_0_2_612 (.A1(n_0_2_584), .A2(n_0_2_588), .ZN(n_0_2_589));
   NAND2_X1 i_0_2_613 (.A1(n_0_48), .A2(\Memory[14] [23]), .ZN(n_0_2_590));
   NAND2_X1 i_0_2_614 (.A1(n_0_49), .A2(\Memory[15] [23]), .ZN(n_0_2_591));
   NAND2_X1 i_0_2_615 (.A1(n_0_34), .A2(\Memory[0] [23]), .ZN(n_0_2_592));
   NAND2_X1 i_0_2_616 (.A1(n_0_43), .A2(\Memory[9] [23]), .ZN(n_0_2_593));
   NAND4_X1 i_0_2_617 (.A1(n_0_2_590), .A2(n_0_2_591), .A3(n_0_2_592), .A4(
      n_0_2_593), .ZN(n_0_2_594));
   NAND2_X1 i_0_2_618 (.A1(n_0_47), .A2(\Memory[13] [23]), .ZN(n_0_2_595));
   NAND2_X1 i_0_2_619 (.A1(n_0_46), .A2(\Memory[12] [23]), .ZN(n_0_2_596));
   NAND2_X1 i_0_2_620 (.A1(n_0_45), .A2(\Memory[11] [23]), .ZN(n_0_2_597));
   NAND3_X1 i_0_2_621 (.A1(n_0_2_595), .A2(n_0_2_596), .A3(n_0_2_597), .ZN(
      n_0_2_598));
   NOR2_X1 i_0_2_622 (.A1(n_0_2_594), .A2(n_0_2_598), .ZN(n_0_2_599));
   NAND3_X1 i_0_2_623 (.A1(n_0_2_580), .A2(n_0_2_589), .A3(n_0_2_599), .ZN(
      dataOut1[23]));
   NAND2_X1 i_0_2_624 (.A1(n_0_38), .A2(\Memory[4] [24]), .ZN(n_0_2_600));
   NAND2_X1 i_0_2_625 (.A1(n_0_41), .A2(\Memory[7] [24]), .ZN(n_0_2_601));
   NAND2_X1 i_0_2_626 (.A1(n_0_37), .A2(\Memory[3] [24]), .ZN(n_0_2_602));
   NAND2_X1 i_0_2_627 (.A1(n_0_36), .A2(\Memory[2] [24]), .ZN(n_0_2_603));
   NAND4_X1 i_0_2_628 (.A1(n_0_2_600), .A2(n_0_2_601), .A3(n_0_2_602), .A4(
      n_0_2_603), .ZN(n_0_2_604));
   INV_X1 i_0_2_629 (.A(n_0_2_604), .ZN(n_0_2_605));
   NAND2_X1 i_0_2_630 (.A1(n_0_50), .A2(\Memory[16] [24]), .ZN(n_0_2_606));
   NAND2_X1 i_0_2_631 (.A1(n_0_40), .A2(\Memory[6] [24]), .ZN(n_0_2_607));
   NAND2_X1 i_0_2_632 (.A1(n_0_39), .A2(\Memory[5] [24]), .ZN(n_0_2_608));
   NAND3_X1 i_0_2_633 (.A1(n_0_2_606), .A2(n_0_2_607), .A3(n_0_2_608), .ZN(
      n_0_2_609));
   NAND2_X1 i_0_2_634 (.A1(n_0_42), .A2(\Memory[8] [24]), .ZN(n_0_2_610));
   NAND2_X1 i_0_2_635 (.A1(n_0_35), .A2(\Memory[1] [24]), .ZN(n_0_2_611));
   NAND2_X1 i_0_2_636 (.A1(n_0_44), .A2(\Memory[10] [24]), .ZN(n_0_2_612));
   NAND3_X1 i_0_2_637 (.A1(n_0_2_610), .A2(n_0_2_611), .A3(n_0_2_612), .ZN(
      n_0_2_613));
   NOR2_X1 i_0_2_638 (.A1(n_0_2_609), .A2(n_0_2_613), .ZN(n_0_2_614));
   NAND2_X1 i_0_2_639 (.A1(n_0_48), .A2(\Memory[14] [24]), .ZN(n_0_2_615));
   NAND2_X1 i_0_2_640 (.A1(n_0_49), .A2(\Memory[15] [24]), .ZN(n_0_2_616));
   NAND2_X1 i_0_2_641 (.A1(n_0_34), .A2(\Memory[0] [24]), .ZN(n_0_2_617));
   NAND2_X1 i_0_2_642 (.A1(n_0_43), .A2(\Memory[9] [24]), .ZN(n_0_2_618));
   NAND4_X1 i_0_2_643 (.A1(n_0_2_615), .A2(n_0_2_616), .A3(n_0_2_617), .A4(
      n_0_2_618), .ZN(n_0_2_619));
   NAND2_X1 i_0_2_644 (.A1(n_0_47), .A2(\Memory[13] [24]), .ZN(n_0_2_620));
   NAND2_X1 i_0_2_645 (.A1(n_0_46), .A2(\Memory[12] [24]), .ZN(n_0_2_621));
   NAND2_X1 i_0_2_646 (.A1(n_0_45), .A2(\Memory[11] [24]), .ZN(n_0_2_622));
   NAND3_X1 i_0_2_647 (.A1(n_0_2_620), .A2(n_0_2_621), .A3(n_0_2_622), .ZN(
      n_0_2_623));
   NOR2_X1 i_0_2_648 (.A1(n_0_2_619), .A2(n_0_2_623), .ZN(n_0_2_624));
   NAND3_X1 i_0_2_649 (.A1(n_0_2_605), .A2(n_0_2_614), .A3(n_0_2_624), .ZN(
      dataOut1[24]));
   NAND2_X1 i_0_2_650 (.A1(n_0_38), .A2(\Memory[4] [25]), .ZN(n_0_2_625));
   NAND2_X1 i_0_2_651 (.A1(n_0_41), .A2(\Memory[7] [25]), .ZN(n_0_2_626));
   NAND2_X1 i_0_2_652 (.A1(n_0_37), .A2(\Memory[3] [25]), .ZN(n_0_2_627));
   NAND2_X1 i_0_2_653 (.A1(n_0_36), .A2(\Memory[2] [25]), .ZN(n_0_2_628));
   NAND4_X1 i_0_2_654 (.A1(n_0_2_625), .A2(n_0_2_626), .A3(n_0_2_627), .A4(
      n_0_2_628), .ZN(n_0_2_629));
   INV_X1 i_0_2_655 (.A(n_0_2_629), .ZN(n_0_2_630));
   NAND2_X1 i_0_2_656 (.A1(n_0_50), .A2(\Memory[16] [25]), .ZN(n_0_2_631));
   NAND2_X1 i_0_2_657 (.A1(n_0_40), .A2(\Memory[6] [25]), .ZN(n_0_2_632));
   NAND2_X1 i_0_2_658 (.A1(n_0_39), .A2(\Memory[5] [25]), .ZN(n_0_2_633));
   NAND3_X1 i_0_2_659 (.A1(n_0_2_631), .A2(n_0_2_632), .A3(n_0_2_633), .ZN(
      n_0_2_634));
   NAND2_X1 i_0_2_660 (.A1(n_0_42), .A2(\Memory[8] [25]), .ZN(n_0_2_635));
   NAND2_X1 i_0_2_661 (.A1(n_0_35), .A2(\Memory[1] [25]), .ZN(n_0_2_636));
   NAND2_X1 i_0_2_662 (.A1(n_0_44), .A2(\Memory[10] [25]), .ZN(n_0_2_637));
   NAND3_X1 i_0_2_663 (.A1(n_0_2_635), .A2(n_0_2_636), .A3(n_0_2_637), .ZN(
      n_0_2_638));
   NOR2_X1 i_0_2_664 (.A1(n_0_2_634), .A2(n_0_2_638), .ZN(n_0_2_639));
   NAND2_X1 i_0_2_665 (.A1(n_0_48), .A2(\Memory[14] [25]), .ZN(n_0_2_640));
   NAND2_X1 i_0_2_666 (.A1(n_0_49), .A2(\Memory[15] [25]), .ZN(n_0_2_641));
   NAND2_X1 i_0_2_667 (.A1(n_0_34), .A2(\Memory[0] [25]), .ZN(n_0_2_642));
   NAND2_X1 i_0_2_668 (.A1(n_0_43), .A2(\Memory[9] [25]), .ZN(n_0_2_643));
   NAND4_X1 i_0_2_669 (.A1(n_0_2_640), .A2(n_0_2_641), .A3(n_0_2_642), .A4(
      n_0_2_643), .ZN(n_0_2_644));
   NAND2_X1 i_0_2_670 (.A1(n_0_47), .A2(\Memory[13] [25]), .ZN(n_0_2_645));
   NAND2_X1 i_0_2_671 (.A1(n_0_46), .A2(\Memory[12] [25]), .ZN(n_0_2_646));
   NAND2_X1 i_0_2_672 (.A1(n_0_45), .A2(\Memory[11] [25]), .ZN(n_0_2_647));
   NAND3_X1 i_0_2_673 (.A1(n_0_2_645), .A2(n_0_2_646), .A3(n_0_2_647), .ZN(
      n_0_2_648));
   NOR2_X1 i_0_2_674 (.A1(n_0_2_644), .A2(n_0_2_648), .ZN(n_0_2_649));
   NAND3_X1 i_0_2_675 (.A1(n_0_2_630), .A2(n_0_2_639), .A3(n_0_2_649), .ZN(
      dataOut1[25]));
   NAND2_X1 i_0_2_676 (.A1(n_0_38), .A2(\Memory[4] [26]), .ZN(n_0_2_650));
   NAND2_X1 i_0_2_677 (.A1(n_0_41), .A2(\Memory[7] [26]), .ZN(n_0_2_651));
   NAND2_X1 i_0_2_678 (.A1(n_0_37), .A2(\Memory[3] [26]), .ZN(n_0_2_652));
   NAND2_X1 i_0_2_679 (.A1(n_0_36), .A2(\Memory[2] [26]), .ZN(n_0_2_653));
   NAND4_X1 i_0_2_680 (.A1(n_0_2_650), .A2(n_0_2_651), .A3(n_0_2_652), .A4(
      n_0_2_653), .ZN(n_0_2_654));
   INV_X1 i_0_2_681 (.A(n_0_2_654), .ZN(n_0_2_655));
   NAND2_X1 i_0_2_682 (.A1(n_0_50), .A2(\Memory[16] [26]), .ZN(n_0_2_656));
   NAND2_X1 i_0_2_683 (.A1(n_0_40), .A2(\Memory[6] [26]), .ZN(n_0_2_657));
   NAND2_X1 i_0_2_684 (.A1(n_0_39), .A2(\Memory[5] [26]), .ZN(n_0_2_658));
   NAND3_X1 i_0_2_685 (.A1(n_0_2_656), .A2(n_0_2_657), .A3(n_0_2_658), .ZN(
      n_0_2_659));
   NAND2_X1 i_0_2_686 (.A1(n_0_42), .A2(\Memory[8] [26]), .ZN(n_0_2_660));
   NAND2_X1 i_0_2_687 (.A1(n_0_35), .A2(\Memory[1] [26]), .ZN(n_0_2_661));
   NAND2_X1 i_0_2_688 (.A1(n_0_44), .A2(\Memory[10] [26]), .ZN(n_0_2_662));
   NAND3_X1 i_0_2_689 (.A1(n_0_2_660), .A2(n_0_2_661), .A3(n_0_2_662), .ZN(
      n_0_2_663));
   NOR2_X1 i_0_2_690 (.A1(n_0_2_659), .A2(n_0_2_663), .ZN(n_0_2_664));
   NAND2_X1 i_0_2_691 (.A1(n_0_48), .A2(\Memory[14] [26]), .ZN(n_0_2_665));
   NAND2_X1 i_0_2_692 (.A1(n_0_49), .A2(\Memory[15] [26]), .ZN(n_0_2_666));
   NAND2_X1 i_0_2_693 (.A1(n_0_34), .A2(\Memory[0] [26]), .ZN(n_0_2_667));
   NAND2_X1 i_0_2_694 (.A1(n_0_43), .A2(\Memory[9] [26]), .ZN(n_0_2_668));
   NAND4_X1 i_0_2_695 (.A1(n_0_2_665), .A2(n_0_2_666), .A3(n_0_2_667), .A4(
      n_0_2_668), .ZN(n_0_2_669));
   NAND2_X1 i_0_2_696 (.A1(n_0_47), .A2(\Memory[13] [26]), .ZN(n_0_2_670));
   NAND2_X1 i_0_2_697 (.A1(n_0_46), .A2(\Memory[12] [26]), .ZN(n_0_2_671));
   NAND2_X1 i_0_2_698 (.A1(n_0_45), .A2(\Memory[11] [26]), .ZN(n_0_2_672));
   NAND3_X1 i_0_2_699 (.A1(n_0_2_670), .A2(n_0_2_671), .A3(n_0_2_672), .ZN(
      n_0_2_673));
   NOR2_X1 i_0_2_700 (.A1(n_0_2_669), .A2(n_0_2_673), .ZN(n_0_2_674));
   NAND3_X1 i_0_2_701 (.A1(n_0_2_655), .A2(n_0_2_664), .A3(n_0_2_674), .ZN(
      dataOut1[26]));
   NAND2_X1 i_0_2_702 (.A1(n_0_38), .A2(\Memory[4] [27]), .ZN(n_0_2_675));
   NAND2_X1 i_0_2_703 (.A1(n_0_41), .A2(\Memory[7] [27]), .ZN(n_0_2_676));
   NAND2_X1 i_0_2_704 (.A1(n_0_37), .A2(\Memory[3] [27]), .ZN(n_0_2_677));
   NAND2_X1 i_0_2_705 (.A1(n_0_36), .A2(\Memory[2] [27]), .ZN(n_0_2_678));
   NAND4_X1 i_0_2_706 (.A1(n_0_2_675), .A2(n_0_2_676), .A3(n_0_2_677), .A4(
      n_0_2_678), .ZN(n_0_2_679));
   INV_X1 i_0_2_707 (.A(n_0_2_679), .ZN(n_0_2_680));
   NAND2_X1 i_0_2_708 (.A1(n_0_50), .A2(\Memory[16] [27]), .ZN(n_0_2_681));
   NAND2_X1 i_0_2_709 (.A1(n_0_40), .A2(\Memory[6] [27]), .ZN(n_0_2_682));
   NAND2_X1 i_0_2_710 (.A1(n_0_39), .A2(\Memory[5] [27]), .ZN(n_0_2_683));
   NAND3_X1 i_0_2_711 (.A1(n_0_2_681), .A2(n_0_2_682), .A3(n_0_2_683), .ZN(
      n_0_2_684));
   NAND2_X1 i_0_2_712 (.A1(n_0_42), .A2(\Memory[8] [27]), .ZN(n_0_2_685));
   NAND2_X1 i_0_2_713 (.A1(n_0_35), .A2(\Memory[1] [27]), .ZN(n_0_2_686));
   NAND2_X1 i_0_2_714 (.A1(n_0_44), .A2(\Memory[10] [27]), .ZN(n_0_2_687));
   NAND3_X1 i_0_2_715 (.A1(n_0_2_685), .A2(n_0_2_686), .A3(n_0_2_687), .ZN(
      n_0_2_688));
   NOR2_X1 i_0_2_716 (.A1(n_0_2_684), .A2(n_0_2_688), .ZN(n_0_2_689));
   NAND2_X1 i_0_2_717 (.A1(n_0_48), .A2(\Memory[14] [27]), .ZN(n_0_2_690));
   NAND2_X1 i_0_2_718 (.A1(n_0_49), .A2(\Memory[15] [27]), .ZN(n_0_2_691));
   NAND2_X1 i_0_2_719 (.A1(n_0_34), .A2(\Memory[0] [27]), .ZN(n_0_2_692));
   NAND2_X1 i_0_2_720 (.A1(n_0_43), .A2(\Memory[9] [27]), .ZN(n_0_2_693));
   NAND4_X1 i_0_2_721 (.A1(n_0_2_690), .A2(n_0_2_691), .A3(n_0_2_692), .A4(
      n_0_2_693), .ZN(n_0_2_694));
   NAND2_X1 i_0_2_722 (.A1(n_0_47), .A2(\Memory[13] [27]), .ZN(n_0_2_695));
   NAND2_X1 i_0_2_723 (.A1(n_0_46), .A2(\Memory[12] [27]), .ZN(n_0_2_696));
   NAND2_X1 i_0_2_724 (.A1(n_0_45), .A2(\Memory[11] [27]), .ZN(n_0_2_697));
   NAND3_X1 i_0_2_725 (.A1(n_0_2_695), .A2(n_0_2_696), .A3(n_0_2_697), .ZN(
      n_0_2_698));
   NOR2_X1 i_0_2_726 (.A1(n_0_2_694), .A2(n_0_2_698), .ZN(n_0_2_699));
   NAND3_X1 i_0_2_727 (.A1(n_0_2_680), .A2(n_0_2_689), .A3(n_0_2_699), .ZN(
      dataOut1[27]));
   NAND2_X1 i_0_2_728 (.A1(n_0_38), .A2(\Memory[4] [28]), .ZN(n_0_2_700));
   NAND2_X1 i_0_2_729 (.A1(n_0_41), .A2(\Memory[7] [28]), .ZN(n_0_2_701));
   NAND2_X1 i_0_2_730 (.A1(n_0_37), .A2(\Memory[3] [28]), .ZN(n_0_2_702));
   NAND2_X1 i_0_2_731 (.A1(n_0_36), .A2(\Memory[2] [28]), .ZN(n_0_2_703));
   NAND4_X1 i_0_2_732 (.A1(n_0_2_700), .A2(n_0_2_701), .A3(n_0_2_702), .A4(
      n_0_2_703), .ZN(n_0_2_704));
   INV_X1 i_0_2_733 (.A(n_0_2_704), .ZN(n_0_2_705));
   NAND2_X1 i_0_2_734 (.A1(n_0_50), .A2(\Memory[16] [28]), .ZN(n_0_2_706));
   NAND2_X1 i_0_2_735 (.A1(n_0_40), .A2(\Memory[6] [28]), .ZN(n_0_2_707));
   NAND2_X1 i_0_2_736 (.A1(n_0_39), .A2(\Memory[5] [28]), .ZN(n_0_2_708));
   NAND3_X1 i_0_2_737 (.A1(n_0_2_706), .A2(n_0_2_707), .A3(n_0_2_708), .ZN(
      n_0_2_709));
   NAND2_X1 i_0_2_738 (.A1(n_0_42), .A2(\Memory[8] [28]), .ZN(n_0_2_710));
   NAND2_X1 i_0_2_739 (.A1(n_0_35), .A2(\Memory[1] [28]), .ZN(n_0_2_711));
   NAND2_X1 i_0_2_740 (.A1(n_0_44), .A2(\Memory[10] [28]), .ZN(n_0_2_712));
   NAND3_X1 i_0_2_741 (.A1(n_0_2_710), .A2(n_0_2_711), .A3(n_0_2_712), .ZN(
      n_0_2_713));
   NOR2_X1 i_0_2_742 (.A1(n_0_2_709), .A2(n_0_2_713), .ZN(n_0_2_714));
   NAND2_X1 i_0_2_743 (.A1(n_0_48), .A2(\Memory[14] [28]), .ZN(n_0_2_715));
   NAND2_X1 i_0_2_744 (.A1(n_0_49), .A2(\Memory[15] [28]), .ZN(n_0_2_716));
   NAND2_X1 i_0_2_745 (.A1(n_0_34), .A2(\Memory[0] [28]), .ZN(n_0_2_717));
   NAND2_X1 i_0_2_746 (.A1(n_0_43), .A2(\Memory[9] [28]), .ZN(n_0_2_718));
   NAND4_X1 i_0_2_747 (.A1(n_0_2_715), .A2(n_0_2_716), .A3(n_0_2_717), .A4(
      n_0_2_718), .ZN(n_0_2_719));
   NAND2_X1 i_0_2_748 (.A1(n_0_47), .A2(\Memory[13] [28]), .ZN(n_0_2_720));
   NAND2_X1 i_0_2_749 (.A1(n_0_46), .A2(\Memory[12] [28]), .ZN(n_0_2_721));
   NAND2_X1 i_0_2_750 (.A1(n_0_45), .A2(\Memory[11] [28]), .ZN(n_0_2_722));
   NAND3_X1 i_0_2_751 (.A1(n_0_2_720), .A2(n_0_2_721), .A3(n_0_2_722), .ZN(
      n_0_2_723));
   NOR2_X1 i_0_2_752 (.A1(n_0_2_719), .A2(n_0_2_723), .ZN(n_0_2_724));
   NAND3_X1 i_0_2_753 (.A1(n_0_2_705), .A2(n_0_2_714), .A3(n_0_2_724), .ZN(
      dataOut1[28]));
   NAND2_X1 i_0_2_754 (.A1(n_0_38), .A2(\Memory[4] [29]), .ZN(n_0_2_725));
   NAND2_X1 i_0_2_755 (.A1(n_0_41), .A2(\Memory[7] [29]), .ZN(n_0_2_726));
   NAND2_X1 i_0_2_756 (.A1(n_0_37), .A2(\Memory[3] [29]), .ZN(n_0_2_727));
   NAND2_X1 i_0_2_757 (.A1(n_0_36), .A2(\Memory[2] [29]), .ZN(n_0_2_728));
   NAND4_X1 i_0_2_758 (.A1(n_0_2_725), .A2(n_0_2_726), .A3(n_0_2_727), .A4(
      n_0_2_728), .ZN(n_0_2_729));
   INV_X1 i_0_2_759 (.A(n_0_2_729), .ZN(n_0_2_730));
   NAND2_X1 i_0_2_760 (.A1(n_0_50), .A2(\Memory[16] [29]), .ZN(n_0_2_731));
   NAND2_X1 i_0_2_761 (.A1(n_0_40), .A2(\Memory[6] [29]), .ZN(n_0_2_732));
   NAND2_X1 i_0_2_762 (.A1(n_0_39), .A2(\Memory[5] [29]), .ZN(n_0_2_733));
   NAND3_X1 i_0_2_763 (.A1(n_0_2_731), .A2(n_0_2_732), .A3(n_0_2_733), .ZN(
      n_0_2_734));
   NAND2_X1 i_0_2_764 (.A1(n_0_42), .A2(\Memory[8] [29]), .ZN(n_0_2_735));
   NAND2_X1 i_0_2_765 (.A1(n_0_35), .A2(\Memory[1] [29]), .ZN(n_0_2_736));
   NAND2_X1 i_0_2_766 (.A1(n_0_44), .A2(\Memory[10] [29]), .ZN(n_0_2_737));
   NAND3_X1 i_0_2_767 (.A1(n_0_2_735), .A2(n_0_2_736), .A3(n_0_2_737), .ZN(
      n_0_2_738));
   NOR2_X1 i_0_2_768 (.A1(n_0_2_734), .A2(n_0_2_738), .ZN(n_0_2_739));
   NAND2_X1 i_0_2_769 (.A1(n_0_48), .A2(\Memory[14] [29]), .ZN(n_0_2_740));
   NAND2_X1 i_0_2_770 (.A1(n_0_49), .A2(\Memory[15] [29]), .ZN(n_0_2_741));
   NAND2_X1 i_0_2_771 (.A1(n_0_34), .A2(\Memory[0] [29]), .ZN(n_0_2_742));
   NAND2_X1 i_0_2_772 (.A1(n_0_43), .A2(\Memory[9] [29]), .ZN(n_0_2_743));
   NAND4_X1 i_0_2_773 (.A1(n_0_2_740), .A2(n_0_2_741), .A3(n_0_2_742), .A4(
      n_0_2_743), .ZN(n_0_2_744));
   NAND2_X1 i_0_2_774 (.A1(n_0_47), .A2(\Memory[13] [29]), .ZN(n_0_2_745));
   NAND2_X1 i_0_2_775 (.A1(n_0_46), .A2(\Memory[12] [29]), .ZN(n_0_2_746));
   NAND2_X1 i_0_2_776 (.A1(n_0_45), .A2(\Memory[11] [29]), .ZN(n_0_2_747));
   NAND3_X1 i_0_2_777 (.A1(n_0_2_745), .A2(n_0_2_746), .A3(n_0_2_747), .ZN(
      n_0_2_748));
   NOR2_X1 i_0_2_778 (.A1(n_0_2_744), .A2(n_0_2_748), .ZN(n_0_2_749));
   NAND3_X1 i_0_2_779 (.A1(n_0_2_730), .A2(n_0_2_739), .A3(n_0_2_749), .ZN(
      dataOut1[29]));
   NAND2_X1 i_0_2_780 (.A1(n_0_38), .A2(\Memory[4] [30]), .ZN(n_0_2_750));
   NAND2_X1 i_0_2_781 (.A1(n_0_41), .A2(\Memory[7] [30]), .ZN(n_0_2_751));
   NAND2_X1 i_0_2_782 (.A1(n_0_37), .A2(\Memory[3] [30]), .ZN(n_0_2_752));
   NAND2_X1 i_0_2_783 (.A1(n_0_36), .A2(\Memory[2] [30]), .ZN(n_0_2_753));
   NAND4_X1 i_0_2_784 (.A1(n_0_2_750), .A2(n_0_2_751), .A3(n_0_2_752), .A4(
      n_0_2_753), .ZN(n_0_2_754));
   INV_X1 i_0_2_785 (.A(n_0_2_754), .ZN(n_0_2_755));
   NAND2_X1 i_0_2_786 (.A1(n_0_50), .A2(\Memory[16] [30]), .ZN(n_0_2_756));
   NAND2_X1 i_0_2_787 (.A1(n_0_40), .A2(\Memory[6] [30]), .ZN(n_0_2_757));
   NAND2_X1 i_0_2_788 (.A1(n_0_39), .A2(\Memory[5] [30]), .ZN(n_0_2_758));
   NAND3_X1 i_0_2_789 (.A1(n_0_2_756), .A2(n_0_2_757), .A3(n_0_2_758), .ZN(
      n_0_2_759));
   NAND2_X1 i_0_2_790 (.A1(n_0_42), .A2(\Memory[8] [30]), .ZN(n_0_2_760));
   NAND2_X1 i_0_2_791 (.A1(n_0_35), .A2(\Memory[1] [30]), .ZN(n_0_2_761));
   NAND2_X1 i_0_2_792 (.A1(n_0_44), .A2(\Memory[10] [30]), .ZN(n_0_2_762));
   NAND3_X1 i_0_2_793 (.A1(n_0_2_760), .A2(n_0_2_761), .A3(n_0_2_762), .ZN(
      n_0_2_763));
   NOR2_X1 i_0_2_794 (.A1(n_0_2_759), .A2(n_0_2_763), .ZN(n_0_2_764));
   NAND2_X1 i_0_2_795 (.A1(n_0_48), .A2(\Memory[14] [30]), .ZN(n_0_2_765));
   NAND2_X1 i_0_2_796 (.A1(n_0_49), .A2(\Memory[15] [30]), .ZN(n_0_2_766));
   NAND2_X1 i_0_2_797 (.A1(n_0_34), .A2(\Memory[0] [30]), .ZN(n_0_2_767));
   NAND2_X1 i_0_2_798 (.A1(n_0_43), .A2(\Memory[9] [30]), .ZN(n_0_2_768));
   NAND4_X1 i_0_2_799 (.A1(n_0_2_765), .A2(n_0_2_766), .A3(n_0_2_767), .A4(
      n_0_2_768), .ZN(n_0_2_769));
   NAND2_X1 i_0_2_800 (.A1(n_0_47), .A2(\Memory[13] [30]), .ZN(n_0_2_770));
   NAND2_X1 i_0_2_801 (.A1(n_0_46), .A2(\Memory[12] [30]), .ZN(n_0_2_771));
   NAND2_X1 i_0_2_802 (.A1(n_0_45), .A2(\Memory[11] [30]), .ZN(n_0_2_772));
   NAND3_X1 i_0_2_803 (.A1(n_0_2_770), .A2(n_0_2_771), .A3(n_0_2_772), .ZN(
      n_0_2_773));
   NOR2_X1 i_0_2_804 (.A1(n_0_2_769), .A2(n_0_2_773), .ZN(n_0_2_774));
   NAND3_X1 i_0_2_805 (.A1(n_0_2_755), .A2(n_0_2_764), .A3(n_0_2_774), .ZN(
      dataOut1[30]));
   NAND2_X1 i_0_2_806 (.A1(n_0_38), .A2(\Memory[4] [31]), .ZN(n_0_2_775));
   NAND2_X1 i_0_2_807 (.A1(n_0_41), .A2(\Memory[7] [31]), .ZN(n_0_2_776));
   NAND2_X1 i_0_2_808 (.A1(n_0_37), .A2(\Memory[3] [31]), .ZN(n_0_2_777));
   NAND2_X1 i_0_2_809 (.A1(n_0_36), .A2(\Memory[2] [31]), .ZN(n_0_2_778));
   NAND4_X1 i_0_2_810 (.A1(n_0_2_775), .A2(n_0_2_776), .A3(n_0_2_777), .A4(
      n_0_2_778), .ZN(n_0_2_779));
   INV_X1 i_0_2_811 (.A(n_0_2_779), .ZN(n_0_2_780));
   NAND2_X1 i_0_2_812 (.A1(n_0_50), .A2(\Memory[16] [31]), .ZN(n_0_2_781));
   NAND2_X1 i_0_2_813 (.A1(n_0_40), .A2(\Memory[6] [31]), .ZN(n_0_2_782));
   NAND2_X1 i_0_2_814 (.A1(n_0_39), .A2(\Memory[5] [31]), .ZN(n_0_2_783));
   NAND3_X1 i_0_2_815 (.A1(n_0_2_781), .A2(n_0_2_782), .A3(n_0_2_783), .ZN(
      n_0_2_784));
   NAND2_X1 i_0_2_816 (.A1(n_0_42), .A2(\Memory[8] [31]), .ZN(n_0_2_785));
   NAND2_X1 i_0_2_817 (.A1(n_0_35), .A2(\Memory[1] [31]), .ZN(n_0_2_786));
   NAND2_X1 i_0_2_818 (.A1(n_0_44), .A2(\Memory[10] [31]), .ZN(n_0_2_787));
   NAND3_X1 i_0_2_819 (.A1(n_0_2_785), .A2(n_0_2_786), .A3(n_0_2_787), .ZN(
      n_0_2_788));
   NOR2_X1 i_0_2_820 (.A1(n_0_2_784), .A2(n_0_2_788), .ZN(n_0_2_789));
   NAND2_X1 i_0_2_821 (.A1(n_0_48), .A2(\Memory[14] [31]), .ZN(n_0_2_790));
   NAND2_X1 i_0_2_822 (.A1(n_0_49), .A2(\Memory[15] [31]), .ZN(n_0_2_791));
   NAND2_X1 i_0_2_823 (.A1(n_0_34), .A2(\Memory[0] [31]), .ZN(n_0_2_792));
   NAND2_X1 i_0_2_824 (.A1(n_0_43), .A2(\Memory[9] [31]), .ZN(n_0_2_793));
   NAND4_X1 i_0_2_825 (.A1(n_0_2_790), .A2(n_0_2_791), .A3(n_0_2_792), .A4(
      n_0_2_793), .ZN(n_0_2_794));
   NAND2_X1 i_0_2_826 (.A1(n_0_47), .A2(\Memory[13] [31]), .ZN(n_0_2_795));
   NAND2_X1 i_0_2_827 (.A1(n_0_46), .A2(\Memory[12] [31]), .ZN(n_0_2_796));
   NAND2_X1 i_0_2_828 (.A1(n_0_45), .A2(\Memory[11] [31]), .ZN(n_0_2_797));
   NAND3_X1 i_0_2_829 (.A1(n_0_2_795), .A2(n_0_2_796), .A3(n_0_2_797), .ZN(
      n_0_2_798));
   NOR2_X1 i_0_2_830 (.A1(n_0_2_794), .A2(n_0_2_798), .ZN(n_0_2_799));
   NAND3_X1 i_0_2_831 (.A1(n_0_2_780), .A2(n_0_2_789), .A3(n_0_2_799), .ZN(
      dataOut1[31]));
   NAND2_X1 i_0_2_832 (.A1(n_0_38), .A2(\Memory[4] [32]), .ZN(n_0_2_800));
   NAND2_X1 i_0_2_833 (.A1(n_0_41), .A2(\Memory[7] [32]), .ZN(n_0_2_801));
   NAND2_X1 i_0_2_834 (.A1(n_0_37), .A2(\Memory[3] [32]), .ZN(n_0_2_802));
   NAND2_X1 i_0_2_835 (.A1(n_0_36), .A2(\Memory[2] [32]), .ZN(n_0_2_803));
   NAND4_X1 i_0_2_836 (.A1(n_0_2_800), .A2(n_0_2_801), .A3(n_0_2_802), .A4(
      n_0_2_803), .ZN(n_0_2_804));
   INV_X1 i_0_2_837 (.A(n_0_2_804), .ZN(n_0_2_805));
   NAND2_X1 i_0_2_838 (.A1(n_0_50), .A2(\Memory[16] [32]), .ZN(n_0_2_806));
   NAND2_X1 i_0_2_839 (.A1(n_0_40), .A2(\Memory[6] [32]), .ZN(n_0_2_807));
   NAND2_X1 i_0_2_840 (.A1(n_0_39), .A2(\Memory[5] [32]), .ZN(n_0_2_808));
   NAND3_X1 i_0_2_841 (.A1(n_0_2_806), .A2(n_0_2_807), .A3(n_0_2_808), .ZN(
      n_0_2_809));
   NAND2_X1 i_0_2_842 (.A1(n_0_42), .A2(\Memory[8] [32]), .ZN(n_0_2_810));
   NAND2_X1 i_0_2_843 (.A1(n_0_35), .A2(\Memory[1] [32]), .ZN(n_0_2_811));
   NAND2_X1 i_0_2_844 (.A1(n_0_44), .A2(\Memory[10] [32]), .ZN(n_0_2_812));
   NAND3_X1 i_0_2_845 (.A1(n_0_2_810), .A2(n_0_2_811), .A3(n_0_2_812), .ZN(
      n_0_2_813));
   NOR2_X1 i_0_2_846 (.A1(n_0_2_809), .A2(n_0_2_813), .ZN(n_0_2_814));
   NAND2_X1 i_0_2_847 (.A1(n_0_48), .A2(\Memory[14] [32]), .ZN(n_0_2_815));
   NAND2_X1 i_0_2_848 (.A1(n_0_49), .A2(\Memory[15] [32]), .ZN(n_0_2_816));
   NAND2_X1 i_0_2_849 (.A1(n_0_34), .A2(\Memory[0] [32]), .ZN(n_0_2_817));
   NAND2_X1 i_0_2_850 (.A1(n_0_43), .A2(\Memory[9] [32]), .ZN(n_0_2_818));
   NAND4_X1 i_0_2_851 (.A1(n_0_2_815), .A2(n_0_2_816), .A3(n_0_2_817), .A4(
      n_0_2_818), .ZN(n_0_2_819));
   NAND2_X1 i_0_2_852 (.A1(n_0_47), .A2(\Memory[13] [32]), .ZN(n_0_2_820));
   NAND2_X1 i_0_2_853 (.A1(n_0_46), .A2(\Memory[12] [32]), .ZN(n_0_2_821));
   NAND2_X1 i_0_2_854 (.A1(n_0_45), .A2(\Memory[11] [32]), .ZN(n_0_2_822));
   NAND3_X1 i_0_2_855 (.A1(n_0_2_820), .A2(n_0_2_821), .A3(n_0_2_822), .ZN(
      n_0_2_823));
   NOR2_X1 i_0_2_856 (.A1(n_0_2_819), .A2(n_0_2_823), .ZN(n_0_2_824));
   NAND3_X1 i_0_2_857 (.A1(n_0_2_805), .A2(n_0_2_814), .A3(n_0_2_824), .ZN(
      dataOut1[32]));
   NAND2_X1 i_0_2_858 (.A1(n_0_38), .A2(\Memory[4] [33]), .ZN(n_0_2_825));
   NAND2_X1 i_0_2_859 (.A1(n_0_41), .A2(\Memory[7] [33]), .ZN(n_0_2_826));
   NAND2_X1 i_0_2_860 (.A1(n_0_37), .A2(\Memory[3] [33]), .ZN(n_0_2_827));
   NAND2_X1 i_0_2_861 (.A1(n_0_36), .A2(\Memory[2] [33]), .ZN(n_0_2_828));
   NAND4_X1 i_0_2_862 (.A1(n_0_2_825), .A2(n_0_2_826), .A3(n_0_2_827), .A4(
      n_0_2_828), .ZN(n_0_2_829));
   INV_X1 i_0_2_863 (.A(n_0_2_829), .ZN(n_0_2_830));
   NAND2_X1 i_0_2_864 (.A1(n_0_50), .A2(\Memory[16] [33]), .ZN(n_0_2_831));
   NAND2_X1 i_0_2_865 (.A1(n_0_40), .A2(\Memory[6] [33]), .ZN(n_0_2_832));
   NAND2_X1 i_0_2_866 (.A1(n_0_39), .A2(\Memory[5] [33]), .ZN(n_0_2_833));
   NAND3_X1 i_0_2_867 (.A1(n_0_2_831), .A2(n_0_2_832), .A3(n_0_2_833), .ZN(
      n_0_2_834));
   NAND2_X1 i_0_2_868 (.A1(n_0_42), .A2(\Memory[8] [33]), .ZN(n_0_2_835));
   NAND2_X1 i_0_2_869 (.A1(n_0_35), .A2(\Memory[1] [33]), .ZN(n_0_2_836));
   NAND2_X1 i_0_2_870 (.A1(n_0_44), .A2(\Memory[10] [33]), .ZN(n_0_2_837));
   NAND3_X1 i_0_2_871 (.A1(n_0_2_835), .A2(n_0_2_836), .A3(n_0_2_837), .ZN(
      n_0_2_838));
   NOR2_X1 i_0_2_872 (.A1(n_0_2_834), .A2(n_0_2_838), .ZN(n_0_2_839));
   NAND2_X1 i_0_2_873 (.A1(n_0_48), .A2(\Memory[14] [33]), .ZN(n_0_2_840));
   NAND2_X1 i_0_2_874 (.A1(n_0_49), .A2(\Memory[15] [33]), .ZN(n_0_2_841));
   NAND2_X1 i_0_2_875 (.A1(n_0_34), .A2(\Memory[0] [33]), .ZN(n_0_2_842));
   NAND2_X1 i_0_2_876 (.A1(n_0_43), .A2(\Memory[9] [33]), .ZN(n_0_2_843));
   NAND4_X1 i_0_2_877 (.A1(n_0_2_840), .A2(n_0_2_841), .A3(n_0_2_842), .A4(
      n_0_2_843), .ZN(n_0_2_844));
   NAND2_X1 i_0_2_878 (.A1(n_0_47), .A2(\Memory[13] [33]), .ZN(n_0_2_845));
   NAND2_X1 i_0_2_879 (.A1(n_0_46), .A2(\Memory[12] [33]), .ZN(n_0_2_846));
   NAND2_X1 i_0_2_880 (.A1(n_0_45), .A2(\Memory[11] [33]), .ZN(n_0_2_847));
   NAND3_X1 i_0_2_881 (.A1(n_0_2_845), .A2(n_0_2_846), .A3(n_0_2_847), .ZN(
      n_0_2_848));
   NOR2_X1 i_0_2_882 (.A1(n_0_2_844), .A2(n_0_2_848), .ZN(n_0_2_849));
   NAND3_X1 i_0_2_883 (.A1(n_0_2_830), .A2(n_0_2_839), .A3(n_0_2_849), .ZN(
      dataOut1[33]));
   NAND2_X1 i_0_2_884 (.A1(n_0_38), .A2(\Memory[4] [34]), .ZN(n_0_2_850));
   NAND2_X1 i_0_2_885 (.A1(n_0_41), .A2(\Memory[7] [34]), .ZN(n_0_2_851));
   NAND2_X1 i_0_2_886 (.A1(n_0_37), .A2(\Memory[3] [34]), .ZN(n_0_2_852));
   NAND2_X1 i_0_2_887 (.A1(n_0_36), .A2(\Memory[2] [34]), .ZN(n_0_2_853));
   NAND4_X1 i_0_2_888 (.A1(n_0_2_850), .A2(n_0_2_851), .A3(n_0_2_852), .A4(
      n_0_2_853), .ZN(n_0_2_854));
   INV_X1 i_0_2_889 (.A(n_0_2_854), .ZN(n_0_2_855));
   NAND2_X1 i_0_2_890 (.A1(n_0_50), .A2(\Memory[16] [34]), .ZN(n_0_2_856));
   NAND2_X1 i_0_2_891 (.A1(n_0_40), .A2(\Memory[6] [34]), .ZN(n_0_2_857));
   NAND2_X1 i_0_2_892 (.A1(n_0_39), .A2(\Memory[5] [34]), .ZN(n_0_2_858));
   NAND3_X1 i_0_2_893 (.A1(n_0_2_856), .A2(n_0_2_857), .A3(n_0_2_858), .ZN(
      n_0_2_859));
   NAND2_X1 i_0_2_894 (.A1(n_0_42), .A2(\Memory[8] [34]), .ZN(n_0_2_860));
   NAND2_X1 i_0_2_895 (.A1(n_0_35), .A2(\Memory[1] [34]), .ZN(n_0_2_861));
   NAND2_X1 i_0_2_896 (.A1(n_0_44), .A2(\Memory[10] [34]), .ZN(n_0_2_862));
   NAND3_X1 i_0_2_897 (.A1(n_0_2_860), .A2(n_0_2_861), .A3(n_0_2_862), .ZN(
      n_0_2_863));
   NOR2_X1 i_0_2_898 (.A1(n_0_2_859), .A2(n_0_2_863), .ZN(n_0_2_864));
   NAND2_X1 i_0_2_899 (.A1(n_0_48), .A2(\Memory[14] [34]), .ZN(n_0_2_865));
   NAND2_X1 i_0_2_900 (.A1(n_0_49), .A2(\Memory[15] [34]), .ZN(n_0_2_866));
   NAND2_X1 i_0_2_901 (.A1(n_0_34), .A2(\Memory[0] [34]), .ZN(n_0_2_867));
   NAND2_X1 i_0_2_902 (.A1(n_0_43), .A2(\Memory[9] [34]), .ZN(n_0_2_868));
   NAND4_X1 i_0_2_903 (.A1(n_0_2_865), .A2(n_0_2_866), .A3(n_0_2_867), .A4(
      n_0_2_868), .ZN(n_0_2_869));
   NAND2_X1 i_0_2_904 (.A1(n_0_47), .A2(\Memory[13] [34]), .ZN(n_0_2_870));
   NAND2_X1 i_0_2_905 (.A1(n_0_46), .A2(\Memory[12] [34]), .ZN(n_0_2_871));
   NAND2_X1 i_0_2_906 (.A1(n_0_45), .A2(\Memory[11] [34]), .ZN(n_0_2_872));
   NAND3_X1 i_0_2_907 (.A1(n_0_2_870), .A2(n_0_2_871), .A3(n_0_2_872), .ZN(
      n_0_2_873));
   NOR2_X1 i_0_2_908 (.A1(n_0_2_869), .A2(n_0_2_873), .ZN(n_0_2_874));
   NAND3_X1 i_0_2_909 (.A1(n_0_2_855), .A2(n_0_2_864), .A3(n_0_2_874), .ZN(
      dataOut1[34]));
   NAND2_X1 i_0_2_910 (.A1(n_0_38), .A2(\Memory[4] [35]), .ZN(n_0_2_875));
   NAND2_X1 i_0_2_911 (.A1(n_0_41), .A2(\Memory[7] [35]), .ZN(n_0_2_876));
   NAND2_X1 i_0_2_912 (.A1(n_0_37), .A2(\Memory[3] [35]), .ZN(n_0_2_877));
   NAND2_X1 i_0_2_913 (.A1(n_0_36), .A2(\Memory[2] [35]), .ZN(n_0_2_878));
   NAND4_X1 i_0_2_914 (.A1(n_0_2_875), .A2(n_0_2_876), .A3(n_0_2_877), .A4(
      n_0_2_878), .ZN(n_0_2_879));
   INV_X1 i_0_2_915 (.A(n_0_2_879), .ZN(n_0_2_880));
   NAND2_X1 i_0_2_916 (.A1(n_0_50), .A2(\Memory[16] [35]), .ZN(n_0_2_881));
   NAND2_X1 i_0_2_917 (.A1(n_0_40), .A2(\Memory[6] [35]), .ZN(n_0_2_882));
   NAND2_X1 i_0_2_918 (.A1(n_0_39), .A2(\Memory[5] [35]), .ZN(n_0_2_883));
   NAND3_X1 i_0_2_919 (.A1(n_0_2_881), .A2(n_0_2_882), .A3(n_0_2_883), .ZN(
      n_0_2_884));
   NAND2_X1 i_0_2_920 (.A1(n_0_42), .A2(\Memory[8] [35]), .ZN(n_0_2_885));
   NAND2_X1 i_0_2_921 (.A1(n_0_35), .A2(\Memory[1] [35]), .ZN(n_0_2_886));
   NAND2_X1 i_0_2_922 (.A1(n_0_44), .A2(\Memory[10] [35]), .ZN(n_0_2_887));
   NAND3_X1 i_0_2_923 (.A1(n_0_2_885), .A2(n_0_2_886), .A3(n_0_2_887), .ZN(
      n_0_2_888));
   NOR2_X1 i_0_2_924 (.A1(n_0_2_884), .A2(n_0_2_888), .ZN(n_0_2_889));
   NAND2_X1 i_0_2_925 (.A1(n_0_48), .A2(\Memory[14] [35]), .ZN(n_0_2_890));
   NAND2_X1 i_0_2_926 (.A1(n_0_49), .A2(\Memory[15] [35]), .ZN(n_0_2_891));
   NAND2_X1 i_0_2_927 (.A1(n_0_34), .A2(\Memory[0] [35]), .ZN(n_0_2_892));
   NAND2_X1 i_0_2_928 (.A1(n_0_43), .A2(\Memory[9] [35]), .ZN(n_0_2_893));
   NAND4_X1 i_0_2_929 (.A1(n_0_2_890), .A2(n_0_2_891), .A3(n_0_2_892), .A4(
      n_0_2_893), .ZN(n_0_2_894));
   NAND2_X1 i_0_2_930 (.A1(n_0_47), .A2(\Memory[13] [35]), .ZN(n_0_2_895));
   NAND2_X1 i_0_2_931 (.A1(n_0_46), .A2(\Memory[12] [35]), .ZN(n_0_2_896));
   NAND2_X1 i_0_2_932 (.A1(n_0_45), .A2(\Memory[11] [35]), .ZN(n_0_2_897));
   NAND3_X1 i_0_2_933 (.A1(n_0_2_895), .A2(n_0_2_896), .A3(n_0_2_897), .ZN(
      n_0_2_898));
   NOR2_X1 i_0_2_934 (.A1(n_0_2_894), .A2(n_0_2_898), .ZN(n_0_2_899));
   NAND3_X1 i_0_2_935 (.A1(n_0_2_880), .A2(n_0_2_889), .A3(n_0_2_899), .ZN(
      dataOut1[35]));
   NAND2_X1 i_0_2_936 (.A1(n_0_38), .A2(\Memory[4] [36]), .ZN(n_0_2_900));
   NAND2_X1 i_0_2_937 (.A1(n_0_41), .A2(\Memory[7] [36]), .ZN(n_0_2_901));
   NAND2_X1 i_0_2_938 (.A1(n_0_37), .A2(\Memory[3] [36]), .ZN(n_0_2_902));
   NAND2_X1 i_0_2_939 (.A1(n_0_36), .A2(\Memory[2] [36]), .ZN(n_0_2_903));
   NAND4_X1 i_0_2_940 (.A1(n_0_2_900), .A2(n_0_2_901), .A3(n_0_2_902), .A4(
      n_0_2_903), .ZN(n_0_2_904));
   INV_X1 i_0_2_941 (.A(n_0_2_904), .ZN(n_0_2_905));
   NAND2_X1 i_0_2_942 (.A1(n_0_50), .A2(\Memory[16] [36]), .ZN(n_0_2_906));
   NAND2_X1 i_0_2_943 (.A1(n_0_40), .A2(\Memory[6] [36]), .ZN(n_0_2_907));
   NAND2_X1 i_0_2_944 (.A1(n_0_39), .A2(\Memory[5] [36]), .ZN(n_0_2_908));
   NAND3_X1 i_0_2_945 (.A1(n_0_2_906), .A2(n_0_2_907), .A3(n_0_2_908), .ZN(
      n_0_2_909));
   NAND2_X1 i_0_2_946 (.A1(n_0_42), .A2(\Memory[8] [36]), .ZN(n_0_2_910));
   NAND2_X1 i_0_2_947 (.A1(n_0_35), .A2(\Memory[1] [36]), .ZN(n_0_2_911));
   NAND2_X1 i_0_2_948 (.A1(n_0_44), .A2(\Memory[10] [36]), .ZN(n_0_2_912));
   NAND3_X1 i_0_2_949 (.A1(n_0_2_910), .A2(n_0_2_911), .A3(n_0_2_912), .ZN(
      n_0_2_913));
   NOR2_X1 i_0_2_950 (.A1(n_0_2_909), .A2(n_0_2_913), .ZN(n_0_2_914));
   NAND2_X1 i_0_2_951 (.A1(n_0_48), .A2(\Memory[14] [36]), .ZN(n_0_2_915));
   NAND2_X1 i_0_2_952 (.A1(n_0_49), .A2(\Memory[15] [36]), .ZN(n_0_2_916));
   NAND2_X1 i_0_2_953 (.A1(n_0_34), .A2(\Memory[0] [36]), .ZN(n_0_2_917));
   NAND2_X1 i_0_2_954 (.A1(n_0_43), .A2(\Memory[9] [36]), .ZN(n_0_2_918));
   NAND4_X1 i_0_2_955 (.A1(n_0_2_915), .A2(n_0_2_916), .A3(n_0_2_917), .A4(
      n_0_2_918), .ZN(n_0_2_919));
   NAND2_X1 i_0_2_956 (.A1(n_0_47), .A2(\Memory[13] [36]), .ZN(n_0_2_920));
   NAND2_X1 i_0_2_957 (.A1(n_0_46), .A2(\Memory[12] [36]), .ZN(n_0_2_921));
   NAND2_X1 i_0_2_958 (.A1(n_0_45), .A2(\Memory[11] [36]), .ZN(n_0_2_922));
   NAND3_X1 i_0_2_959 (.A1(n_0_2_920), .A2(n_0_2_921), .A3(n_0_2_922), .ZN(
      n_0_2_923));
   NOR2_X1 i_0_2_960 (.A1(n_0_2_919), .A2(n_0_2_923), .ZN(n_0_2_924));
   NAND3_X1 i_0_2_961 (.A1(n_0_2_905), .A2(n_0_2_914), .A3(n_0_2_924), .ZN(
      dataOut1[36]));
   NAND2_X1 i_0_2_962 (.A1(n_0_38), .A2(\Memory[4] [37]), .ZN(n_0_2_925));
   NAND2_X1 i_0_2_963 (.A1(n_0_41), .A2(\Memory[7] [37]), .ZN(n_0_2_926));
   NAND2_X1 i_0_2_964 (.A1(n_0_37), .A2(\Memory[3] [37]), .ZN(n_0_2_927));
   NAND2_X1 i_0_2_965 (.A1(n_0_36), .A2(\Memory[2] [37]), .ZN(n_0_2_928));
   NAND4_X1 i_0_2_966 (.A1(n_0_2_925), .A2(n_0_2_926), .A3(n_0_2_927), .A4(
      n_0_2_928), .ZN(n_0_2_929));
   INV_X1 i_0_2_967 (.A(n_0_2_929), .ZN(n_0_2_930));
   NAND2_X1 i_0_2_968 (.A1(n_0_50), .A2(\Memory[16] [37]), .ZN(n_0_2_931));
   NAND2_X1 i_0_2_969 (.A1(n_0_40), .A2(\Memory[6] [37]), .ZN(n_0_2_932));
   NAND2_X1 i_0_2_970 (.A1(n_0_39), .A2(\Memory[5] [37]), .ZN(n_0_2_933));
   NAND3_X1 i_0_2_971 (.A1(n_0_2_931), .A2(n_0_2_932), .A3(n_0_2_933), .ZN(
      n_0_2_934));
   NAND2_X1 i_0_2_972 (.A1(n_0_42), .A2(\Memory[8] [37]), .ZN(n_0_2_935));
   NAND2_X1 i_0_2_973 (.A1(n_0_35), .A2(\Memory[1] [37]), .ZN(n_0_2_936));
   NAND2_X1 i_0_2_974 (.A1(n_0_44), .A2(\Memory[10] [37]), .ZN(n_0_2_937));
   NAND3_X1 i_0_2_975 (.A1(n_0_2_935), .A2(n_0_2_936), .A3(n_0_2_937), .ZN(
      n_0_2_938));
   NOR2_X1 i_0_2_976 (.A1(n_0_2_934), .A2(n_0_2_938), .ZN(n_0_2_939));
   NAND2_X1 i_0_2_977 (.A1(n_0_48), .A2(\Memory[14] [37]), .ZN(n_0_2_940));
   NAND2_X1 i_0_2_978 (.A1(n_0_49), .A2(\Memory[15] [37]), .ZN(n_0_2_941));
   NAND2_X1 i_0_2_979 (.A1(n_0_34), .A2(\Memory[0] [37]), .ZN(n_0_2_942));
   NAND2_X1 i_0_2_980 (.A1(n_0_43), .A2(\Memory[9] [37]), .ZN(n_0_2_943));
   NAND4_X1 i_0_2_981 (.A1(n_0_2_940), .A2(n_0_2_941), .A3(n_0_2_942), .A4(
      n_0_2_943), .ZN(n_0_2_944));
   NAND2_X1 i_0_2_982 (.A1(n_0_47), .A2(\Memory[13] [37]), .ZN(n_0_2_945));
   NAND2_X1 i_0_2_983 (.A1(n_0_46), .A2(\Memory[12] [37]), .ZN(n_0_2_946));
   NAND2_X1 i_0_2_984 (.A1(n_0_45), .A2(\Memory[11] [37]), .ZN(n_0_2_947));
   NAND3_X1 i_0_2_985 (.A1(n_0_2_945), .A2(n_0_2_946), .A3(n_0_2_947), .ZN(
      n_0_2_948));
   NOR2_X1 i_0_2_986 (.A1(n_0_2_944), .A2(n_0_2_948), .ZN(n_0_2_949));
   NAND3_X1 i_0_2_987 (.A1(n_0_2_930), .A2(n_0_2_939), .A3(n_0_2_949), .ZN(
      dataOut1[37]));
   NAND2_X1 i_0_2_988 (.A1(n_0_38), .A2(\Memory[4] [38]), .ZN(n_0_2_950));
   NAND2_X1 i_0_2_989 (.A1(n_0_41), .A2(\Memory[7] [38]), .ZN(n_0_2_951));
   NAND2_X1 i_0_2_990 (.A1(n_0_37), .A2(\Memory[3] [38]), .ZN(n_0_2_952));
   NAND2_X1 i_0_2_991 (.A1(n_0_36), .A2(\Memory[2] [38]), .ZN(n_0_2_953));
   NAND4_X1 i_0_2_992 (.A1(n_0_2_950), .A2(n_0_2_951), .A3(n_0_2_952), .A4(
      n_0_2_953), .ZN(n_0_2_954));
   INV_X1 i_0_2_993 (.A(n_0_2_954), .ZN(n_0_2_955));
   NAND2_X1 i_0_2_994 (.A1(n_0_50), .A2(\Memory[16] [38]), .ZN(n_0_2_956));
   NAND2_X1 i_0_2_995 (.A1(n_0_40), .A2(\Memory[6] [38]), .ZN(n_0_2_957));
   NAND2_X1 i_0_2_996 (.A1(n_0_39), .A2(\Memory[5] [38]), .ZN(n_0_2_958));
   NAND3_X1 i_0_2_997 (.A1(n_0_2_956), .A2(n_0_2_957), .A3(n_0_2_958), .ZN(
      n_0_2_959));
   NAND2_X1 i_0_2_998 (.A1(n_0_42), .A2(\Memory[8] [38]), .ZN(n_0_2_960));
   NAND2_X1 i_0_2_999 (.A1(n_0_35), .A2(\Memory[1] [38]), .ZN(n_0_2_961));
   NAND2_X1 i_0_2_1000 (.A1(n_0_44), .A2(\Memory[10] [38]), .ZN(n_0_2_962));
   NAND3_X1 i_0_2_1001 (.A1(n_0_2_960), .A2(n_0_2_961), .A3(n_0_2_962), .ZN(
      n_0_2_963));
   NOR2_X1 i_0_2_1002 (.A1(n_0_2_959), .A2(n_0_2_963), .ZN(n_0_2_964));
   NAND2_X1 i_0_2_1003 (.A1(n_0_48), .A2(\Memory[14] [38]), .ZN(n_0_2_965));
   NAND2_X1 i_0_2_1004 (.A1(n_0_49), .A2(\Memory[15] [38]), .ZN(n_0_2_966));
   NAND2_X1 i_0_2_1005 (.A1(n_0_34), .A2(\Memory[0] [38]), .ZN(n_0_2_967));
   NAND2_X1 i_0_2_1006 (.A1(n_0_43), .A2(\Memory[9] [38]), .ZN(n_0_2_968));
   NAND4_X1 i_0_2_1007 (.A1(n_0_2_965), .A2(n_0_2_966), .A3(n_0_2_967), .A4(
      n_0_2_968), .ZN(n_0_2_969));
   NAND2_X1 i_0_2_1008 (.A1(n_0_47), .A2(\Memory[13] [38]), .ZN(n_0_2_970));
   NAND2_X1 i_0_2_1009 (.A1(n_0_46), .A2(\Memory[12] [38]), .ZN(n_0_2_971));
   NAND2_X1 i_0_2_1010 (.A1(n_0_45), .A2(\Memory[11] [38]), .ZN(n_0_2_972));
   NAND3_X1 i_0_2_1011 (.A1(n_0_2_970), .A2(n_0_2_971), .A3(n_0_2_972), .ZN(
      n_0_2_973));
   NOR2_X1 i_0_2_1012 (.A1(n_0_2_969), .A2(n_0_2_973), .ZN(n_0_2_974));
   NAND3_X1 i_0_2_1013 (.A1(n_0_2_955), .A2(n_0_2_964), .A3(n_0_2_974), .ZN(
      dataOut1[38]));
   NAND2_X1 i_0_2_1014 (.A1(n_0_38), .A2(\Memory[4] [39]), .ZN(n_0_2_975));
   NAND2_X1 i_0_2_1015 (.A1(n_0_41), .A2(\Memory[7] [39]), .ZN(n_0_2_976));
   NAND2_X1 i_0_2_1016 (.A1(n_0_37), .A2(\Memory[3] [39]), .ZN(n_0_2_977));
   NAND2_X1 i_0_2_1017 (.A1(n_0_36), .A2(\Memory[2] [39]), .ZN(n_0_2_978));
   NAND4_X1 i_0_2_1018 (.A1(n_0_2_975), .A2(n_0_2_976), .A3(n_0_2_977), .A4(
      n_0_2_978), .ZN(n_0_2_979));
   INV_X1 i_0_2_1019 (.A(n_0_2_979), .ZN(n_0_2_980));
   NAND2_X1 i_0_2_1020 (.A1(n_0_50), .A2(\Memory[16] [39]), .ZN(n_0_2_981));
   NAND2_X1 i_0_2_1021 (.A1(n_0_40), .A2(\Memory[6] [39]), .ZN(n_0_2_982));
   NAND2_X1 i_0_2_1022 (.A1(n_0_39), .A2(\Memory[5] [39]), .ZN(n_0_2_983));
   NAND3_X1 i_0_2_1023 (.A1(n_0_2_981), .A2(n_0_2_982), .A3(n_0_2_983), .ZN(
      n_0_2_984));
   NAND2_X1 i_0_2_1024 (.A1(n_0_42), .A2(\Memory[8] [39]), .ZN(n_0_2_985));
   NAND2_X1 i_0_2_1025 (.A1(n_0_35), .A2(\Memory[1] [39]), .ZN(n_0_2_986));
   NAND2_X1 i_0_2_1026 (.A1(n_0_44), .A2(\Memory[10] [39]), .ZN(n_0_2_987));
   NAND3_X1 i_0_2_1027 (.A1(n_0_2_985), .A2(n_0_2_986), .A3(n_0_2_987), .ZN(
      n_0_2_988));
   NOR2_X1 i_0_2_1028 (.A1(n_0_2_984), .A2(n_0_2_988), .ZN(n_0_2_989));
   NAND2_X1 i_0_2_1029 (.A1(n_0_48), .A2(\Memory[14] [39]), .ZN(n_0_2_990));
   NAND2_X1 i_0_2_1030 (.A1(n_0_49), .A2(\Memory[15] [39]), .ZN(n_0_2_991));
   NAND2_X1 i_0_2_1031 (.A1(n_0_34), .A2(\Memory[0] [39]), .ZN(n_0_2_992));
   NAND2_X1 i_0_2_1032 (.A1(n_0_43), .A2(\Memory[9] [39]), .ZN(n_0_2_993));
   NAND4_X1 i_0_2_1033 (.A1(n_0_2_990), .A2(n_0_2_991), .A3(n_0_2_992), .A4(
      n_0_2_993), .ZN(n_0_2_994));
   NAND2_X1 i_0_2_1034 (.A1(n_0_47), .A2(\Memory[13] [39]), .ZN(n_0_2_995));
   NAND2_X1 i_0_2_1035 (.A1(n_0_46), .A2(\Memory[12] [39]), .ZN(n_0_2_996));
   NAND2_X1 i_0_2_1036 (.A1(n_0_45), .A2(\Memory[11] [39]), .ZN(n_0_2_997));
   NAND3_X1 i_0_2_1037 (.A1(n_0_2_995), .A2(n_0_2_996), .A3(n_0_2_997), .ZN(
      n_0_2_998));
   NOR2_X1 i_0_2_1038 (.A1(n_0_2_994), .A2(n_0_2_998), .ZN(n_0_2_999));
   NAND3_X1 i_0_2_1039 (.A1(n_0_2_980), .A2(n_0_2_989), .A3(n_0_2_999), .ZN(
      dataOut1[39]));
   NAND2_X1 i_0_2_1040 (.A1(n_0_38), .A2(\Memory[4] [40]), .ZN(n_0_2_1000));
   NAND2_X1 i_0_2_1041 (.A1(n_0_41), .A2(\Memory[7] [40]), .ZN(n_0_2_1001));
   NAND2_X1 i_0_2_1042 (.A1(n_0_37), .A2(\Memory[3] [40]), .ZN(n_0_2_1002));
   NAND2_X1 i_0_2_1043 (.A1(n_0_36), .A2(\Memory[2] [40]), .ZN(n_0_2_1003));
   NAND4_X1 i_0_2_1044 (.A1(n_0_2_1000), .A2(n_0_2_1001), .A3(n_0_2_1002), 
      .A4(n_0_2_1003), .ZN(n_0_2_1004));
   INV_X1 i_0_2_1045 (.A(n_0_2_1004), .ZN(n_0_2_1005));
   NAND2_X1 i_0_2_1046 (.A1(n_0_50), .A2(\Memory[16] [40]), .ZN(n_0_2_1006));
   NAND2_X1 i_0_2_1047 (.A1(n_0_40), .A2(\Memory[6] [40]), .ZN(n_0_2_1007));
   NAND2_X1 i_0_2_1048 (.A1(n_0_39), .A2(\Memory[5] [40]), .ZN(n_0_2_1008));
   NAND3_X1 i_0_2_1049 (.A1(n_0_2_1006), .A2(n_0_2_1007), .A3(n_0_2_1008), 
      .ZN(n_0_2_1009));
   NAND2_X1 i_0_2_1050 (.A1(n_0_42), .A2(\Memory[8] [40]), .ZN(n_0_2_1010));
   NAND2_X1 i_0_2_1051 (.A1(n_0_35), .A2(\Memory[1] [40]), .ZN(n_0_2_1011));
   NAND2_X1 i_0_2_1052 (.A1(n_0_44), .A2(\Memory[10] [40]), .ZN(n_0_2_1012));
   NAND3_X1 i_0_2_1053 (.A1(n_0_2_1010), .A2(n_0_2_1011), .A3(n_0_2_1012), 
      .ZN(n_0_2_1013));
   NOR2_X1 i_0_2_1054 (.A1(n_0_2_1009), .A2(n_0_2_1013), .ZN(n_0_2_1014));
   NAND2_X1 i_0_2_1055 (.A1(n_0_48), .A2(\Memory[14] [40]), .ZN(n_0_2_1015));
   NAND2_X1 i_0_2_1056 (.A1(n_0_49), .A2(\Memory[15] [40]), .ZN(n_0_2_1016));
   NAND2_X1 i_0_2_1057 (.A1(n_0_34), .A2(\Memory[0] [40]), .ZN(n_0_2_1017));
   NAND2_X1 i_0_2_1058 (.A1(n_0_43), .A2(\Memory[9] [40]), .ZN(n_0_2_1018));
   NAND4_X1 i_0_2_1059 (.A1(n_0_2_1015), .A2(n_0_2_1016), .A3(n_0_2_1017), 
      .A4(n_0_2_1018), .ZN(n_0_2_1019));
   NAND2_X1 i_0_2_1060 (.A1(n_0_47), .A2(\Memory[13] [40]), .ZN(n_0_2_1020));
   NAND2_X1 i_0_2_1061 (.A1(n_0_46), .A2(\Memory[12] [40]), .ZN(n_0_2_1021));
   NAND2_X1 i_0_2_1062 (.A1(n_0_45), .A2(\Memory[11] [40]), .ZN(n_0_2_1022));
   NAND3_X1 i_0_2_1063 (.A1(n_0_2_1020), .A2(n_0_2_1021), .A3(n_0_2_1022), 
      .ZN(n_0_2_1023));
   NOR2_X1 i_0_2_1064 (.A1(n_0_2_1019), .A2(n_0_2_1023), .ZN(n_0_2_1024));
   NAND3_X1 i_0_2_1065 (.A1(n_0_2_1005), .A2(n_0_2_1014), .A3(n_0_2_1024), 
      .ZN(dataOut1[40]));
   NAND2_X1 i_0_2_1066 (.A1(n_0_38), .A2(\Memory[4] [41]), .ZN(n_0_2_1025));
   NAND2_X1 i_0_2_1067 (.A1(n_0_41), .A2(\Memory[7] [41]), .ZN(n_0_2_1026));
   NAND2_X1 i_0_2_1068 (.A1(n_0_37), .A2(\Memory[3] [41]), .ZN(n_0_2_1027));
   NAND2_X1 i_0_2_1069 (.A1(n_0_36), .A2(\Memory[2] [41]), .ZN(n_0_2_1028));
   NAND4_X1 i_0_2_1070 (.A1(n_0_2_1025), .A2(n_0_2_1026), .A3(n_0_2_1027), 
      .A4(n_0_2_1028), .ZN(n_0_2_1029));
   INV_X1 i_0_2_1071 (.A(n_0_2_1029), .ZN(n_0_2_1030));
   NAND2_X1 i_0_2_1072 (.A1(n_0_50), .A2(\Memory[16] [41]), .ZN(n_0_2_1031));
   NAND2_X1 i_0_2_1073 (.A1(n_0_40), .A2(\Memory[6] [41]), .ZN(n_0_2_1032));
   NAND2_X1 i_0_2_1074 (.A1(n_0_39), .A2(\Memory[5] [41]), .ZN(n_0_2_1033));
   NAND3_X1 i_0_2_1075 (.A1(n_0_2_1031), .A2(n_0_2_1032), .A3(n_0_2_1033), 
      .ZN(n_0_2_1034));
   NAND2_X1 i_0_2_1076 (.A1(n_0_42), .A2(\Memory[8] [41]), .ZN(n_0_2_1035));
   NAND2_X1 i_0_2_1077 (.A1(n_0_35), .A2(\Memory[1] [41]), .ZN(n_0_2_1036));
   NAND2_X1 i_0_2_1078 (.A1(n_0_44), .A2(\Memory[10] [41]), .ZN(n_0_2_1037));
   NAND3_X1 i_0_2_1079 (.A1(n_0_2_1035), .A2(n_0_2_1036), .A3(n_0_2_1037), 
      .ZN(n_0_2_1038));
   NOR2_X1 i_0_2_1080 (.A1(n_0_2_1034), .A2(n_0_2_1038), .ZN(n_0_2_1039));
   NAND2_X1 i_0_2_1081 (.A1(n_0_48), .A2(\Memory[14] [41]), .ZN(n_0_2_1040));
   NAND2_X1 i_0_2_1082 (.A1(n_0_49), .A2(\Memory[15] [41]), .ZN(n_0_2_1041));
   NAND2_X1 i_0_2_1083 (.A1(n_0_34), .A2(\Memory[0] [41]), .ZN(n_0_2_1042));
   NAND2_X1 i_0_2_1084 (.A1(n_0_43), .A2(\Memory[9] [41]), .ZN(n_0_2_1043));
   NAND4_X1 i_0_2_1085 (.A1(n_0_2_1040), .A2(n_0_2_1041), .A3(n_0_2_1042), 
      .A4(n_0_2_1043), .ZN(n_0_2_1044));
   NAND2_X1 i_0_2_1086 (.A1(n_0_47), .A2(\Memory[13] [41]), .ZN(n_0_2_1045));
   NAND2_X1 i_0_2_1087 (.A1(n_0_46), .A2(\Memory[12] [41]), .ZN(n_0_2_1046));
   NAND2_X1 i_0_2_1088 (.A1(n_0_45), .A2(\Memory[11] [41]), .ZN(n_0_2_1047));
   NAND3_X1 i_0_2_1089 (.A1(n_0_2_1045), .A2(n_0_2_1046), .A3(n_0_2_1047), 
      .ZN(n_0_2_1048));
   NOR2_X1 i_0_2_1090 (.A1(n_0_2_1044), .A2(n_0_2_1048), .ZN(n_0_2_1049));
   NAND3_X1 i_0_2_1091 (.A1(n_0_2_1030), .A2(n_0_2_1039), .A3(n_0_2_1049), 
      .ZN(dataOut1[41]));
   NAND2_X1 i_0_2_1092 (.A1(n_0_38), .A2(\Memory[4] [42]), .ZN(n_0_2_1050));
   NAND2_X1 i_0_2_1093 (.A1(n_0_41), .A2(\Memory[7] [42]), .ZN(n_0_2_1051));
   NAND2_X1 i_0_2_1094 (.A1(n_0_37), .A2(\Memory[3] [42]), .ZN(n_0_2_1052));
   NAND2_X1 i_0_2_1095 (.A1(n_0_36), .A2(\Memory[2] [42]), .ZN(n_0_2_1053));
   NAND4_X1 i_0_2_1096 (.A1(n_0_2_1050), .A2(n_0_2_1051), .A3(n_0_2_1052), 
      .A4(n_0_2_1053), .ZN(n_0_2_1054));
   INV_X1 i_0_2_1097 (.A(n_0_2_1054), .ZN(n_0_2_1055));
   NAND2_X1 i_0_2_1098 (.A1(n_0_50), .A2(\Memory[16] [42]), .ZN(n_0_2_1056));
   NAND2_X1 i_0_2_1099 (.A1(n_0_40), .A2(\Memory[6] [42]), .ZN(n_0_2_1057));
   NAND2_X1 i_0_2_1100 (.A1(n_0_39), .A2(\Memory[5] [42]), .ZN(n_0_2_1058));
   NAND3_X1 i_0_2_1101 (.A1(n_0_2_1056), .A2(n_0_2_1057), .A3(n_0_2_1058), 
      .ZN(n_0_2_1059));
   NAND2_X1 i_0_2_1102 (.A1(n_0_42), .A2(\Memory[8] [42]), .ZN(n_0_2_1060));
   NAND2_X1 i_0_2_1103 (.A1(n_0_35), .A2(\Memory[1] [42]), .ZN(n_0_2_1061));
   NAND2_X1 i_0_2_1104 (.A1(n_0_44), .A2(\Memory[10] [42]), .ZN(n_0_2_1062));
   NAND3_X1 i_0_2_1105 (.A1(n_0_2_1060), .A2(n_0_2_1061), .A3(n_0_2_1062), 
      .ZN(n_0_2_1063));
   NOR2_X1 i_0_2_1106 (.A1(n_0_2_1059), .A2(n_0_2_1063), .ZN(n_0_2_1064));
   NAND2_X1 i_0_2_1107 (.A1(n_0_48), .A2(\Memory[14] [42]), .ZN(n_0_2_1065));
   NAND2_X1 i_0_2_1108 (.A1(n_0_49), .A2(\Memory[15] [42]), .ZN(n_0_2_1066));
   NAND2_X1 i_0_2_1109 (.A1(n_0_34), .A2(\Memory[0] [42]), .ZN(n_0_2_1067));
   NAND2_X1 i_0_2_1110 (.A1(n_0_43), .A2(\Memory[9] [42]), .ZN(n_0_2_1068));
   NAND4_X1 i_0_2_1111 (.A1(n_0_2_1065), .A2(n_0_2_1066), .A3(n_0_2_1067), 
      .A4(n_0_2_1068), .ZN(n_0_2_1069));
   NAND2_X1 i_0_2_1112 (.A1(n_0_47), .A2(\Memory[13] [42]), .ZN(n_0_2_1070));
   NAND2_X1 i_0_2_1113 (.A1(n_0_46), .A2(\Memory[12] [42]), .ZN(n_0_2_1071));
   NAND2_X1 i_0_2_1114 (.A1(n_0_45), .A2(\Memory[11] [42]), .ZN(n_0_2_1072));
   NAND3_X1 i_0_2_1115 (.A1(n_0_2_1070), .A2(n_0_2_1071), .A3(n_0_2_1072), 
      .ZN(n_0_2_1073));
   NOR2_X1 i_0_2_1116 (.A1(n_0_2_1069), .A2(n_0_2_1073), .ZN(n_0_2_1074));
   NAND3_X1 i_0_2_1117 (.A1(n_0_2_1055), .A2(n_0_2_1064), .A3(n_0_2_1074), 
      .ZN(dataOut1[42]));
   NAND2_X1 i_0_2_1118 (.A1(n_0_38), .A2(\Memory[4] [43]), .ZN(n_0_2_1075));
   NAND2_X1 i_0_2_1119 (.A1(n_0_41), .A2(\Memory[7] [43]), .ZN(n_0_2_1076));
   NAND2_X1 i_0_2_1120 (.A1(n_0_37), .A2(\Memory[3] [43]), .ZN(n_0_2_1077));
   NAND2_X1 i_0_2_1121 (.A1(n_0_36), .A2(\Memory[2] [43]), .ZN(n_0_2_1078));
   NAND4_X1 i_0_2_1122 (.A1(n_0_2_1075), .A2(n_0_2_1076), .A3(n_0_2_1077), 
      .A4(n_0_2_1078), .ZN(n_0_2_1079));
   INV_X1 i_0_2_1123 (.A(n_0_2_1079), .ZN(n_0_2_1080));
   NAND2_X1 i_0_2_1124 (.A1(n_0_50), .A2(\Memory[16] [43]), .ZN(n_0_2_1081));
   NAND2_X1 i_0_2_1125 (.A1(n_0_40), .A2(\Memory[6] [43]), .ZN(n_0_2_1082));
   NAND2_X1 i_0_2_1126 (.A1(n_0_39), .A2(\Memory[5] [43]), .ZN(n_0_2_1083));
   NAND3_X1 i_0_2_1127 (.A1(n_0_2_1081), .A2(n_0_2_1082), .A3(n_0_2_1083), 
      .ZN(n_0_2_1084));
   NAND2_X1 i_0_2_1128 (.A1(n_0_42), .A2(\Memory[8] [43]), .ZN(n_0_2_1085));
   NAND2_X1 i_0_2_1129 (.A1(n_0_35), .A2(\Memory[1] [43]), .ZN(n_0_2_1086));
   NAND2_X1 i_0_2_1130 (.A1(n_0_44), .A2(\Memory[10] [43]), .ZN(n_0_2_1087));
   NAND3_X1 i_0_2_1131 (.A1(n_0_2_1085), .A2(n_0_2_1086), .A3(n_0_2_1087), 
      .ZN(n_0_2_1088));
   NOR2_X1 i_0_2_1132 (.A1(n_0_2_1084), .A2(n_0_2_1088), .ZN(n_0_2_1089));
   NAND2_X1 i_0_2_1133 (.A1(n_0_48), .A2(\Memory[14] [43]), .ZN(n_0_2_1090));
   NAND2_X1 i_0_2_1134 (.A1(n_0_49), .A2(\Memory[15] [43]), .ZN(n_0_2_1091));
   NAND2_X1 i_0_2_1135 (.A1(n_0_34), .A2(\Memory[0] [43]), .ZN(n_0_2_1092));
   NAND2_X1 i_0_2_1136 (.A1(n_0_43), .A2(\Memory[9] [43]), .ZN(n_0_2_1093));
   NAND4_X1 i_0_2_1137 (.A1(n_0_2_1090), .A2(n_0_2_1091), .A3(n_0_2_1092), 
      .A4(n_0_2_1093), .ZN(n_0_2_1094));
   NAND2_X1 i_0_2_1138 (.A1(n_0_47), .A2(\Memory[13] [43]), .ZN(n_0_2_1095));
   NAND2_X1 i_0_2_1139 (.A1(n_0_46), .A2(\Memory[12] [43]), .ZN(n_0_2_1096));
   NAND2_X1 i_0_2_1140 (.A1(n_0_45), .A2(\Memory[11] [43]), .ZN(n_0_2_1097));
   NAND3_X1 i_0_2_1141 (.A1(n_0_2_1095), .A2(n_0_2_1096), .A3(n_0_2_1097), 
      .ZN(n_0_2_1098));
   NOR2_X1 i_0_2_1142 (.A1(n_0_2_1094), .A2(n_0_2_1098), .ZN(n_0_2_1099));
   NAND3_X1 i_0_2_1143 (.A1(n_0_2_1080), .A2(n_0_2_1089), .A3(n_0_2_1099), 
      .ZN(dataOut1[43]));
   NAND2_X1 i_0_2_1144 (.A1(n_0_38), .A2(\Memory[4] [44]), .ZN(n_0_2_1100));
   NAND2_X1 i_0_2_1145 (.A1(n_0_41), .A2(\Memory[7] [44]), .ZN(n_0_2_1101));
   NAND2_X1 i_0_2_1146 (.A1(n_0_37), .A2(\Memory[3] [44]), .ZN(n_0_2_1102));
   NAND2_X1 i_0_2_1147 (.A1(n_0_36), .A2(\Memory[2] [44]), .ZN(n_0_2_1103));
   NAND4_X1 i_0_2_1148 (.A1(n_0_2_1100), .A2(n_0_2_1101), .A3(n_0_2_1102), 
      .A4(n_0_2_1103), .ZN(n_0_2_1104));
   INV_X1 i_0_2_1149 (.A(n_0_2_1104), .ZN(n_0_2_1105));
   NAND2_X1 i_0_2_1150 (.A1(n_0_50), .A2(\Memory[16] [44]), .ZN(n_0_2_1106));
   NAND2_X1 i_0_2_1151 (.A1(n_0_40), .A2(\Memory[6] [44]), .ZN(n_0_2_1107));
   NAND2_X1 i_0_2_1152 (.A1(n_0_39), .A2(\Memory[5] [44]), .ZN(n_0_2_1108));
   NAND3_X1 i_0_2_1153 (.A1(n_0_2_1106), .A2(n_0_2_1107), .A3(n_0_2_1108), 
      .ZN(n_0_2_1109));
   NAND2_X1 i_0_2_1154 (.A1(n_0_42), .A2(\Memory[8] [44]), .ZN(n_0_2_1110));
   NAND2_X1 i_0_2_1155 (.A1(n_0_35), .A2(\Memory[1] [44]), .ZN(n_0_2_1111));
   NAND2_X1 i_0_2_1156 (.A1(n_0_44), .A2(\Memory[10] [44]), .ZN(n_0_2_1112));
   NAND3_X1 i_0_2_1157 (.A1(n_0_2_1110), .A2(n_0_2_1111), .A3(n_0_2_1112), 
      .ZN(n_0_2_1113));
   NOR2_X1 i_0_2_1158 (.A1(n_0_2_1109), .A2(n_0_2_1113), .ZN(n_0_2_1114));
   NAND2_X1 i_0_2_1159 (.A1(n_0_48), .A2(\Memory[14] [44]), .ZN(n_0_2_1115));
   NAND2_X1 i_0_2_1160 (.A1(n_0_49), .A2(\Memory[15] [44]), .ZN(n_0_2_1116));
   NAND2_X1 i_0_2_1161 (.A1(n_0_34), .A2(\Memory[0] [44]), .ZN(n_0_2_1117));
   NAND2_X1 i_0_2_1162 (.A1(n_0_43), .A2(\Memory[9] [44]), .ZN(n_0_2_1118));
   NAND4_X1 i_0_2_1163 (.A1(n_0_2_1115), .A2(n_0_2_1116), .A3(n_0_2_1117), 
      .A4(n_0_2_1118), .ZN(n_0_2_1119));
   NAND2_X1 i_0_2_1164 (.A1(n_0_47), .A2(\Memory[13] [44]), .ZN(n_0_2_1120));
   NAND2_X1 i_0_2_1165 (.A1(n_0_46), .A2(\Memory[12] [44]), .ZN(n_0_2_1121));
   NAND2_X1 i_0_2_1166 (.A1(n_0_45), .A2(\Memory[11] [44]), .ZN(n_0_2_1122));
   NAND3_X1 i_0_2_1167 (.A1(n_0_2_1120), .A2(n_0_2_1121), .A3(n_0_2_1122), 
      .ZN(n_0_2_1123));
   NOR2_X1 i_0_2_1168 (.A1(n_0_2_1119), .A2(n_0_2_1123), .ZN(n_0_2_1124));
   NAND3_X1 i_0_2_1169 (.A1(n_0_2_1105), .A2(n_0_2_1114), .A3(n_0_2_1124), 
      .ZN(dataOut1[44]));
   NAND2_X1 i_0_2_1170 (.A1(n_0_38), .A2(\Memory[4] [45]), .ZN(n_0_2_1125));
   NAND2_X1 i_0_2_1171 (.A1(n_0_41), .A2(\Memory[7] [45]), .ZN(n_0_2_1126));
   NAND2_X1 i_0_2_1172 (.A1(n_0_37), .A2(\Memory[3] [45]), .ZN(n_0_2_1127));
   NAND2_X1 i_0_2_1173 (.A1(n_0_36), .A2(\Memory[2] [45]), .ZN(n_0_2_1128));
   NAND4_X1 i_0_2_1174 (.A1(n_0_2_1125), .A2(n_0_2_1126), .A3(n_0_2_1127), 
      .A4(n_0_2_1128), .ZN(n_0_2_1129));
   INV_X1 i_0_2_1175 (.A(n_0_2_1129), .ZN(n_0_2_1130));
   NAND2_X1 i_0_2_1176 (.A1(n_0_50), .A2(\Memory[16] [45]), .ZN(n_0_2_1131));
   NAND2_X1 i_0_2_1177 (.A1(n_0_40), .A2(\Memory[6] [45]), .ZN(n_0_2_1132));
   NAND2_X1 i_0_2_1178 (.A1(n_0_39), .A2(\Memory[5] [45]), .ZN(n_0_2_1133));
   NAND3_X1 i_0_2_1179 (.A1(n_0_2_1131), .A2(n_0_2_1132), .A3(n_0_2_1133), 
      .ZN(n_0_2_1134));
   NAND2_X1 i_0_2_1180 (.A1(n_0_42), .A2(\Memory[8] [45]), .ZN(n_0_2_1135));
   NAND2_X1 i_0_2_1181 (.A1(n_0_35), .A2(\Memory[1] [45]), .ZN(n_0_2_1136));
   NAND2_X1 i_0_2_1182 (.A1(n_0_44), .A2(\Memory[10] [45]), .ZN(n_0_2_1137));
   NAND3_X1 i_0_2_1183 (.A1(n_0_2_1135), .A2(n_0_2_1136), .A3(n_0_2_1137), 
      .ZN(n_0_2_1138));
   NOR2_X1 i_0_2_1184 (.A1(n_0_2_1134), .A2(n_0_2_1138), .ZN(n_0_2_1139));
   NAND2_X1 i_0_2_1185 (.A1(n_0_48), .A2(\Memory[14] [45]), .ZN(n_0_2_1140));
   NAND2_X1 i_0_2_1186 (.A1(n_0_49), .A2(\Memory[15] [45]), .ZN(n_0_2_1141));
   NAND2_X1 i_0_2_1187 (.A1(n_0_34), .A2(\Memory[0] [45]), .ZN(n_0_2_1142));
   NAND2_X1 i_0_2_1188 (.A1(n_0_43), .A2(\Memory[9] [45]), .ZN(n_0_2_1143));
   NAND4_X1 i_0_2_1189 (.A1(n_0_2_1140), .A2(n_0_2_1141), .A3(n_0_2_1142), 
      .A4(n_0_2_1143), .ZN(n_0_2_1144));
   NAND2_X1 i_0_2_1190 (.A1(n_0_47), .A2(\Memory[13] [45]), .ZN(n_0_2_1145));
   NAND2_X1 i_0_2_1191 (.A1(n_0_46), .A2(\Memory[12] [45]), .ZN(n_0_2_1146));
   NAND2_X1 i_0_2_1192 (.A1(n_0_45), .A2(\Memory[11] [45]), .ZN(n_0_2_1147));
   NAND3_X1 i_0_2_1193 (.A1(n_0_2_1145), .A2(n_0_2_1146), .A3(n_0_2_1147), 
      .ZN(n_0_2_1148));
   NOR2_X1 i_0_2_1194 (.A1(n_0_2_1144), .A2(n_0_2_1148), .ZN(n_0_2_1149));
   NAND3_X1 i_0_2_1195 (.A1(n_0_2_1130), .A2(n_0_2_1139), .A3(n_0_2_1149), 
      .ZN(dataOut1[45]));
   NAND2_X1 i_0_2_1196 (.A1(n_0_38), .A2(\Memory[4] [46]), .ZN(n_0_2_1150));
   NAND2_X1 i_0_2_1197 (.A1(n_0_41), .A2(\Memory[7] [46]), .ZN(n_0_2_1151));
   NAND2_X1 i_0_2_1198 (.A1(n_0_37), .A2(\Memory[3] [46]), .ZN(n_0_2_1152));
   NAND2_X1 i_0_2_1199 (.A1(n_0_36), .A2(\Memory[2] [46]), .ZN(n_0_2_1153));
   NAND4_X1 i_0_2_1200 (.A1(n_0_2_1150), .A2(n_0_2_1151), .A3(n_0_2_1152), 
      .A4(n_0_2_1153), .ZN(n_0_2_1154));
   INV_X1 i_0_2_1201 (.A(n_0_2_1154), .ZN(n_0_2_1155));
   NAND2_X1 i_0_2_1202 (.A1(n_0_50), .A2(\Memory[16] [46]), .ZN(n_0_2_1156));
   NAND2_X1 i_0_2_1203 (.A1(n_0_40), .A2(\Memory[6] [46]), .ZN(n_0_2_1157));
   NAND2_X1 i_0_2_1204 (.A1(n_0_39), .A2(\Memory[5] [46]), .ZN(n_0_2_1158));
   NAND3_X1 i_0_2_1205 (.A1(n_0_2_1156), .A2(n_0_2_1157), .A3(n_0_2_1158), 
      .ZN(n_0_2_1159));
   NAND2_X1 i_0_2_1206 (.A1(n_0_42), .A2(\Memory[8] [46]), .ZN(n_0_2_1160));
   NAND2_X1 i_0_2_1207 (.A1(n_0_35), .A2(\Memory[1] [46]), .ZN(n_0_2_1161));
   NAND2_X1 i_0_2_1208 (.A1(n_0_44), .A2(\Memory[10] [46]), .ZN(n_0_2_1162));
   NAND3_X1 i_0_2_1209 (.A1(n_0_2_1160), .A2(n_0_2_1161), .A3(n_0_2_1162), 
      .ZN(n_0_2_1163));
   NOR2_X1 i_0_2_1210 (.A1(n_0_2_1159), .A2(n_0_2_1163), .ZN(n_0_2_1164));
   NAND2_X1 i_0_2_1211 (.A1(n_0_48), .A2(\Memory[14] [46]), .ZN(n_0_2_1165));
   NAND2_X1 i_0_2_1212 (.A1(n_0_49), .A2(\Memory[15] [46]), .ZN(n_0_2_1166));
   NAND2_X1 i_0_2_1213 (.A1(n_0_34), .A2(\Memory[0] [46]), .ZN(n_0_2_1167));
   NAND2_X1 i_0_2_1214 (.A1(n_0_43), .A2(\Memory[9] [46]), .ZN(n_0_2_1168));
   NAND4_X1 i_0_2_1215 (.A1(n_0_2_1165), .A2(n_0_2_1166), .A3(n_0_2_1167), 
      .A4(n_0_2_1168), .ZN(n_0_2_1169));
   NAND2_X1 i_0_2_1216 (.A1(n_0_47), .A2(\Memory[13] [46]), .ZN(n_0_2_1170));
   NAND2_X1 i_0_2_1217 (.A1(n_0_46), .A2(\Memory[12] [46]), .ZN(n_0_2_1171));
   NAND2_X1 i_0_2_1218 (.A1(n_0_45), .A2(\Memory[11] [46]), .ZN(n_0_2_1172));
   NAND3_X1 i_0_2_1219 (.A1(n_0_2_1170), .A2(n_0_2_1171), .A3(n_0_2_1172), 
      .ZN(n_0_2_1173));
   NOR2_X1 i_0_2_1220 (.A1(n_0_2_1169), .A2(n_0_2_1173), .ZN(n_0_2_1174));
   NAND3_X1 i_0_2_1221 (.A1(n_0_2_1155), .A2(n_0_2_1164), .A3(n_0_2_1174), 
      .ZN(dataOut1[46]));
   NAND2_X1 i_0_2_1222 (.A1(n_0_38), .A2(\Memory[4] [47]), .ZN(n_0_2_1175));
   NAND2_X1 i_0_2_1223 (.A1(n_0_41), .A2(\Memory[7] [47]), .ZN(n_0_2_1176));
   NAND2_X1 i_0_2_1224 (.A1(n_0_37), .A2(\Memory[3] [47]), .ZN(n_0_2_1177));
   NAND2_X1 i_0_2_1225 (.A1(n_0_36), .A2(\Memory[2] [47]), .ZN(n_0_2_1178));
   NAND4_X1 i_0_2_1226 (.A1(n_0_2_1175), .A2(n_0_2_1176), .A3(n_0_2_1177), 
      .A4(n_0_2_1178), .ZN(n_0_2_1179));
   INV_X1 i_0_2_1227 (.A(n_0_2_1179), .ZN(n_0_2_1180));
   NAND2_X1 i_0_2_1228 (.A1(n_0_50), .A2(\Memory[16] [47]), .ZN(n_0_2_1181));
   NAND2_X1 i_0_2_1229 (.A1(n_0_40), .A2(\Memory[6] [47]), .ZN(n_0_2_1182));
   NAND2_X1 i_0_2_1230 (.A1(n_0_39), .A2(\Memory[5] [47]), .ZN(n_0_2_1183));
   NAND3_X1 i_0_2_1231 (.A1(n_0_2_1181), .A2(n_0_2_1182), .A3(n_0_2_1183), 
      .ZN(n_0_2_1184));
   NAND2_X1 i_0_2_1232 (.A1(n_0_42), .A2(\Memory[8] [47]), .ZN(n_0_2_1185));
   NAND2_X1 i_0_2_1233 (.A1(n_0_35), .A2(\Memory[1] [47]), .ZN(n_0_2_1186));
   NAND2_X1 i_0_2_1234 (.A1(n_0_44), .A2(\Memory[10] [47]), .ZN(n_0_2_1187));
   NAND3_X1 i_0_2_1235 (.A1(n_0_2_1185), .A2(n_0_2_1186), .A3(n_0_2_1187), 
      .ZN(n_0_2_1188));
   NOR2_X1 i_0_2_1236 (.A1(n_0_2_1184), .A2(n_0_2_1188), .ZN(n_0_2_1189));
   NAND2_X1 i_0_2_1237 (.A1(n_0_48), .A2(\Memory[14] [47]), .ZN(n_0_2_1190));
   NAND2_X1 i_0_2_1238 (.A1(n_0_49), .A2(\Memory[15] [47]), .ZN(n_0_2_1191));
   NAND2_X1 i_0_2_1239 (.A1(n_0_34), .A2(\Memory[0] [47]), .ZN(n_0_2_1192));
   NAND2_X1 i_0_2_1240 (.A1(n_0_43), .A2(\Memory[9] [47]), .ZN(n_0_2_1193));
   NAND4_X1 i_0_2_1241 (.A1(n_0_2_1190), .A2(n_0_2_1191), .A3(n_0_2_1192), 
      .A4(n_0_2_1193), .ZN(n_0_2_1194));
   NAND2_X1 i_0_2_1242 (.A1(n_0_47), .A2(\Memory[13] [47]), .ZN(n_0_2_1195));
   NAND2_X1 i_0_2_1243 (.A1(n_0_46), .A2(\Memory[12] [47]), .ZN(n_0_2_1196));
   NAND2_X1 i_0_2_1244 (.A1(n_0_45), .A2(\Memory[11] [47]), .ZN(n_0_2_1197));
   NAND3_X1 i_0_2_1245 (.A1(n_0_2_1195), .A2(n_0_2_1196), .A3(n_0_2_1197), 
      .ZN(n_0_2_1198));
   NOR2_X1 i_0_2_1246 (.A1(n_0_2_1194), .A2(n_0_2_1198), .ZN(n_0_2_1199));
   NAND3_X1 i_0_2_1247 (.A1(n_0_2_1180), .A2(n_0_2_1189), .A3(n_0_2_1199), 
      .ZN(dataOut1[47]));
   NAND2_X1 i_0_2_1248 (.A1(n_0_38), .A2(\Memory[4] [48]), .ZN(n_0_2_1200));
   NAND2_X1 i_0_2_1249 (.A1(n_0_41), .A2(\Memory[7] [48]), .ZN(n_0_2_1201));
   NAND2_X1 i_0_2_1250 (.A1(n_0_37), .A2(\Memory[3] [48]), .ZN(n_0_2_1202));
   NAND2_X1 i_0_2_1251 (.A1(n_0_36), .A2(\Memory[2] [48]), .ZN(n_0_2_1203));
   NAND4_X1 i_0_2_1252 (.A1(n_0_2_1200), .A2(n_0_2_1201), .A3(n_0_2_1202), 
      .A4(n_0_2_1203), .ZN(n_0_2_1204));
   INV_X1 i_0_2_1253 (.A(n_0_2_1204), .ZN(n_0_2_1205));
   NAND2_X1 i_0_2_1254 (.A1(n_0_50), .A2(\Memory[16] [48]), .ZN(n_0_2_1206));
   NAND2_X1 i_0_2_1255 (.A1(n_0_40), .A2(\Memory[6] [48]), .ZN(n_0_2_1207));
   NAND2_X1 i_0_2_1256 (.A1(n_0_39), .A2(\Memory[5] [48]), .ZN(n_0_2_1208));
   NAND3_X1 i_0_2_1257 (.A1(n_0_2_1206), .A2(n_0_2_1207), .A3(n_0_2_1208), 
      .ZN(n_0_2_1209));
   NAND2_X1 i_0_2_1258 (.A1(n_0_42), .A2(\Memory[8] [48]), .ZN(n_0_2_1210));
   NAND2_X1 i_0_2_1259 (.A1(n_0_35), .A2(\Memory[1] [48]), .ZN(n_0_2_1211));
   NAND2_X1 i_0_2_1260 (.A1(n_0_44), .A2(\Memory[10] [48]), .ZN(n_0_2_1212));
   NAND3_X1 i_0_2_1261 (.A1(n_0_2_1210), .A2(n_0_2_1211), .A3(n_0_2_1212), 
      .ZN(n_0_2_1213));
   NOR2_X1 i_0_2_1262 (.A1(n_0_2_1209), .A2(n_0_2_1213), .ZN(n_0_2_1214));
   NAND2_X1 i_0_2_1263 (.A1(n_0_48), .A2(\Memory[14] [48]), .ZN(n_0_2_1215));
   NAND2_X1 i_0_2_1264 (.A1(n_0_49), .A2(\Memory[15] [48]), .ZN(n_0_2_1216));
   NAND2_X1 i_0_2_1265 (.A1(n_0_34), .A2(\Memory[0] [48]), .ZN(n_0_2_1217));
   NAND2_X1 i_0_2_1266 (.A1(n_0_43), .A2(\Memory[9] [48]), .ZN(n_0_2_1218));
   NAND4_X1 i_0_2_1267 (.A1(n_0_2_1215), .A2(n_0_2_1216), .A3(n_0_2_1217), 
      .A4(n_0_2_1218), .ZN(n_0_2_1219));
   NAND2_X1 i_0_2_1268 (.A1(n_0_47), .A2(\Memory[13] [48]), .ZN(n_0_2_1220));
   NAND2_X1 i_0_2_1269 (.A1(n_0_46), .A2(\Memory[12] [48]), .ZN(n_0_2_1221));
   NAND2_X1 i_0_2_1270 (.A1(n_0_45), .A2(\Memory[11] [48]), .ZN(n_0_2_1222));
   NAND3_X1 i_0_2_1271 (.A1(n_0_2_1220), .A2(n_0_2_1221), .A3(n_0_2_1222), 
      .ZN(n_0_2_1223));
   NOR2_X1 i_0_2_1272 (.A1(n_0_2_1219), .A2(n_0_2_1223), .ZN(n_0_2_1224));
   NAND3_X1 i_0_2_1273 (.A1(n_0_2_1205), .A2(n_0_2_1214), .A3(n_0_2_1224), 
      .ZN(dataOut1[48]));
   NAND2_X1 i_0_2_1274 (.A1(n_0_38), .A2(\Memory[4] [49]), .ZN(n_0_2_1225));
   NAND2_X1 i_0_2_1275 (.A1(n_0_41), .A2(\Memory[7] [49]), .ZN(n_0_2_1226));
   NAND2_X1 i_0_2_1276 (.A1(n_0_37), .A2(\Memory[3] [49]), .ZN(n_0_2_1227));
   NAND2_X1 i_0_2_1277 (.A1(n_0_36), .A2(\Memory[2] [49]), .ZN(n_0_2_1228));
   NAND4_X1 i_0_2_1278 (.A1(n_0_2_1225), .A2(n_0_2_1226), .A3(n_0_2_1227), 
      .A4(n_0_2_1228), .ZN(n_0_2_1229));
   INV_X1 i_0_2_1279 (.A(n_0_2_1229), .ZN(n_0_2_1230));
   NAND2_X1 i_0_2_1280 (.A1(n_0_50), .A2(\Memory[16] [49]), .ZN(n_0_2_1231));
   NAND2_X1 i_0_2_1281 (.A1(n_0_40), .A2(\Memory[6] [49]), .ZN(n_0_2_1232));
   NAND2_X1 i_0_2_1282 (.A1(n_0_39), .A2(\Memory[5] [49]), .ZN(n_0_2_1233));
   NAND3_X1 i_0_2_1283 (.A1(n_0_2_1231), .A2(n_0_2_1232), .A3(n_0_2_1233), 
      .ZN(n_0_2_1234));
   NAND2_X1 i_0_2_1284 (.A1(n_0_42), .A2(\Memory[8] [49]), .ZN(n_0_2_1235));
   NAND2_X1 i_0_2_1285 (.A1(n_0_35), .A2(\Memory[1] [49]), .ZN(n_0_2_1236));
   NAND2_X1 i_0_2_1286 (.A1(n_0_44), .A2(\Memory[10] [49]), .ZN(n_0_2_1237));
   NAND3_X1 i_0_2_1287 (.A1(n_0_2_1235), .A2(n_0_2_1236), .A3(n_0_2_1237), 
      .ZN(n_0_2_1238));
   NOR2_X1 i_0_2_1288 (.A1(n_0_2_1234), .A2(n_0_2_1238), .ZN(n_0_2_1239));
   NAND2_X1 i_0_2_1289 (.A1(n_0_48), .A2(\Memory[14] [49]), .ZN(n_0_2_1240));
   NAND2_X1 i_0_2_1290 (.A1(n_0_49), .A2(\Memory[15] [49]), .ZN(n_0_2_1241));
   NAND2_X1 i_0_2_1291 (.A1(n_0_34), .A2(\Memory[0] [49]), .ZN(n_0_2_1242));
   NAND2_X1 i_0_2_1292 (.A1(n_0_43), .A2(\Memory[9] [49]), .ZN(n_0_2_1243));
   NAND4_X1 i_0_2_1293 (.A1(n_0_2_1240), .A2(n_0_2_1241), .A3(n_0_2_1242), 
      .A4(n_0_2_1243), .ZN(n_0_2_1244));
   NAND2_X1 i_0_2_1294 (.A1(n_0_47), .A2(\Memory[13] [49]), .ZN(n_0_2_1245));
   NAND2_X1 i_0_2_1295 (.A1(n_0_46), .A2(\Memory[12] [49]), .ZN(n_0_2_1246));
   NAND2_X1 i_0_2_1296 (.A1(n_0_45), .A2(\Memory[11] [49]), .ZN(n_0_2_1247));
   NAND3_X1 i_0_2_1297 (.A1(n_0_2_1245), .A2(n_0_2_1246), .A3(n_0_2_1247), 
      .ZN(n_0_2_1248));
   NOR2_X1 i_0_2_1298 (.A1(n_0_2_1244), .A2(n_0_2_1248), .ZN(n_0_2_1249));
   NAND3_X1 i_0_2_1299 (.A1(n_0_2_1230), .A2(n_0_2_1239), .A3(n_0_2_1249), 
      .ZN(dataOut1[49]));
   NAND2_X1 i_0_2_1300 (.A1(n_0_38), .A2(\Memory[4] [50]), .ZN(n_0_2_1250));
   NAND2_X1 i_0_2_1301 (.A1(n_0_41), .A2(\Memory[7] [50]), .ZN(n_0_2_1251));
   NAND2_X1 i_0_2_1302 (.A1(n_0_37), .A2(\Memory[3] [50]), .ZN(n_0_2_1252));
   NAND2_X1 i_0_2_1303 (.A1(n_0_36), .A2(\Memory[2] [50]), .ZN(n_0_2_1253));
   NAND4_X1 i_0_2_1304 (.A1(n_0_2_1250), .A2(n_0_2_1251), .A3(n_0_2_1252), 
      .A4(n_0_2_1253), .ZN(n_0_2_1254));
   INV_X1 i_0_2_1305 (.A(n_0_2_1254), .ZN(n_0_2_1255));
   NAND2_X1 i_0_2_1306 (.A1(n_0_50), .A2(\Memory[16] [50]), .ZN(n_0_2_1256));
   NAND2_X1 i_0_2_1307 (.A1(n_0_40), .A2(\Memory[6] [50]), .ZN(n_0_2_1257));
   NAND2_X1 i_0_2_1308 (.A1(n_0_39), .A2(\Memory[5] [50]), .ZN(n_0_2_1258));
   NAND3_X1 i_0_2_1309 (.A1(n_0_2_1256), .A2(n_0_2_1257), .A3(n_0_2_1258), 
      .ZN(n_0_2_1259));
   NAND2_X1 i_0_2_1310 (.A1(n_0_42), .A2(\Memory[8] [50]), .ZN(n_0_2_1260));
   NAND2_X1 i_0_2_1311 (.A1(n_0_35), .A2(\Memory[1] [50]), .ZN(n_0_2_1261));
   NAND2_X1 i_0_2_1312 (.A1(n_0_44), .A2(\Memory[10] [50]), .ZN(n_0_2_1262));
   NAND3_X1 i_0_2_1313 (.A1(n_0_2_1260), .A2(n_0_2_1261), .A3(n_0_2_1262), 
      .ZN(n_0_2_1263));
   NOR2_X1 i_0_2_1314 (.A1(n_0_2_1259), .A2(n_0_2_1263), .ZN(n_0_2_1264));
   NAND2_X1 i_0_2_1315 (.A1(n_0_48), .A2(\Memory[14] [50]), .ZN(n_0_2_1265));
   NAND2_X1 i_0_2_1316 (.A1(n_0_49), .A2(\Memory[15] [50]), .ZN(n_0_2_1266));
   NAND2_X1 i_0_2_1317 (.A1(n_0_34), .A2(\Memory[0] [50]), .ZN(n_0_2_1267));
   NAND2_X1 i_0_2_1318 (.A1(n_0_43), .A2(\Memory[9] [50]), .ZN(n_0_2_1268));
   NAND4_X1 i_0_2_1319 (.A1(n_0_2_1265), .A2(n_0_2_1266), .A3(n_0_2_1267), 
      .A4(n_0_2_1268), .ZN(n_0_2_1269));
   NAND2_X1 i_0_2_1320 (.A1(n_0_47), .A2(\Memory[13] [50]), .ZN(n_0_2_1270));
   NAND2_X1 i_0_2_1321 (.A1(n_0_46), .A2(\Memory[12] [50]), .ZN(n_0_2_1271));
   NAND2_X1 i_0_2_1322 (.A1(n_0_45), .A2(\Memory[11] [50]), .ZN(n_0_2_1272));
   NAND3_X1 i_0_2_1323 (.A1(n_0_2_1270), .A2(n_0_2_1271), .A3(n_0_2_1272), 
      .ZN(n_0_2_1273));
   NOR2_X1 i_0_2_1324 (.A1(n_0_2_1269), .A2(n_0_2_1273), .ZN(n_0_2_1274));
   NAND3_X1 i_0_2_1325 (.A1(n_0_2_1255), .A2(n_0_2_1264), .A3(n_0_2_1274), 
      .ZN(dataOut1[50]));
   NAND2_X1 i_0_2_1326 (.A1(n_0_38), .A2(\Memory[4] [51]), .ZN(n_0_2_1275));
   NAND2_X1 i_0_2_1327 (.A1(n_0_41), .A2(\Memory[7] [51]), .ZN(n_0_2_1276));
   NAND2_X1 i_0_2_1328 (.A1(n_0_37), .A2(\Memory[3] [51]), .ZN(n_0_2_1277));
   NAND2_X1 i_0_2_1329 (.A1(n_0_36), .A2(\Memory[2] [51]), .ZN(n_0_2_1278));
   NAND4_X1 i_0_2_1330 (.A1(n_0_2_1275), .A2(n_0_2_1276), .A3(n_0_2_1277), 
      .A4(n_0_2_1278), .ZN(n_0_2_1279));
   INV_X1 i_0_2_1331 (.A(n_0_2_1279), .ZN(n_0_2_1280));
   NAND2_X1 i_0_2_1332 (.A1(n_0_50), .A2(\Memory[16] [51]), .ZN(n_0_2_1281));
   NAND2_X1 i_0_2_1333 (.A1(n_0_40), .A2(\Memory[6] [51]), .ZN(n_0_2_1282));
   NAND2_X1 i_0_2_1334 (.A1(n_0_39), .A2(\Memory[5] [51]), .ZN(n_0_2_1283));
   NAND3_X1 i_0_2_1335 (.A1(n_0_2_1281), .A2(n_0_2_1282), .A3(n_0_2_1283), 
      .ZN(n_0_2_1284));
   NAND2_X1 i_0_2_1336 (.A1(n_0_42), .A2(\Memory[8] [51]), .ZN(n_0_2_1285));
   NAND2_X1 i_0_2_1337 (.A1(n_0_35), .A2(\Memory[1] [51]), .ZN(n_0_2_1286));
   NAND2_X1 i_0_2_1338 (.A1(n_0_44), .A2(\Memory[10] [51]), .ZN(n_0_2_1287));
   NAND3_X1 i_0_2_1339 (.A1(n_0_2_1285), .A2(n_0_2_1286), .A3(n_0_2_1287), 
      .ZN(n_0_2_1288));
   NOR2_X1 i_0_2_1340 (.A1(n_0_2_1284), .A2(n_0_2_1288), .ZN(n_0_2_1289));
   NAND2_X1 i_0_2_1341 (.A1(n_0_48), .A2(\Memory[14] [51]), .ZN(n_0_2_1290));
   NAND2_X1 i_0_2_1342 (.A1(n_0_49), .A2(\Memory[15] [51]), .ZN(n_0_2_1291));
   NAND2_X1 i_0_2_1343 (.A1(n_0_34), .A2(\Memory[0] [51]), .ZN(n_0_2_1292));
   NAND2_X1 i_0_2_1344 (.A1(n_0_43), .A2(\Memory[9] [51]), .ZN(n_0_2_1293));
   NAND4_X1 i_0_2_1345 (.A1(n_0_2_1290), .A2(n_0_2_1291), .A3(n_0_2_1292), 
      .A4(n_0_2_1293), .ZN(n_0_2_1294));
   NAND2_X1 i_0_2_1346 (.A1(n_0_47), .A2(\Memory[13] [51]), .ZN(n_0_2_1295));
   NAND2_X1 i_0_2_1347 (.A1(n_0_46), .A2(\Memory[12] [51]), .ZN(n_0_2_1296));
   NAND2_X1 i_0_2_1348 (.A1(n_0_45), .A2(\Memory[11] [51]), .ZN(n_0_2_1297));
   NAND3_X1 i_0_2_1349 (.A1(n_0_2_1295), .A2(n_0_2_1296), .A3(n_0_2_1297), 
      .ZN(n_0_2_1298));
   NOR2_X1 i_0_2_1350 (.A1(n_0_2_1294), .A2(n_0_2_1298), .ZN(n_0_2_1299));
   NAND3_X1 i_0_2_1351 (.A1(n_0_2_1280), .A2(n_0_2_1289), .A3(n_0_2_1299), 
      .ZN(dataOut1[51]));
   NAND2_X1 i_0_2_1352 (.A1(n_0_38), .A2(\Memory[4] [52]), .ZN(n_0_2_1300));
   NAND2_X1 i_0_2_1353 (.A1(n_0_41), .A2(\Memory[7] [52]), .ZN(n_0_2_1301));
   NAND2_X1 i_0_2_1354 (.A1(n_0_37), .A2(\Memory[3] [52]), .ZN(n_0_2_1302));
   NAND2_X1 i_0_2_1355 (.A1(n_0_36), .A2(\Memory[2] [52]), .ZN(n_0_2_1303));
   NAND4_X1 i_0_2_1356 (.A1(n_0_2_1300), .A2(n_0_2_1301), .A3(n_0_2_1302), 
      .A4(n_0_2_1303), .ZN(n_0_2_1304));
   INV_X1 i_0_2_1357 (.A(n_0_2_1304), .ZN(n_0_2_1305));
   NAND2_X1 i_0_2_1358 (.A1(n_0_50), .A2(\Memory[16] [52]), .ZN(n_0_2_1306));
   NAND2_X1 i_0_2_1359 (.A1(n_0_40), .A2(\Memory[6] [52]), .ZN(n_0_2_1307));
   NAND2_X1 i_0_2_1360 (.A1(n_0_39), .A2(\Memory[5] [52]), .ZN(n_0_2_1308));
   NAND3_X1 i_0_2_1361 (.A1(n_0_2_1306), .A2(n_0_2_1307), .A3(n_0_2_1308), 
      .ZN(n_0_2_1309));
   NAND2_X1 i_0_2_1362 (.A1(n_0_42), .A2(\Memory[8] [52]), .ZN(n_0_2_1310));
   NAND2_X1 i_0_2_1363 (.A1(n_0_35), .A2(\Memory[1] [52]), .ZN(n_0_2_1311));
   NAND2_X1 i_0_2_1364 (.A1(n_0_44), .A2(\Memory[10] [52]), .ZN(n_0_2_1312));
   NAND3_X1 i_0_2_1365 (.A1(n_0_2_1310), .A2(n_0_2_1311), .A3(n_0_2_1312), 
      .ZN(n_0_2_1313));
   NOR2_X1 i_0_2_1366 (.A1(n_0_2_1309), .A2(n_0_2_1313), .ZN(n_0_2_1314));
   NAND2_X1 i_0_2_1367 (.A1(n_0_48), .A2(\Memory[14] [52]), .ZN(n_0_2_1315));
   NAND2_X1 i_0_2_1368 (.A1(n_0_49), .A2(\Memory[15] [52]), .ZN(n_0_2_1316));
   NAND2_X1 i_0_2_1369 (.A1(n_0_34), .A2(\Memory[0] [52]), .ZN(n_0_2_1317));
   NAND2_X1 i_0_2_1370 (.A1(n_0_43), .A2(\Memory[9] [52]), .ZN(n_0_2_1318));
   NAND4_X1 i_0_2_1371 (.A1(n_0_2_1315), .A2(n_0_2_1316), .A3(n_0_2_1317), 
      .A4(n_0_2_1318), .ZN(n_0_2_1319));
   NAND2_X1 i_0_2_1372 (.A1(n_0_47), .A2(\Memory[13] [52]), .ZN(n_0_2_1320));
   NAND2_X1 i_0_2_1373 (.A1(n_0_46), .A2(\Memory[12] [52]), .ZN(n_0_2_1321));
   NAND2_X1 i_0_2_1374 (.A1(n_0_45), .A2(\Memory[11] [52]), .ZN(n_0_2_1322));
   NAND3_X1 i_0_2_1375 (.A1(n_0_2_1320), .A2(n_0_2_1321), .A3(n_0_2_1322), 
      .ZN(n_0_2_1323));
   NOR2_X1 i_0_2_1376 (.A1(n_0_2_1319), .A2(n_0_2_1323), .ZN(n_0_2_1324));
   NAND3_X1 i_0_2_1377 (.A1(n_0_2_1305), .A2(n_0_2_1314), .A3(n_0_2_1324), 
      .ZN(dataOut1[52]));
   NAND2_X1 i_0_2_1378 (.A1(n_0_38), .A2(\Memory[4] [53]), .ZN(n_0_2_1325));
   NAND2_X1 i_0_2_1379 (.A1(n_0_41), .A2(\Memory[7] [53]), .ZN(n_0_2_1326));
   NAND2_X1 i_0_2_1380 (.A1(n_0_37), .A2(\Memory[3] [53]), .ZN(n_0_2_1327));
   NAND2_X1 i_0_2_1381 (.A1(n_0_36), .A2(\Memory[2] [53]), .ZN(n_0_2_1328));
   NAND4_X1 i_0_2_1382 (.A1(n_0_2_1325), .A2(n_0_2_1326), .A3(n_0_2_1327), 
      .A4(n_0_2_1328), .ZN(n_0_2_1329));
   INV_X1 i_0_2_1383 (.A(n_0_2_1329), .ZN(n_0_2_1330));
   NAND2_X1 i_0_2_1384 (.A1(n_0_50), .A2(\Memory[16] [53]), .ZN(n_0_2_1331));
   NAND2_X1 i_0_2_1385 (.A1(n_0_40), .A2(\Memory[6] [53]), .ZN(n_0_2_1332));
   NAND2_X1 i_0_2_1386 (.A1(n_0_39), .A2(\Memory[5] [53]), .ZN(n_0_2_1333));
   NAND3_X1 i_0_2_1387 (.A1(n_0_2_1331), .A2(n_0_2_1332), .A3(n_0_2_1333), 
      .ZN(n_0_2_1334));
   NAND2_X1 i_0_2_1388 (.A1(n_0_42), .A2(\Memory[8] [53]), .ZN(n_0_2_1335));
   NAND2_X1 i_0_2_1389 (.A1(n_0_35), .A2(\Memory[1] [53]), .ZN(n_0_2_1336));
   NAND2_X1 i_0_2_1390 (.A1(n_0_44), .A2(\Memory[10] [53]), .ZN(n_0_2_1337));
   NAND3_X1 i_0_2_1391 (.A1(n_0_2_1335), .A2(n_0_2_1336), .A3(n_0_2_1337), 
      .ZN(n_0_2_1338));
   NOR2_X1 i_0_2_1392 (.A1(n_0_2_1334), .A2(n_0_2_1338), .ZN(n_0_2_1339));
   NAND2_X1 i_0_2_1393 (.A1(n_0_48), .A2(\Memory[14] [53]), .ZN(n_0_2_1340));
   NAND2_X1 i_0_2_1394 (.A1(n_0_49), .A2(\Memory[15] [53]), .ZN(n_0_2_1341));
   NAND2_X1 i_0_2_1395 (.A1(n_0_34), .A2(\Memory[0] [53]), .ZN(n_0_2_1342));
   NAND2_X1 i_0_2_1396 (.A1(n_0_43), .A2(\Memory[9] [53]), .ZN(n_0_2_1343));
   NAND4_X1 i_0_2_1397 (.A1(n_0_2_1340), .A2(n_0_2_1341), .A3(n_0_2_1342), 
      .A4(n_0_2_1343), .ZN(n_0_2_1344));
   NAND2_X1 i_0_2_1398 (.A1(n_0_47), .A2(\Memory[13] [53]), .ZN(n_0_2_1345));
   NAND2_X1 i_0_2_1399 (.A1(n_0_46), .A2(\Memory[12] [53]), .ZN(n_0_2_1346));
   NAND2_X1 i_0_2_1400 (.A1(n_0_45), .A2(\Memory[11] [53]), .ZN(n_0_2_1347));
   NAND3_X1 i_0_2_1401 (.A1(n_0_2_1345), .A2(n_0_2_1346), .A3(n_0_2_1347), 
      .ZN(n_0_2_1348));
   NOR2_X1 i_0_2_1402 (.A1(n_0_2_1344), .A2(n_0_2_1348), .ZN(n_0_2_1349));
   NAND3_X1 i_0_2_1403 (.A1(n_0_2_1330), .A2(n_0_2_1339), .A3(n_0_2_1349), 
      .ZN(dataOut1[53]));
   NAND2_X1 i_0_2_1404 (.A1(n_0_38), .A2(\Memory[4] [54]), .ZN(n_0_2_1350));
   NAND2_X1 i_0_2_1405 (.A1(n_0_41), .A2(\Memory[7] [54]), .ZN(n_0_2_1351));
   NAND2_X1 i_0_2_1406 (.A1(n_0_37), .A2(\Memory[3] [54]), .ZN(n_0_2_1352));
   NAND2_X1 i_0_2_1407 (.A1(n_0_36), .A2(\Memory[2] [54]), .ZN(n_0_2_1353));
   NAND4_X1 i_0_2_1408 (.A1(n_0_2_1350), .A2(n_0_2_1351), .A3(n_0_2_1352), 
      .A4(n_0_2_1353), .ZN(n_0_2_1354));
   INV_X1 i_0_2_1409 (.A(n_0_2_1354), .ZN(n_0_2_1355));
   NAND2_X1 i_0_2_1410 (.A1(n_0_50), .A2(\Memory[16] [54]), .ZN(n_0_2_1356));
   NAND2_X1 i_0_2_1411 (.A1(n_0_40), .A2(\Memory[6] [54]), .ZN(n_0_2_1357));
   NAND2_X1 i_0_2_1412 (.A1(n_0_39), .A2(\Memory[5] [54]), .ZN(n_0_2_1358));
   NAND3_X1 i_0_2_1413 (.A1(n_0_2_1356), .A2(n_0_2_1357), .A3(n_0_2_1358), 
      .ZN(n_0_2_1359));
   NAND2_X1 i_0_2_1414 (.A1(n_0_42), .A2(\Memory[8] [54]), .ZN(n_0_2_1360));
   NAND2_X1 i_0_2_1415 (.A1(n_0_35), .A2(\Memory[1] [54]), .ZN(n_0_2_1361));
   NAND2_X1 i_0_2_1416 (.A1(n_0_44), .A2(\Memory[10] [54]), .ZN(n_0_2_1362));
   NAND3_X1 i_0_2_1417 (.A1(n_0_2_1360), .A2(n_0_2_1361), .A3(n_0_2_1362), 
      .ZN(n_0_2_1363));
   NOR2_X1 i_0_2_1418 (.A1(n_0_2_1359), .A2(n_0_2_1363), .ZN(n_0_2_1364));
   NAND2_X1 i_0_2_1419 (.A1(n_0_48), .A2(\Memory[14] [54]), .ZN(n_0_2_1365));
   NAND2_X1 i_0_2_1420 (.A1(n_0_49), .A2(\Memory[15] [54]), .ZN(n_0_2_1366));
   NAND2_X1 i_0_2_1421 (.A1(n_0_34), .A2(\Memory[0] [54]), .ZN(n_0_2_1367));
   NAND2_X1 i_0_2_1422 (.A1(n_0_43), .A2(\Memory[9] [54]), .ZN(n_0_2_1368));
   NAND4_X1 i_0_2_1423 (.A1(n_0_2_1365), .A2(n_0_2_1366), .A3(n_0_2_1367), 
      .A4(n_0_2_1368), .ZN(n_0_2_1369));
   NAND2_X1 i_0_2_1424 (.A1(n_0_47), .A2(\Memory[13] [54]), .ZN(n_0_2_1370));
   NAND2_X1 i_0_2_1425 (.A1(n_0_46), .A2(\Memory[12] [54]), .ZN(n_0_2_1371));
   NAND2_X1 i_0_2_1426 (.A1(n_0_45), .A2(\Memory[11] [54]), .ZN(n_0_2_1372));
   NAND3_X1 i_0_2_1427 (.A1(n_0_2_1370), .A2(n_0_2_1371), .A3(n_0_2_1372), 
      .ZN(n_0_2_1373));
   NOR2_X1 i_0_2_1428 (.A1(n_0_2_1369), .A2(n_0_2_1373), .ZN(n_0_2_1374));
   NAND3_X1 i_0_2_1429 (.A1(n_0_2_1355), .A2(n_0_2_1364), .A3(n_0_2_1374), 
      .ZN(dataOut1[54]));
   NAND2_X1 i_0_2_1430 (.A1(n_0_38), .A2(\Memory[4] [55]), .ZN(n_0_2_1375));
   NAND2_X1 i_0_2_1431 (.A1(n_0_41), .A2(\Memory[7] [55]), .ZN(n_0_2_1376));
   NAND2_X1 i_0_2_1432 (.A1(n_0_37), .A2(\Memory[3] [55]), .ZN(n_0_2_1377));
   NAND2_X1 i_0_2_1433 (.A1(n_0_36), .A2(\Memory[2] [55]), .ZN(n_0_2_1378));
   NAND4_X1 i_0_2_1434 (.A1(n_0_2_1375), .A2(n_0_2_1376), .A3(n_0_2_1377), 
      .A4(n_0_2_1378), .ZN(n_0_2_1379));
   INV_X1 i_0_2_1435 (.A(n_0_2_1379), .ZN(n_0_2_1380));
   NAND2_X1 i_0_2_1436 (.A1(n_0_50), .A2(\Memory[16] [55]), .ZN(n_0_2_1381));
   NAND2_X1 i_0_2_1437 (.A1(n_0_40), .A2(\Memory[6] [55]), .ZN(n_0_2_1382));
   NAND2_X1 i_0_2_1438 (.A1(n_0_39), .A2(\Memory[5] [55]), .ZN(n_0_2_1383));
   NAND3_X1 i_0_2_1439 (.A1(n_0_2_1381), .A2(n_0_2_1382), .A3(n_0_2_1383), 
      .ZN(n_0_2_1384));
   NAND2_X1 i_0_2_1440 (.A1(n_0_42), .A2(\Memory[8] [55]), .ZN(n_0_2_1385));
   NAND2_X1 i_0_2_1441 (.A1(n_0_35), .A2(\Memory[1] [55]), .ZN(n_0_2_1386));
   NAND2_X1 i_0_2_1442 (.A1(n_0_44), .A2(\Memory[10] [55]), .ZN(n_0_2_1387));
   NAND3_X1 i_0_2_1443 (.A1(n_0_2_1385), .A2(n_0_2_1386), .A3(n_0_2_1387), 
      .ZN(n_0_2_1388));
   NOR2_X1 i_0_2_1444 (.A1(n_0_2_1384), .A2(n_0_2_1388), .ZN(n_0_2_1389));
   NAND2_X1 i_0_2_1445 (.A1(n_0_48), .A2(\Memory[14] [55]), .ZN(n_0_2_1390));
   NAND2_X1 i_0_2_1446 (.A1(n_0_49), .A2(\Memory[15] [55]), .ZN(n_0_2_1391));
   NAND2_X1 i_0_2_1447 (.A1(n_0_34), .A2(\Memory[0] [55]), .ZN(n_0_2_1392));
   NAND2_X1 i_0_2_1448 (.A1(n_0_43), .A2(\Memory[9] [55]), .ZN(n_0_2_1393));
   NAND4_X1 i_0_2_1449 (.A1(n_0_2_1390), .A2(n_0_2_1391), .A3(n_0_2_1392), 
      .A4(n_0_2_1393), .ZN(n_0_2_1394));
   NAND2_X1 i_0_2_1450 (.A1(n_0_47), .A2(\Memory[13] [55]), .ZN(n_0_2_1395));
   NAND2_X1 i_0_2_1451 (.A1(n_0_46), .A2(\Memory[12] [55]), .ZN(n_0_2_1396));
   NAND2_X1 i_0_2_1452 (.A1(n_0_45), .A2(\Memory[11] [55]), .ZN(n_0_2_1397));
   NAND3_X1 i_0_2_1453 (.A1(n_0_2_1395), .A2(n_0_2_1396), .A3(n_0_2_1397), 
      .ZN(n_0_2_1398));
   NOR2_X1 i_0_2_1454 (.A1(n_0_2_1394), .A2(n_0_2_1398), .ZN(n_0_2_1399));
   NAND3_X1 i_0_2_1455 (.A1(n_0_2_1380), .A2(n_0_2_1389), .A3(n_0_2_1399), 
      .ZN(dataOut1[55]));
   NAND2_X1 i_0_2_1456 (.A1(n_0_38), .A2(\Memory[4] [56]), .ZN(n_0_2_1400));
   NAND2_X1 i_0_2_1457 (.A1(n_0_41), .A2(\Memory[7] [56]), .ZN(n_0_2_1401));
   NAND2_X1 i_0_2_1458 (.A1(n_0_37), .A2(\Memory[3] [56]), .ZN(n_0_2_1402));
   NAND2_X1 i_0_2_1459 (.A1(n_0_36), .A2(\Memory[2] [56]), .ZN(n_0_2_1403));
   NAND4_X1 i_0_2_1460 (.A1(n_0_2_1400), .A2(n_0_2_1401), .A3(n_0_2_1402), 
      .A4(n_0_2_1403), .ZN(n_0_2_1404));
   INV_X1 i_0_2_1461 (.A(n_0_2_1404), .ZN(n_0_2_1405));
   NAND2_X1 i_0_2_1462 (.A1(n_0_50), .A2(\Memory[16] [56]), .ZN(n_0_2_1406));
   NAND2_X1 i_0_2_1463 (.A1(n_0_40), .A2(\Memory[6] [56]), .ZN(n_0_2_1407));
   NAND2_X1 i_0_2_1464 (.A1(n_0_39), .A2(\Memory[5] [56]), .ZN(n_0_2_1408));
   NAND3_X1 i_0_2_1465 (.A1(n_0_2_1406), .A2(n_0_2_1407), .A3(n_0_2_1408), 
      .ZN(n_0_2_1409));
   NAND2_X1 i_0_2_1466 (.A1(n_0_42), .A2(\Memory[8] [56]), .ZN(n_0_2_1410));
   NAND2_X1 i_0_2_1467 (.A1(n_0_35), .A2(\Memory[1] [56]), .ZN(n_0_2_1411));
   NAND2_X1 i_0_2_1468 (.A1(n_0_44), .A2(\Memory[10] [56]), .ZN(n_0_2_1412));
   NAND3_X1 i_0_2_1469 (.A1(n_0_2_1410), .A2(n_0_2_1411), .A3(n_0_2_1412), 
      .ZN(n_0_2_1413));
   NOR2_X1 i_0_2_1470 (.A1(n_0_2_1409), .A2(n_0_2_1413), .ZN(n_0_2_1414));
   NAND2_X1 i_0_2_1471 (.A1(n_0_48), .A2(\Memory[14] [56]), .ZN(n_0_2_1415));
   NAND2_X1 i_0_2_1472 (.A1(n_0_49), .A2(\Memory[15] [56]), .ZN(n_0_2_1416));
   NAND2_X1 i_0_2_1473 (.A1(n_0_34), .A2(\Memory[0] [56]), .ZN(n_0_2_1417));
   NAND2_X1 i_0_2_1474 (.A1(n_0_43), .A2(\Memory[9] [56]), .ZN(n_0_2_1418));
   NAND4_X1 i_0_2_1475 (.A1(n_0_2_1415), .A2(n_0_2_1416), .A3(n_0_2_1417), 
      .A4(n_0_2_1418), .ZN(n_0_2_1419));
   NAND2_X1 i_0_2_1476 (.A1(n_0_47), .A2(\Memory[13] [56]), .ZN(n_0_2_1420));
   NAND2_X1 i_0_2_1477 (.A1(n_0_46), .A2(\Memory[12] [56]), .ZN(n_0_2_1421));
   NAND2_X1 i_0_2_1478 (.A1(n_0_45), .A2(\Memory[11] [56]), .ZN(n_0_2_1422));
   NAND3_X1 i_0_2_1479 (.A1(n_0_2_1420), .A2(n_0_2_1421), .A3(n_0_2_1422), 
      .ZN(n_0_2_1423));
   NOR2_X1 i_0_2_1480 (.A1(n_0_2_1419), .A2(n_0_2_1423), .ZN(n_0_2_1424));
   NAND3_X1 i_0_2_1481 (.A1(n_0_2_1405), .A2(n_0_2_1414), .A3(n_0_2_1424), 
      .ZN(dataOut1[56]));
   NAND2_X1 i_0_2_1482 (.A1(n_0_38), .A2(\Memory[4] [57]), .ZN(n_0_2_1425));
   NAND2_X1 i_0_2_1483 (.A1(n_0_41), .A2(\Memory[7] [57]), .ZN(n_0_2_1426));
   NAND2_X1 i_0_2_1484 (.A1(n_0_37), .A2(\Memory[3] [57]), .ZN(n_0_2_1427));
   NAND2_X1 i_0_2_1485 (.A1(n_0_36), .A2(\Memory[2] [57]), .ZN(n_0_2_1428));
   NAND4_X1 i_0_2_1486 (.A1(n_0_2_1425), .A2(n_0_2_1426), .A3(n_0_2_1427), 
      .A4(n_0_2_1428), .ZN(n_0_2_1429));
   INV_X1 i_0_2_1487 (.A(n_0_2_1429), .ZN(n_0_2_1430));
   NAND2_X1 i_0_2_1488 (.A1(n_0_50), .A2(\Memory[16] [57]), .ZN(n_0_2_1431));
   NAND2_X1 i_0_2_1489 (.A1(n_0_40), .A2(\Memory[6] [57]), .ZN(n_0_2_1432));
   NAND2_X1 i_0_2_1490 (.A1(n_0_39), .A2(\Memory[5] [57]), .ZN(n_0_2_1433));
   NAND3_X1 i_0_2_1491 (.A1(n_0_2_1431), .A2(n_0_2_1432), .A3(n_0_2_1433), 
      .ZN(n_0_2_1434));
   NAND2_X1 i_0_2_1492 (.A1(n_0_42), .A2(\Memory[8] [57]), .ZN(n_0_2_1435));
   NAND2_X1 i_0_2_1493 (.A1(n_0_35), .A2(\Memory[1] [57]), .ZN(n_0_2_1436));
   NAND2_X1 i_0_2_1494 (.A1(n_0_44), .A2(\Memory[10] [57]), .ZN(n_0_2_1437));
   NAND3_X1 i_0_2_1495 (.A1(n_0_2_1435), .A2(n_0_2_1436), .A3(n_0_2_1437), 
      .ZN(n_0_2_1438));
   NOR2_X1 i_0_2_1496 (.A1(n_0_2_1434), .A2(n_0_2_1438), .ZN(n_0_2_1439));
   NAND2_X1 i_0_2_1497 (.A1(n_0_48), .A2(\Memory[14] [57]), .ZN(n_0_2_1440));
   NAND2_X1 i_0_2_1498 (.A1(n_0_49), .A2(\Memory[15] [57]), .ZN(n_0_2_1441));
   NAND2_X1 i_0_2_1499 (.A1(n_0_34), .A2(\Memory[0] [57]), .ZN(n_0_2_1442));
   NAND2_X1 i_0_2_1500 (.A1(n_0_43), .A2(\Memory[9] [57]), .ZN(n_0_2_1443));
   NAND4_X1 i_0_2_1501 (.A1(n_0_2_1440), .A2(n_0_2_1441), .A3(n_0_2_1442), 
      .A4(n_0_2_1443), .ZN(n_0_2_1444));
   NAND2_X1 i_0_2_1502 (.A1(n_0_47), .A2(\Memory[13] [57]), .ZN(n_0_2_1445));
   NAND2_X1 i_0_2_1503 (.A1(n_0_46), .A2(\Memory[12] [57]), .ZN(n_0_2_1446));
   NAND2_X1 i_0_2_1504 (.A1(n_0_45), .A2(\Memory[11] [57]), .ZN(n_0_2_1447));
   NAND3_X1 i_0_2_1505 (.A1(n_0_2_1445), .A2(n_0_2_1446), .A3(n_0_2_1447), 
      .ZN(n_0_2_1448));
   NOR2_X1 i_0_2_1506 (.A1(n_0_2_1444), .A2(n_0_2_1448), .ZN(n_0_2_1449));
   NAND3_X1 i_0_2_1507 (.A1(n_0_2_1430), .A2(n_0_2_1439), .A3(n_0_2_1449), 
      .ZN(dataOut1[57]));
   NAND2_X1 i_0_2_1508 (.A1(n_0_38), .A2(\Memory[4] [58]), .ZN(n_0_2_1450));
   NAND2_X1 i_0_2_1509 (.A1(n_0_41), .A2(\Memory[7] [58]), .ZN(n_0_2_1451));
   NAND2_X1 i_0_2_1510 (.A1(n_0_37), .A2(\Memory[3] [58]), .ZN(n_0_2_1452));
   NAND2_X1 i_0_2_1511 (.A1(n_0_36), .A2(\Memory[2] [58]), .ZN(n_0_2_1453));
   NAND4_X1 i_0_2_1512 (.A1(n_0_2_1450), .A2(n_0_2_1451), .A3(n_0_2_1452), 
      .A4(n_0_2_1453), .ZN(n_0_2_1454));
   INV_X1 i_0_2_1513 (.A(n_0_2_1454), .ZN(n_0_2_1455));
   NAND2_X1 i_0_2_1514 (.A1(n_0_50), .A2(\Memory[16] [58]), .ZN(n_0_2_1456));
   NAND2_X1 i_0_2_1515 (.A1(n_0_40), .A2(\Memory[6] [58]), .ZN(n_0_2_1457));
   NAND2_X1 i_0_2_1516 (.A1(n_0_39), .A2(\Memory[5] [58]), .ZN(n_0_2_1458));
   NAND3_X1 i_0_2_1517 (.A1(n_0_2_1456), .A2(n_0_2_1457), .A3(n_0_2_1458), 
      .ZN(n_0_2_1459));
   NAND2_X1 i_0_2_1518 (.A1(n_0_42), .A2(\Memory[8] [58]), .ZN(n_0_2_1460));
   NAND2_X1 i_0_2_1519 (.A1(n_0_35), .A2(\Memory[1] [58]), .ZN(n_0_2_1461));
   NAND2_X1 i_0_2_1520 (.A1(n_0_44), .A2(\Memory[10] [58]), .ZN(n_0_2_1462));
   NAND3_X1 i_0_2_1521 (.A1(n_0_2_1460), .A2(n_0_2_1461), .A3(n_0_2_1462), 
      .ZN(n_0_2_1463));
   NOR2_X1 i_0_2_1522 (.A1(n_0_2_1459), .A2(n_0_2_1463), .ZN(n_0_2_1464));
   NAND2_X1 i_0_2_1523 (.A1(n_0_48), .A2(\Memory[14] [58]), .ZN(n_0_2_1465));
   NAND2_X1 i_0_2_1524 (.A1(n_0_49), .A2(\Memory[15] [58]), .ZN(n_0_2_1466));
   NAND2_X1 i_0_2_1525 (.A1(n_0_34), .A2(\Memory[0] [58]), .ZN(n_0_2_1467));
   NAND2_X1 i_0_2_1526 (.A1(n_0_43), .A2(\Memory[9] [58]), .ZN(n_0_2_1468));
   NAND4_X1 i_0_2_1527 (.A1(n_0_2_1465), .A2(n_0_2_1466), .A3(n_0_2_1467), 
      .A4(n_0_2_1468), .ZN(n_0_2_1469));
   NAND2_X1 i_0_2_1528 (.A1(n_0_47), .A2(\Memory[13] [58]), .ZN(n_0_2_1470));
   NAND2_X1 i_0_2_1529 (.A1(n_0_46), .A2(\Memory[12] [58]), .ZN(n_0_2_1471));
   NAND2_X1 i_0_2_1530 (.A1(n_0_45), .A2(\Memory[11] [58]), .ZN(n_0_2_1472));
   NAND3_X1 i_0_2_1531 (.A1(n_0_2_1470), .A2(n_0_2_1471), .A3(n_0_2_1472), 
      .ZN(n_0_2_1473));
   NOR2_X1 i_0_2_1532 (.A1(n_0_2_1469), .A2(n_0_2_1473), .ZN(n_0_2_1474));
   NAND3_X1 i_0_2_1533 (.A1(n_0_2_1455), .A2(n_0_2_1464), .A3(n_0_2_1474), 
      .ZN(dataOut1[58]));
   NAND2_X1 i_0_2_1534 (.A1(n_0_38), .A2(\Memory[4] [59]), .ZN(n_0_2_1475));
   NAND2_X1 i_0_2_1535 (.A1(n_0_41), .A2(\Memory[7] [59]), .ZN(n_0_2_1476));
   NAND2_X1 i_0_2_1536 (.A1(n_0_37), .A2(\Memory[3] [59]), .ZN(n_0_2_1477));
   NAND2_X1 i_0_2_1537 (.A1(n_0_36), .A2(\Memory[2] [59]), .ZN(n_0_2_1478));
   NAND4_X1 i_0_2_1538 (.A1(n_0_2_1475), .A2(n_0_2_1476), .A3(n_0_2_1477), 
      .A4(n_0_2_1478), .ZN(n_0_2_1479));
   INV_X1 i_0_2_1539 (.A(n_0_2_1479), .ZN(n_0_2_1480));
   NAND2_X1 i_0_2_1540 (.A1(n_0_50), .A2(\Memory[16] [59]), .ZN(n_0_2_1481));
   NAND2_X1 i_0_2_1541 (.A1(n_0_40), .A2(\Memory[6] [59]), .ZN(n_0_2_1482));
   NAND2_X1 i_0_2_1542 (.A1(n_0_39), .A2(\Memory[5] [59]), .ZN(n_0_2_1483));
   NAND3_X1 i_0_2_1543 (.A1(n_0_2_1481), .A2(n_0_2_1482), .A3(n_0_2_1483), 
      .ZN(n_0_2_1484));
   NAND2_X1 i_0_2_1544 (.A1(n_0_42), .A2(\Memory[8] [59]), .ZN(n_0_2_1485));
   NAND2_X1 i_0_2_1545 (.A1(n_0_35), .A2(\Memory[1] [59]), .ZN(n_0_2_1486));
   NAND2_X1 i_0_2_1546 (.A1(n_0_44), .A2(\Memory[10] [59]), .ZN(n_0_2_1487));
   NAND3_X1 i_0_2_1547 (.A1(n_0_2_1485), .A2(n_0_2_1486), .A3(n_0_2_1487), 
      .ZN(n_0_2_1488));
   NOR2_X1 i_0_2_1548 (.A1(n_0_2_1484), .A2(n_0_2_1488), .ZN(n_0_2_1489));
   NAND2_X1 i_0_2_1549 (.A1(n_0_48), .A2(\Memory[14] [59]), .ZN(n_0_2_1490));
   NAND2_X1 i_0_2_1550 (.A1(n_0_49), .A2(\Memory[15] [59]), .ZN(n_0_2_1491));
   NAND2_X1 i_0_2_1551 (.A1(n_0_34), .A2(\Memory[0] [59]), .ZN(n_0_2_1492));
   NAND2_X1 i_0_2_1552 (.A1(n_0_43), .A2(\Memory[9] [59]), .ZN(n_0_2_1493));
   NAND4_X1 i_0_2_1553 (.A1(n_0_2_1490), .A2(n_0_2_1491), .A3(n_0_2_1492), 
      .A4(n_0_2_1493), .ZN(n_0_2_1494));
   NAND2_X1 i_0_2_1554 (.A1(n_0_47), .A2(\Memory[13] [59]), .ZN(n_0_2_1495));
   NAND2_X1 i_0_2_1555 (.A1(n_0_46), .A2(\Memory[12] [59]), .ZN(n_0_2_1496));
   NAND2_X1 i_0_2_1556 (.A1(n_0_45), .A2(\Memory[11] [59]), .ZN(n_0_2_1497));
   NAND3_X1 i_0_2_1557 (.A1(n_0_2_1495), .A2(n_0_2_1496), .A3(n_0_2_1497), 
      .ZN(n_0_2_1498));
   NOR2_X1 i_0_2_1558 (.A1(n_0_2_1494), .A2(n_0_2_1498), .ZN(n_0_2_1499));
   NAND3_X1 i_0_2_1559 (.A1(n_0_2_1480), .A2(n_0_2_1489), .A3(n_0_2_1499), 
      .ZN(dataOut1[59]));
   NAND2_X1 i_0_2_1560 (.A1(n_0_38), .A2(\Memory[4] [60]), .ZN(n_0_2_1500));
   NAND2_X1 i_0_2_1561 (.A1(n_0_41), .A2(\Memory[7] [60]), .ZN(n_0_2_1501));
   NAND2_X1 i_0_2_1562 (.A1(n_0_37), .A2(\Memory[3] [60]), .ZN(n_0_2_1502));
   NAND2_X1 i_0_2_1563 (.A1(n_0_36), .A2(\Memory[2] [60]), .ZN(n_0_2_1503));
   NAND4_X1 i_0_2_1564 (.A1(n_0_2_1500), .A2(n_0_2_1501), .A3(n_0_2_1502), 
      .A4(n_0_2_1503), .ZN(n_0_2_1504));
   INV_X1 i_0_2_1565 (.A(n_0_2_1504), .ZN(n_0_2_1505));
   NAND2_X1 i_0_2_1566 (.A1(n_0_50), .A2(\Memory[16] [60]), .ZN(n_0_2_1506));
   NAND2_X1 i_0_2_1567 (.A1(n_0_40), .A2(\Memory[6] [60]), .ZN(n_0_2_1507));
   NAND2_X1 i_0_2_1568 (.A1(n_0_39), .A2(\Memory[5] [60]), .ZN(n_0_2_1508));
   NAND3_X1 i_0_2_1569 (.A1(n_0_2_1506), .A2(n_0_2_1507), .A3(n_0_2_1508), 
      .ZN(n_0_2_1509));
   NAND2_X1 i_0_2_1570 (.A1(n_0_42), .A2(\Memory[8] [60]), .ZN(n_0_2_1510));
   NAND2_X1 i_0_2_1571 (.A1(n_0_35), .A2(\Memory[1] [60]), .ZN(n_0_2_1511));
   NAND2_X1 i_0_2_1572 (.A1(n_0_44), .A2(\Memory[10] [60]), .ZN(n_0_2_1512));
   NAND3_X1 i_0_2_1573 (.A1(n_0_2_1510), .A2(n_0_2_1511), .A3(n_0_2_1512), 
      .ZN(n_0_2_1513));
   NOR2_X1 i_0_2_1574 (.A1(n_0_2_1509), .A2(n_0_2_1513), .ZN(n_0_2_1514));
   NAND2_X1 i_0_2_1575 (.A1(n_0_48), .A2(\Memory[14] [60]), .ZN(n_0_2_1515));
   NAND2_X1 i_0_2_1576 (.A1(n_0_49), .A2(\Memory[15] [60]), .ZN(n_0_2_1516));
   NAND2_X1 i_0_2_1577 (.A1(n_0_34), .A2(\Memory[0] [60]), .ZN(n_0_2_1517));
   NAND2_X1 i_0_2_1578 (.A1(n_0_43), .A2(\Memory[9] [60]), .ZN(n_0_2_1518));
   NAND4_X1 i_0_2_1579 (.A1(n_0_2_1515), .A2(n_0_2_1516), .A3(n_0_2_1517), 
      .A4(n_0_2_1518), .ZN(n_0_2_1519));
   NAND2_X1 i_0_2_1580 (.A1(n_0_47), .A2(\Memory[13] [60]), .ZN(n_0_2_1520));
   NAND2_X1 i_0_2_1581 (.A1(n_0_46), .A2(\Memory[12] [60]), .ZN(n_0_2_1521));
   NAND2_X1 i_0_2_1582 (.A1(n_0_45), .A2(\Memory[11] [60]), .ZN(n_0_2_1522));
   NAND3_X1 i_0_2_1583 (.A1(n_0_2_1520), .A2(n_0_2_1521), .A3(n_0_2_1522), 
      .ZN(n_0_2_1523));
   NOR2_X1 i_0_2_1584 (.A1(n_0_2_1519), .A2(n_0_2_1523), .ZN(n_0_2_1524));
   NAND3_X1 i_0_2_1585 (.A1(n_0_2_1505), .A2(n_0_2_1514), .A3(n_0_2_1524), 
      .ZN(dataOut1[60]));
   NAND2_X1 i_0_2_1586 (.A1(n_0_38), .A2(\Memory[4] [61]), .ZN(n_0_2_1525));
   NAND2_X1 i_0_2_1587 (.A1(n_0_41), .A2(\Memory[7] [61]), .ZN(n_0_2_1526));
   NAND2_X1 i_0_2_1588 (.A1(n_0_37), .A2(\Memory[3] [61]), .ZN(n_0_2_1527));
   NAND2_X1 i_0_2_1589 (.A1(n_0_36), .A2(\Memory[2] [61]), .ZN(n_0_2_1528));
   NAND4_X1 i_0_2_1590 (.A1(n_0_2_1525), .A2(n_0_2_1526), .A3(n_0_2_1527), 
      .A4(n_0_2_1528), .ZN(n_0_2_1529));
   INV_X1 i_0_2_1591 (.A(n_0_2_1529), .ZN(n_0_2_1530));
   NAND2_X1 i_0_2_1592 (.A1(n_0_50), .A2(\Memory[16] [61]), .ZN(n_0_2_1531));
   NAND2_X1 i_0_2_1593 (.A1(n_0_40), .A2(\Memory[6] [61]), .ZN(n_0_2_1532));
   NAND2_X1 i_0_2_1594 (.A1(n_0_39), .A2(\Memory[5] [61]), .ZN(n_0_2_1533));
   NAND3_X1 i_0_2_1595 (.A1(n_0_2_1531), .A2(n_0_2_1532), .A3(n_0_2_1533), 
      .ZN(n_0_2_1534));
   NAND2_X1 i_0_2_1596 (.A1(n_0_42), .A2(\Memory[8] [61]), .ZN(n_0_2_1535));
   NAND2_X1 i_0_2_1597 (.A1(n_0_35), .A2(\Memory[1] [61]), .ZN(n_0_2_1536));
   NAND2_X1 i_0_2_1598 (.A1(n_0_44), .A2(\Memory[10] [61]), .ZN(n_0_2_1537));
   NAND3_X1 i_0_2_1599 (.A1(n_0_2_1535), .A2(n_0_2_1536), .A3(n_0_2_1537), 
      .ZN(n_0_2_1538));
   NOR2_X1 i_0_2_1600 (.A1(n_0_2_1534), .A2(n_0_2_1538), .ZN(n_0_2_1539));
   NAND2_X1 i_0_2_1601 (.A1(n_0_48), .A2(\Memory[14] [61]), .ZN(n_0_2_1540));
   NAND2_X1 i_0_2_1602 (.A1(n_0_49), .A2(\Memory[15] [61]), .ZN(n_0_2_1541));
   NAND2_X1 i_0_2_1603 (.A1(n_0_34), .A2(\Memory[0] [61]), .ZN(n_0_2_1542));
   NAND2_X1 i_0_2_1604 (.A1(n_0_43), .A2(\Memory[9] [61]), .ZN(n_0_2_1543));
   NAND4_X1 i_0_2_1605 (.A1(n_0_2_1540), .A2(n_0_2_1541), .A3(n_0_2_1542), 
      .A4(n_0_2_1543), .ZN(n_0_2_1544));
   NAND2_X1 i_0_2_1606 (.A1(n_0_47), .A2(\Memory[13] [61]), .ZN(n_0_2_1545));
   NAND2_X1 i_0_2_1607 (.A1(n_0_46), .A2(\Memory[12] [61]), .ZN(n_0_2_1546));
   NAND2_X1 i_0_2_1608 (.A1(n_0_45), .A2(\Memory[11] [61]), .ZN(n_0_2_1547));
   NAND3_X1 i_0_2_1609 (.A1(n_0_2_1545), .A2(n_0_2_1546), .A3(n_0_2_1547), 
      .ZN(n_0_2_1548));
   NOR2_X1 i_0_2_1610 (.A1(n_0_2_1544), .A2(n_0_2_1548), .ZN(n_0_2_1549));
   NAND3_X1 i_0_2_1611 (.A1(n_0_2_1530), .A2(n_0_2_1539), .A3(n_0_2_1549), 
      .ZN(dataOut1[61]));
   NAND2_X1 i_0_2_1612 (.A1(n_0_38), .A2(\Memory[4] [62]), .ZN(n_0_2_1550));
   NAND2_X1 i_0_2_1613 (.A1(n_0_41), .A2(\Memory[7] [62]), .ZN(n_0_2_1551));
   NAND2_X1 i_0_2_1614 (.A1(n_0_37), .A2(\Memory[3] [62]), .ZN(n_0_2_1552));
   NAND2_X1 i_0_2_1615 (.A1(n_0_36), .A2(\Memory[2] [62]), .ZN(n_0_2_1553));
   NAND4_X1 i_0_2_1616 (.A1(n_0_2_1550), .A2(n_0_2_1551), .A3(n_0_2_1552), 
      .A4(n_0_2_1553), .ZN(n_0_2_1554));
   INV_X1 i_0_2_1617 (.A(n_0_2_1554), .ZN(n_0_2_1555));
   NAND2_X1 i_0_2_1618 (.A1(n_0_50), .A2(\Memory[16] [62]), .ZN(n_0_2_1556));
   NAND2_X1 i_0_2_1619 (.A1(n_0_40), .A2(\Memory[6] [62]), .ZN(n_0_2_1557));
   NAND2_X1 i_0_2_1620 (.A1(n_0_39), .A2(\Memory[5] [62]), .ZN(n_0_2_1558));
   NAND3_X1 i_0_2_1621 (.A1(n_0_2_1556), .A2(n_0_2_1557), .A3(n_0_2_1558), 
      .ZN(n_0_2_1559));
   NAND2_X1 i_0_2_1622 (.A1(n_0_42), .A2(\Memory[8] [62]), .ZN(n_0_2_1560));
   NAND2_X1 i_0_2_1623 (.A1(n_0_35), .A2(\Memory[1] [62]), .ZN(n_0_2_1561));
   NAND2_X1 i_0_2_1624 (.A1(n_0_44), .A2(\Memory[10] [62]), .ZN(n_0_2_1562));
   NAND3_X1 i_0_2_1625 (.A1(n_0_2_1560), .A2(n_0_2_1561), .A3(n_0_2_1562), 
      .ZN(n_0_2_1563));
   NOR2_X1 i_0_2_1626 (.A1(n_0_2_1559), .A2(n_0_2_1563), .ZN(n_0_2_1564));
   NAND2_X1 i_0_2_1627 (.A1(n_0_48), .A2(\Memory[14] [62]), .ZN(n_0_2_1565));
   NAND2_X1 i_0_2_1628 (.A1(n_0_49), .A2(\Memory[15] [62]), .ZN(n_0_2_1566));
   NAND2_X1 i_0_2_1629 (.A1(n_0_34), .A2(\Memory[0] [62]), .ZN(n_0_2_1567));
   NAND2_X1 i_0_2_1630 (.A1(n_0_43), .A2(\Memory[9] [62]), .ZN(n_0_2_1568));
   NAND4_X1 i_0_2_1631 (.A1(n_0_2_1565), .A2(n_0_2_1566), .A3(n_0_2_1567), 
      .A4(n_0_2_1568), .ZN(n_0_2_1569));
   NAND2_X1 i_0_2_1632 (.A1(n_0_47), .A2(\Memory[13] [62]), .ZN(n_0_2_1570));
   NAND2_X1 i_0_2_1633 (.A1(n_0_46), .A2(\Memory[12] [62]), .ZN(n_0_2_1571));
   NAND2_X1 i_0_2_1634 (.A1(n_0_45), .A2(\Memory[11] [62]), .ZN(n_0_2_1572));
   NAND3_X1 i_0_2_1635 (.A1(n_0_2_1570), .A2(n_0_2_1571), .A3(n_0_2_1572), 
      .ZN(n_0_2_1573));
   NOR2_X1 i_0_2_1636 (.A1(n_0_2_1569), .A2(n_0_2_1573), .ZN(n_0_2_1574));
   NAND3_X1 i_0_2_1637 (.A1(n_0_2_1555), .A2(n_0_2_1564), .A3(n_0_2_1574), 
      .ZN(dataOut1[62]));
   NAND2_X1 i_0_2_1638 (.A1(n_0_38), .A2(\Memory[4] [63]), .ZN(n_0_2_1575));
   NAND2_X1 i_0_2_1639 (.A1(n_0_41), .A2(\Memory[7] [63]), .ZN(n_0_2_1576));
   NAND2_X1 i_0_2_1640 (.A1(n_0_37), .A2(\Memory[3] [63]), .ZN(n_0_2_1577));
   NAND2_X1 i_0_2_1641 (.A1(n_0_36), .A2(\Memory[2] [63]), .ZN(n_0_2_1578));
   NAND4_X1 i_0_2_1642 (.A1(n_0_2_1575), .A2(n_0_2_1576), .A3(n_0_2_1577), 
      .A4(n_0_2_1578), .ZN(n_0_2_1579));
   INV_X1 i_0_2_1643 (.A(n_0_2_1579), .ZN(n_0_2_1580));
   NAND2_X1 i_0_2_1644 (.A1(n_0_50), .A2(\Memory[16] [63]), .ZN(n_0_2_1581));
   NAND2_X1 i_0_2_1645 (.A1(n_0_40), .A2(\Memory[6] [63]), .ZN(n_0_2_1582));
   NAND2_X1 i_0_2_1646 (.A1(n_0_39), .A2(\Memory[5] [63]), .ZN(n_0_2_1583));
   NAND3_X1 i_0_2_1647 (.A1(n_0_2_1581), .A2(n_0_2_1582), .A3(n_0_2_1583), 
      .ZN(n_0_2_1584));
   NAND2_X1 i_0_2_1648 (.A1(n_0_42), .A2(\Memory[8] [63]), .ZN(n_0_2_1585));
   NAND2_X1 i_0_2_1649 (.A1(n_0_35), .A2(\Memory[1] [63]), .ZN(n_0_2_1586));
   NAND2_X1 i_0_2_1650 (.A1(n_0_44), .A2(\Memory[10] [63]), .ZN(n_0_2_1587));
   NAND3_X1 i_0_2_1651 (.A1(n_0_2_1585), .A2(n_0_2_1586), .A3(n_0_2_1587), 
      .ZN(n_0_2_1588));
   NOR2_X1 i_0_2_1652 (.A1(n_0_2_1584), .A2(n_0_2_1588), .ZN(n_0_2_1589));
   NAND2_X1 i_0_2_1653 (.A1(n_0_48), .A2(\Memory[14] [63]), .ZN(n_0_2_1590));
   NAND2_X1 i_0_2_1654 (.A1(n_0_49), .A2(\Memory[15] [63]), .ZN(n_0_2_1591));
   NAND2_X1 i_0_2_1655 (.A1(n_0_34), .A2(\Memory[0] [63]), .ZN(n_0_2_1592));
   NAND2_X1 i_0_2_1656 (.A1(n_0_43), .A2(\Memory[9] [63]), .ZN(n_0_2_1593));
   NAND4_X1 i_0_2_1657 (.A1(n_0_2_1590), .A2(n_0_2_1591), .A3(n_0_2_1592), 
      .A4(n_0_2_1593), .ZN(n_0_2_1594));
   NAND2_X1 i_0_2_1658 (.A1(n_0_47), .A2(\Memory[13] [63]), .ZN(n_0_2_1595));
   NAND2_X1 i_0_2_1659 (.A1(n_0_46), .A2(\Memory[12] [63]), .ZN(n_0_2_1596));
   NAND2_X1 i_0_2_1660 (.A1(n_0_45), .A2(\Memory[11] [63]), .ZN(n_0_2_1597));
   NAND3_X1 i_0_2_1661 (.A1(n_0_2_1595), .A2(n_0_2_1596), .A3(n_0_2_1597), 
      .ZN(n_0_2_1598));
   NOR2_X1 i_0_2_1662 (.A1(n_0_2_1594), .A2(n_0_2_1598), .ZN(n_0_2_1599));
   NAND3_X1 i_0_2_1663 (.A1(n_0_2_1580), .A2(n_0_2_1589), .A3(n_0_2_1599), 
      .ZN(dataOut1[63]));
   INV_X1 i_0_3_0 (.A(n_0_3_0), .ZN(n_0_51));
   NAND3_X1 i_0_3_1 (.A1(n_0_3_12), .A2(n_0_3_8), .A3(n_0_3_22), .ZN(n_0_3_0));
   INV_X1 i_0_3_2 (.A(n_0_3_1), .ZN(n_0_52));
   NAND3_X1 i_0_3_3 (.A1(n_0_3_12), .A2(n_0_3_8), .A3(address_RD2[0]), .ZN(
      n_0_3_1));
   INV_X1 i_0_3_4 (.A(n_0_3_2), .ZN(n_0_53));
   NAND4_X1 i_0_3_5 (.A1(n_0_3_8), .A2(n_0_3_26), .A3(address_RD2[1]), .A4(
      n_0_3_22), .ZN(n_0_3_2));
   INV_X1 i_0_3_6 (.A(n_0_3_3), .ZN(n_0_54));
   NAND4_X1 i_0_3_7 (.A1(n_0_3_8), .A2(n_0_3_26), .A3(address_RD2[1]), .A4(
      address_RD2[0]), .ZN(n_0_3_3));
   INV_X1 i_0_3_8 (.A(n_0_3_4), .ZN(n_0_55));
   NAND4_X1 i_0_3_9 (.A1(n_0_3_8), .A2(address_RD2[2]), .A3(n_0_3_25), .A4(
      n_0_3_22), .ZN(n_0_3_4));
   INV_X1 i_0_3_10 (.A(n_0_3_5), .ZN(n_0_56));
   NAND4_X1 i_0_3_11 (.A1(n_0_3_8), .A2(address_RD2[2]), .A3(n_0_3_25), .A4(
      address_RD2[0]), .ZN(n_0_3_5));
   INV_X1 i_0_3_12 (.A(n_0_3_6), .ZN(n_0_57));
   NAND4_X1 i_0_3_13 (.A1(n_0_3_8), .A2(address_RD2[2]), .A3(address_RD2[1]), 
      .A4(n_0_3_22), .ZN(n_0_3_6));
   INV_X1 i_0_3_14 (.A(n_0_3_7), .ZN(n_0_58));
   NAND4_X1 i_0_3_15 (.A1(n_0_3_8), .A2(address_RD2[2]), .A3(address_RD2[1]), 
      .A4(address_RD2[0]), .ZN(n_0_3_7));
   INV_X1 i_0_3_16 (.A(n_0_3_9), .ZN(n_0_3_8));
   NAND2_X1 i_0_3_17 (.A1(n_0_3_20), .A2(n_0_3_23), .ZN(n_0_3_9));
   INV_X1 i_0_3_18 (.A(n_0_3_10), .ZN(n_0_59));
   NAND3_X1 i_0_3_19 (.A1(n_0_3_12), .A2(n_0_3_17), .A3(n_0_3_22), .ZN(n_0_3_10));
   INV_X1 i_0_3_20 (.A(n_0_3_11), .ZN(n_0_60));
   NAND3_X1 i_0_3_21 (.A1(n_0_3_12), .A2(n_0_3_17), .A3(address_RD2[0]), 
      .ZN(n_0_3_11));
   INV_X1 i_0_3_22 (.A(n_0_3_24), .ZN(n_0_3_12));
   INV_X1 i_0_3_23 (.A(n_0_3_13), .ZN(n_0_61));
   NAND4_X1 i_0_3_24 (.A1(n_0_3_17), .A2(n_0_3_26), .A3(address_RD2[1]), 
      .A4(n_0_3_22), .ZN(n_0_3_13));
   INV_X1 i_0_3_25 (.A(n_0_3_14), .ZN(n_0_62));
   NAND4_X1 i_0_3_26 (.A1(n_0_3_17), .A2(n_0_3_26), .A3(address_RD2[1]), 
      .A4(address_RD2[0]), .ZN(n_0_3_14));
   INV_X1 i_0_3_27 (.A(n_0_3_15), .ZN(n_0_63));
   NAND4_X1 i_0_3_28 (.A1(n_0_3_17), .A2(address_RD2[2]), .A3(n_0_3_25), 
      .A4(n_0_3_22), .ZN(n_0_3_15));
   INV_X1 i_0_3_29 (.A(n_0_3_16), .ZN(n_0_64));
   NAND4_X1 i_0_3_30 (.A1(n_0_3_17), .A2(address_RD2[2]), .A3(n_0_3_25), 
      .A4(address_RD2[0]), .ZN(n_0_3_16));
   INV_X1 i_0_3_31 (.A(n_0_3_18), .ZN(n_0_3_17));
   NAND2_X1 i_0_3_32 (.A1(n_0_3_20), .A2(address_RD2[3]), .ZN(n_0_3_18));
   NOR2_X1 i_0_3_33 (.A1(n_0_3_19), .A2(address_RD2[0]), .ZN(n_0_65));
   NOR2_X1 i_0_3_34 (.A1(n_0_3_19), .A2(n_0_3_22), .ZN(n_0_66));
   NAND4_X1 i_0_3_35 (.A1(n_0_3_20), .A2(address_RD2[3]), .A3(address_RD2[2]), 
      .A4(address_RD2[1]), .ZN(n_0_3_19));
   INV_X1 i_0_3_36 (.A(address_RD2[4]), .ZN(n_0_3_20));
   NOR2_X1 i_0_3_37 (.A1(n_0_3_21), .A2(n_0_3_24), .ZN(n_0_67));
   NAND3_X1 i_0_3_38 (.A1(n_0_3_23), .A2(n_0_3_22), .A3(address_RD2[4]), 
      .ZN(n_0_3_21));
   INV_X1 i_0_3_39 (.A(address_RD2[0]), .ZN(n_0_3_22));
   INV_X1 i_0_3_40 (.A(address_RD2[3]), .ZN(n_0_3_23));
   NAND2_X1 i_0_3_41 (.A1(n_0_3_26), .A2(n_0_3_25), .ZN(n_0_3_24));
   INV_X1 i_0_3_42 (.A(address_RD2[1]), .ZN(n_0_3_25));
   INV_X1 i_0_3_43 (.A(address_RD2[2]), .ZN(n_0_3_26));
   NAND2_X1 i_0_4_0 (.A1(n_0_55), .A2(\Memory[4] [0]), .ZN(n_0_4_0));
   NAND2_X1 i_0_4_1 (.A1(n_0_58), .A2(\Memory[7] [0]), .ZN(n_0_4_1));
   NAND2_X1 i_0_4_2 (.A1(n_0_54), .A2(\Memory[3] [0]), .ZN(n_0_4_2));
   NAND2_X1 i_0_4_3 (.A1(n_0_53), .A2(\Memory[2] [0]), .ZN(n_0_4_3));
   NAND4_X1 i_0_4_4 (.A1(n_0_4_0), .A2(n_0_4_1), .A3(n_0_4_2), .A4(n_0_4_3), 
      .ZN(n_0_4_4));
   INV_X1 i_0_4_5 (.A(n_0_4_4), .ZN(n_0_4_5));
   NAND2_X1 i_0_4_6 (.A1(n_0_67), .A2(\Memory[16] [0]), .ZN(n_0_4_6));
   NAND2_X1 i_0_4_7 (.A1(n_0_57), .A2(\Memory[6] [0]), .ZN(n_0_4_7));
   NAND2_X1 i_0_4_8 (.A1(n_0_56), .A2(\Memory[5] [0]), .ZN(n_0_4_8));
   NAND3_X1 i_0_4_9 (.A1(n_0_4_6), .A2(n_0_4_7), .A3(n_0_4_8), .ZN(n_0_4_9));
   NAND2_X1 i_0_4_10 (.A1(n_0_59), .A2(\Memory[8] [0]), .ZN(n_0_4_10));
   NAND2_X1 i_0_4_11 (.A1(n_0_52), .A2(\Memory[1] [0]), .ZN(n_0_4_11));
   NAND2_X1 i_0_4_12 (.A1(n_0_61), .A2(\Memory[10] [0]), .ZN(n_0_4_12));
   NAND3_X1 i_0_4_13 (.A1(n_0_4_10), .A2(n_0_4_11), .A3(n_0_4_12), .ZN(n_0_4_13));
   NOR2_X1 i_0_4_14 (.A1(n_0_4_9), .A2(n_0_4_13), .ZN(n_0_4_14));
   NAND2_X1 i_0_4_15 (.A1(n_0_65), .A2(\Memory[14] [0]), .ZN(n_0_4_15));
   NAND2_X1 i_0_4_16 (.A1(n_0_66), .A2(\Memory[15] [0]), .ZN(n_0_4_16));
   NAND2_X1 i_0_4_17 (.A1(n_0_51), .A2(\Memory[0] [0]), .ZN(n_0_4_17));
   NAND2_X1 i_0_4_18 (.A1(n_0_60), .A2(\Memory[9] [0]), .ZN(n_0_4_18));
   NAND4_X1 i_0_4_19 (.A1(n_0_4_15), .A2(n_0_4_16), .A3(n_0_4_17), .A4(n_0_4_18), 
      .ZN(n_0_4_19));
   NAND2_X1 i_0_4_20 (.A1(n_0_64), .A2(\Memory[13] [0]), .ZN(n_0_4_20));
   NAND2_X1 i_0_4_21 (.A1(n_0_63), .A2(\Memory[12] [0]), .ZN(n_0_4_21));
   NAND2_X1 i_0_4_22 (.A1(n_0_62), .A2(\Memory[11] [0]), .ZN(n_0_4_22));
   NAND3_X1 i_0_4_23 (.A1(n_0_4_20), .A2(n_0_4_21), .A3(n_0_4_22), .ZN(n_0_4_23));
   NOR2_X1 i_0_4_24 (.A1(n_0_4_19), .A2(n_0_4_23), .ZN(n_0_4_24));
   NAND3_X1 i_0_4_25 (.A1(n_0_4_5), .A2(n_0_4_14), .A3(n_0_4_24), .ZN(
      dataOut2[0]));
   NAND2_X1 i_0_4_26 (.A1(n_0_55), .A2(\Memory[4] [1]), .ZN(n_0_4_25));
   NAND2_X1 i_0_4_27 (.A1(n_0_58), .A2(\Memory[7] [1]), .ZN(n_0_4_26));
   NAND2_X1 i_0_4_28 (.A1(n_0_54), .A2(\Memory[3] [1]), .ZN(n_0_4_27));
   NAND2_X1 i_0_4_29 (.A1(n_0_53), .A2(\Memory[2] [1]), .ZN(n_0_4_28));
   NAND4_X1 i_0_4_30 (.A1(n_0_4_25), .A2(n_0_4_26), .A3(n_0_4_27), .A4(n_0_4_28), 
      .ZN(n_0_4_29));
   INV_X1 i_0_4_31 (.A(n_0_4_29), .ZN(n_0_4_30));
   NAND2_X1 i_0_4_32 (.A1(n_0_67), .A2(\Memory[16] [1]), .ZN(n_0_4_31));
   NAND2_X1 i_0_4_33 (.A1(n_0_57), .A2(\Memory[6] [1]), .ZN(n_0_4_32));
   NAND2_X1 i_0_4_34 (.A1(n_0_56), .A2(\Memory[5] [1]), .ZN(n_0_4_33));
   NAND3_X1 i_0_4_35 (.A1(n_0_4_31), .A2(n_0_4_32), .A3(n_0_4_33), .ZN(n_0_4_34));
   NAND2_X1 i_0_4_36 (.A1(n_0_59), .A2(\Memory[8] [1]), .ZN(n_0_4_35));
   NAND2_X1 i_0_4_37 (.A1(n_0_52), .A2(\Memory[1] [1]), .ZN(n_0_4_36));
   NAND2_X1 i_0_4_38 (.A1(n_0_61), .A2(\Memory[10] [1]), .ZN(n_0_4_37));
   NAND3_X1 i_0_4_39 (.A1(n_0_4_35), .A2(n_0_4_36), .A3(n_0_4_37), .ZN(n_0_4_38));
   NOR2_X1 i_0_4_40 (.A1(n_0_4_34), .A2(n_0_4_38), .ZN(n_0_4_39));
   NAND2_X1 i_0_4_41 (.A1(n_0_65), .A2(\Memory[14] [1]), .ZN(n_0_4_40));
   NAND2_X1 i_0_4_42 (.A1(n_0_66), .A2(\Memory[15] [1]), .ZN(n_0_4_41));
   NAND2_X1 i_0_4_43 (.A1(n_0_51), .A2(\Memory[0] [1]), .ZN(n_0_4_42));
   NAND2_X1 i_0_4_44 (.A1(n_0_60), .A2(\Memory[9] [1]), .ZN(n_0_4_43));
   NAND4_X1 i_0_4_45 (.A1(n_0_4_40), .A2(n_0_4_41), .A3(n_0_4_42), .A4(n_0_4_43), 
      .ZN(n_0_4_44));
   NAND2_X1 i_0_4_46 (.A1(n_0_64), .A2(\Memory[13] [1]), .ZN(n_0_4_45));
   NAND2_X1 i_0_4_47 (.A1(n_0_63), .A2(\Memory[12] [1]), .ZN(n_0_4_46));
   NAND2_X1 i_0_4_48 (.A1(n_0_62), .A2(\Memory[11] [1]), .ZN(n_0_4_47));
   NAND3_X1 i_0_4_49 (.A1(n_0_4_45), .A2(n_0_4_46), .A3(n_0_4_47), .ZN(n_0_4_48));
   NOR2_X1 i_0_4_50 (.A1(n_0_4_44), .A2(n_0_4_48), .ZN(n_0_4_49));
   NAND3_X1 i_0_4_51 (.A1(n_0_4_30), .A2(n_0_4_39), .A3(n_0_4_49), .ZN(
      dataOut2[1]));
   NAND2_X1 i_0_4_52 (.A1(n_0_55), .A2(\Memory[4] [2]), .ZN(n_0_4_50));
   NAND2_X1 i_0_4_53 (.A1(n_0_58), .A2(\Memory[7] [2]), .ZN(n_0_4_51));
   NAND2_X1 i_0_4_54 (.A1(n_0_54), .A2(\Memory[3] [2]), .ZN(n_0_4_52));
   NAND2_X1 i_0_4_55 (.A1(n_0_53), .A2(\Memory[2] [2]), .ZN(n_0_4_53));
   NAND4_X1 i_0_4_56 (.A1(n_0_4_50), .A2(n_0_4_51), .A3(n_0_4_52), .A4(n_0_4_53), 
      .ZN(n_0_4_54));
   INV_X1 i_0_4_57 (.A(n_0_4_54), .ZN(n_0_4_55));
   NAND2_X1 i_0_4_58 (.A1(n_0_67), .A2(\Memory[16] [2]), .ZN(n_0_4_56));
   NAND2_X1 i_0_4_59 (.A1(n_0_57), .A2(\Memory[6] [2]), .ZN(n_0_4_57));
   NAND2_X1 i_0_4_60 (.A1(n_0_56), .A2(\Memory[5] [2]), .ZN(n_0_4_58));
   NAND3_X1 i_0_4_61 (.A1(n_0_4_56), .A2(n_0_4_57), .A3(n_0_4_58), .ZN(n_0_4_59));
   NAND2_X1 i_0_4_62 (.A1(n_0_59), .A2(\Memory[8] [2]), .ZN(n_0_4_60));
   NAND2_X1 i_0_4_63 (.A1(n_0_52), .A2(\Memory[1] [2]), .ZN(n_0_4_61));
   NAND2_X1 i_0_4_64 (.A1(n_0_61), .A2(\Memory[10] [2]), .ZN(n_0_4_62));
   NAND3_X1 i_0_4_65 (.A1(n_0_4_60), .A2(n_0_4_61), .A3(n_0_4_62), .ZN(n_0_4_63));
   NOR2_X1 i_0_4_66 (.A1(n_0_4_59), .A2(n_0_4_63), .ZN(n_0_4_64));
   NAND2_X1 i_0_4_67 (.A1(n_0_65), .A2(\Memory[14] [2]), .ZN(n_0_4_65));
   NAND2_X1 i_0_4_68 (.A1(n_0_66), .A2(\Memory[15] [2]), .ZN(n_0_4_66));
   NAND2_X1 i_0_4_69 (.A1(n_0_51), .A2(\Memory[0] [2]), .ZN(n_0_4_67));
   NAND2_X1 i_0_4_70 (.A1(n_0_60), .A2(\Memory[9] [2]), .ZN(n_0_4_68));
   NAND4_X1 i_0_4_71 (.A1(n_0_4_65), .A2(n_0_4_66), .A3(n_0_4_67), .A4(n_0_4_68), 
      .ZN(n_0_4_69));
   NAND2_X1 i_0_4_72 (.A1(n_0_64), .A2(\Memory[13] [2]), .ZN(n_0_4_70));
   NAND2_X1 i_0_4_73 (.A1(n_0_63), .A2(\Memory[12] [2]), .ZN(n_0_4_71));
   NAND2_X1 i_0_4_74 (.A1(n_0_62), .A2(\Memory[11] [2]), .ZN(n_0_4_72));
   NAND3_X1 i_0_4_75 (.A1(n_0_4_70), .A2(n_0_4_71), .A3(n_0_4_72), .ZN(n_0_4_73));
   NOR2_X1 i_0_4_76 (.A1(n_0_4_69), .A2(n_0_4_73), .ZN(n_0_4_74));
   NAND3_X1 i_0_4_77 (.A1(n_0_4_55), .A2(n_0_4_64), .A3(n_0_4_74), .ZN(
      dataOut2[2]));
   NAND2_X1 i_0_4_78 (.A1(n_0_55), .A2(\Memory[4] [3]), .ZN(n_0_4_75));
   NAND2_X1 i_0_4_79 (.A1(n_0_58), .A2(\Memory[7] [3]), .ZN(n_0_4_76));
   NAND2_X1 i_0_4_80 (.A1(n_0_54), .A2(\Memory[3] [3]), .ZN(n_0_4_77));
   NAND2_X1 i_0_4_81 (.A1(n_0_53), .A2(\Memory[2] [3]), .ZN(n_0_4_78));
   NAND4_X1 i_0_4_82 (.A1(n_0_4_75), .A2(n_0_4_76), .A3(n_0_4_77), .A4(n_0_4_78), 
      .ZN(n_0_4_79));
   INV_X1 i_0_4_83 (.A(n_0_4_79), .ZN(n_0_4_80));
   NAND2_X1 i_0_4_84 (.A1(n_0_67), .A2(\Memory[16] [3]), .ZN(n_0_4_81));
   NAND2_X1 i_0_4_85 (.A1(n_0_57), .A2(\Memory[6] [3]), .ZN(n_0_4_82));
   NAND2_X1 i_0_4_86 (.A1(n_0_56), .A2(\Memory[5] [3]), .ZN(n_0_4_83));
   NAND3_X1 i_0_4_87 (.A1(n_0_4_81), .A2(n_0_4_82), .A3(n_0_4_83), .ZN(n_0_4_84));
   NAND2_X1 i_0_4_88 (.A1(n_0_59), .A2(\Memory[8] [3]), .ZN(n_0_4_85));
   NAND2_X1 i_0_4_89 (.A1(n_0_52), .A2(\Memory[1] [3]), .ZN(n_0_4_86));
   NAND2_X1 i_0_4_90 (.A1(n_0_61), .A2(\Memory[10] [3]), .ZN(n_0_4_87));
   NAND3_X1 i_0_4_91 (.A1(n_0_4_85), .A2(n_0_4_86), .A3(n_0_4_87), .ZN(n_0_4_88));
   NOR2_X1 i_0_4_92 (.A1(n_0_4_84), .A2(n_0_4_88), .ZN(n_0_4_89));
   NAND2_X1 i_0_4_93 (.A1(n_0_65), .A2(\Memory[14] [3]), .ZN(n_0_4_90));
   NAND2_X1 i_0_4_94 (.A1(n_0_66), .A2(\Memory[15] [3]), .ZN(n_0_4_91));
   NAND2_X1 i_0_4_95 (.A1(n_0_51), .A2(\Memory[0] [3]), .ZN(n_0_4_92));
   NAND2_X1 i_0_4_96 (.A1(n_0_60), .A2(\Memory[9] [3]), .ZN(n_0_4_93));
   NAND4_X1 i_0_4_97 (.A1(n_0_4_90), .A2(n_0_4_91), .A3(n_0_4_92), .A4(n_0_4_93), 
      .ZN(n_0_4_94));
   NAND2_X1 i_0_4_98 (.A1(n_0_64), .A2(\Memory[13] [3]), .ZN(n_0_4_95));
   NAND2_X1 i_0_4_99 (.A1(n_0_63), .A2(\Memory[12] [3]), .ZN(n_0_4_96));
   NAND2_X1 i_0_4_100 (.A1(n_0_62), .A2(\Memory[11] [3]), .ZN(n_0_4_97));
   NAND3_X1 i_0_4_101 (.A1(n_0_4_95), .A2(n_0_4_96), .A3(n_0_4_97), .ZN(n_0_4_98));
   NOR2_X1 i_0_4_102 (.A1(n_0_4_94), .A2(n_0_4_98), .ZN(n_0_4_99));
   NAND3_X1 i_0_4_103 (.A1(n_0_4_80), .A2(n_0_4_89), .A3(n_0_4_99), .ZN(
      dataOut2[3]));
   NAND2_X1 i_0_4_104 (.A1(n_0_55), .A2(\Memory[4] [4]), .ZN(n_0_4_100));
   NAND2_X1 i_0_4_105 (.A1(n_0_58), .A2(\Memory[7] [4]), .ZN(n_0_4_101));
   NAND2_X1 i_0_4_106 (.A1(n_0_54), .A2(\Memory[3] [4]), .ZN(n_0_4_102));
   NAND2_X1 i_0_4_107 (.A1(n_0_53), .A2(\Memory[2] [4]), .ZN(n_0_4_103));
   NAND4_X1 i_0_4_108 (.A1(n_0_4_100), .A2(n_0_4_101), .A3(n_0_4_102), .A4(
      n_0_4_103), .ZN(n_0_4_104));
   INV_X1 i_0_4_109 (.A(n_0_4_104), .ZN(n_0_4_105));
   NAND2_X1 i_0_4_110 (.A1(n_0_67), .A2(\Memory[16] [4]), .ZN(n_0_4_106));
   NAND2_X1 i_0_4_111 (.A1(n_0_57), .A2(\Memory[6] [4]), .ZN(n_0_4_107));
   NAND2_X1 i_0_4_112 (.A1(n_0_56), .A2(\Memory[5] [4]), .ZN(n_0_4_108));
   NAND3_X1 i_0_4_113 (.A1(n_0_4_106), .A2(n_0_4_107), .A3(n_0_4_108), .ZN(
      n_0_4_109));
   NAND2_X1 i_0_4_114 (.A1(n_0_59), .A2(\Memory[8] [4]), .ZN(n_0_4_110));
   NAND2_X1 i_0_4_115 (.A1(n_0_52), .A2(\Memory[1] [4]), .ZN(n_0_4_111));
   NAND2_X1 i_0_4_116 (.A1(n_0_61), .A2(\Memory[10] [4]), .ZN(n_0_4_112));
   NAND3_X1 i_0_4_117 (.A1(n_0_4_110), .A2(n_0_4_111), .A3(n_0_4_112), .ZN(
      n_0_4_113));
   NOR2_X1 i_0_4_118 (.A1(n_0_4_109), .A2(n_0_4_113), .ZN(n_0_4_114));
   NAND2_X1 i_0_4_119 (.A1(n_0_65), .A2(\Memory[14] [4]), .ZN(n_0_4_115));
   NAND2_X1 i_0_4_120 (.A1(n_0_66), .A2(\Memory[15] [4]), .ZN(n_0_4_116));
   NAND2_X1 i_0_4_121 (.A1(n_0_51), .A2(\Memory[0] [4]), .ZN(n_0_4_117));
   NAND2_X1 i_0_4_122 (.A1(n_0_60), .A2(\Memory[9] [4]), .ZN(n_0_4_118));
   NAND4_X1 i_0_4_123 (.A1(n_0_4_115), .A2(n_0_4_116), .A3(n_0_4_117), .A4(
      n_0_4_118), .ZN(n_0_4_119));
   NAND2_X1 i_0_4_124 (.A1(n_0_64), .A2(\Memory[13] [4]), .ZN(n_0_4_120));
   NAND2_X1 i_0_4_125 (.A1(n_0_63), .A2(\Memory[12] [4]), .ZN(n_0_4_121));
   NAND2_X1 i_0_4_126 (.A1(n_0_62), .A2(\Memory[11] [4]), .ZN(n_0_4_122));
   NAND3_X1 i_0_4_127 (.A1(n_0_4_120), .A2(n_0_4_121), .A3(n_0_4_122), .ZN(
      n_0_4_123));
   NOR2_X1 i_0_4_128 (.A1(n_0_4_119), .A2(n_0_4_123), .ZN(n_0_4_124));
   NAND3_X1 i_0_4_129 (.A1(n_0_4_105), .A2(n_0_4_114), .A3(n_0_4_124), .ZN(
      dataOut2[4]));
   NAND2_X1 i_0_4_130 (.A1(n_0_55), .A2(\Memory[4] [5]), .ZN(n_0_4_125));
   NAND2_X1 i_0_4_131 (.A1(n_0_58), .A2(\Memory[7] [5]), .ZN(n_0_4_126));
   NAND2_X1 i_0_4_132 (.A1(n_0_54), .A2(\Memory[3] [5]), .ZN(n_0_4_127));
   NAND2_X1 i_0_4_133 (.A1(n_0_53), .A2(\Memory[2] [5]), .ZN(n_0_4_128));
   NAND4_X1 i_0_4_134 (.A1(n_0_4_125), .A2(n_0_4_126), .A3(n_0_4_127), .A4(
      n_0_4_128), .ZN(n_0_4_129));
   INV_X1 i_0_4_135 (.A(n_0_4_129), .ZN(n_0_4_130));
   NAND2_X1 i_0_4_136 (.A1(n_0_67), .A2(\Memory[16] [5]), .ZN(n_0_4_131));
   NAND2_X1 i_0_4_137 (.A1(n_0_57), .A2(\Memory[6] [5]), .ZN(n_0_4_132));
   NAND2_X1 i_0_4_138 (.A1(n_0_56), .A2(\Memory[5] [5]), .ZN(n_0_4_133));
   NAND3_X1 i_0_4_139 (.A1(n_0_4_131), .A2(n_0_4_132), .A3(n_0_4_133), .ZN(
      n_0_4_134));
   NAND2_X1 i_0_4_140 (.A1(n_0_59), .A2(\Memory[8] [5]), .ZN(n_0_4_135));
   NAND2_X1 i_0_4_141 (.A1(n_0_52), .A2(\Memory[1] [5]), .ZN(n_0_4_136));
   NAND2_X1 i_0_4_142 (.A1(n_0_61), .A2(\Memory[10] [5]), .ZN(n_0_4_137));
   NAND3_X1 i_0_4_143 (.A1(n_0_4_135), .A2(n_0_4_136), .A3(n_0_4_137), .ZN(
      n_0_4_138));
   NOR2_X1 i_0_4_144 (.A1(n_0_4_134), .A2(n_0_4_138), .ZN(n_0_4_139));
   NAND2_X1 i_0_4_145 (.A1(n_0_65), .A2(\Memory[14] [5]), .ZN(n_0_4_140));
   NAND2_X1 i_0_4_146 (.A1(n_0_66), .A2(\Memory[15] [5]), .ZN(n_0_4_141));
   NAND2_X1 i_0_4_147 (.A1(n_0_51), .A2(\Memory[0] [5]), .ZN(n_0_4_142));
   NAND2_X1 i_0_4_148 (.A1(n_0_60), .A2(\Memory[9] [5]), .ZN(n_0_4_143));
   NAND4_X1 i_0_4_149 (.A1(n_0_4_140), .A2(n_0_4_141), .A3(n_0_4_142), .A4(
      n_0_4_143), .ZN(n_0_4_144));
   NAND2_X1 i_0_4_150 (.A1(n_0_64), .A2(\Memory[13] [5]), .ZN(n_0_4_145));
   NAND2_X1 i_0_4_151 (.A1(n_0_63), .A2(\Memory[12] [5]), .ZN(n_0_4_146));
   NAND2_X1 i_0_4_152 (.A1(n_0_62), .A2(\Memory[11] [5]), .ZN(n_0_4_147));
   NAND3_X1 i_0_4_153 (.A1(n_0_4_145), .A2(n_0_4_146), .A3(n_0_4_147), .ZN(
      n_0_4_148));
   NOR2_X1 i_0_4_154 (.A1(n_0_4_144), .A2(n_0_4_148), .ZN(n_0_4_149));
   NAND3_X1 i_0_4_155 (.A1(n_0_4_130), .A2(n_0_4_139), .A3(n_0_4_149), .ZN(
      dataOut2[5]));
   NAND2_X1 i_0_4_156 (.A1(n_0_55), .A2(\Memory[4] [6]), .ZN(n_0_4_150));
   NAND2_X1 i_0_4_157 (.A1(n_0_58), .A2(\Memory[7] [6]), .ZN(n_0_4_151));
   NAND2_X1 i_0_4_158 (.A1(n_0_54), .A2(\Memory[3] [6]), .ZN(n_0_4_152));
   NAND2_X1 i_0_4_159 (.A1(n_0_53), .A2(\Memory[2] [6]), .ZN(n_0_4_153));
   NAND4_X1 i_0_4_160 (.A1(n_0_4_150), .A2(n_0_4_151), .A3(n_0_4_152), .A4(
      n_0_4_153), .ZN(n_0_4_154));
   INV_X1 i_0_4_161 (.A(n_0_4_154), .ZN(n_0_4_155));
   NAND2_X1 i_0_4_162 (.A1(n_0_67), .A2(\Memory[16] [6]), .ZN(n_0_4_156));
   NAND2_X1 i_0_4_163 (.A1(n_0_57), .A2(\Memory[6] [6]), .ZN(n_0_4_157));
   NAND2_X1 i_0_4_164 (.A1(n_0_56), .A2(\Memory[5] [6]), .ZN(n_0_4_158));
   NAND3_X1 i_0_4_165 (.A1(n_0_4_156), .A2(n_0_4_157), .A3(n_0_4_158), .ZN(
      n_0_4_159));
   NAND2_X1 i_0_4_166 (.A1(n_0_59), .A2(\Memory[8] [6]), .ZN(n_0_4_160));
   NAND2_X1 i_0_4_167 (.A1(n_0_52), .A2(\Memory[1] [6]), .ZN(n_0_4_161));
   NAND2_X1 i_0_4_168 (.A1(n_0_61), .A2(\Memory[10] [6]), .ZN(n_0_4_162));
   NAND3_X1 i_0_4_169 (.A1(n_0_4_160), .A2(n_0_4_161), .A3(n_0_4_162), .ZN(
      n_0_4_163));
   NOR2_X1 i_0_4_170 (.A1(n_0_4_159), .A2(n_0_4_163), .ZN(n_0_4_164));
   NAND2_X1 i_0_4_171 (.A1(n_0_65), .A2(\Memory[14] [6]), .ZN(n_0_4_165));
   NAND2_X1 i_0_4_172 (.A1(n_0_66), .A2(\Memory[15] [6]), .ZN(n_0_4_166));
   NAND2_X1 i_0_4_173 (.A1(n_0_51), .A2(\Memory[0] [6]), .ZN(n_0_4_167));
   NAND2_X1 i_0_4_174 (.A1(n_0_60), .A2(\Memory[9] [6]), .ZN(n_0_4_168));
   NAND4_X1 i_0_4_175 (.A1(n_0_4_165), .A2(n_0_4_166), .A3(n_0_4_167), .A4(
      n_0_4_168), .ZN(n_0_4_169));
   NAND2_X1 i_0_4_176 (.A1(n_0_64), .A2(\Memory[13] [6]), .ZN(n_0_4_170));
   NAND2_X1 i_0_4_177 (.A1(n_0_63), .A2(\Memory[12] [6]), .ZN(n_0_4_171));
   NAND2_X1 i_0_4_178 (.A1(n_0_62), .A2(\Memory[11] [6]), .ZN(n_0_4_172));
   NAND3_X1 i_0_4_179 (.A1(n_0_4_170), .A2(n_0_4_171), .A3(n_0_4_172), .ZN(
      n_0_4_173));
   NOR2_X1 i_0_4_180 (.A1(n_0_4_169), .A2(n_0_4_173), .ZN(n_0_4_174));
   NAND3_X1 i_0_4_181 (.A1(n_0_4_155), .A2(n_0_4_164), .A3(n_0_4_174), .ZN(
      dataOut2[6]));
   NAND2_X1 i_0_4_182 (.A1(n_0_55), .A2(\Memory[4] [7]), .ZN(n_0_4_175));
   NAND2_X1 i_0_4_183 (.A1(n_0_58), .A2(\Memory[7] [7]), .ZN(n_0_4_176));
   NAND2_X1 i_0_4_184 (.A1(n_0_54), .A2(\Memory[3] [7]), .ZN(n_0_4_177));
   NAND2_X1 i_0_4_185 (.A1(n_0_53), .A2(\Memory[2] [7]), .ZN(n_0_4_178));
   NAND4_X1 i_0_4_186 (.A1(n_0_4_175), .A2(n_0_4_176), .A3(n_0_4_177), .A4(
      n_0_4_178), .ZN(n_0_4_179));
   INV_X1 i_0_4_187 (.A(n_0_4_179), .ZN(n_0_4_180));
   NAND2_X1 i_0_4_188 (.A1(n_0_67), .A2(\Memory[16] [7]), .ZN(n_0_4_181));
   NAND2_X1 i_0_4_189 (.A1(n_0_57), .A2(\Memory[6] [7]), .ZN(n_0_4_182));
   NAND2_X1 i_0_4_190 (.A1(n_0_56), .A2(\Memory[5] [7]), .ZN(n_0_4_183));
   NAND3_X1 i_0_4_191 (.A1(n_0_4_181), .A2(n_0_4_182), .A3(n_0_4_183), .ZN(
      n_0_4_184));
   NAND2_X1 i_0_4_192 (.A1(n_0_59), .A2(\Memory[8] [7]), .ZN(n_0_4_185));
   NAND2_X1 i_0_4_193 (.A1(n_0_52), .A2(\Memory[1] [7]), .ZN(n_0_4_186));
   NAND2_X1 i_0_4_194 (.A1(n_0_61), .A2(\Memory[10] [7]), .ZN(n_0_4_187));
   NAND3_X1 i_0_4_195 (.A1(n_0_4_185), .A2(n_0_4_186), .A3(n_0_4_187), .ZN(
      n_0_4_188));
   NOR2_X1 i_0_4_196 (.A1(n_0_4_184), .A2(n_0_4_188), .ZN(n_0_4_189));
   NAND2_X1 i_0_4_197 (.A1(n_0_65), .A2(\Memory[14] [7]), .ZN(n_0_4_190));
   NAND2_X1 i_0_4_198 (.A1(n_0_66), .A2(\Memory[15] [7]), .ZN(n_0_4_191));
   NAND2_X1 i_0_4_199 (.A1(n_0_51), .A2(\Memory[0] [7]), .ZN(n_0_4_192));
   NAND2_X1 i_0_4_200 (.A1(n_0_60), .A2(\Memory[9] [7]), .ZN(n_0_4_193));
   NAND4_X1 i_0_4_201 (.A1(n_0_4_190), .A2(n_0_4_191), .A3(n_0_4_192), .A4(
      n_0_4_193), .ZN(n_0_4_194));
   NAND2_X1 i_0_4_202 (.A1(n_0_64), .A2(\Memory[13] [7]), .ZN(n_0_4_195));
   NAND2_X1 i_0_4_203 (.A1(n_0_63), .A2(\Memory[12] [7]), .ZN(n_0_4_196));
   NAND2_X1 i_0_4_204 (.A1(n_0_62), .A2(\Memory[11] [7]), .ZN(n_0_4_197));
   NAND3_X1 i_0_4_205 (.A1(n_0_4_195), .A2(n_0_4_196), .A3(n_0_4_197), .ZN(
      n_0_4_198));
   NOR2_X1 i_0_4_206 (.A1(n_0_4_194), .A2(n_0_4_198), .ZN(n_0_4_199));
   NAND3_X1 i_0_4_207 (.A1(n_0_4_180), .A2(n_0_4_189), .A3(n_0_4_199), .ZN(
      dataOut2[7]));
   NAND2_X1 i_0_4_208 (.A1(n_0_55), .A2(\Memory[4] [8]), .ZN(n_0_4_200));
   NAND2_X1 i_0_4_209 (.A1(n_0_58), .A2(\Memory[7] [8]), .ZN(n_0_4_201));
   NAND2_X1 i_0_4_210 (.A1(n_0_54), .A2(\Memory[3] [8]), .ZN(n_0_4_202));
   NAND2_X1 i_0_4_211 (.A1(n_0_53), .A2(\Memory[2] [8]), .ZN(n_0_4_203));
   NAND4_X1 i_0_4_212 (.A1(n_0_4_200), .A2(n_0_4_201), .A3(n_0_4_202), .A4(
      n_0_4_203), .ZN(n_0_4_204));
   INV_X1 i_0_4_213 (.A(n_0_4_204), .ZN(n_0_4_205));
   NAND2_X1 i_0_4_214 (.A1(n_0_67), .A2(\Memory[16] [8]), .ZN(n_0_4_206));
   NAND2_X1 i_0_4_215 (.A1(n_0_57), .A2(\Memory[6] [8]), .ZN(n_0_4_207));
   NAND2_X1 i_0_4_216 (.A1(n_0_56), .A2(\Memory[5] [8]), .ZN(n_0_4_208));
   NAND3_X1 i_0_4_217 (.A1(n_0_4_206), .A2(n_0_4_207), .A3(n_0_4_208), .ZN(
      n_0_4_209));
   NAND2_X1 i_0_4_218 (.A1(n_0_59), .A2(\Memory[8] [8]), .ZN(n_0_4_210));
   NAND2_X1 i_0_4_219 (.A1(n_0_52), .A2(\Memory[1] [8]), .ZN(n_0_4_211));
   NAND2_X1 i_0_4_220 (.A1(n_0_61), .A2(\Memory[10] [8]), .ZN(n_0_4_212));
   NAND3_X1 i_0_4_221 (.A1(n_0_4_210), .A2(n_0_4_211), .A3(n_0_4_212), .ZN(
      n_0_4_213));
   NOR2_X1 i_0_4_222 (.A1(n_0_4_209), .A2(n_0_4_213), .ZN(n_0_4_214));
   NAND2_X1 i_0_4_223 (.A1(n_0_65), .A2(\Memory[14] [8]), .ZN(n_0_4_215));
   NAND2_X1 i_0_4_224 (.A1(n_0_66), .A2(\Memory[15] [8]), .ZN(n_0_4_216));
   NAND2_X1 i_0_4_225 (.A1(n_0_51), .A2(\Memory[0] [8]), .ZN(n_0_4_217));
   NAND2_X1 i_0_4_226 (.A1(n_0_60), .A2(\Memory[9] [8]), .ZN(n_0_4_218));
   NAND4_X1 i_0_4_227 (.A1(n_0_4_215), .A2(n_0_4_216), .A3(n_0_4_217), .A4(
      n_0_4_218), .ZN(n_0_4_219));
   NAND2_X1 i_0_4_228 (.A1(n_0_64), .A2(\Memory[13] [8]), .ZN(n_0_4_220));
   NAND2_X1 i_0_4_229 (.A1(n_0_63), .A2(\Memory[12] [8]), .ZN(n_0_4_221));
   NAND2_X1 i_0_4_230 (.A1(n_0_62), .A2(\Memory[11] [8]), .ZN(n_0_4_222));
   NAND3_X1 i_0_4_231 (.A1(n_0_4_220), .A2(n_0_4_221), .A3(n_0_4_222), .ZN(
      n_0_4_223));
   NOR2_X1 i_0_4_232 (.A1(n_0_4_219), .A2(n_0_4_223), .ZN(n_0_4_224));
   NAND3_X1 i_0_4_233 (.A1(n_0_4_205), .A2(n_0_4_214), .A3(n_0_4_224), .ZN(
      dataOut2[8]));
   NAND2_X1 i_0_4_234 (.A1(n_0_55), .A2(\Memory[4] [9]), .ZN(n_0_4_225));
   NAND2_X1 i_0_4_235 (.A1(n_0_58), .A2(\Memory[7] [9]), .ZN(n_0_4_226));
   NAND2_X1 i_0_4_236 (.A1(n_0_54), .A2(\Memory[3] [9]), .ZN(n_0_4_227));
   NAND2_X1 i_0_4_237 (.A1(n_0_53), .A2(\Memory[2] [9]), .ZN(n_0_4_228));
   NAND4_X1 i_0_4_238 (.A1(n_0_4_225), .A2(n_0_4_226), .A3(n_0_4_227), .A4(
      n_0_4_228), .ZN(n_0_4_229));
   INV_X1 i_0_4_239 (.A(n_0_4_229), .ZN(n_0_4_230));
   NAND2_X1 i_0_4_240 (.A1(n_0_67), .A2(\Memory[16] [9]), .ZN(n_0_4_231));
   NAND2_X1 i_0_4_241 (.A1(n_0_57), .A2(\Memory[6] [9]), .ZN(n_0_4_232));
   NAND2_X1 i_0_4_242 (.A1(n_0_56), .A2(\Memory[5] [9]), .ZN(n_0_4_233));
   NAND3_X1 i_0_4_243 (.A1(n_0_4_231), .A2(n_0_4_232), .A3(n_0_4_233), .ZN(
      n_0_4_234));
   NAND2_X1 i_0_4_244 (.A1(n_0_59), .A2(\Memory[8] [9]), .ZN(n_0_4_235));
   NAND2_X1 i_0_4_245 (.A1(n_0_52), .A2(\Memory[1] [9]), .ZN(n_0_4_236));
   NAND2_X1 i_0_4_246 (.A1(n_0_61), .A2(\Memory[10] [9]), .ZN(n_0_4_237));
   NAND3_X1 i_0_4_247 (.A1(n_0_4_235), .A2(n_0_4_236), .A3(n_0_4_237), .ZN(
      n_0_4_238));
   NOR2_X1 i_0_4_248 (.A1(n_0_4_234), .A2(n_0_4_238), .ZN(n_0_4_239));
   NAND2_X1 i_0_4_249 (.A1(n_0_65), .A2(\Memory[14] [9]), .ZN(n_0_4_240));
   NAND2_X1 i_0_4_250 (.A1(n_0_66), .A2(\Memory[15] [9]), .ZN(n_0_4_241));
   NAND2_X1 i_0_4_251 (.A1(n_0_51), .A2(\Memory[0] [9]), .ZN(n_0_4_242));
   NAND2_X1 i_0_4_252 (.A1(n_0_60), .A2(\Memory[9] [9]), .ZN(n_0_4_243));
   NAND4_X1 i_0_4_253 (.A1(n_0_4_240), .A2(n_0_4_241), .A3(n_0_4_242), .A4(
      n_0_4_243), .ZN(n_0_4_244));
   NAND2_X1 i_0_4_254 (.A1(n_0_64), .A2(\Memory[13] [9]), .ZN(n_0_4_245));
   NAND2_X1 i_0_4_255 (.A1(n_0_63), .A2(\Memory[12] [9]), .ZN(n_0_4_246));
   NAND2_X1 i_0_4_256 (.A1(n_0_62), .A2(\Memory[11] [9]), .ZN(n_0_4_247));
   NAND3_X1 i_0_4_257 (.A1(n_0_4_245), .A2(n_0_4_246), .A3(n_0_4_247), .ZN(
      n_0_4_248));
   NOR2_X1 i_0_4_258 (.A1(n_0_4_244), .A2(n_0_4_248), .ZN(n_0_4_249));
   NAND3_X1 i_0_4_259 (.A1(n_0_4_230), .A2(n_0_4_239), .A3(n_0_4_249), .ZN(
      dataOut2[9]));
   NAND2_X1 i_0_4_260 (.A1(n_0_55), .A2(\Memory[4] [10]), .ZN(n_0_4_250));
   NAND2_X1 i_0_4_261 (.A1(n_0_58), .A2(\Memory[7] [10]), .ZN(n_0_4_251));
   NAND2_X1 i_0_4_262 (.A1(n_0_54), .A2(\Memory[3] [10]), .ZN(n_0_4_252));
   NAND2_X1 i_0_4_263 (.A1(n_0_53), .A2(\Memory[2] [10]), .ZN(n_0_4_253));
   NAND4_X1 i_0_4_264 (.A1(n_0_4_250), .A2(n_0_4_251), .A3(n_0_4_252), .A4(
      n_0_4_253), .ZN(n_0_4_254));
   INV_X1 i_0_4_265 (.A(n_0_4_254), .ZN(n_0_4_255));
   NAND2_X1 i_0_4_266 (.A1(n_0_67), .A2(\Memory[16] [10]), .ZN(n_0_4_256));
   NAND2_X1 i_0_4_267 (.A1(n_0_57), .A2(\Memory[6] [10]), .ZN(n_0_4_257));
   NAND2_X1 i_0_4_268 (.A1(n_0_56), .A2(\Memory[5] [10]), .ZN(n_0_4_258));
   NAND3_X1 i_0_4_269 (.A1(n_0_4_256), .A2(n_0_4_257), .A3(n_0_4_258), .ZN(
      n_0_4_259));
   NAND2_X1 i_0_4_270 (.A1(n_0_59), .A2(\Memory[8] [10]), .ZN(n_0_4_260));
   NAND2_X1 i_0_4_271 (.A1(n_0_52), .A2(\Memory[1] [10]), .ZN(n_0_4_261));
   NAND2_X1 i_0_4_272 (.A1(n_0_61), .A2(\Memory[10] [10]), .ZN(n_0_4_262));
   NAND3_X1 i_0_4_273 (.A1(n_0_4_260), .A2(n_0_4_261), .A3(n_0_4_262), .ZN(
      n_0_4_263));
   NOR2_X1 i_0_4_274 (.A1(n_0_4_259), .A2(n_0_4_263), .ZN(n_0_4_264));
   NAND2_X1 i_0_4_275 (.A1(n_0_65), .A2(\Memory[14] [10]), .ZN(n_0_4_265));
   NAND2_X1 i_0_4_276 (.A1(n_0_66), .A2(\Memory[15] [10]), .ZN(n_0_4_266));
   NAND2_X1 i_0_4_277 (.A1(n_0_51), .A2(\Memory[0] [10]), .ZN(n_0_4_267));
   NAND2_X1 i_0_4_278 (.A1(n_0_60), .A2(\Memory[9] [10]), .ZN(n_0_4_268));
   NAND4_X1 i_0_4_279 (.A1(n_0_4_265), .A2(n_0_4_266), .A3(n_0_4_267), .A4(
      n_0_4_268), .ZN(n_0_4_269));
   NAND2_X1 i_0_4_280 (.A1(n_0_64), .A2(\Memory[13] [10]), .ZN(n_0_4_270));
   NAND2_X1 i_0_4_281 (.A1(n_0_63), .A2(\Memory[12] [10]), .ZN(n_0_4_271));
   NAND2_X1 i_0_4_282 (.A1(n_0_62), .A2(\Memory[11] [10]), .ZN(n_0_4_272));
   NAND3_X1 i_0_4_283 (.A1(n_0_4_270), .A2(n_0_4_271), .A3(n_0_4_272), .ZN(
      n_0_4_273));
   NOR2_X1 i_0_4_284 (.A1(n_0_4_269), .A2(n_0_4_273), .ZN(n_0_4_274));
   NAND3_X1 i_0_4_285 (.A1(n_0_4_255), .A2(n_0_4_264), .A3(n_0_4_274), .ZN(
      dataOut2[10]));
   NAND2_X1 i_0_4_286 (.A1(n_0_55), .A2(\Memory[4] [11]), .ZN(n_0_4_275));
   NAND2_X1 i_0_4_287 (.A1(n_0_58), .A2(\Memory[7] [11]), .ZN(n_0_4_276));
   NAND2_X1 i_0_4_288 (.A1(n_0_54), .A2(\Memory[3] [11]), .ZN(n_0_4_277));
   NAND2_X1 i_0_4_289 (.A1(n_0_53), .A2(\Memory[2] [11]), .ZN(n_0_4_278));
   NAND4_X1 i_0_4_290 (.A1(n_0_4_275), .A2(n_0_4_276), .A3(n_0_4_277), .A4(
      n_0_4_278), .ZN(n_0_4_279));
   INV_X1 i_0_4_291 (.A(n_0_4_279), .ZN(n_0_4_280));
   NAND2_X1 i_0_4_292 (.A1(n_0_67), .A2(\Memory[16] [11]), .ZN(n_0_4_281));
   NAND2_X1 i_0_4_293 (.A1(n_0_57), .A2(\Memory[6] [11]), .ZN(n_0_4_282));
   NAND2_X1 i_0_4_294 (.A1(n_0_56), .A2(\Memory[5] [11]), .ZN(n_0_4_283));
   NAND3_X1 i_0_4_295 (.A1(n_0_4_281), .A2(n_0_4_282), .A3(n_0_4_283), .ZN(
      n_0_4_284));
   NAND2_X1 i_0_4_296 (.A1(n_0_59), .A2(\Memory[8] [11]), .ZN(n_0_4_285));
   NAND2_X1 i_0_4_297 (.A1(n_0_52), .A2(\Memory[1] [11]), .ZN(n_0_4_286));
   NAND2_X1 i_0_4_298 (.A1(n_0_61), .A2(\Memory[10] [11]), .ZN(n_0_4_287));
   NAND3_X1 i_0_4_299 (.A1(n_0_4_285), .A2(n_0_4_286), .A3(n_0_4_287), .ZN(
      n_0_4_288));
   NOR2_X1 i_0_4_300 (.A1(n_0_4_284), .A2(n_0_4_288), .ZN(n_0_4_289));
   NAND2_X1 i_0_4_301 (.A1(n_0_65), .A2(\Memory[14] [11]), .ZN(n_0_4_290));
   NAND2_X1 i_0_4_302 (.A1(n_0_66), .A2(\Memory[15] [11]), .ZN(n_0_4_291));
   NAND2_X1 i_0_4_303 (.A1(n_0_51), .A2(\Memory[0] [11]), .ZN(n_0_4_292));
   NAND2_X1 i_0_4_304 (.A1(n_0_60), .A2(\Memory[9] [11]), .ZN(n_0_4_293));
   NAND4_X1 i_0_4_305 (.A1(n_0_4_290), .A2(n_0_4_291), .A3(n_0_4_292), .A4(
      n_0_4_293), .ZN(n_0_4_294));
   NAND2_X1 i_0_4_306 (.A1(n_0_64), .A2(\Memory[13] [11]), .ZN(n_0_4_295));
   NAND2_X1 i_0_4_307 (.A1(n_0_63), .A2(\Memory[12] [11]), .ZN(n_0_4_296));
   NAND2_X1 i_0_4_308 (.A1(n_0_62), .A2(\Memory[11] [11]), .ZN(n_0_4_297));
   NAND3_X1 i_0_4_309 (.A1(n_0_4_295), .A2(n_0_4_296), .A3(n_0_4_297), .ZN(
      n_0_4_298));
   NOR2_X1 i_0_4_310 (.A1(n_0_4_294), .A2(n_0_4_298), .ZN(n_0_4_299));
   NAND3_X1 i_0_4_311 (.A1(n_0_4_280), .A2(n_0_4_289), .A3(n_0_4_299), .ZN(
      dataOut2[11]));
   NAND2_X1 i_0_4_312 (.A1(n_0_55), .A2(\Memory[4] [12]), .ZN(n_0_4_300));
   NAND2_X1 i_0_4_313 (.A1(n_0_58), .A2(\Memory[7] [12]), .ZN(n_0_4_301));
   NAND2_X1 i_0_4_314 (.A1(n_0_54), .A2(\Memory[3] [12]), .ZN(n_0_4_302));
   NAND2_X1 i_0_4_315 (.A1(n_0_53), .A2(\Memory[2] [12]), .ZN(n_0_4_303));
   NAND4_X1 i_0_4_316 (.A1(n_0_4_300), .A2(n_0_4_301), .A3(n_0_4_302), .A4(
      n_0_4_303), .ZN(n_0_4_304));
   INV_X1 i_0_4_317 (.A(n_0_4_304), .ZN(n_0_4_305));
   NAND2_X1 i_0_4_318 (.A1(n_0_67), .A2(\Memory[16] [12]), .ZN(n_0_4_306));
   NAND2_X1 i_0_4_319 (.A1(n_0_57), .A2(\Memory[6] [12]), .ZN(n_0_4_307));
   NAND2_X1 i_0_4_320 (.A1(n_0_56), .A2(\Memory[5] [12]), .ZN(n_0_4_308));
   NAND3_X1 i_0_4_321 (.A1(n_0_4_306), .A2(n_0_4_307), .A3(n_0_4_308), .ZN(
      n_0_4_309));
   NAND2_X1 i_0_4_322 (.A1(n_0_59), .A2(\Memory[8] [12]), .ZN(n_0_4_310));
   NAND2_X1 i_0_4_323 (.A1(n_0_52), .A2(\Memory[1] [12]), .ZN(n_0_4_311));
   NAND2_X1 i_0_4_324 (.A1(n_0_61), .A2(\Memory[10] [12]), .ZN(n_0_4_312));
   NAND3_X1 i_0_4_325 (.A1(n_0_4_310), .A2(n_0_4_311), .A3(n_0_4_312), .ZN(
      n_0_4_313));
   NOR2_X1 i_0_4_326 (.A1(n_0_4_309), .A2(n_0_4_313), .ZN(n_0_4_314));
   NAND2_X1 i_0_4_327 (.A1(n_0_65), .A2(\Memory[14] [12]), .ZN(n_0_4_315));
   NAND2_X1 i_0_4_328 (.A1(n_0_66), .A2(\Memory[15] [12]), .ZN(n_0_4_316));
   NAND2_X1 i_0_4_329 (.A1(n_0_51), .A2(\Memory[0] [12]), .ZN(n_0_4_317));
   NAND2_X1 i_0_4_330 (.A1(n_0_60), .A2(\Memory[9] [12]), .ZN(n_0_4_318));
   NAND4_X1 i_0_4_331 (.A1(n_0_4_315), .A2(n_0_4_316), .A3(n_0_4_317), .A4(
      n_0_4_318), .ZN(n_0_4_319));
   NAND2_X1 i_0_4_332 (.A1(n_0_64), .A2(\Memory[13] [12]), .ZN(n_0_4_320));
   NAND2_X1 i_0_4_333 (.A1(n_0_63), .A2(\Memory[12] [12]), .ZN(n_0_4_321));
   NAND2_X1 i_0_4_334 (.A1(n_0_62), .A2(\Memory[11] [12]), .ZN(n_0_4_322));
   NAND3_X1 i_0_4_335 (.A1(n_0_4_320), .A2(n_0_4_321), .A3(n_0_4_322), .ZN(
      n_0_4_323));
   NOR2_X1 i_0_4_336 (.A1(n_0_4_319), .A2(n_0_4_323), .ZN(n_0_4_324));
   NAND3_X1 i_0_4_337 (.A1(n_0_4_305), .A2(n_0_4_314), .A3(n_0_4_324), .ZN(
      dataOut2[12]));
   NAND2_X1 i_0_4_338 (.A1(n_0_55), .A2(\Memory[4] [13]), .ZN(n_0_4_325));
   NAND2_X1 i_0_4_339 (.A1(n_0_58), .A2(\Memory[7] [13]), .ZN(n_0_4_326));
   NAND2_X1 i_0_4_340 (.A1(n_0_54), .A2(\Memory[3] [13]), .ZN(n_0_4_327));
   NAND2_X1 i_0_4_341 (.A1(n_0_53), .A2(\Memory[2] [13]), .ZN(n_0_4_328));
   NAND4_X1 i_0_4_342 (.A1(n_0_4_325), .A2(n_0_4_326), .A3(n_0_4_327), .A4(
      n_0_4_328), .ZN(n_0_4_329));
   INV_X1 i_0_4_343 (.A(n_0_4_329), .ZN(n_0_4_330));
   NAND2_X1 i_0_4_344 (.A1(n_0_67), .A2(\Memory[16] [13]), .ZN(n_0_4_331));
   NAND2_X1 i_0_4_345 (.A1(n_0_57), .A2(\Memory[6] [13]), .ZN(n_0_4_332));
   NAND2_X1 i_0_4_346 (.A1(n_0_56), .A2(\Memory[5] [13]), .ZN(n_0_4_333));
   NAND3_X1 i_0_4_347 (.A1(n_0_4_331), .A2(n_0_4_332), .A3(n_0_4_333), .ZN(
      n_0_4_334));
   NAND2_X1 i_0_4_348 (.A1(n_0_59), .A2(\Memory[8] [13]), .ZN(n_0_4_335));
   NAND2_X1 i_0_4_349 (.A1(n_0_52), .A2(\Memory[1] [13]), .ZN(n_0_4_336));
   NAND2_X1 i_0_4_350 (.A1(n_0_61), .A2(\Memory[10] [13]), .ZN(n_0_4_337));
   NAND3_X1 i_0_4_351 (.A1(n_0_4_335), .A2(n_0_4_336), .A3(n_0_4_337), .ZN(
      n_0_4_338));
   NOR2_X1 i_0_4_352 (.A1(n_0_4_334), .A2(n_0_4_338), .ZN(n_0_4_339));
   NAND2_X1 i_0_4_353 (.A1(n_0_65), .A2(\Memory[14] [13]), .ZN(n_0_4_340));
   NAND2_X1 i_0_4_354 (.A1(n_0_66), .A2(\Memory[15] [13]), .ZN(n_0_4_341));
   NAND2_X1 i_0_4_355 (.A1(n_0_51), .A2(\Memory[0] [13]), .ZN(n_0_4_342));
   NAND2_X1 i_0_4_356 (.A1(n_0_60), .A2(\Memory[9] [13]), .ZN(n_0_4_343));
   NAND4_X1 i_0_4_357 (.A1(n_0_4_340), .A2(n_0_4_341), .A3(n_0_4_342), .A4(
      n_0_4_343), .ZN(n_0_4_344));
   NAND2_X1 i_0_4_358 (.A1(n_0_64), .A2(\Memory[13] [13]), .ZN(n_0_4_345));
   NAND2_X1 i_0_4_359 (.A1(n_0_63), .A2(\Memory[12] [13]), .ZN(n_0_4_346));
   NAND2_X1 i_0_4_360 (.A1(n_0_62), .A2(\Memory[11] [13]), .ZN(n_0_4_347));
   NAND3_X1 i_0_4_361 (.A1(n_0_4_345), .A2(n_0_4_346), .A3(n_0_4_347), .ZN(
      n_0_4_348));
   NOR2_X1 i_0_4_362 (.A1(n_0_4_344), .A2(n_0_4_348), .ZN(n_0_4_349));
   NAND3_X1 i_0_4_363 (.A1(n_0_4_330), .A2(n_0_4_339), .A3(n_0_4_349), .ZN(
      dataOut2[13]));
   NAND2_X1 i_0_4_364 (.A1(n_0_55), .A2(\Memory[4] [14]), .ZN(n_0_4_350));
   NAND2_X1 i_0_4_365 (.A1(n_0_58), .A2(\Memory[7] [14]), .ZN(n_0_4_351));
   NAND2_X1 i_0_4_366 (.A1(n_0_54), .A2(\Memory[3] [14]), .ZN(n_0_4_352));
   NAND2_X1 i_0_4_367 (.A1(n_0_53), .A2(\Memory[2] [14]), .ZN(n_0_4_353));
   NAND4_X1 i_0_4_368 (.A1(n_0_4_350), .A2(n_0_4_351), .A3(n_0_4_352), .A4(
      n_0_4_353), .ZN(n_0_4_354));
   INV_X1 i_0_4_369 (.A(n_0_4_354), .ZN(n_0_4_355));
   NAND2_X1 i_0_4_370 (.A1(n_0_67), .A2(\Memory[16] [14]), .ZN(n_0_4_356));
   NAND2_X1 i_0_4_371 (.A1(n_0_57), .A2(\Memory[6] [14]), .ZN(n_0_4_357));
   NAND2_X1 i_0_4_372 (.A1(n_0_56), .A2(\Memory[5] [14]), .ZN(n_0_4_358));
   NAND3_X1 i_0_4_373 (.A1(n_0_4_356), .A2(n_0_4_357), .A3(n_0_4_358), .ZN(
      n_0_4_359));
   NAND2_X1 i_0_4_374 (.A1(n_0_59), .A2(\Memory[8] [14]), .ZN(n_0_4_360));
   NAND2_X1 i_0_4_375 (.A1(n_0_52), .A2(\Memory[1] [14]), .ZN(n_0_4_361));
   NAND2_X1 i_0_4_376 (.A1(n_0_61), .A2(\Memory[10] [14]), .ZN(n_0_4_362));
   NAND3_X1 i_0_4_377 (.A1(n_0_4_360), .A2(n_0_4_361), .A3(n_0_4_362), .ZN(
      n_0_4_363));
   NOR2_X1 i_0_4_378 (.A1(n_0_4_359), .A2(n_0_4_363), .ZN(n_0_4_364));
   NAND2_X1 i_0_4_379 (.A1(n_0_65), .A2(\Memory[14] [14]), .ZN(n_0_4_365));
   NAND2_X1 i_0_4_380 (.A1(n_0_66), .A2(\Memory[15] [14]), .ZN(n_0_4_366));
   NAND2_X1 i_0_4_381 (.A1(n_0_51), .A2(\Memory[0] [14]), .ZN(n_0_4_367));
   NAND2_X1 i_0_4_382 (.A1(n_0_60), .A2(\Memory[9] [14]), .ZN(n_0_4_368));
   NAND4_X1 i_0_4_383 (.A1(n_0_4_365), .A2(n_0_4_366), .A3(n_0_4_367), .A4(
      n_0_4_368), .ZN(n_0_4_369));
   NAND2_X1 i_0_4_384 (.A1(n_0_64), .A2(\Memory[13] [14]), .ZN(n_0_4_370));
   NAND2_X1 i_0_4_385 (.A1(n_0_63), .A2(\Memory[12] [14]), .ZN(n_0_4_371));
   NAND2_X1 i_0_4_386 (.A1(n_0_62), .A2(\Memory[11] [14]), .ZN(n_0_4_372));
   NAND3_X1 i_0_4_387 (.A1(n_0_4_370), .A2(n_0_4_371), .A3(n_0_4_372), .ZN(
      n_0_4_373));
   NOR2_X1 i_0_4_388 (.A1(n_0_4_369), .A2(n_0_4_373), .ZN(n_0_4_374));
   NAND3_X1 i_0_4_389 (.A1(n_0_4_355), .A2(n_0_4_364), .A3(n_0_4_374), .ZN(
      dataOut2[14]));
   NAND2_X1 i_0_4_390 (.A1(n_0_55), .A2(\Memory[4] [15]), .ZN(n_0_4_375));
   NAND2_X1 i_0_4_391 (.A1(n_0_58), .A2(\Memory[7] [15]), .ZN(n_0_4_376));
   NAND2_X1 i_0_4_392 (.A1(n_0_54), .A2(\Memory[3] [15]), .ZN(n_0_4_377));
   NAND2_X1 i_0_4_393 (.A1(n_0_53), .A2(\Memory[2] [15]), .ZN(n_0_4_378));
   NAND4_X1 i_0_4_394 (.A1(n_0_4_375), .A2(n_0_4_376), .A3(n_0_4_377), .A4(
      n_0_4_378), .ZN(n_0_4_379));
   INV_X1 i_0_4_395 (.A(n_0_4_379), .ZN(n_0_4_380));
   NAND2_X1 i_0_4_396 (.A1(n_0_67), .A2(\Memory[16] [15]), .ZN(n_0_4_381));
   NAND2_X1 i_0_4_397 (.A1(n_0_57), .A2(\Memory[6] [15]), .ZN(n_0_4_382));
   NAND2_X1 i_0_4_398 (.A1(n_0_56), .A2(\Memory[5] [15]), .ZN(n_0_4_383));
   NAND3_X1 i_0_4_399 (.A1(n_0_4_381), .A2(n_0_4_382), .A3(n_0_4_383), .ZN(
      n_0_4_384));
   NAND2_X1 i_0_4_400 (.A1(n_0_59), .A2(\Memory[8] [15]), .ZN(n_0_4_385));
   NAND2_X1 i_0_4_401 (.A1(n_0_52), .A2(\Memory[1] [15]), .ZN(n_0_4_386));
   NAND2_X1 i_0_4_402 (.A1(n_0_61), .A2(\Memory[10] [15]), .ZN(n_0_4_387));
   NAND3_X1 i_0_4_403 (.A1(n_0_4_385), .A2(n_0_4_386), .A3(n_0_4_387), .ZN(
      n_0_4_388));
   NOR2_X1 i_0_4_404 (.A1(n_0_4_384), .A2(n_0_4_388), .ZN(n_0_4_389));
   NAND2_X1 i_0_4_405 (.A1(n_0_65), .A2(\Memory[14] [15]), .ZN(n_0_4_390));
   NAND2_X1 i_0_4_406 (.A1(n_0_66), .A2(\Memory[15] [15]), .ZN(n_0_4_391));
   NAND2_X1 i_0_4_407 (.A1(n_0_51), .A2(\Memory[0] [15]), .ZN(n_0_4_392));
   NAND2_X1 i_0_4_408 (.A1(n_0_60), .A2(\Memory[9] [15]), .ZN(n_0_4_393));
   NAND4_X1 i_0_4_409 (.A1(n_0_4_390), .A2(n_0_4_391), .A3(n_0_4_392), .A4(
      n_0_4_393), .ZN(n_0_4_394));
   NAND2_X1 i_0_4_410 (.A1(n_0_64), .A2(\Memory[13] [15]), .ZN(n_0_4_395));
   NAND2_X1 i_0_4_411 (.A1(n_0_63), .A2(\Memory[12] [15]), .ZN(n_0_4_396));
   NAND2_X1 i_0_4_412 (.A1(n_0_62), .A2(\Memory[11] [15]), .ZN(n_0_4_397));
   NAND3_X1 i_0_4_413 (.A1(n_0_4_395), .A2(n_0_4_396), .A3(n_0_4_397), .ZN(
      n_0_4_398));
   NOR2_X1 i_0_4_414 (.A1(n_0_4_394), .A2(n_0_4_398), .ZN(n_0_4_399));
   NAND3_X1 i_0_4_415 (.A1(n_0_4_380), .A2(n_0_4_389), .A3(n_0_4_399), .ZN(
      dataOut2[15]));
   NAND2_X1 i_0_4_416 (.A1(n_0_55), .A2(\Memory[4] [16]), .ZN(n_0_4_400));
   NAND2_X1 i_0_4_417 (.A1(n_0_58), .A2(\Memory[7] [16]), .ZN(n_0_4_401));
   NAND2_X1 i_0_4_418 (.A1(n_0_54), .A2(\Memory[3] [16]), .ZN(n_0_4_402));
   NAND2_X1 i_0_4_419 (.A1(n_0_53), .A2(\Memory[2] [16]), .ZN(n_0_4_403));
   NAND4_X1 i_0_4_420 (.A1(n_0_4_400), .A2(n_0_4_401), .A3(n_0_4_402), .A4(
      n_0_4_403), .ZN(n_0_4_404));
   INV_X1 i_0_4_421 (.A(n_0_4_404), .ZN(n_0_4_405));
   NAND2_X1 i_0_4_422 (.A1(n_0_67), .A2(\Memory[16] [16]), .ZN(n_0_4_406));
   NAND2_X1 i_0_4_423 (.A1(n_0_57), .A2(\Memory[6] [16]), .ZN(n_0_4_407));
   NAND2_X1 i_0_4_424 (.A1(n_0_56), .A2(\Memory[5] [16]), .ZN(n_0_4_408));
   NAND3_X1 i_0_4_425 (.A1(n_0_4_406), .A2(n_0_4_407), .A3(n_0_4_408), .ZN(
      n_0_4_409));
   NAND2_X1 i_0_4_426 (.A1(n_0_59), .A2(\Memory[8] [16]), .ZN(n_0_4_410));
   NAND2_X1 i_0_4_427 (.A1(n_0_52), .A2(\Memory[1] [16]), .ZN(n_0_4_411));
   NAND2_X1 i_0_4_428 (.A1(n_0_61), .A2(\Memory[10] [16]), .ZN(n_0_4_412));
   NAND3_X1 i_0_4_429 (.A1(n_0_4_410), .A2(n_0_4_411), .A3(n_0_4_412), .ZN(
      n_0_4_413));
   NOR2_X1 i_0_4_430 (.A1(n_0_4_409), .A2(n_0_4_413), .ZN(n_0_4_414));
   NAND2_X1 i_0_4_431 (.A1(n_0_65), .A2(\Memory[14] [16]), .ZN(n_0_4_415));
   NAND2_X1 i_0_4_432 (.A1(n_0_66), .A2(\Memory[15] [16]), .ZN(n_0_4_416));
   NAND2_X1 i_0_4_433 (.A1(n_0_51), .A2(\Memory[0] [16]), .ZN(n_0_4_417));
   NAND2_X1 i_0_4_434 (.A1(n_0_60), .A2(\Memory[9] [16]), .ZN(n_0_4_418));
   NAND4_X1 i_0_4_435 (.A1(n_0_4_415), .A2(n_0_4_416), .A3(n_0_4_417), .A4(
      n_0_4_418), .ZN(n_0_4_419));
   NAND2_X1 i_0_4_436 (.A1(n_0_64), .A2(\Memory[13] [16]), .ZN(n_0_4_420));
   NAND2_X1 i_0_4_437 (.A1(n_0_63), .A2(\Memory[12] [16]), .ZN(n_0_4_421));
   NAND2_X1 i_0_4_438 (.A1(n_0_62), .A2(\Memory[11] [16]), .ZN(n_0_4_422));
   NAND3_X1 i_0_4_439 (.A1(n_0_4_420), .A2(n_0_4_421), .A3(n_0_4_422), .ZN(
      n_0_4_423));
   NOR2_X1 i_0_4_440 (.A1(n_0_4_419), .A2(n_0_4_423), .ZN(n_0_4_424));
   NAND3_X1 i_0_4_441 (.A1(n_0_4_405), .A2(n_0_4_414), .A3(n_0_4_424), .ZN(
      dataOut2[16]));
   NAND2_X1 i_0_4_442 (.A1(n_0_55), .A2(\Memory[4] [17]), .ZN(n_0_4_425));
   NAND2_X1 i_0_4_443 (.A1(n_0_58), .A2(\Memory[7] [17]), .ZN(n_0_4_426));
   NAND2_X1 i_0_4_444 (.A1(n_0_54), .A2(\Memory[3] [17]), .ZN(n_0_4_427));
   NAND2_X1 i_0_4_445 (.A1(n_0_53), .A2(\Memory[2] [17]), .ZN(n_0_4_428));
   NAND4_X1 i_0_4_446 (.A1(n_0_4_425), .A2(n_0_4_426), .A3(n_0_4_427), .A4(
      n_0_4_428), .ZN(n_0_4_429));
   INV_X1 i_0_4_447 (.A(n_0_4_429), .ZN(n_0_4_430));
   NAND2_X1 i_0_4_448 (.A1(n_0_67), .A2(\Memory[16] [17]), .ZN(n_0_4_431));
   NAND2_X1 i_0_4_449 (.A1(n_0_57), .A2(\Memory[6] [17]), .ZN(n_0_4_432));
   NAND2_X1 i_0_4_450 (.A1(n_0_56), .A2(\Memory[5] [17]), .ZN(n_0_4_433));
   NAND3_X1 i_0_4_451 (.A1(n_0_4_431), .A2(n_0_4_432), .A3(n_0_4_433), .ZN(
      n_0_4_434));
   NAND2_X1 i_0_4_452 (.A1(n_0_59), .A2(\Memory[8] [17]), .ZN(n_0_4_435));
   NAND2_X1 i_0_4_453 (.A1(n_0_52), .A2(\Memory[1] [17]), .ZN(n_0_4_436));
   NAND2_X1 i_0_4_454 (.A1(n_0_61), .A2(\Memory[10] [17]), .ZN(n_0_4_437));
   NAND3_X1 i_0_4_455 (.A1(n_0_4_435), .A2(n_0_4_436), .A3(n_0_4_437), .ZN(
      n_0_4_438));
   NOR2_X1 i_0_4_456 (.A1(n_0_4_434), .A2(n_0_4_438), .ZN(n_0_4_439));
   NAND2_X1 i_0_4_457 (.A1(n_0_65), .A2(\Memory[14] [17]), .ZN(n_0_4_440));
   NAND2_X1 i_0_4_458 (.A1(n_0_66), .A2(\Memory[15] [17]), .ZN(n_0_4_441));
   NAND2_X1 i_0_4_459 (.A1(n_0_51), .A2(\Memory[0] [17]), .ZN(n_0_4_442));
   NAND2_X1 i_0_4_460 (.A1(n_0_60), .A2(\Memory[9] [17]), .ZN(n_0_4_443));
   NAND4_X1 i_0_4_461 (.A1(n_0_4_440), .A2(n_0_4_441), .A3(n_0_4_442), .A4(
      n_0_4_443), .ZN(n_0_4_444));
   NAND2_X1 i_0_4_462 (.A1(n_0_64), .A2(\Memory[13] [17]), .ZN(n_0_4_445));
   NAND2_X1 i_0_4_463 (.A1(n_0_63), .A2(\Memory[12] [17]), .ZN(n_0_4_446));
   NAND2_X1 i_0_4_464 (.A1(n_0_62), .A2(\Memory[11] [17]), .ZN(n_0_4_447));
   NAND3_X1 i_0_4_465 (.A1(n_0_4_445), .A2(n_0_4_446), .A3(n_0_4_447), .ZN(
      n_0_4_448));
   NOR2_X1 i_0_4_466 (.A1(n_0_4_444), .A2(n_0_4_448), .ZN(n_0_4_449));
   NAND3_X1 i_0_4_467 (.A1(n_0_4_430), .A2(n_0_4_439), .A3(n_0_4_449), .ZN(
      dataOut2[17]));
   NAND2_X1 i_0_4_468 (.A1(n_0_55), .A2(\Memory[4] [18]), .ZN(n_0_4_450));
   NAND2_X1 i_0_4_469 (.A1(n_0_58), .A2(\Memory[7] [18]), .ZN(n_0_4_451));
   NAND2_X1 i_0_4_470 (.A1(n_0_54), .A2(\Memory[3] [18]), .ZN(n_0_4_452));
   NAND2_X1 i_0_4_471 (.A1(n_0_53), .A2(\Memory[2] [18]), .ZN(n_0_4_453));
   NAND4_X1 i_0_4_472 (.A1(n_0_4_450), .A2(n_0_4_451), .A3(n_0_4_452), .A4(
      n_0_4_453), .ZN(n_0_4_454));
   INV_X1 i_0_4_473 (.A(n_0_4_454), .ZN(n_0_4_455));
   NAND2_X1 i_0_4_474 (.A1(n_0_67), .A2(\Memory[16] [18]), .ZN(n_0_4_456));
   NAND2_X1 i_0_4_475 (.A1(n_0_57), .A2(\Memory[6] [18]), .ZN(n_0_4_457));
   NAND2_X1 i_0_4_476 (.A1(n_0_56), .A2(\Memory[5] [18]), .ZN(n_0_4_458));
   NAND3_X1 i_0_4_477 (.A1(n_0_4_456), .A2(n_0_4_457), .A3(n_0_4_458), .ZN(
      n_0_4_459));
   NAND2_X1 i_0_4_478 (.A1(n_0_59), .A2(\Memory[8] [18]), .ZN(n_0_4_460));
   NAND2_X1 i_0_4_479 (.A1(n_0_52), .A2(\Memory[1] [18]), .ZN(n_0_4_461));
   NAND2_X1 i_0_4_480 (.A1(n_0_61), .A2(\Memory[10] [18]), .ZN(n_0_4_462));
   NAND3_X1 i_0_4_481 (.A1(n_0_4_460), .A2(n_0_4_461), .A3(n_0_4_462), .ZN(
      n_0_4_463));
   NOR2_X1 i_0_4_482 (.A1(n_0_4_459), .A2(n_0_4_463), .ZN(n_0_4_464));
   NAND2_X1 i_0_4_483 (.A1(n_0_65), .A2(\Memory[14] [18]), .ZN(n_0_4_465));
   NAND2_X1 i_0_4_484 (.A1(n_0_66), .A2(\Memory[15] [18]), .ZN(n_0_4_466));
   NAND2_X1 i_0_4_485 (.A1(n_0_51), .A2(\Memory[0] [18]), .ZN(n_0_4_467));
   NAND2_X1 i_0_4_486 (.A1(n_0_60), .A2(\Memory[9] [18]), .ZN(n_0_4_468));
   NAND4_X1 i_0_4_487 (.A1(n_0_4_465), .A2(n_0_4_466), .A3(n_0_4_467), .A4(
      n_0_4_468), .ZN(n_0_4_469));
   NAND2_X1 i_0_4_488 (.A1(n_0_64), .A2(\Memory[13] [18]), .ZN(n_0_4_470));
   NAND2_X1 i_0_4_489 (.A1(n_0_63), .A2(\Memory[12] [18]), .ZN(n_0_4_471));
   NAND2_X1 i_0_4_490 (.A1(n_0_62), .A2(\Memory[11] [18]), .ZN(n_0_4_472));
   NAND3_X1 i_0_4_491 (.A1(n_0_4_470), .A2(n_0_4_471), .A3(n_0_4_472), .ZN(
      n_0_4_473));
   NOR2_X1 i_0_4_492 (.A1(n_0_4_469), .A2(n_0_4_473), .ZN(n_0_4_474));
   NAND3_X1 i_0_4_493 (.A1(n_0_4_455), .A2(n_0_4_464), .A3(n_0_4_474), .ZN(
      dataOut2[18]));
   NAND2_X1 i_0_4_494 (.A1(n_0_55), .A2(\Memory[4] [19]), .ZN(n_0_4_475));
   NAND2_X1 i_0_4_495 (.A1(n_0_58), .A2(\Memory[7] [19]), .ZN(n_0_4_476));
   NAND2_X1 i_0_4_496 (.A1(n_0_54), .A2(\Memory[3] [19]), .ZN(n_0_4_477));
   NAND2_X1 i_0_4_497 (.A1(n_0_53), .A2(\Memory[2] [19]), .ZN(n_0_4_478));
   NAND4_X1 i_0_4_498 (.A1(n_0_4_475), .A2(n_0_4_476), .A3(n_0_4_477), .A4(
      n_0_4_478), .ZN(n_0_4_479));
   INV_X1 i_0_4_499 (.A(n_0_4_479), .ZN(n_0_4_480));
   NAND2_X1 i_0_4_500 (.A1(n_0_67), .A2(\Memory[16] [19]), .ZN(n_0_4_481));
   NAND2_X1 i_0_4_501 (.A1(n_0_57), .A2(\Memory[6] [19]), .ZN(n_0_4_482));
   NAND2_X1 i_0_4_502 (.A1(n_0_56), .A2(\Memory[5] [19]), .ZN(n_0_4_483));
   NAND3_X1 i_0_4_503 (.A1(n_0_4_481), .A2(n_0_4_482), .A3(n_0_4_483), .ZN(
      n_0_4_484));
   NAND2_X1 i_0_4_504 (.A1(n_0_59), .A2(\Memory[8] [19]), .ZN(n_0_4_485));
   NAND2_X1 i_0_4_505 (.A1(n_0_52), .A2(\Memory[1] [19]), .ZN(n_0_4_486));
   NAND2_X1 i_0_4_506 (.A1(n_0_61), .A2(\Memory[10] [19]), .ZN(n_0_4_487));
   NAND3_X1 i_0_4_507 (.A1(n_0_4_485), .A2(n_0_4_486), .A3(n_0_4_487), .ZN(
      n_0_4_488));
   NOR2_X1 i_0_4_508 (.A1(n_0_4_484), .A2(n_0_4_488), .ZN(n_0_4_489));
   NAND2_X1 i_0_4_509 (.A1(n_0_65), .A2(\Memory[14] [19]), .ZN(n_0_4_490));
   NAND2_X1 i_0_4_510 (.A1(n_0_66), .A2(\Memory[15] [19]), .ZN(n_0_4_491));
   NAND2_X1 i_0_4_511 (.A1(n_0_51), .A2(\Memory[0] [19]), .ZN(n_0_4_492));
   NAND2_X1 i_0_4_512 (.A1(n_0_60), .A2(\Memory[9] [19]), .ZN(n_0_4_493));
   NAND4_X1 i_0_4_513 (.A1(n_0_4_490), .A2(n_0_4_491), .A3(n_0_4_492), .A4(
      n_0_4_493), .ZN(n_0_4_494));
   NAND2_X1 i_0_4_514 (.A1(n_0_64), .A2(\Memory[13] [19]), .ZN(n_0_4_495));
   NAND2_X1 i_0_4_515 (.A1(n_0_63), .A2(\Memory[12] [19]), .ZN(n_0_4_496));
   NAND2_X1 i_0_4_516 (.A1(n_0_62), .A2(\Memory[11] [19]), .ZN(n_0_4_497));
   NAND3_X1 i_0_4_517 (.A1(n_0_4_495), .A2(n_0_4_496), .A3(n_0_4_497), .ZN(
      n_0_4_498));
   NOR2_X1 i_0_4_518 (.A1(n_0_4_494), .A2(n_0_4_498), .ZN(n_0_4_499));
   NAND3_X1 i_0_4_519 (.A1(n_0_4_480), .A2(n_0_4_489), .A3(n_0_4_499), .ZN(
      dataOut2[19]));
   NAND2_X1 i_0_4_520 (.A1(n_0_55), .A2(\Memory[4] [20]), .ZN(n_0_4_500));
   NAND2_X1 i_0_4_521 (.A1(n_0_58), .A2(\Memory[7] [20]), .ZN(n_0_4_501));
   NAND2_X1 i_0_4_522 (.A1(n_0_54), .A2(\Memory[3] [20]), .ZN(n_0_4_502));
   NAND2_X1 i_0_4_523 (.A1(n_0_53), .A2(\Memory[2] [20]), .ZN(n_0_4_503));
   NAND4_X1 i_0_4_524 (.A1(n_0_4_500), .A2(n_0_4_501), .A3(n_0_4_502), .A4(
      n_0_4_503), .ZN(n_0_4_504));
   INV_X1 i_0_4_525 (.A(n_0_4_504), .ZN(n_0_4_505));
   NAND2_X1 i_0_4_526 (.A1(n_0_67), .A2(\Memory[16] [20]), .ZN(n_0_4_506));
   NAND2_X1 i_0_4_527 (.A1(n_0_57), .A2(\Memory[6] [20]), .ZN(n_0_4_507));
   NAND2_X1 i_0_4_528 (.A1(n_0_56), .A2(\Memory[5] [20]), .ZN(n_0_4_508));
   NAND3_X1 i_0_4_529 (.A1(n_0_4_506), .A2(n_0_4_507), .A3(n_0_4_508), .ZN(
      n_0_4_509));
   NAND2_X1 i_0_4_530 (.A1(n_0_59), .A2(\Memory[8] [20]), .ZN(n_0_4_510));
   NAND2_X1 i_0_4_531 (.A1(n_0_52), .A2(\Memory[1] [20]), .ZN(n_0_4_511));
   NAND2_X1 i_0_4_532 (.A1(n_0_61), .A2(\Memory[10] [20]), .ZN(n_0_4_512));
   NAND3_X1 i_0_4_533 (.A1(n_0_4_510), .A2(n_0_4_511), .A3(n_0_4_512), .ZN(
      n_0_4_513));
   NOR2_X1 i_0_4_534 (.A1(n_0_4_509), .A2(n_0_4_513), .ZN(n_0_4_514));
   NAND2_X1 i_0_4_535 (.A1(n_0_65), .A2(\Memory[14] [20]), .ZN(n_0_4_515));
   NAND2_X1 i_0_4_536 (.A1(n_0_66), .A2(\Memory[15] [20]), .ZN(n_0_4_516));
   NAND2_X1 i_0_4_537 (.A1(n_0_51), .A2(\Memory[0] [20]), .ZN(n_0_4_517));
   NAND2_X1 i_0_4_538 (.A1(n_0_60), .A2(\Memory[9] [20]), .ZN(n_0_4_518));
   NAND4_X1 i_0_4_539 (.A1(n_0_4_515), .A2(n_0_4_516), .A3(n_0_4_517), .A4(
      n_0_4_518), .ZN(n_0_4_519));
   NAND2_X1 i_0_4_540 (.A1(n_0_64), .A2(\Memory[13] [20]), .ZN(n_0_4_520));
   NAND2_X1 i_0_4_541 (.A1(n_0_63), .A2(\Memory[12] [20]), .ZN(n_0_4_521));
   NAND2_X1 i_0_4_542 (.A1(n_0_62), .A2(\Memory[11] [20]), .ZN(n_0_4_522));
   NAND3_X1 i_0_4_543 (.A1(n_0_4_520), .A2(n_0_4_521), .A3(n_0_4_522), .ZN(
      n_0_4_523));
   NOR2_X1 i_0_4_544 (.A1(n_0_4_519), .A2(n_0_4_523), .ZN(n_0_4_524));
   NAND3_X1 i_0_4_545 (.A1(n_0_4_505), .A2(n_0_4_514), .A3(n_0_4_524), .ZN(
      dataOut2[20]));
   NAND2_X1 i_0_4_546 (.A1(n_0_55), .A2(\Memory[4] [21]), .ZN(n_0_4_525));
   NAND2_X1 i_0_4_547 (.A1(n_0_58), .A2(\Memory[7] [21]), .ZN(n_0_4_526));
   NAND2_X1 i_0_4_548 (.A1(n_0_54), .A2(\Memory[3] [21]), .ZN(n_0_4_527));
   NAND2_X1 i_0_4_549 (.A1(n_0_53), .A2(\Memory[2] [21]), .ZN(n_0_4_528));
   NAND4_X1 i_0_4_550 (.A1(n_0_4_525), .A2(n_0_4_526), .A3(n_0_4_527), .A4(
      n_0_4_528), .ZN(n_0_4_529));
   INV_X1 i_0_4_551 (.A(n_0_4_529), .ZN(n_0_4_530));
   NAND2_X1 i_0_4_552 (.A1(n_0_67), .A2(\Memory[16] [21]), .ZN(n_0_4_531));
   NAND2_X1 i_0_4_553 (.A1(n_0_57), .A2(\Memory[6] [21]), .ZN(n_0_4_532));
   NAND2_X1 i_0_4_554 (.A1(n_0_56), .A2(\Memory[5] [21]), .ZN(n_0_4_533));
   NAND3_X1 i_0_4_555 (.A1(n_0_4_531), .A2(n_0_4_532), .A3(n_0_4_533), .ZN(
      n_0_4_534));
   NAND2_X1 i_0_4_556 (.A1(n_0_59), .A2(\Memory[8] [21]), .ZN(n_0_4_535));
   NAND2_X1 i_0_4_557 (.A1(n_0_52), .A2(\Memory[1] [21]), .ZN(n_0_4_536));
   NAND2_X1 i_0_4_558 (.A1(n_0_61), .A2(\Memory[10] [21]), .ZN(n_0_4_537));
   NAND3_X1 i_0_4_559 (.A1(n_0_4_535), .A2(n_0_4_536), .A3(n_0_4_537), .ZN(
      n_0_4_538));
   NOR2_X1 i_0_4_560 (.A1(n_0_4_534), .A2(n_0_4_538), .ZN(n_0_4_539));
   NAND2_X1 i_0_4_561 (.A1(n_0_65), .A2(\Memory[14] [21]), .ZN(n_0_4_540));
   NAND2_X1 i_0_4_562 (.A1(n_0_66), .A2(\Memory[15] [21]), .ZN(n_0_4_541));
   NAND2_X1 i_0_4_563 (.A1(n_0_51), .A2(\Memory[0] [21]), .ZN(n_0_4_542));
   NAND2_X1 i_0_4_564 (.A1(n_0_60), .A2(\Memory[9] [21]), .ZN(n_0_4_543));
   NAND4_X1 i_0_4_565 (.A1(n_0_4_540), .A2(n_0_4_541), .A3(n_0_4_542), .A4(
      n_0_4_543), .ZN(n_0_4_544));
   NAND2_X1 i_0_4_566 (.A1(n_0_64), .A2(\Memory[13] [21]), .ZN(n_0_4_545));
   NAND2_X1 i_0_4_567 (.A1(n_0_63), .A2(\Memory[12] [21]), .ZN(n_0_4_546));
   NAND2_X1 i_0_4_568 (.A1(n_0_62), .A2(\Memory[11] [21]), .ZN(n_0_4_547));
   NAND3_X1 i_0_4_569 (.A1(n_0_4_545), .A2(n_0_4_546), .A3(n_0_4_547), .ZN(
      n_0_4_548));
   NOR2_X1 i_0_4_570 (.A1(n_0_4_544), .A2(n_0_4_548), .ZN(n_0_4_549));
   NAND3_X1 i_0_4_571 (.A1(n_0_4_530), .A2(n_0_4_539), .A3(n_0_4_549), .ZN(
      dataOut2[21]));
   NAND2_X1 i_0_4_572 (.A1(n_0_55), .A2(\Memory[4] [22]), .ZN(n_0_4_550));
   NAND2_X1 i_0_4_573 (.A1(n_0_58), .A2(\Memory[7] [22]), .ZN(n_0_4_551));
   NAND2_X1 i_0_4_574 (.A1(n_0_54), .A2(\Memory[3] [22]), .ZN(n_0_4_552));
   NAND2_X1 i_0_4_575 (.A1(n_0_53), .A2(\Memory[2] [22]), .ZN(n_0_4_553));
   NAND4_X1 i_0_4_576 (.A1(n_0_4_550), .A2(n_0_4_551), .A3(n_0_4_552), .A4(
      n_0_4_553), .ZN(n_0_4_554));
   INV_X1 i_0_4_577 (.A(n_0_4_554), .ZN(n_0_4_555));
   NAND2_X1 i_0_4_578 (.A1(n_0_67), .A2(\Memory[16] [22]), .ZN(n_0_4_556));
   NAND2_X1 i_0_4_579 (.A1(n_0_57), .A2(\Memory[6] [22]), .ZN(n_0_4_557));
   NAND2_X1 i_0_4_580 (.A1(n_0_56), .A2(\Memory[5] [22]), .ZN(n_0_4_558));
   NAND3_X1 i_0_4_581 (.A1(n_0_4_556), .A2(n_0_4_557), .A3(n_0_4_558), .ZN(
      n_0_4_559));
   NAND2_X1 i_0_4_582 (.A1(n_0_59), .A2(\Memory[8] [22]), .ZN(n_0_4_560));
   NAND2_X1 i_0_4_583 (.A1(n_0_52), .A2(\Memory[1] [22]), .ZN(n_0_4_561));
   NAND2_X1 i_0_4_584 (.A1(n_0_61), .A2(\Memory[10] [22]), .ZN(n_0_4_562));
   NAND3_X1 i_0_4_585 (.A1(n_0_4_560), .A2(n_0_4_561), .A3(n_0_4_562), .ZN(
      n_0_4_563));
   NOR2_X1 i_0_4_586 (.A1(n_0_4_559), .A2(n_0_4_563), .ZN(n_0_4_564));
   NAND2_X1 i_0_4_587 (.A1(n_0_65), .A2(\Memory[14] [22]), .ZN(n_0_4_565));
   NAND2_X1 i_0_4_588 (.A1(n_0_66), .A2(\Memory[15] [22]), .ZN(n_0_4_566));
   NAND2_X1 i_0_4_589 (.A1(n_0_51), .A2(\Memory[0] [22]), .ZN(n_0_4_567));
   NAND2_X1 i_0_4_590 (.A1(n_0_60), .A2(\Memory[9] [22]), .ZN(n_0_4_568));
   NAND4_X1 i_0_4_591 (.A1(n_0_4_565), .A2(n_0_4_566), .A3(n_0_4_567), .A4(
      n_0_4_568), .ZN(n_0_4_569));
   NAND2_X1 i_0_4_592 (.A1(n_0_64), .A2(\Memory[13] [22]), .ZN(n_0_4_570));
   NAND2_X1 i_0_4_593 (.A1(n_0_63), .A2(\Memory[12] [22]), .ZN(n_0_4_571));
   NAND2_X1 i_0_4_594 (.A1(n_0_62), .A2(\Memory[11] [22]), .ZN(n_0_4_572));
   NAND3_X1 i_0_4_595 (.A1(n_0_4_570), .A2(n_0_4_571), .A3(n_0_4_572), .ZN(
      n_0_4_573));
   NOR2_X1 i_0_4_596 (.A1(n_0_4_569), .A2(n_0_4_573), .ZN(n_0_4_574));
   NAND3_X1 i_0_4_597 (.A1(n_0_4_555), .A2(n_0_4_564), .A3(n_0_4_574), .ZN(
      dataOut2[22]));
   NAND2_X1 i_0_4_598 (.A1(n_0_55), .A2(\Memory[4] [23]), .ZN(n_0_4_575));
   NAND2_X1 i_0_4_599 (.A1(n_0_58), .A2(\Memory[7] [23]), .ZN(n_0_4_576));
   NAND2_X1 i_0_4_600 (.A1(n_0_54), .A2(\Memory[3] [23]), .ZN(n_0_4_577));
   NAND2_X1 i_0_4_601 (.A1(n_0_53), .A2(\Memory[2] [23]), .ZN(n_0_4_578));
   NAND4_X1 i_0_4_602 (.A1(n_0_4_575), .A2(n_0_4_576), .A3(n_0_4_577), .A4(
      n_0_4_578), .ZN(n_0_4_579));
   INV_X1 i_0_4_603 (.A(n_0_4_579), .ZN(n_0_4_580));
   NAND2_X1 i_0_4_604 (.A1(n_0_67), .A2(\Memory[16] [23]), .ZN(n_0_4_581));
   NAND2_X1 i_0_4_605 (.A1(n_0_57), .A2(\Memory[6] [23]), .ZN(n_0_4_582));
   NAND2_X1 i_0_4_606 (.A1(n_0_56), .A2(\Memory[5] [23]), .ZN(n_0_4_583));
   NAND3_X1 i_0_4_607 (.A1(n_0_4_581), .A2(n_0_4_582), .A3(n_0_4_583), .ZN(
      n_0_4_584));
   NAND2_X1 i_0_4_608 (.A1(n_0_59), .A2(\Memory[8] [23]), .ZN(n_0_4_585));
   NAND2_X1 i_0_4_609 (.A1(n_0_52), .A2(\Memory[1] [23]), .ZN(n_0_4_586));
   NAND2_X1 i_0_4_610 (.A1(n_0_61), .A2(\Memory[10] [23]), .ZN(n_0_4_587));
   NAND3_X1 i_0_4_611 (.A1(n_0_4_585), .A2(n_0_4_586), .A3(n_0_4_587), .ZN(
      n_0_4_588));
   NOR2_X1 i_0_4_612 (.A1(n_0_4_584), .A2(n_0_4_588), .ZN(n_0_4_589));
   NAND2_X1 i_0_4_613 (.A1(n_0_65), .A2(\Memory[14] [23]), .ZN(n_0_4_590));
   NAND2_X1 i_0_4_614 (.A1(n_0_66), .A2(\Memory[15] [23]), .ZN(n_0_4_591));
   NAND2_X1 i_0_4_615 (.A1(n_0_51), .A2(\Memory[0] [23]), .ZN(n_0_4_592));
   NAND2_X1 i_0_4_616 (.A1(n_0_60), .A2(\Memory[9] [23]), .ZN(n_0_4_593));
   NAND4_X1 i_0_4_617 (.A1(n_0_4_590), .A2(n_0_4_591), .A3(n_0_4_592), .A4(
      n_0_4_593), .ZN(n_0_4_594));
   NAND2_X1 i_0_4_618 (.A1(n_0_64), .A2(\Memory[13] [23]), .ZN(n_0_4_595));
   NAND2_X1 i_0_4_619 (.A1(n_0_63), .A2(\Memory[12] [23]), .ZN(n_0_4_596));
   NAND2_X1 i_0_4_620 (.A1(n_0_62), .A2(\Memory[11] [23]), .ZN(n_0_4_597));
   NAND3_X1 i_0_4_621 (.A1(n_0_4_595), .A2(n_0_4_596), .A3(n_0_4_597), .ZN(
      n_0_4_598));
   NOR2_X1 i_0_4_622 (.A1(n_0_4_594), .A2(n_0_4_598), .ZN(n_0_4_599));
   NAND3_X1 i_0_4_623 (.A1(n_0_4_580), .A2(n_0_4_589), .A3(n_0_4_599), .ZN(
      dataOut2[23]));
   NAND2_X1 i_0_4_624 (.A1(n_0_55), .A2(\Memory[4] [24]), .ZN(n_0_4_600));
   NAND2_X1 i_0_4_625 (.A1(n_0_58), .A2(\Memory[7] [24]), .ZN(n_0_4_601));
   NAND2_X1 i_0_4_626 (.A1(n_0_54), .A2(\Memory[3] [24]), .ZN(n_0_4_602));
   NAND2_X1 i_0_4_627 (.A1(n_0_53), .A2(\Memory[2] [24]), .ZN(n_0_4_603));
   NAND4_X1 i_0_4_628 (.A1(n_0_4_600), .A2(n_0_4_601), .A3(n_0_4_602), .A4(
      n_0_4_603), .ZN(n_0_4_604));
   INV_X1 i_0_4_629 (.A(n_0_4_604), .ZN(n_0_4_605));
   NAND2_X1 i_0_4_630 (.A1(n_0_67), .A2(\Memory[16] [24]), .ZN(n_0_4_606));
   NAND2_X1 i_0_4_631 (.A1(n_0_57), .A2(\Memory[6] [24]), .ZN(n_0_4_607));
   NAND2_X1 i_0_4_632 (.A1(n_0_56), .A2(\Memory[5] [24]), .ZN(n_0_4_608));
   NAND3_X1 i_0_4_633 (.A1(n_0_4_606), .A2(n_0_4_607), .A3(n_0_4_608), .ZN(
      n_0_4_609));
   NAND2_X1 i_0_4_634 (.A1(n_0_59), .A2(\Memory[8] [24]), .ZN(n_0_4_610));
   NAND2_X1 i_0_4_635 (.A1(n_0_52), .A2(\Memory[1] [24]), .ZN(n_0_4_611));
   NAND2_X1 i_0_4_636 (.A1(n_0_61), .A2(\Memory[10] [24]), .ZN(n_0_4_612));
   NAND3_X1 i_0_4_637 (.A1(n_0_4_610), .A2(n_0_4_611), .A3(n_0_4_612), .ZN(
      n_0_4_613));
   NOR2_X1 i_0_4_638 (.A1(n_0_4_609), .A2(n_0_4_613), .ZN(n_0_4_614));
   NAND2_X1 i_0_4_639 (.A1(n_0_65), .A2(\Memory[14] [24]), .ZN(n_0_4_615));
   NAND2_X1 i_0_4_640 (.A1(n_0_66), .A2(\Memory[15] [24]), .ZN(n_0_4_616));
   NAND2_X1 i_0_4_641 (.A1(n_0_51), .A2(\Memory[0] [24]), .ZN(n_0_4_617));
   NAND2_X1 i_0_4_642 (.A1(n_0_60), .A2(\Memory[9] [24]), .ZN(n_0_4_618));
   NAND4_X1 i_0_4_643 (.A1(n_0_4_615), .A2(n_0_4_616), .A3(n_0_4_617), .A4(
      n_0_4_618), .ZN(n_0_4_619));
   NAND2_X1 i_0_4_644 (.A1(n_0_64), .A2(\Memory[13] [24]), .ZN(n_0_4_620));
   NAND2_X1 i_0_4_645 (.A1(n_0_63), .A2(\Memory[12] [24]), .ZN(n_0_4_621));
   NAND2_X1 i_0_4_646 (.A1(n_0_62), .A2(\Memory[11] [24]), .ZN(n_0_4_622));
   NAND3_X1 i_0_4_647 (.A1(n_0_4_620), .A2(n_0_4_621), .A3(n_0_4_622), .ZN(
      n_0_4_623));
   NOR2_X1 i_0_4_648 (.A1(n_0_4_619), .A2(n_0_4_623), .ZN(n_0_4_624));
   NAND3_X1 i_0_4_649 (.A1(n_0_4_605), .A2(n_0_4_614), .A3(n_0_4_624), .ZN(
      dataOut2[24]));
   NAND2_X1 i_0_4_650 (.A1(n_0_55), .A2(\Memory[4] [25]), .ZN(n_0_4_625));
   NAND2_X1 i_0_4_651 (.A1(n_0_58), .A2(\Memory[7] [25]), .ZN(n_0_4_626));
   NAND2_X1 i_0_4_652 (.A1(n_0_54), .A2(\Memory[3] [25]), .ZN(n_0_4_627));
   NAND2_X1 i_0_4_653 (.A1(n_0_53), .A2(\Memory[2] [25]), .ZN(n_0_4_628));
   NAND4_X1 i_0_4_654 (.A1(n_0_4_625), .A2(n_0_4_626), .A3(n_0_4_627), .A4(
      n_0_4_628), .ZN(n_0_4_629));
   INV_X1 i_0_4_655 (.A(n_0_4_629), .ZN(n_0_4_630));
   NAND2_X1 i_0_4_656 (.A1(n_0_67), .A2(\Memory[16] [25]), .ZN(n_0_4_631));
   NAND2_X1 i_0_4_657 (.A1(n_0_57), .A2(\Memory[6] [25]), .ZN(n_0_4_632));
   NAND2_X1 i_0_4_658 (.A1(n_0_56), .A2(\Memory[5] [25]), .ZN(n_0_4_633));
   NAND3_X1 i_0_4_659 (.A1(n_0_4_631), .A2(n_0_4_632), .A3(n_0_4_633), .ZN(
      n_0_4_634));
   NAND2_X1 i_0_4_660 (.A1(n_0_59), .A2(\Memory[8] [25]), .ZN(n_0_4_635));
   NAND2_X1 i_0_4_661 (.A1(n_0_52), .A2(\Memory[1] [25]), .ZN(n_0_4_636));
   NAND2_X1 i_0_4_662 (.A1(n_0_61), .A2(\Memory[10] [25]), .ZN(n_0_4_637));
   NAND3_X1 i_0_4_663 (.A1(n_0_4_635), .A2(n_0_4_636), .A3(n_0_4_637), .ZN(
      n_0_4_638));
   NOR2_X1 i_0_4_664 (.A1(n_0_4_634), .A2(n_0_4_638), .ZN(n_0_4_639));
   NAND2_X1 i_0_4_665 (.A1(n_0_65), .A2(\Memory[14] [25]), .ZN(n_0_4_640));
   NAND2_X1 i_0_4_666 (.A1(n_0_66), .A2(\Memory[15] [25]), .ZN(n_0_4_641));
   NAND2_X1 i_0_4_667 (.A1(n_0_51), .A2(\Memory[0] [25]), .ZN(n_0_4_642));
   NAND2_X1 i_0_4_668 (.A1(n_0_60), .A2(\Memory[9] [25]), .ZN(n_0_4_643));
   NAND4_X1 i_0_4_669 (.A1(n_0_4_640), .A2(n_0_4_641), .A3(n_0_4_642), .A4(
      n_0_4_643), .ZN(n_0_4_644));
   NAND2_X1 i_0_4_670 (.A1(n_0_64), .A2(\Memory[13] [25]), .ZN(n_0_4_645));
   NAND2_X1 i_0_4_671 (.A1(n_0_63), .A2(\Memory[12] [25]), .ZN(n_0_4_646));
   NAND2_X1 i_0_4_672 (.A1(n_0_62), .A2(\Memory[11] [25]), .ZN(n_0_4_647));
   NAND3_X1 i_0_4_673 (.A1(n_0_4_645), .A2(n_0_4_646), .A3(n_0_4_647), .ZN(
      n_0_4_648));
   NOR2_X1 i_0_4_674 (.A1(n_0_4_644), .A2(n_0_4_648), .ZN(n_0_4_649));
   NAND3_X1 i_0_4_675 (.A1(n_0_4_630), .A2(n_0_4_639), .A3(n_0_4_649), .ZN(
      dataOut2[25]));
   NAND2_X1 i_0_4_676 (.A1(n_0_55), .A2(\Memory[4] [26]), .ZN(n_0_4_650));
   NAND2_X1 i_0_4_677 (.A1(n_0_58), .A2(\Memory[7] [26]), .ZN(n_0_4_651));
   NAND2_X1 i_0_4_678 (.A1(n_0_54), .A2(\Memory[3] [26]), .ZN(n_0_4_652));
   NAND2_X1 i_0_4_679 (.A1(n_0_53), .A2(\Memory[2] [26]), .ZN(n_0_4_653));
   NAND4_X1 i_0_4_680 (.A1(n_0_4_650), .A2(n_0_4_651), .A3(n_0_4_652), .A4(
      n_0_4_653), .ZN(n_0_4_654));
   INV_X1 i_0_4_681 (.A(n_0_4_654), .ZN(n_0_4_655));
   NAND2_X1 i_0_4_682 (.A1(n_0_67), .A2(\Memory[16] [26]), .ZN(n_0_4_656));
   NAND2_X1 i_0_4_683 (.A1(n_0_57), .A2(\Memory[6] [26]), .ZN(n_0_4_657));
   NAND2_X1 i_0_4_684 (.A1(n_0_56), .A2(\Memory[5] [26]), .ZN(n_0_4_658));
   NAND3_X1 i_0_4_685 (.A1(n_0_4_656), .A2(n_0_4_657), .A3(n_0_4_658), .ZN(
      n_0_4_659));
   NAND2_X1 i_0_4_686 (.A1(n_0_59), .A2(\Memory[8] [26]), .ZN(n_0_4_660));
   NAND2_X1 i_0_4_687 (.A1(n_0_52), .A2(\Memory[1] [26]), .ZN(n_0_4_661));
   NAND2_X1 i_0_4_688 (.A1(n_0_61), .A2(\Memory[10] [26]), .ZN(n_0_4_662));
   NAND3_X1 i_0_4_689 (.A1(n_0_4_660), .A2(n_0_4_661), .A3(n_0_4_662), .ZN(
      n_0_4_663));
   NOR2_X1 i_0_4_690 (.A1(n_0_4_659), .A2(n_0_4_663), .ZN(n_0_4_664));
   NAND2_X1 i_0_4_691 (.A1(n_0_65), .A2(\Memory[14] [26]), .ZN(n_0_4_665));
   NAND2_X1 i_0_4_692 (.A1(n_0_66), .A2(\Memory[15] [26]), .ZN(n_0_4_666));
   NAND2_X1 i_0_4_693 (.A1(n_0_51), .A2(\Memory[0] [26]), .ZN(n_0_4_667));
   NAND2_X1 i_0_4_694 (.A1(n_0_60), .A2(\Memory[9] [26]), .ZN(n_0_4_668));
   NAND4_X1 i_0_4_695 (.A1(n_0_4_665), .A2(n_0_4_666), .A3(n_0_4_667), .A4(
      n_0_4_668), .ZN(n_0_4_669));
   NAND2_X1 i_0_4_696 (.A1(n_0_64), .A2(\Memory[13] [26]), .ZN(n_0_4_670));
   NAND2_X1 i_0_4_697 (.A1(n_0_63), .A2(\Memory[12] [26]), .ZN(n_0_4_671));
   NAND2_X1 i_0_4_698 (.A1(n_0_62), .A2(\Memory[11] [26]), .ZN(n_0_4_672));
   NAND3_X1 i_0_4_699 (.A1(n_0_4_670), .A2(n_0_4_671), .A3(n_0_4_672), .ZN(
      n_0_4_673));
   NOR2_X1 i_0_4_700 (.A1(n_0_4_669), .A2(n_0_4_673), .ZN(n_0_4_674));
   NAND3_X1 i_0_4_701 (.A1(n_0_4_655), .A2(n_0_4_664), .A3(n_0_4_674), .ZN(
      dataOut2[26]));
   NAND2_X1 i_0_4_702 (.A1(n_0_55), .A2(\Memory[4] [27]), .ZN(n_0_4_675));
   NAND2_X1 i_0_4_703 (.A1(n_0_58), .A2(\Memory[7] [27]), .ZN(n_0_4_676));
   NAND2_X1 i_0_4_704 (.A1(n_0_54), .A2(\Memory[3] [27]), .ZN(n_0_4_677));
   NAND2_X1 i_0_4_705 (.A1(n_0_53), .A2(\Memory[2] [27]), .ZN(n_0_4_678));
   NAND4_X1 i_0_4_706 (.A1(n_0_4_675), .A2(n_0_4_676), .A3(n_0_4_677), .A4(
      n_0_4_678), .ZN(n_0_4_679));
   INV_X1 i_0_4_707 (.A(n_0_4_679), .ZN(n_0_4_680));
   NAND2_X1 i_0_4_708 (.A1(n_0_67), .A2(\Memory[16] [27]), .ZN(n_0_4_681));
   NAND2_X1 i_0_4_709 (.A1(n_0_57), .A2(\Memory[6] [27]), .ZN(n_0_4_682));
   NAND2_X1 i_0_4_710 (.A1(n_0_56), .A2(\Memory[5] [27]), .ZN(n_0_4_683));
   NAND3_X1 i_0_4_711 (.A1(n_0_4_681), .A2(n_0_4_682), .A3(n_0_4_683), .ZN(
      n_0_4_684));
   NAND2_X1 i_0_4_712 (.A1(n_0_59), .A2(\Memory[8] [27]), .ZN(n_0_4_685));
   NAND2_X1 i_0_4_713 (.A1(n_0_52), .A2(\Memory[1] [27]), .ZN(n_0_4_686));
   NAND2_X1 i_0_4_714 (.A1(n_0_61), .A2(\Memory[10] [27]), .ZN(n_0_4_687));
   NAND3_X1 i_0_4_715 (.A1(n_0_4_685), .A2(n_0_4_686), .A3(n_0_4_687), .ZN(
      n_0_4_688));
   NOR2_X1 i_0_4_716 (.A1(n_0_4_684), .A2(n_0_4_688), .ZN(n_0_4_689));
   NAND2_X1 i_0_4_717 (.A1(n_0_65), .A2(\Memory[14] [27]), .ZN(n_0_4_690));
   NAND2_X1 i_0_4_718 (.A1(n_0_66), .A2(\Memory[15] [27]), .ZN(n_0_4_691));
   NAND2_X1 i_0_4_719 (.A1(n_0_51), .A2(\Memory[0] [27]), .ZN(n_0_4_692));
   NAND2_X1 i_0_4_720 (.A1(n_0_60), .A2(\Memory[9] [27]), .ZN(n_0_4_693));
   NAND4_X1 i_0_4_721 (.A1(n_0_4_690), .A2(n_0_4_691), .A3(n_0_4_692), .A4(
      n_0_4_693), .ZN(n_0_4_694));
   NAND2_X1 i_0_4_722 (.A1(n_0_64), .A2(\Memory[13] [27]), .ZN(n_0_4_695));
   NAND2_X1 i_0_4_723 (.A1(n_0_63), .A2(\Memory[12] [27]), .ZN(n_0_4_696));
   NAND2_X1 i_0_4_724 (.A1(n_0_62), .A2(\Memory[11] [27]), .ZN(n_0_4_697));
   NAND3_X1 i_0_4_725 (.A1(n_0_4_695), .A2(n_0_4_696), .A3(n_0_4_697), .ZN(
      n_0_4_698));
   NOR2_X1 i_0_4_726 (.A1(n_0_4_694), .A2(n_0_4_698), .ZN(n_0_4_699));
   NAND3_X1 i_0_4_727 (.A1(n_0_4_680), .A2(n_0_4_689), .A3(n_0_4_699), .ZN(
      dataOut2[27]));
   NAND2_X1 i_0_4_728 (.A1(n_0_55), .A2(\Memory[4] [28]), .ZN(n_0_4_700));
   NAND2_X1 i_0_4_729 (.A1(n_0_58), .A2(\Memory[7] [28]), .ZN(n_0_4_701));
   NAND2_X1 i_0_4_730 (.A1(n_0_54), .A2(\Memory[3] [28]), .ZN(n_0_4_702));
   NAND2_X1 i_0_4_731 (.A1(n_0_53), .A2(\Memory[2] [28]), .ZN(n_0_4_703));
   NAND4_X1 i_0_4_732 (.A1(n_0_4_700), .A2(n_0_4_701), .A3(n_0_4_702), .A4(
      n_0_4_703), .ZN(n_0_4_704));
   INV_X1 i_0_4_733 (.A(n_0_4_704), .ZN(n_0_4_705));
   NAND2_X1 i_0_4_734 (.A1(n_0_67), .A2(\Memory[16] [28]), .ZN(n_0_4_706));
   NAND2_X1 i_0_4_735 (.A1(n_0_57), .A2(\Memory[6] [28]), .ZN(n_0_4_707));
   NAND2_X1 i_0_4_736 (.A1(n_0_56), .A2(\Memory[5] [28]), .ZN(n_0_4_708));
   NAND3_X1 i_0_4_737 (.A1(n_0_4_706), .A2(n_0_4_707), .A3(n_0_4_708), .ZN(
      n_0_4_709));
   NAND2_X1 i_0_4_738 (.A1(n_0_59), .A2(\Memory[8] [28]), .ZN(n_0_4_710));
   NAND2_X1 i_0_4_739 (.A1(n_0_52), .A2(\Memory[1] [28]), .ZN(n_0_4_711));
   NAND2_X1 i_0_4_740 (.A1(n_0_61), .A2(\Memory[10] [28]), .ZN(n_0_4_712));
   NAND3_X1 i_0_4_741 (.A1(n_0_4_710), .A2(n_0_4_711), .A3(n_0_4_712), .ZN(
      n_0_4_713));
   NOR2_X1 i_0_4_742 (.A1(n_0_4_709), .A2(n_0_4_713), .ZN(n_0_4_714));
   NAND2_X1 i_0_4_743 (.A1(n_0_65), .A2(\Memory[14] [28]), .ZN(n_0_4_715));
   NAND2_X1 i_0_4_744 (.A1(n_0_66), .A2(\Memory[15] [28]), .ZN(n_0_4_716));
   NAND2_X1 i_0_4_745 (.A1(n_0_51), .A2(\Memory[0] [28]), .ZN(n_0_4_717));
   NAND2_X1 i_0_4_746 (.A1(n_0_60), .A2(\Memory[9] [28]), .ZN(n_0_4_718));
   NAND4_X1 i_0_4_747 (.A1(n_0_4_715), .A2(n_0_4_716), .A3(n_0_4_717), .A4(
      n_0_4_718), .ZN(n_0_4_719));
   NAND2_X1 i_0_4_748 (.A1(n_0_64), .A2(\Memory[13] [28]), .ZN(n_0_4_720));
   NAND2_X1 i_0_4_749 (.A1(n_0_63), .A2(\Memory[12] [28]), .ZN(n_0_4_721));
   NAND2_X1 i_0_4_750 (.A1(n_0_62), .A2(\Memory[11] [28]), .ZN(n_0_4_722));
   NAND3_X1 i_0_4_751 (.A1(n_0_4_720), .A2(n_0_4_721), .A3(n_0_4_722), .ZN(
      n_0_4_723));
   NOR2_X1 i_0_4_752 (.A1(n_0_4_719), .A2(n_0_4_723), .ZN(n_0_4_724));
   NAND3_X1 i_0_4_753 (.A1(n_0_4_705), .A2(n_0_4_714), .A3(n_0_4_724), .ZN(
      dataOut2[28]));
   NAND2_X1 i_0_4_754 (.A1(n_0_55), .A2(\Memory[4] [29]), .ZN(n_0_4_725));
   NAND2_X1 i_0_4_755 (.A1(n_0_58), .A2(\Memory[7] [29]), .ZN(n_0_4_726));
   NAND2_X1 i_0_4_756 (.A1(n_0_54), .A2(\Memory[3] [29]), .ZN(n_0_4_727));
   NAND2_X1 i_0_4_757 (.A1(n_0_53), .A2(\Memory[2] [29]), .ZN(n_0_4_728));
   NAND4_X1 i_0_4_758 (.A1(n_0_4_725), .A2(n_0_4_726), .A3(n_0_4_727), .A4(
      n_0_4_728), .ZN(n_0_4_729));
   INV_X1 i_0_4_759 (.A(n_0_4_729), .ZN(n_0_4_730));
   NAND2_X1 i_0_4_760 (.A1(n_0_67), .A2(\Memory[16] [29]), .ZN(n_0_4_731));
   NAND2_X1 i_0_4_761 (.A1(n_0_57), .A2(\Memory[6] [29]), .ZN(n_0_4_732));
   NAND2_X1 i_0_4_762 (.A1(n_0_56), .A2(\Memory[5] [29]), .ZN(n_0_4_733));
   NAND3_X1 i_0_4_763 (.A1(n_0_4_731), .A2(n_0_4_732), .A3(n_0_4_733), .ZN(
      n_0_4_734));
   NAND2_X1 i_0_4_764 (.A1(n_0_59), .A2(\Memory[8] [29]), .ZN(n_0_4_735));
   NAND2_X1 i_0_4_765 (.A1(n_0_52), .A2(\Memory[1] [29]), .ZN(n_0_4_736));
   NAND2_X1 i_0_4_766 (.A1(n_0_61), .A2(\Memory[10] [29]), .ZN(n_0_4_737));
   NAND3_X1 i_0_4_767 (.A1(n_0_4_735), .A2(n_0_4_736), .A3(n_0_4_737), .ZN(
      n_0_4_738));
   NOR2_X1 i_0_4_768 (.A1(n_0_4_734), .A2(n_0_4_738), .ZN(n_0_4_739));
   NAND2_X1 i_0_4_769 (.A1(n_0_65), .A2(\Memory[14] [29]), .ZN(n_0_4_740));
   NAND2_X1 i_0_4_770 (.A1(n_0_66), .A2(\Memory[15] [29]), .ZN(n_0_4_741));
   NAND2_X1 i_0_4_771 (.A1(n_0_51), .A2(\Memory[0] [29]), .ZN(n_0_4_742));
   NAND2_X1 i_0_4_772 (.A1(n_0_60), .A2(\Memory[9] [29]), .ZN(n_0_4_743));
   NAND4_X1 i_0_4_773 (.A1(n_0_4_740), .A2(n_0_4_741), .A3(n_0_4_742), .A4(
      n_0_4_743), .ZN(n_0_4_744));
   NAND2_X1 i_0_4_774 (.A1(n_0_64), .A2(\Memory[13] [29]), .ZN(n_0_4_745));
   NAND2_X1 i_0_4_775 (.A1(n_0_63), .A2(\Memory[12] [29]), .ZN(n_0_4_746));
   NAND2_X1 i_0_4_776 (.A1(n_0_62), .A2(\Memory[11] [29]), .ZN(n_0_4_747));
   NAND3_X1 i_0_4_777 (.A1(n_0_4_745), .A2(n_0_4_746), .A3(n_0_4_747), .ZN(
      n_0_4_748));
   NOR2_X1 i_0_4_778 (.A1(n_0_4_744), .A2(n_0_4_748), .ZN(n_0_4_749));
   NAND3_X1 i_0_4_779 (.A1(n_0_4_730), .A2(n_0_4_739), .A3(n_0_4_749), .ZN(
      dataOut2[29]));
   NAND2_X1 i_0_4_780 (.A1(n_0_55), .A2(\Memory[4] [30]), .ZN(n_0_4_750));
   NAND2_X1 i_0_4_781 (.A1(n_0_58), .A2(\Memory[7] [30]), .ZN(n_0_4_751));
   NAND2_X1 i_0_4_782 (.A1(n_0_54), .A2(\Memory[3] [30]), .ZN(n_0_4_752));
   NAND2_X1 i_0_4_783 (.A1(n_0_53), .A2(\Memory[2] [30]), .ZN(n_0_4_753));
   NAND4_X1 i_0_4_784 (.A1(n_0_4_750), .A2(n_0_4_751), .A3(n_0_4_752), .A4(
      n_0_4_753), .ZN(n_0_4_754));
   INV_X1 i_0_4_785 (.A(n_0_4_754), .ZN(n_0_4_755));
   NAND2_X1 i_0_4_786 (.A1(n_0_67), .A2(\Memory[16] [30]), .ZN(n_0_4_756));
   NAND2_X1 i_0_4_787 (.A1(n_0_57), .A2(\Memory[6] [30]), .ZN(n_0_4_757));
   NAND2_X1 i_0_4_788 (.A1(n_0_56), .A2(\Memory[5] [30]), .ZN(n_0_4_758));
   NAND3_X1 i_0_4_789 (.A1(n_0_4_756), .A2(n_0_4_757), .A3(n_0_4_758), .ZN(
      n_0_4_759));
   NAND2_X1 i_0_4_790 (.A1(n_0_59), .A2(\Memory[8] [30]), .ZN(n_0_4_760));
   NAND2_X1 i_0_4_791 (.A1(n_0_52), .A2(\Memory[1] [30]), .ZN(n_0_4_761));
   NAND2_X1 i_0_4_792 (.A1(n_0_61), .A2(\Memory[10] [30]), .ZN(n_0_4_762));
   NAND3_X1 i_0_4_793 (.A1(n_0_4_760), .A2(n_0_4_761), .A3(n_0_4_762), .ZN(
      n_0_4_763));
   NOR2_X1 i_0_4_794 (.A1(n_0_4_759), .A2(n_0_4_763), .ZN(n_0_4_764));
   NAND2_X1 i_0_4_795 (.A1(n_0_65), .A2(\Memory[14] [30]), .ZN(n_0_4_765));
   NAND2_X1 i_0_4_796 (.A1(n_0_66), .A2(\Memory[15] [30]), .ZN(n_0_4_766));
   NAND2_X1 i_0_4_797 (.A1(n_0_51), .A2(\Memory[0] [30]), .ZN(n_0_4_767));
   NAND2_X1 i_0_4_798 (.A1(n_0_60), .A2(\Memory[9] [30]), .ZN(n_0_4_768));
   NAND4_X1 i_0_4_799 (.A1(n_0_4_765), .A2(n_0_4_766), .A3(n_0_4_767), .A4(
      n_0_4_768), .ZN(n_0_4_769));
   NAND2_X1 i_0_4_800 (.A1(n_0_64), .A2(\Memory[13] [30]), .ZN(n_0_4_770));
   NAND2_X1 i_0_4_801 (.A1(n_0_63), .A2(\Memory[12] [30]), .ZN(n_0_4_771));
   NAND2_X1 i_0_4_802 (.A1(n_0_62), .A2(\Memory[11] [30]), .ZN(n_0_4_772));
   NAND3_X1 i_0_4_803 (.A1(n_0_4_770), .A2(n_0_4_771), .A3(n_0_4_772), .ZN(
      n_0_4_773));
   NOR2_X1 i_0_4_804 (.A1(n_0_4_769), .A2(n_0_4_773), .ZN(n_0_4_774));
   NAND3_X1 i_0_4_805 (.A1(n_0_4_755), .A2(n_0_4_764), .A3(n_0_4_774), .ZN(
      dataOut2[30]));
   NAND2_X1 i_0_4_806 (.A1(n_0_55), .A2(\Memory[4] [31]), .ZN(n_0_4_775));
   NAND2_X1 i_0_4_807 (.A1(n_0_58), .A2(\Memory[7] [31]), .ZN(n_0_4_776));
   NAND2_X1 i_0_4_808 (.A1(n_0_54), .A2(\Memory[3] [31]), .ZN(n_0_4_777));
   NAND2_X1 i_0_4_809 (.A1(n_0_53), .A2(\Memory[2] [31]), .ZN(n_0_4_778));
   NAND4_X1 i_0_4_810 (.A1(n_0_4_775), .A2(n_0_4_776), .A3(n_0_4_777), .A4(
      n_0_4_778), .ZN(n_0_4_779));
   INV_X1 i_0_4_811 (.A(n_0_4_779), .ZN(n_0_4_780));
   NAND2_X1 i_0_4_812 (.A1(n_0_67), .A2(\Memory[16] [31]), .ZN(n_0_4_781));
   NAND2_X1 i_0_4_813 (.A1(n_0_57), .A2(\Memory[6] [31]), .ZN(n_0_4_782));
   NAND2_X1 i_0_4_814 (.A1(n_0_56), .A2(\Memory[5] [31]), .ZN(n_0_4_783));
   NAND3_X1 i_0_4_815 (.A1(n_0_4_781), .A2(n_0_4_782), .A3(n_0_4_783), .ZN(
      n_0_4_784));
   NAND2_X1 i_0_4_816 (.A1(n_0_59), .A2(\Memory[8] [31]), .ZN(n_0_4_785));
   NAND2_X1 i_0_4_817 (.A1(n_0_52), .A2(\Memory[1] [31]), .ZN(n_0_4_786));
   NAND2_X1 i_0_4_818 (.A1(n_0_61), .A2(\Memory[10] [31]), .ZN(n_0_4_787));
   NAND3_X1 i_0_4_819 (.A1(n_0_4_785), .A2(n_0_4_786), .A3(n_0_4_787), .ZN(
      n_0_4_788));
   NOR2_X1 i_0_4_820 (.A1(n_0_4_784), .A2(n_0_4_788), .ZN(n_0_4_789));
   NAND2_X1 i_0_4_821 (.A1(n_0_65), .A2(\Memory[14] [31]), .ZN(n_0_4_790));
   NAND2_X1 i_0_4_822 (.A1(n_0_66), .A2(\Memory[15] [31]), .ZN(n_0_4_791));
   NAND2_X1 i_0_4_823 (.A1(n_0_51), .A2(\Memory[0] [31]), .ZN(n_0_4_792));
   NAND2_X1 i_0_4_824 (.A1(n_0_60), .A2(\Memory[9] [31]), .ZN(n_0_4_793));
   NAND4_X1 i_0_4_825 (.A1(n_0_4_790), .A2(n_0_4_791), .A3(n_0_4_792), .A4(
      n_0_4_793), .ZN(n_0_4_794));
   NAND2_X1 i_0_4_826 (.A1(n_0_64), .A2(\Memory[13] [31]), .ZN(n_0_4_795));
   NAND2_X1 i_0_4_827 (.A1(n_0_63), .A2(\Memory[12] [31]), .ZN(n_0_4_796));
   NAND2_X1 i_0_4_828 (.A1(n_0_62), .A2(\Memory[11] [31]), .ZN(n_0_4_797));
   NAND3_X1 i_0_4_829 (.A1(n_0_4_795), .A2(n_0_4_796), .A3(n_0_4_797), .ZN(
      n_0_4_798));
   NOR2_X1 i_0_4_830 (.A1(n_0_4_794), .A2(n_0_4_798), .ZN(n_0_4_799));
   NAND3_X1 i_0_4_831 (.A1(n_0_4_780), .A2(n_0_4_789), .A3(n_0_4_799), .ZN(
      dataOut2[31]));
   NAND2_X1 i_0_4_832 (.A1(n_0_55), .A2(\Memory[4] [32]), .ZN(n_0_4_800));
   NAND2_X1 i_0_4_833 (.A1(n_0_58), .A2(\Memory[7] [32]), .ZN(n_0_4_801));
   NAND2_X1 i_0_4_834 (.A1(n_0_54), .A2(\Memory[3] [32]), .ZN(n_0_4_802));
   NAND2_X1 i_0_4_835 (.A1(n_0_53), .A2(\Memory[2] [32]), .ZN(n_0_4_803));
   NAND4_X1 i_0_4_836 (.A1(n_0_4_800), .A2(n_0_4_801), .A3(n_0_4_802), .A4(
      n_0_4_803), .ZN(n_0_4_804));
   INV_X1 i_0_4_837 (.A(n_0_4_804), .ZN(n_0_4_805));
   NAND2_X1 i_0_4_838 (.A1(n_0_67), .A2(\Memory[16] [32]), .ZN(n_0_4_806));
   NAND2_X1 i_0_4_839 (.A1(n_0_57), .A2(\Memory[6] [32]), .ZN(n_0_4_807));
   NAND2_X1 i_0_4_840 (.A1(n_0_56), .A2(\Memory[5] [32]), .ZN(n_0_4_808));
   NAND3_X1 i_0_4_841 (.A1(n_0_4_806), .A2(n_0_4_807), .A3(n_0_4_808), .ZN(
      n_0_4_809));
   NAND2_X1 i_0_4_842 (.A1(n_0_59), .A2(\Memory[8] [32]), .ZN(n_0_4_810));
   NAND2_X1 i_0_4_843 (.A1(n_0_52), .A2(\Memory[1] [32]), .ZN(n_0_4_811));
   NAND2_X1 i_0_4_844 (.A1(n_0_61), .A2(\Memory[10] [32]), .ZN(n_0_4_812));
   NAND3_X1 i_0_4_845 (.A1(n_0_4_810), .A2(n_0_4_811), .A3(n_0_4_812), .ZN(
      n_0_4_813));
   NOR2_X1 i_0_4_846 (.A1(n_0_4_809), .A2(n_0_4_813), .ZN(n_0_4_814));
   NAND2_X1 i_0_4_847 (.A1(n_0_65), .A2(\Memory[14] [32]), .ZN(n_0_4_815));
   NAND2_X1 i_0_4_848 (.A1(n_0_66), .A2(\Memory[15] [32]), .ZN(n_0_4_816));
   NAND2_X1 i_0_4_849 (.A1(n_0_51), .A2(\Memory[0] [32]), .ZN(n_0_4_817));
   NAND2_X1 i_0_4_850 (.A1(n_0_60), .A2(\Memory[9] [32]), .ZN(n_0_4_818));
   NAND4_X1 i_0_4_851 (.A1(n_0_4_815), .A2(n_0_4_816), .A3(n_0_4_817), .A4(
      n_0_4_818), .ZN(n_0_4_819));
   NAND2_X1 i_0_4_852 (.A1(n_0_64), .A2(\Memory[13] [32]), .ZN(n_0_4_820));
   NAND2_X1 i_0_4_853 (.A1(n_0_63), .A2(\Memory[12] [32]), .ZN(n_0_4_821));
   NAND2_X1 i_0_4_854 (.A1(n_0_62), .A2(\Memory[11] [32]), .ZN(n_0_4_822));
   NAND3_X1 i_0_4_855 (.A1(n_0_4_820), .A2(n_0_4_821), .A3(n_0_4_822), .ZN(
      n_0_4_823));
   NOR2_X1 i_0_4_856 (.A1(n_0_4_819), .A2(n_0_4_823), .ZN(n_0_4_824));
   NAND3_X1 i_0_4_857 (.A1(n_0_4_805), .A2(n_0_4_814), .A3(n_0_4_824), .ZN(
      dataOut2[32]));
   NAND2_X1 i_0_4_858 (.A1(n_0_55), .A2(\Memory[4] [33]), .ZN(n_0_4_825));
   NAND2_X1 i_0_4_859 (.A1(n_0_58), .A2(\Memory[7] [33]), .ZN(n_0_4_826));
   NAND2_X1 i_0_4_860 (.A1(n_0_54), .A2(\Memory[3] [33]), .ZN(n_0_4_827));
   NAND2_X1 i_0_4_861 (.A1(n_0_53), .A2(\Memory[2] [33]), .ZN(n_0_4_828));
   NAND4_X1 i_0_4_862 (.A1(n_0_4_825), .A2(n_0_4_826), .A3(n_0_4_827), .A4(
      n_0_4_828), .ZN(n_0_4_829));
   INV_X1 i_0_4_863 (.A(n_0_4_829), .ZN(n_0_4_830));
   NAND2_X1 i_0_4_864 (.A1(n_0_67), .A2(\Memory[16] [33]), .ZN(n_0_4_831));
   NAND2_X1 i_0_4_865 (.A1(n_0_57), .A2(\Memory[6] [33]), .ZN(n_0_4_832));
   NAND2_X1 i_0_4_866 (.A1(n_0_56), .A2(\Memory[5] [33]), .ZN(n_0_4_833));
   NAND3_X1 i_0_4_867 (.A1(n_0_4_831), .A2(n_0_4_832), .A3(n_0_4_833), .ZN(
      n_0_4_834));
   NAND2_X1 i_0_4_868 (.A1(n_0_59), .A2(\Memory[8] [33]), .ZN(n_0_4_835));
   NAND2_X1 i_0_4_869 (.A1(n_0_52), .A2(\Memory[1] [33]), .ZN(n_0_4_836));
   NAND2_X1 i_0_4_870 (.A1(n_0_61), .A2(\Memory[10] [33]), .ZN(n_0_4_837));
   NAND3_X1 i_0_4_871 (.A1(n_0_4_835), .A2(n_0_4_836), .A3(n_0_4_837), .ZN(
      n_0_4_838));
   NOR2_X1 i_0_4_872 (.A1(n_0_4_834), .A2(n_0_4_838), .ZN(n_0_4_839));
   NAND2_X1 i_0_4_873 (.A1(n_0_65), .A2(\Memory[14] [33]), .ZN(n_0_4_840));
   NAND2_X1 i_0_4_874 (.A1(n_0_66), .A2(\Memory[15] [33]), .ZN(n_0_4_841));
   NAND2_X1 i_0_4_875 (.A1(n_0_51), .A2(\Memory[0] [33]), .ZN(n_0_4_842));
   NAND2_X1 i_0_4_876 (.A1(n_0_60), .A2(\Memory[9] [33]), .ZN(n_0_4_843));
   NAND4_X1 i_0_4_877 (.A1(n_0_4_840), .A2(n_0_4_841), .A3(n_0_4_842), .A4(
      n_0_4_843), .ZN(n_0_4_844));
   NAND2_X1 i_0_4_878 (.A1(n_0_64), .A2(\Memory[13] [33]), .ZN(n_0_4_845));
   NAND2_X1 i_0_4_879 (.A1(n_0_63), .A2(\Memory[12] [33]), .ZN(n_0_4_846));
   NAND2_X1 i_0_4_880 (.A1(n_0_62), .A2(\Memory[11] [33]), .ZN(n_0_4_847));
   NAND3_X1 i_0_4_881 (.A1(n_0_4_845), .A2(n_0_4_846), .A3(n_0_4_847), .ZN(
      n_0_4_848));
   NOR2_X1 i_0_4_882 (.A1(n_0_4_844), .A2(n_0_4_848), .ZN(n_0_4_849));
   NAND3_X1 i_0_4_883 (.A1(n_0_4_830), .A2(n_0_4_839), .A3(n_0_4_849), .ZN(
      dataOut2[33]));
   NAND2_X1 i_0_4_884 (.A1(n_0_55), .A2(\Memory[4] [34]), .ZN(n_0_4_850));
   NAND2_X1 i_0_4_885 (.A1(n_0_58), .A2(\Memory[7] [34]), .ZN(n_0_4_851));
   NAND2_X1 i_0_4_886 (.A1(n_0_54), .A2(\Memory[3] [34]), .ZN(n_0_4_852));
   NAND2_X1 i_0_4_887 (.A1(n_0_53), .A2(\Memory[2] [34]), .ZN(n_0_4_853));
   NAND4_X1 i_0_4_888 (.A1(n_0_4_850), .A2(n_0_4_851), .A3(n_0_4_852), .A4(
      n_0_4_853), .ZN(n_0_4_854));
   INV_X1 i_0_4_889 (.A(n_0_4_854), .ZN(n_0_4_855));
   NAND2_X1 i_0_4_890 (.A1(n_0_67), .A2(\Memory[16] [34]), .ZN(n_0_4_856));
   NAND2_X1 i_0_4_891 (.A1(n_0_57), .A2(\Memory[6] [34]), .ZN(n_0_4_857));
   NAND2_X1 i_0_4_892 (.A1(n_0_56), .A2(\Memory[5] [34]), .ZN(n_0_4_858));
   NAND3_X1 i_0_4_893 (.A1(n_0_4_856), .A2(n_0_4_857), .A3(n_0_4_858), .ZN(
      n_0_4_859));
   NAND2_X1 i_0_4_894 (.A1(n_0_59), .A2(\Memory[8] [34]), .ZN(n_0_4_860));
   NAND2_X1 i_0_4_895 (.A1(n_0_52), .A2(\Memory[1] [34]), .ZN(n_0_4_861));
   NAND2_X1 i_0_4_896 (.A1(n_0_61), .A2(\Memory[10] [34]), .ZN(n_0_4_862));
   NAND3_X1 i_0_4_897 (.A1(n_0_4_860), .A2(n_0_4_861), .A3(n_0_4_862), .ZN(
      n_0_4_863));
   NOR2_X1 i_0_4_898 (.A1(n_0_4_859), .A2(n_0_4_863), .ZN(n_0_4_864));
   NAND2_X1 i_0_4_899 (.A1(n_0_65), .A2(\Memory[14] [34]), .ZN(n_0_4_865));
   NAND2_X1 i_0_4_900 (.A1(n_0_66), .A2(\Memory[15] [34]), .ZN(n_0_4_866));
   NAND2_X1 i_0_4_901 (.A1(n_0_51), .A2(\Memory[0] [34]), .ZN(n_0_4_867));
   NAND2_X1 i_0_4_902 (.A1(n_0_60), .A2(\Memory[9] [34]), .ZN(n_0_4_868));
   NAND4_X1 i_0_4_903 (.A1(n_0_4_865), .A2(n_0_4_866), .A3(n_0_4_867), .A4(
      n_0_4_868), .ZN(n_0_4_869));
   NAND2_X1 i_0_4_904 (.A1(n_0_64), .A2(\Memory[13] [34]), .ZN(n_0_4_870));
   NAND2_X1 i_0_4_905 (.A1(n_0_63), .A2(\Memory[12] [34]), .ZN(n_0_4_871));
   NAND2_X1 i_0_4_906 (.A1(n_0_62), .A2(\Memory[11] [34]), .ZN(n_0_4_872));
   NAND3_X1 i_0_4_907 (.A1(n_0_4_870), .A2(n_0_4_871), .A3(n_0_4_872), .ZN(
      n_0_4_873));
   NOR2_X1 i_0_4_908 (.A1(n_0_4_869), .A2(n_0_4_873), .ZN(n_0_4_874));
   NAND3_X1 i_0_4_909 (.A1(n_0_4_855), .A2(n_0_4_864), .A3(n_0_4_874), .ZN(
      dataOut2[34]));
   NAND2_X1 i_0_4_910 (.A1(n_0_55), .A2(\Memory[4] [35]), .ZN(n_0_4_875));
   NAND2_X1 i_0_4_911 (.A1(n_0_58), .A2(\Memory[7] [35]), .ZN(n_0_4_876));
   NAND2_X1 i_0_4_912 (.A1(n_0_54), .A2(\Memory[3] [35]), .ZN(n_0_4_877));
   NAND2_X1 i_0_4_913 (.A1(n_0_53), .A2(\Memory[2] [35]), .ZN(n_0_4_878));
   NAND4_X1 i_0_4_914 (.A1(n_0_4_875), .A2(n_0_4_876), .A3(n_0_4_877), .A4(
      n_0_4_878), .ZN(n_0_4_879));
   INV_X1 i_0_4_915 (.A(n_0_4_879), .ZN(n_0_4_880));
   NAND2_X1 i_0_4_916 (.A1(n_0_67), .A2(\Memory[16] [35]), .ZN(n_0_4_881));
   NAND2_X1 i_0_4_917 (.A1(n_0_57), .A2(\Memory[6] [35]), .ZN(n_0_4_882));
   NAND2_X1 i_0_4_918 (.A1(n_0_56), .A2(\Memory[5] [35]), .ZN(n_0_4_883));
   NAND3_X1 i_0_4_919 (.A1(n_0_4_881), .A2(n_0_4_882), .A3(n_0_4_883), .ZN(
      n_0_4_884));
   NAND2_X1 i_0_4_920 (.A1(n_0_59), .A2(\Memory[8] [35]), .ZN(n_0_4_885));
   NAND2_X1 i_0_4_921 (.A1(n_0_52), .A2(\Memory[1] [35]), .ZN(n_0_4_886));
   NAND2_X1 i_0_4_922 (.A1(n_0_61), .A2(\Memory[10] [35]), .ZN(n_0_4_887));
   NAND3_X1 i_0_4_923 (.A1(n_0_4_885), .A2(n_0_4_886), .A3(n_0_4_887), .ZN(
      n_0_4_888));
   NOR2_X1 i_0_4_924 (.A1(n_0_4_884), .A2(n_0_4_888), .ZN(n_0_4_889));
   NAND2_X1 i_0_4_925 (.A1(n_0_65), .A2(\Memory[14] [35]), .ZN(n_0_4_890));
   NAND2_X1 i_0_4_926 (.A1(n_0_66), .A2(\Memory[15] [35]), .ZN(n_0_4_891));
   NAND2_X1 i_0_4_927 (.A1(n_0_51), .A2(\Memory[0] [35]), .ZN(n_0_4_892));
   NAND2_X1 i_0_4_928 (.A1(n_0_60), .A2(\Memory[9] [35]), .ZN(n_0_4_893));
   NAND4_X1 i_0_4_929 (.A1(n_0_4_890), .A2(n_0_4_891), .A3(n_0_4_892), .A4(
      n_0_4_893), .ZN(n_0_4_894));
   NAND2_X1 i_0_4_930 (.A1(n_0_64), .A2(\Memory[13] [35]), .ZN(n_0_4_895));
   NAND2_X1 i_0_4_931 (.A1(n_0_63), .A2(\Memory[12] [35]), .ZN(n_0_4_896));
   NAND2_X1 i_0_4_932 (.A1(n_0_62), .A2(\Memory[11] [35]), .ZN(n_0_4_897));
   NAND3_X1 i_0_4_933 (.A1(n_0_4_895), .A2(n_0_4_896), .A3(n_0_4_897), .ZN(
      n_0_4_898));
   NOR2_X1 i_0_4_934 (.A1(n_0_4_894), .A2(n_0_4_898), .ZN(n_0_4_899));
   NAND3_X1 i_0_4_935 (.A1(n_0_4_880), .A2(n_0_4_889), .A3(n_0_4_899), .ZN(
      dataOut2[35]));
   NAND2_X1 i_0_4_936 (.A1(n_0_55), .A2(\Memory[4] [36]), .ZN(n_0_4_900));
   NAND2_X1 i_0_4_937 (.A1(n_0_58), .A2(\Memory[7] [36]), .ZN(n_0_4_901));
   NAND2_X1 i_0_4_938 (.A1(n_0_54), .A2(\Memory[3] [36]), .ZN(n_0_4_902));
   NAND2_X1 i_0_4_939 (.A1(n_0_53), .A2(\Memory[2] [36]), .ZN(n_0_4_903));
   NAND4_X1 i_0_4_940 (.A1(n_0_4_900), .A2(n_0_4_901), .A3(n_0_4_902), .A4(
      n_0_4_903), .ZN(n_0_4_904));
   INV_X1 i_0_4_941 (.A(n_0_4_904), .ZN(n_0_4_905));
   NAND2_X1 i_0_4_942 (.A1(n_0_67), .A2(\Memory[16] [36]), .ZN(n_0_4_906));
   NAND2_X1 i_0_4_943 (.A1(n_0_57), .A2(\Memory[6] [36]), .ZN(n_0_4_907));
   NAND2_X1 i_0_4_944 (.A1(n_0_56), .A2(\Memory[5] [36]), .ZN(n_0_4_908));
   NAND3_X1 i_0_4_945 (.A1(n_0_4_906), .A2(n_0_4_907), .A3(n_0_4_908), .ZN(
      n_0_4_909));
   NAND2_X1 i_0_4_946 (.A1(n_0_59), .A2(\Memory[8] [36]), .ZN(n_0_4_910));
   NAND2_X1 i_0_4_947 (.A1(n_0_52), .A2(\Memory[1] [36]), .ZN(n_0_4_911));
   NAND2_X1 i_0_4_948 (.A1(n_0_61), .A2(\Memory[10] [36]), .ZN(n_0_4_912));
   NAND3_X1 i_0_4_949 (.A1(n_0_4_910), .A2(n_0_4_911), .A3(n_0_4_912), .ZN(
      n_0_4_913));
   NOR2_X1 i_0_4_950 (.A1(n_0_4_909), .A2(n_0_4_913), .ZN(n_0_4_914));
   NAND2_X1 i_0_4_951 (.A1(n_0_65), .A2(\Memory[14] [36]), .ZN(n_0_4_915));
   NAND2_X1 i_0_4_952 (.A1(n_0_66), .A2(\Memory[15] [36]), .ZN(n_0_4_916));
   NAND2_X1 i_0_4_953 (.A1(n_0_51), .A2(\Memory[0] [36]), .ZN(n_0_4_917));
   NAND2_X1 i_0_4_954 (.A1(n_0_60), .A2(\Memory[9] [36]), .ZN(n_0_4_918));
   NAND4_X1 i_0_4_955 (.A1(n_0_4_915), .A2(n_0_4_916), .A3(n_0_4_917), .A4(
      n_0_4_918), .ZN(n_0_4_919));
   NAND2_X1 i_0_4_956 (.A1(n_0_64), .A2(\Memory[13] [36]), .ZN(n_0_4_920));
   NAND2_X1 i_0_4_957 (.A1(n_0_63), .A2(\Memory[12] [36]), .ZN(n_0_4_921));
   NAND2_X1 i_0_4_958 (.A1(n_0_62), .A2(\Memory[11] [36]), .ZN(n_0_4_922));
   NAND3_X1 i_0_4_959 (.A1(n_0_4_920), .A2(n_0_4_921), .A3(n_0_4_922), .ZN(
      n_0_4_923));
   NOR2_X1 i_0_4_960 (.A1(n_0_4_919), .A2(n_0_4_923), .ZN(n_0_4_924));
   NAND3_X1 i_0_4_961 (.A1(n_0_4_905), .A2(n_0_4_914), .A3(n_0_4_924), .ZN(
      dataOut2[36]));
   NAND2_X1 i_0_4_962 (.A1(n_0_55), .A2(\Memory[4] [37]), .ZN(n_0_4_925));
   NAND2_X1 i_0_4_963 (.A1(n_0_58), .A2(\Memory[7] [37]), .ZN(n_0_4_926));
   NAND2_X1 i_0_4_964 (.A1(n_0_54), .A2(\Memory[3] [37]), .ZN(n_0_4_927));
   NAND2_X1 i_0_4_965 (.A1(n_0_53), .A2(\Memory[2] [37]), .ZN(n_0_4_928));
   NAND4_X1 i_0_4_966 (.A1(n_0_4_925), .A2(n_0_4_926), .A3(n_0_4_927), .A4(
      n_0_4_928), .ZN(n_0_4_929));
   INV_X1 i_0_4_967 (.A(n_0_4_929), .ZN(n_0_4_930));
   NAND2_X1 i_0_4_968 (.A1(n_0_67), .A2(\Memory[16] [37]), .ZN(n_0_4_931));
   NAND2_X1 i_0_4_969 (.A1(n_0_57), .A2(\Memory[6] [37]), .ZN(n_0_4_932));
   NAND2_X1 i_0_4_970 (.A1(n_0_56), .A2(\Memory[5] [37]), .ZN(n_0_4_933));
   NAND3_X1 i_0_4_971 (.A1(n_0_4_931), .A2(n_0_4_932), .A3(n_0_4_933), .ZN(
      n_0_4_934));
   NAND2_X1 i_0_4_972 (.A1(n_0_59), .A2(\Memory[8] [37]), .ZN(n_0_4_935));
   NAND2_X1 i_0_4_973 (.A1(n_0_52), .A2(\Memory[1] [37]), .ZN(n_0_4_936));
   NAND2_X1 i_0_4_974 (.A1(n_0_61), .A2(\Memory[10] [37]), .ZN(n_0_4_937));
   NAND3_X1 i_0_4_975 (.A1(n_0_4_935), .A2(n_0_4_936), .A3(n_0_4_937), .ZN(
      n_0_4_938));
   NOR2_X1 i_0_4_976 (.A1(n_0_4_934), .A2(n_0_4_938), .ZN(n_0_4_939));
   NAND2_X1 i_0_4_977 (.A1(n_0_65), .A2(\Memory[14] [37]), .ZN(n_0_4_940));
   NAND2_X1 i_0_4_978 (.A1(n_0_66), .A2(\Memory[15] [37]), .ZN(n_0_4_941));
   NAND2_X1 i_0_4_979 (.A1(n_0_51), .A2(\Memory[0] [37]), .ZN(n_0_4_942));
   NAND2_X1 i_0_4_980 (.A1(n_0_60), .A2(\Memory[9] [37]), .ZN(n_0_4_943));
   NAND4_X1 i_0_4_981 (.A1(n_0_4_940), .A2(n_0_4_941), .A3(n_0_4_942), .A4(
      n_0_4_943), .ZN(n_0_4_944));
   NAND2_X1 i_0_4_982 (.A1(n_0_64), .A2(\Memory[13] [37]), .ZN(n_0_4_945));
   NAND2_X1 i_0_4_983 (.A1(n_0_63), .A2(\Memory[12] [37]), .ZN(n_0_4_946));
   NAND2_X1 i_0_4_984 (.A1(n_0_62), .A2(\Memory[11] [37]), .ZN(n_0_4_947));
   NAND3_X1 i_0_4_985 (.A1(n_0_4_945), .A2(n_0_4_946), .A3(n_0_4_947), .ZN(
      n_0_4_948));
   NOR2_X1 i_0_4_986 (.A1(n_0_4_944), .A2(n_0_4_948), .ZN(n_0_4_949));
   NAND3_X1 i_0_4_987 (.A1(n_0_4_930), .A2(n_0_4_939), .A3(n_0_4_949), .ZN(
      dataOut2[37]));
   NAND2_X1 i_0_4_988 (.A1(n_0_55), .A2(\Memory[4] [38]), .ZN(n_0_4_950));
   NAND2_X1 i_0_4_989 (.A1(n_0_58), .A2(\Memory[7] [38]), .ZN(n_0_4_951));
   NAND2_X1 i_0_4_990 (.A1(n_0_54), .A2(\Memory[3] [38]), .ZN(n_0_4_952));
   NAND2_X1 i_0_4_991 (.A1(n_0_53), .A2(\Memory[2] [38]), .ZN(n_0_4_953));
   NAND4_X1 i_0_4_992 (.A1(n_0_4_950), .A2(n_0_4_951), .A3(n_0_4_952), .A4(
      n_0_4_953), .ZN(n_0_4_954));
   INV_X1 i_0_4_993 (.A(n_0_4_954), .ZN(n_0_4_955));
   NAND2_X1 i_0_4_994 (.A1(n_0_67), .A2(\Memory[16] [38]), .ZN(n_0_4_956));
   NAND2_X1 i_0_4_995 (.A1(n_0_57), .A2(\Memory[6] [38]), .ZN(n_0_4_957));
   NAND2_X1 i_0_4_996 (.A1(n_0_56), .A2(\Memory[5] [38]), .ZN(n_0_4_958));
   NAND3_X1 i_0_4_997 (.A1(n_0_4_956), .A2(n_0_4_957), .A3(n_0_4_958), .ZN(
      n_0_4_959));
   NAND2_X1 i_0_4_998 (.A1(n_0_59), .A2(\Memory[8] [38]), .ZN(n_0_4_960));
   NAND2_X1 i_0_4_999 (.A1(n_0_52), .A2(\Memory[1] [38]), .ZN(n_0_4_961));
   NAND2_X1 i_0_4_1000 (.A1(n_0_61), .A2(\Memory[10] [38]), .ZN(n_0_4_962));
   NAND3_X1 i_0_4_1001 (.A1(n_0_4_960), .A2(n_0_4_961), .A3(n_0_4_962), .ZN(
      n_0_4_963));
   NOR2_X1 i_0_4_1002 (.A1(n_0_4_959), .A2(n_0_4_963), .ZN(n_0_4_964));
   NAND2_X1 i_0_4_1003 (.A1(n_0_65), .A2(\Memory[14] [38]), .ZN(n_0_4_965));
   NAND2_X1 i_0_4_1004 (.A1(n_0_66), .A2(\Memory[15] [38]), .ZN(n_0_4_966));
   NAND2_X1 i_0_4_1005 (.A1(n_0_51), .A2(\Memory[0] [38]), .ZN(n_0_4_967));
   NAND2_X1 i_0_4_1006 (.A1(n_0_60), .A2(\Memory[9] [38]), .ZN(n_0_4_968));
   NAND4_X1 i_0_4_1007 (.A1(n_0_4_965), .A2(n_0_4_966), .A3(n_0_4_967), .A4(
      n_0_4_968), .ZN(n_0_4_969));
   NAND2_X1 i_0_4_1008 (.A1(n_0_64), .A2(\Memory[13] [38]), .ZN(n_0_4_970));
   NAND2_X1 i_0_4_1009 (.A1(n_0_63), .A2(\Memory[12] [38]), .ZN(n_0_4_971));
   NAND2_X1 i_0_4_1010 (.A1(n_0_62), .A2(\Memory[11] [38]), .ZN(n_0_4_972));
   NAND3_X1 i_0_4_1011 (.A1(n_0_4_970), .A2(n_0_4_971), .A3(n_0_4_972), .ZN(
      n_0_4_973));
   NOR2_X1 i_0_4_1012 (.A1(n_0_4_969), .A2(n_0_4_973), .ZN(n_0_4_974));
   NAND3_X1 i_0_4_1013 (.A1(n_0_4_955), .A2(n_0_4_964), .A3(n_0_4_974), .ZN(
      dataOut2[38]));
   NAND2_X1 i_0_4_1014 (.A1(n_0_55), .A2(\Memory[4] [39]), .ZN(n_0_4_975));
   NAND2_X1 i_0_4_1015 (.A1(n_0_58), .A2(\Memory[7] [39]), .ZN(n_0_4_976));
   NAND2_X1 i_0_4_1016 (.A1(n_0_54), .A2(\Memory[3] [39]), .ZN(n_0_4_977));
   NAND2_X1 i_0_4_1017 (.A1(n_0_53), .A2(\Memory[2] [39]), .ZN(n_0_4_978));
   NAND4_X1 i_0_4_1018 (.A1(n_0_4_975), .A2(n_0_4_976), .A3(n_0_4_977), .A4(
      n_0_4_978), .ZN(n_0_4_979));
   INV_X1 i_0_4_1019 (.A(n_0_4_979), .ZN(n_0_4_980));
   NAND2_X1 i_0_4_1020 (.A1(n_0_67), .A2(\Memory[16] [39]), .ZN(n_0_4_981));
   NAND2_X1 i_0_4_1021 (.A1(n_0_57), .A2(\Memory[6] [39]), .ZN(n_0_4_982));
   NAND2_X1 i_0_4_1022 (.A1(n_0_56), .A2(\Memory[5] [39]), .ZN(n_0_4_983));
   NAND3_X1 i_0_4_1023 (.A1(n_0_4_981), .A2(n_0_4_982), .A3(n_0_4_983), .ZN(
      n_0_4_984));
   NAND2_X1 i_0_4_1024 (.A1(n_0_59), .A2(\Memory[8] [39]), .ZN(n_0_4_985));
   NAND2_X1 i_0_4_1025 (.A1(n_0_52), .A2(\Memory[1] [39]), .ZN(n_0_4_986));
   NAND2_X1 i_0_4_1026 (.A1(n_0_61), .A2(\Memory[10] [39]), .ZN(n_0_4_987));
   NAND3_X1 i_0_4_1027 (.A1(n_0_4_985), .A2(n_0_4_986), .A3(n_0_4_987), .ZN(
      n_0_4_988));
   NOR2_X1 i_0_4_1028 (.A1(n_0_4_984), .A2(n_0_4_988), .ZN(n_0_4_989));
   NAND2_X1 i_0_4_1029 (.A1(n_0_65), .A2(\Memory[14] [39]), .ZN(n_0_4_990));
   NAND2_X1 i_0_4_1030 (.A1(n_0_66), .A2(\Memory[15] [39]), .ZN(n_0_4_991));
   NAND2_X1 i_0_4_1031 (.A1(n_0_51), .A2(\Memory[0] [39]), .ZN(n_0_4_992));
   NAND2_X1 i_0_4_1032 (.A1(n_0_60), .A2(\Memory[9] [39]), .ZN(n_0_4_993));
   NAND4_X1 i_0_4_1033 (.A1(n_0_4_990), .A2(n_0_4_991), .A3(n_0_4_992), .A4(
      n_0_4_993), .ZN(n_0_4_994));
   NAND2_X1 i_0_4_1034 (.A1(n_0_64), .A2(\Memory[13] [39]), .ZN(n_0_4_995));
   NAND2_X1 i_0_4_1035 (.A1(n_0_63), .A2(\Memory[12] [39]), .ZN(n_0_4_996));
   NAND2_X1 i_0_4_1036 (.A1(n_0_62), .A2(\Memory[11] [39]), .ZN(n_0_4_997));
   NAND3_X1 i_0_4_1037 (.A1(n_0_4_995), .A2(n_0_4_996), .A3(n_0_4_997), .ZN(
      n_0_4_998));
   NOR2_X1 i_0_4_1038 (.A1(n_0_4_994), .A2(n_0_4_998), .ZN(n_0_4_999));
   NAND3_X1 i_0_4_1039 (.A1(n_0_4_980), .A2(n_0_4_989), .A3(n_0_4_999), .ZN(
      dataOut2[39]));
   NAND2_X1 i_0_4_1040 (.A1(n_0_55), .A2(\Memory[4] [40]), .ZN(n_0_4_1000));
   NAND2_X1 i_0_4_1041 (.A1(n_0_58), .A2(\Memory[7] [40]), .ZN(n_0_4_1001));
   NAND2_X1 i_0_4_1042 (.A1(n_0_54), .A2(\Memory[3] [40]), .ZN(n_0_4_1002));
   NAND2_X1 i_0_4_1043 (.A1(n_0_53), .A2(\Memory[2] [40]), .ZN(n_0_4_1003));
   NAND4_X1 i_0_4_1044 (.A1(n_0_4_1000), .A2(n_0_4_1001), .A3(n_0_4_1002), 
      .A4(n_0_4_1003), .ZN(n_0_4_1004));
   INV_X1 i_0_4_1045 (.A(n_0_4_1004), .ZN(n_0_4_1005));
   NAND2_X1 i_0_4_1046 (.A1(n_0_67), .A2(\Memory[16] [40]), .ZN(n_0_4_1006));
   NAND2_X1 i_0_4_1047 (.A1(n_0_57), .A2(\Memory[6] [40]), .ZN(n_0_4_1007));
   NAND2_X1 i_0_4_1048 (.A1(n_0_56), .A2(\Memory[5] [40]), .ZN(n_0_4_1008));
   NAND3_X1 i_0_4_1049 (.A1(n_0_4_1006), .A2(n_0_4_1007), .A3(n_0_4_1008), 
      .ZN(n_0_4_1009));
   NAND2_X1 i_0_4_1050 (.A1(n_0_59), .A2(\Memory[8] [40]), .ZN(n_0_4_1010));
   NAND2_X1 i_0_4_1051 (.A1(n_0_52), .A2(\Memory[1] [40]), .ZN(n_0_4_1011));
   NAND2_X1 i_0_4_1052 (.A1(n_0_61), .A2(\Memory[10] [40]), .ZN(n_0_4_1012));
   NAND3_X1 i_0_4_1053 (.A1(n_0_4_1010), .A2(n_0_4_1011), .A3(n_0_4_1012), 
      .ZN(n_0_4_1013));
   NOR2_X1 i_0_4_1054 (.A1(n_0_4_1009), .A2(n_0_4_1013), .ZN(n_0_4_1014));
   NAND2_X1 i_0_4_1055 (.A1(n_0_65), .A2(\Memory[14] [40]), .ZN(n_0_4_1015));
   NAND2_X1 i_0_4_1056 (.A1(n_0_66), .A2(\Memory[15] [40]), .ZN(n_0_4_1016));
   NAND2_X1 i_0_4_1057 (.A1(n_0_51), .A2(\Memory[0] [40]), .ZN(n_0_4_1017));
   NAND2_X1 i_0_4_1058 (.A1(n_0_60), .A2(\Memory[9] [40]), .ZN(n_0_4_1018));
   NAND4_X1 i_0_4_1059 (.A1(n_0_4_1015), .A2(n_0_4_1016), .A3(n_0_4_1017), 
      .A4(n_0_4_1018), .ZN(n_0_4_1019));
   NAND2_X1 i_0_4_1060 (.A1(n_0_64), .A2(\Memory[13] [40]), .ZN(n_0_4_1020));
   NAND2_X1 i_0_4_1061 (.A1(n_0_63), .A2(\Memory[12] [40]), .ZN(n_0_4_1021));
   NAND2_X1 i_0_4_1062 (.A1(n_0_62), .A2(\Memory[11] [40]), .ZN(n_0_4_1022));
   NAND3_X1 i_0_4_1063 (.A1(n_0_4_1020), .A2(n_0_4_1021), .A3(n_0_4_1022), 
      .ZN(n_0_4_1023));
   NOR2_X1 i_0_4_1064 (.A1(n_0_4_1019), .A2(n_0_4_1023), .ZN(n_0_4_1024));
   NAND3_X1 i_0_4_1065 (.A1(n_0_4_1005), .A2(n_0_4_1014), .A3(n_0_4_1024), 
      .ZN(dataOut2[40]));
   NAND2_X1 i_0_4_1066 (.A1(n_0_55), .A2(\Memory[4] [41]), .ZN(n_0_4_1025));
   NAND2_X1 i_0_4_1067 (.A1(n_0_58), .A2(\Memory[7] [41]), .ZN(n_0_4_1026));
   NAND2_X1 i_0_4_1068 (.A1(n_0_54), .A2(\Memory[3] [41]), .ZN(n_0_4_1027));
   NAND2_X1 i_0_4_1069 (.A1(n_0_53), .A2(\Memory[2] [41]), .ZN(n_0_4_1028));
   NAND4_X1 i_0_4_1070 (.A1(n_0_4_1025), .A2(n_0_4_1026), .A3(n_0_4_1027), 
      .A4(n_0_4_1028), .ZN(n_0_4_1029));
   INV_X1 i_0_4_1071 (.A(n_0_4_1029), .ZN(n_0_4_1030));
   NAND2_X1 i_0_4_1072 (.A1(n_0_67), .A2(\Memory[16] [41]), .ZN(n_0_4_1031));
   NAND2_X1 i_0_4_1073 (.A1(n_0_57), .A2(\Memory[6] [41]), .ZN(n_0_4_1032));
   NAND2_X1 i_0_4_1074 (.A1(n_0_56), .A2(\Memory[5] [41]), .ZN(n_0_4_1033));
   NAND3_X1 i_0_4_1075 (.A1(n_0_4_1031), .A2(n_0_4_1032), .A3(n_0_4_1033), 
      .ZN(n_0_4_1034));
   NAND2_X1 i_0_4_1076 (.A1(n_0_59), .A2(\Memory[8] [41]), .ZN(n_0_4_1035));
   NAND2_X1 i_0_4_1077 (.A1(n_0_52), .A2(\Memory[1] [41]), .ZN(n_0_4_1036));
   NAND2_X1 i_0_4_1078 (.A1(n_0_61), .A2(\Memory[10] [41]), .ZN(n_0_4_1037));
   NAND3_X1 i_0_4_1079 (.A1(n_0_4_1035), .A2(n_0_4_1036), .A3(n_0_4_1037), 
      .ZN(n_0_4_1038));
   NOR2_X1 i_0_4_1080 (.A1(n_0_4_1034), .A2(n_0_4_1038), .ZN(n_0_4_1039));
   NAND2_X1 i_0_4_1081 (.A1(n_0_65), .A2(\Memory[14] [41]), .ZN(n_0_4_1040));
   NAND2_X1 i_0_4_1082 (.A1(n_0_66), .A2(\Memory[15] [41]), .ZN(n_0_4_1041));
   NAND2_X1 i_0_4_1083 (.A1(n_0_51), .A2(\Memory[0] [41]), .ZN(n_0_4_1042));
   NAND2_X1 i_0_4_1084 (.A1(n_0_60), .A2(\Memory[9] [41]), .ZN(n_0_4_1043));
   NAND4_X1 i_0_4_1085 (.A1(n_0_4_1040), .A2(n_0_4_1041), .A3(n_0_4_1042), 
      .A4(n_0_4_1043), .ZN(n_0_4_1044));
   NAND2_X1 i_0_4_1086 (.A1(n_0_64), .A2(\Memory[13] [41]), .ZN(n_0_4_1045));
   NAND2_X1 i_0_4_1087 (.A1(n_0_63), .A2(\Memory[12] [41]), .ZN(n_0_4_1046));
   NAND2_X1 i_0_4_1088 (.A1(n_0_62), .A2(\Memory[11] [41]), .ZN(n_0_4_1047));
   NAND3_X1 i_0_4_1089 (.A1(n_0_4_1045), .A2(n_0_4_1046), .A3(n_0_4_1047), 
      .ZN(n_0_4_1048));
   NOR2_X1 i_0_4_1090 (.A1(n_0_4_1044), .A2(n_0_4_1048), .ZN(n_0_4_1049));
   NAND3_X1 i_0_4_1091 (.A1(n_0_4_1030), .A2(n_0_4_1039), .A3(n_0_4_1049), 
      .ZN(dataOut2[41]));
   NAND2_X1 i_0_4_1092 (.A1(n_0_55), .A2(\Memory[4] [42]), .ZN(n_0_4_1050));
   NAND2_X1 i_0_4_1093 (.A1(n_0_58), .A2(\Memory[7] [42]), .ZN(n_0_4_1051));
   NAND2_X1 i_0_4_1094 (.A1(n_0_54), .A2(\Memory[3] [42]), .ZN(n_0_4_1052));
   NAND2_X1 i_0_4_1095 (.A1(n_0_53), .A2(\Memory[2] [42]), .ZN(n_0_4_1053));
   NAND4_X1 i_0_4_1096 (.A1(n_0_4_1050), .A2(n_0_4_1051), .A3(n_0_4_1052), 
      .A4(n_0_4_1053), .ZN(n_0_4_1054));
   INV_X1 i_0_4_1097 (.A(n_0_4_1054), .ZN(n_0_4_1055));
   NAND2_X1 i_0_4_1098 (.A1(n_0_67), .A2(\Memory[16] [42]), .ZN(n_0_4_1056));
   NAND2_X1 i_0_4_1099 (.A1(n_0_57), .A2(\Memory[6] [42]), .ZN(n_0_4_1057));
   NAND2_X1 i_0_4_1100 (.A1(n_0_56), .A2(\Memory[5] [42]), .ZN(n_0_4_1058));
   NAND3_X1 i_0_4_1101 (.A1(n_0_4_1056), .A2(n_0_4_1057), .A3(n_0_4_1058), 
      .ZN(n_0_4_1059));
   NAND2_X1 i_0_4_1102 (.A1(n_0_59), .A2(\Memory[8] [42]), .ZN(n_0_4_1060));
   NAND2_X1 i_0_4_1103 (.A1(n_0_52), .A2(\Memory[1] [42]), .ZN(n_0_4_1061));
   NAND2_X1 i_0_4_1104 (.A1(n_0_61), .A2(\Memory[10] [42]), .ZN(n_0_4_1062));
   NAND3_X1 i_0_4_1105 (.A1(n_0_4_1060), .A2(n_0_4_1061), .A3(n_0_4_1062), 
      .ZN(n_0_4_1063));
   NOR2_X1 i_0_4_1106 (.A1(n_0_4_1059), .A2(n_0_4_1063), .ZN(n_0_4_1064));
   NAND2_X1 i_0_4_1107 (.A1(n_0_65), .A2(\Memory[14] [42]), .ZN(n_0_4_1065));
   NAND2_X1 i_0_4_1108 (.A1(n_0_66), .A2(\Memory[15] [42]), .ZN(n_0_4_1066));
   NAND2_X1 i_0_4_1109 (.A1(n_0_51), .A2(\Memory[0] [42]), .ZN(n_0_4_1067));
   NAND2_X1 i_0_4_1110 (.A1(n_0_60), .A2(\Memory[9] [42]), .ZN(n_0_4_1068));
   NAND4_X1 i_0_4_1111 (.A1(n_0_4_1065), .A2(n_0_4_1066), .A3(n_0_4_1067), 
      .A4(n_0_4_1068), .ZN(n_0_4_1069));
   NAND2_X1 i_0_4_1112 (.A1(n_0_64), .A2(\Memory[13] [42]), .ZN(n_0_4_1070));
   NAND2_X1 i_0_4_1113 (.A1(n_0_63), .A2(\Memory[12] [42]), .ZN(n_0_4_1071));
   NAND2_X1 i_0_4_1114 (.A1(n_0_62), .A2(\Memory[11] [42]), .ZN(n_0_4_1072));
   NAND3_X1 i_0_4_1115 (.A1(n_0_4_1070), .A2(n_0_4_1071), .A3(n_0_4_1072), 
      .ZN(n_0_4_1073));
   NOR2_X1 i_0_4_1116 (.A1(n_0_4_1069), .A2(n_0_4_1073), .ZN(n_0_4_1074));
   NAND3_X1 i_0_4_1117 (.A1(n_0_4_1055), .A2(n_0_4_1064), .A3(n_0_4_1074), 
      .ZN(dataOut2[42]));
   NAND2_X1 i_0_4_1118 (.A1(n_0_55), .A2(\Memory[4] [43]), .ZN(n_0_4_1075));
   NAND2_X1 i_0_4_1119 (.A1(n_0_58), .A2(\Memory[7] [43]), .ZN(n_0_4_1076));
   NAND2_X1 i_0_4_1120 (.A1(n_0_54), .A2(\Memory[3] [43]), .ZN(n_0_4_1077));
   NAND2_X1 i_0_4_1121 (.A1(n_0_53), .A2(\Memory[2] [43]), .ZN(n_0_4_1078));
   NAND4_X1 i_0_4_1122 (.A1(n_0_4_1075), .A2(n_0_4_1076), .A3(n_0_4_1077), 
      .A4(n_0_4_1078), .ZN(n_0_4_1079));
   INV_X1 i_0_4_1123 (.A(n_0_4_1079), .ZN(n_0_4_1080));
   NAND2_X1 i_0_4_1124 (.A1(n_0_67), .A2(\Memory[16] [43]), .ZN(n_0_4_1081));
   NAND2_X1 i_0_4_1125 (.A1(n_0_57), .A2(\Memory[6] [43]), .ZN(n_0_4_1082));
   NAND2_X1 i_0_4_1126 (.A1(n_0_56), .A2(\Memory[5] [43]), .ZN(n_0_4_1083));
   NAND3_X1 i_0_4_1127 (.A1(n_0_4_1081), .A2(n_0_4_1082), .A3(n_0_4_1083), 
      .ZN(n_0_4_1084));
   NAND2_X1 i_0_4_1128 (.A1(n_0_59), .A2(\Memory[8] [43]), .ZN(n_0_4_1085));
   NAND2_X1 i_0_4_1129 (.A1(n_0_52), .A2(\Memory[1] [43]), .ZN(n_0_4_1086));
   NAND2_X1 i_0_4_1130 (.A1(n_0_61), .A2(\Memory[10] [43]), .ZN(n_0_4_1087));
   NAND3_X1 i_0_4_1131 (.A1(n_0_4_1085), .A2(n_0_4_1086), .A3(n_0_4_1087), 
      .ZN(n_0_4_1088));
   NOR2_X1 i_0_4_1132 (.A1(n_0_4_1084), .A2(n_0_4_1088), .ZN(n_0_4_1089));
   NAND2_X1 i_0_4_1133 (.A1(n_0_65), .A2(\Memory[14] [43]), .ZN(n_0_4_1090));
   NAND2_X1 i_0_4_1134 (.A1(n_0_66), .A2(\Memory[15] [43]), .ZN(n_0_4_1091));
   NAND2_X1 i_0_4_1135 (.A1(n_0_51), .A2(\Memory[0] [43]), .ZN(n_0_4_1092));
   NAND2_X1 i_0_4_1136 (.A1(n_0_60), .A2(\Memory[9] [43]), .ZN(n_0_4_1093));
   NAND4_X1 i_0_4_1137 (.A1(n_0_4_1090), .A2(n_0_4_1091), .A3(n_0_4_1092), 
      .A4(n_0_4_1093), .ZN(n_0_4_1094));
   NAND2_X1 i_0_4_1138 (.A1(n_0_64), .A2(\Memory[13] [43]), .ZN(n_0_4_1095));
   NAND2_X1 i_0_4_1139 (.A1(n_0_63), .A2(\Memory[12] [43]), .ZN(n_0_4_1096));
   NAND2_X1 i_0_4_1140 (.A1(n_0_62), .A2(\Memory[11] [43]), .ZN(n_0_4_1097));
   NAND3_X1 i_0_4_1141 (.A1(n_0_4_1095), .A2(n_0_4_1096), .A3(n_0_4_1097), 
      .ZN(n_0_4_1098));
   NOR2_X1 i_0_4_1142 (.A1(n_0_4_1094), .A2(n_0_4_1098), .ZN(n_0_4_1099));
   NAND3_X1 i_0_4_1143 (.A1(n_0_4_1080), .A2(n_0_4_1089), .A3(n_0_4_1099), 
      .ZN(dataOut2[43]));
   NAND2_X1 i_0_4_1144 (.A1(n_0_55), .A2(\Memory[4] [44]), .ZN(n_0_4_1100));
   NAND2_X1 i_0_4_1145 (.A1(n_0_58), .A2(\Memory[7] [44]), .ZN(n_0_4_1101));
   NAND2_X1 i_0_4_1146 (.A1(n_0_54), .A2(\Memory[3] [44]), .ZN(n_0_4_1102));
   NAND2_X1 i_0_4_1147 (.A1(n_0_53), .A2(\Memory[2] [44]), .ZN(n_0_4_1103));
   NAND4_X1 i_0_4_1148 (.A1(n_0_4_1100), .A2(n_0_4_1101), .A3(n_0_4_1102), 
      .A4(n_0_4_1103), .ZN(n_0_4_1104));
   INV_X1 i_0_4_1149 (.A(n_0_4_1104), .ZN(n_0_4_1105));
   NAND2_X1 i_0_4_1150 (.A1(n_0_67), .A2(\Memory[16] [44]), .ZN(n_0_4_1106));
   NAND2_X1 i_0_4_1151 (.A1(n_0_57), .A2(\Memory[6] [44]), .ZN(n_0_4_1107));
   NAND2_X1 i_0_4_1152 (.A1(n_0_56), .A2(\Memory[5] [44]), .ZN(n_0_4_1108));
   NAND3_X1 i_0_4_1153 (.A1(n_0_4_1106), .A2(n_0_4_1107), .A3(n_0_4_1108), 
      .ZN(n_0_4_1109));
   NAND2_X1 i_0_4_1154 (.A1(n_0_59), .A2(\Memory[8] [44]), .ZN(n_0_4_1110));
   NAND2_X1 i_0_4_1155 (.A1(n_0_52), .A2(\Memory[1] [44]), .ZN(n_0_4_1111));
   NAND2_X1 i_0_4_1156 (.A1(n_0_61), .A2(\Memory[10] [44]), .ZN(n_0_4_1112));
   NAND3_X1 i_0_4_1157 (.A1(n_0_4_1110), .A2(n_0_4_1111), .A3(n_0_4_1112), 
      .ZN(n_0_4_1113));
   NOR2_X1 i_0_4_1158 (.A1(n_0_4_1109), .A2(n_0_4_1113), .ZN(n_0_4_1114));
   NAND2_X1 i_0_4_1159 (.A1(n_0_65), .A2(\Memory[14] [44]), .ZN(n_0_4_1115));
   NAND2_X1 i_0_4_1160 (.A1(n_0_66), .A2(\Memory[15] [44]), .ZN(n_0_4_1116));
   NAND2_X1 i_0_4_1161 (.A1(n_0_51), .A2(\Memory[0] [44]), .ZN(n_0_4_1117));
   NAND2_X1 i_0_4_1162 (.A1(n_0_60), .A2(\Memory[9] [44]), .ZN(n_0_4_1118));
   NAND4_X1 i_0_4_1163 (.A1(n_0_4_1115), .A2(n_0_4_1116), .A3(n_0_4_1117), 
      .A4(n_0_4_1118), .ZN(n_0_4_1119));
   NAND2_X1 i_0_4_1164 (.A1(n_0_64), .A2(\Memory[13] [44]), .ZN(n_0_4_1120));
   NAND2_X1 i_0_4_1165 (.A1(n_0_63), .A2(\Memory[12] [44]), .ZN(n_0_4_1121));
   NAND2_X1 i_0_4_1166 (.A1(n_0_62), .A2(\Memory[11] [44]), .ZN(n_0_4_1122));
   NAND3_X1 i_0_4_1167 (.A1(n_0_4_1120), .A2(n_0_4_1121), .A3(n_0_4_1122), 
      .ZN(n_0_4_1123));
   NOR2_X1 i_0_4_1168 (.A1(n_0_4_1119), .A2(n_0_4_1123), .ZN(n_0_4_1124));
   NAND3_X1 i_0_4_1169 (.A1(n_0_4_1105), .A2(n_0_4_1114), .A3(n_0_4_1124), 
      .ZN(dataOut2[44]));
   NAND2_X1 i_0_4_1170 (.A1(n_0_55), .A2(\Memory[4] [45]), .ZN(n_0_4_1125));
   NAND2_X1 i_0_4_1171 (.A1(n_0_58), .A2(\Memory[7] [45]), .ZN(n_0_4_1126));
   NAND2_X1 i_0_4_1172 (.A1(n_0_54), .A2(\Memory[3] [45]), .ZN(n_0_4_1127));
   NAND2_X1 i_0_4_1173 (.A1(n_0_53), .A2(\Memory[2] [45]), .ZN(n_0_4_1128));
   NAND4_X1 i_0_4_1174 (.A1(n_0_4_1125), .A2(n_0_4_1126), .A3(n_0_4_1127), 
      .A4(n_0_4_1128), .ZN(n_0_4_1129));
   INV_X1 i_0_4_1175 (.A(n_0_4_1129), .ZN(n_0_4_1130));
   NAND2_X1 i_0_4_1176 (.A1(n_0_67), .A2(\Memory[16] [45]), .ZN(n_0_4_1131));
   NAND2_X1 i_0_4_1177 (.A1(n_0_57), .A2(\Memory[6] [45]), .ZN(n_0_4_1132));
   NAND2_X1 i_0_4_1178 (.A1(n_0_56), .A2(\Memory[5] [45]), .ZN(n_0_4_1133));
   NAND3_X1 i_0_4_1179 (.A1(n_0_4_1131), .A2(n_0_4_1132), .A3(n_0_4_1133), 
      .ZN(n_0_4_1134));
   NAND2_X1 i_0_4_1180 (.A1(n_0_59), .A2(\Memory[8] [45]), .ZN(n_0_4_1135));
   NAND2_X1 i_0_4_1181 (.A1(n_0_52), .A2(\Memory[1] [45]), .ZN(n_0_4_1136));
   NAND2_X1 i_0_4_1182 (.A1(n_0_61), .A2(\Memory[10] [45]), .ZN(n_0_4_1137));
   NAND3_X1 i_0_4_1183 (.A1(n_0_4_1135), .A2(n_0_4_1136), .A3(n_0_4_1137), 
      .ZN(n_0_4_1138));
   NOR2_X1 i_0_4_1184 (.A1(n_0_4_1134), .A2(n_0_4_1138), .ZN(n_0_4_1139));
   NAND2_X1 i_0_4_1185 (.A1(n_0_65), .A2(\Memory[14] [45]), .ZN(n_0_4_1140));
   NAND2_X1 i_0_4_1186 (.A1(n_0_66), .A2(\Memory[15] [45]), .ZN(n_0_4_1141));
   NAND2_X1 i_0_4_1187 (.A1(n_0_51), .A2(\Memory[0] [45]), .ZN(n_0_4_1142));
   NAND2_X1 i_0_4_1188 (.A1(n_0_60), .A2(\Memory[9] [45]), .ZN(n_0_4_1143));
   NAND4_X1 i_0_4_1189 (.A1(n_0_4_1140), .A2(n_0_4_1141), .A3(n_0_4_1142), 
      .A4(n_0_4_1143), .ZN(n_0_4_1144));
   NAND2_X1 i_0_4_1190 (.A1(n_0_64), .A2(\Memory[13] [45]), .ZN(n_0_4_1145));
   NAND2_X1 i_0_4_1191 (.A1(n_0_63), .A2(\Memory[12] [45]), .ZN(n_0_4_1146));
   NAND2_X1 i_0_4_1192 (.A1(n_0_62), .A2(\Memory[11] [45]), .ZN(n_0_4_1147));
   NAND3_X1 i_0_4_1193 (.A1(n_0_4_1145), .A2(n_0_4_1146), .A3(n_0_4_1147), 
      .ZN(n_0_4_1148));
   NOR2_X1 i_0_4_1194 (.A1(n_0_4_1144), .A2(n_0_4_1148), .ZN(n_0_4_1149));
   NAND3_X1 i_0_4_1195 (.A1(n_0_4_1130), .A2(n_0_4_1139), .A3(n_0_4_1149), 
      .ZN(dataOut2[45]));
   NAND2_X1 i_0_4_1196 (.A1(n_0_55), .A2(\Memory[4] [46]), .ZN(n_0_4_1150));
   NAND2_X1 i_0_4_1197 (.A1(n_0_58), .A2(\Memory[7] [46]), .ZN(n_0_4_1151));
   NAND2_X1 i_0_4_1198 (.A1(n_0_54), .A2(\Memory[3] [46]), .ZN(n_0_4_1152));
   NAND2_X1 i_0_4_1199 (.A1(n_0_53), .A2(\Memory[2] [46]), .ZN(n_0_4_1153));
   NAND4_X1 i_0_4_1200 (.A1(n_0_4_1150), .A2(n_0_4_1151), .A3(n_0_4_1152), 
      .A4(n_0_4_1153), .ZN(n_0_4_1154));
   INV_X1 i_0_4_1201 (.A(n_0_4_1154), .ZN(n_0_4_1155));
   NAND2_X1 i_0_4_1202 (.A1(n_0_67), .A2(\Memory[16] [46]), .ZN(n_0_4_1156));
   NAND2_X1 i_0_4_1203 (.A1(n_0_57), .A2(\Memory[6] [46]), .ZN(n_0_4_1157));
   NAND2_X1 i_0_4_1204 (.A1(n_0_56), .A2(\Memory[5] [46]), .ZN(n_0_4_1158));
   NAND3_X1 i_0_4_1205 (.A1(n_0_4_1156), .A2(n_0_4_1157), .A3(n_0_4_1158), 
      .ZN(n_0_4_1159));
   NAND2_X1 i_0_4_1206 (.A1(n_0_59), .A2(\Memory[8] [46]), .ZN(n_0_4_1160));
   NAND2_X1 i_0_4_1207 (.A1(n_0_52), .A2(\Memory[1] [46]), .ZN(n_0_4_1161));
   NAND2_X1 i_0_4_1208 (.A1(n_0_61), .A2(\Memory[10] [46]), .ZN(n_0_4_1162));
   NAND3_X1 i_0_4_1209 (.A1(n_0_4_1160), .A2(n_0_4_1161), .A3(n_0_4_1162), 
      .ZN(n_0_4_1163));
   NOR2_X1 i_0_4_1210 (.A1(n_0_4_1159), .A2(n_0_4_1163), .ZN(n_0_4_1164));
   NAND2_X1 i_0_4_1211 (.A1(n_0_65), .A2(\Memory[14] [46]), .ZN(n_0_4_1165));
   NAND2_X1 i_0_4_1212 (.A1(n_0_66), .A2(\Memory[15] [46]), .ZN(n_0_4_1166));
   NAND2_X1 i_0_4_1213 (.A1(n_0_51), .A2(\Memory[0] [46]), .ZN(n_0_4_1167));
   NAND2_X1 i_0_4_1214 (.A1(n_0_60), .A2(\Memory[9] [46]), .ZN(n_0_4_1168));
   NAND4_X1 i_0_4_1215 (.A1(n_0_4_1165), .A2(n_0_4_1166), .A3(n_0_4_1167), 
      .A4(n_0_4_1168), .ZN(n_0_4_1169));
   NAND2_X1 i_0_4_1216 (.A1(n_0_64), .A2(\Memory[13] [46]), .ZN(n_0_4_1170));
   NAND2_X1 i_0_4_1217 (.A1(n_0_63), .A2(\Memory[12] [46]), .ZN(n_0_4_1171));
   NAND2_X1 i_0_4_1218 (.A1(n_0_62), .A2(\Memory[11] [46]), .ZN(n_0_4_1172));
   NAND3_X1 i_0_4_1219 (.A1(n_0_4_1170), .A2(n_0_4_1171), .A3(n_0_4_1172), 
      .ZN(n_0_4_1173));
   NOR2_X1 i_0_4_1220 (.A1(n_0_4_1169), .A2(n_0_4_1173), .ZN(n_0_4_1174));
   NAND3_X1 i_0_4_1221 (.A1(n_0_4_1155), .A2(n_0_4_1164), .A3(n_0_4_1174), 
      .ZN(dataOut2[46]));
   NAND2_X1 i_0_4_1222 (.A1(n_0_55), .A2(\Memory[4] [47]), .ZN(n_0_4_1175));
   NAND2_X1 i_0_4_1223 (.A1(n_0_58), .A2(\Memory[7] [47]), .ZN(n_0_4_1176));
   NAND2_X1 i_0_4_1224 (.A1(n_0_54), .A2(\Memory[3] [47]), .ZN(n_0_4_1177));
   NAND2_X1 i_0_4_1225 (.A1(n_0_53), .A2(\Memory[2] [47]), .ZN(n_0_4_1178));
   NAND4_X1 i_0_4_1226 (.A1(n_0_4_1175), .A2(n_0_4_1176), .A3(n_0_4_1177), 
      .A4(n_0_4_1178), .ZN(n_0_4_1179));
   INV_X1 i_0_4_1227 (.A(n_0_4_1179), .ZN(n_0_4_1180));
   NAND2_X1 i_0_4_1228 (.A1(n_0_67), .A2(\Memory[16] [47]), .ZN(n_0_4_1181));
   NAND2_X1 i_0_4_1229 (.A1(n_0_57), .A2(\Memory[6] [47]), .ZN(n_0_4_1182));
   NAND2_X1 i_0_4_1230 (.A1(n_0_56), .A2(\Memory[5] [47]), .ZN(n_0_4_1183));
   NAND3_X1 i_0_4_1231 (.A1(n_0_4_1181), .A2(n_0_4_1182), .A3(n_0_4_1183), 
      .ZN(n_0_4_1184));
   NAND2_X1 i_0_4_1232 (.A1(n_0_59), .A2(\Memory[8] [47]), .ZN(n_0_4_1185));
   NAND2_X1 i_0_4_1233 (.A1(n_0_52), .A2(\Memory[1] [47]), .ZN(n_0_4_1186));
   NAND2_X1 i_0_4_1234 (.A1(n_0_61), .A2(\Memory[10] [47]), .ZN(n_0_4_1187));
   NAND3_X1 i_0_4_1235 (.A1(n_0_4_1185), .A2(n_0_4_1186), .A3(n_0_4_1187), 
      .ZN(n_0_4_1188));
   NOR2_X1 i_0_4_1236 (.A1(n_0_4_1184), .A2(n_0_4_1188), .ZN(n_0_4_1189));
   NAND2_X1 i_0_4_1237 (.A1(n_0_65), .A2(\Memory[14] [47]), .ZN(n_0_4_1190));
   NAND2_X1 i_0_4_1238 (.A1(n_0_66), .A2(\Memory[15] [47]), .ZN(n_0_4_1191));
   NAND2_X1 i_0_4_1239 (.A1(n_0_51), .A2(\Memory[0] [47]), .ZN(n_0_4_1192));
   NAND2_X1 i_0_4_1240 (.A1(n_0_60), .A2(\Memory[9] [47]), .ZN(n_0_4_1193));
   NAND4_X1 i_0_4_1241 (.A1(n_0_4_1190), .A2(n_0_4_1191), .A3(n_0_4_1192), 
      .A4(n_0_4_1193), .ZN(n_0_4_1194));
   NAND2_X1 i_0_4_1242 (.A1(n_0_64), .A2(\Memory[13] [47]), .ZN(n_0_4_1195));
   NAND2_X1 i_0_4_1243 (.A1(n_0_63), .A2(\Memory[12] [47]), .ZN(n_0_4_1196));
   NAND2_X1 i_0_4_1244 (.A1(n_0_62), .A2(\Memory[11] [47]), .ZN(n_0_4_1197));
   NAND3_X1 i_0_4_1245 (.A1(n_0_4_1195), .A2(n_0_4_1196), .A3(n_0_4_1197), 
      .ZN(n_0_4_1198));
   NOR2_X1 i_0_4_1246 (.A1(n_0_4_1194), .A2(n_0_4_1198), .ZN(n_0_4_1199));
   NAND3_X1 i_0_4_1247 (.A1(n_0_4_1180), .A2(n_0_4_1189), .A3(n_0_4_1199), 
      .ZN(dataOut2[47]));
   NAND2_X1 i_0_4_1248 (.A1(n_0_55), .A2(\Memory[4] [48]), .ZN(n_0_4_1200));
   NAND2_X1 i_0_4_1249 (.A1(n_0_58), .A2(\Memory[7] [48]), .ZN(n_0_4_1201));
   NAND2_X1 i_0_4_1250 (.A1(n_0_54), .A2(\Memory[3] [48]), .ZN(n_0_4_1202));
   NAND2_X1 i_0_4_1251 (.A1(n_0_53), .A2(\Memory[2] [48]), .ZN(n_0_4_1203));
   NAND4_X1 i_0_4_1252 (.A1(n_0_4_1200), .A2(n_0_4_1201), .A3(n_0_4_1202), 
      .A4(n_0_4_1203), .ZN(n_0_4_1204));
   INV_X1 i_0_4_1253 (.A(n_0_4_1204), .ZN(n_0_4_1205));
   NAND2_X1 i_0_4_1254 (.A1(n_0_67), .A2(\Memory[16] [48]), .ZN(n_0_4_1206));
   NAND2_X1 i_0_4_1255 (.A1(n_0_57), .A2(\Memory[6] [48]), .ZN(n_0_4_1207));
   NAND2_X1 i_0_4_1256 (.A1(n_0_56), .A2(\Memory[5] [48]), .ZN(n_0_4_1208));
   NAND3_X1 i_0_4_1257 (.A1(n_0_4_1206), .A2(n_0_4_1207), .A3(n_0_4_1208), 
      .ZN(n_0_4_1209));
   NAND2_X1 i_0_4_1258 (.A1(n_0_59), .A2(\Memory[8] [48]), .ZN(n_0_4_1210));
   NAND2_X1 i_0_4_1259 (.A1(n_0_52), .A2(\Memory[1] [48]), .ZN(n_0_4_1211));
   NAND2_X1 i_0_4_1260 (.A1(n_0_61), .A2(\Memory[10] [48]), .ZN(n_0_4_1212));
   NAND3_X1 i_0_4_1261 (.A1(n_0_4_1210), .A2(n_0_4_1211), .A3(n_0_4_1212), 
      .ZN(n_0_4_1213));
   NOR2_X1 i_0_4_1262 (.A1(n_0_4_1209), .A2(n_0_4_1213), .ZN(n_0_4_1214));
   NAND2_X1 i_0_4_1263 (.A1(n_0_65), .A2(\Memory[14] [48]), .ZN(n_0_4_1215));
   NAND2_X1 i_0_4_1264 (.A1(n_0_66), .A2(\Memory[15] [48]), .ZN(n_0_4_1216));
   NAND2_X1 i_0_4_1265 (.A1(n_0_51), .A2(\Memory[0] [48]), .ZN(n_0_4_1217));
   NAND2_X1 i_0_4_1266 (.A1(n_0_60), .A2(\Memory[9] [48]), .ZN(n_0_4_1218));
   NAND4_X1 i_0_4_1267 (.A1(n_0_4_1215), .A2(n_0_4_1216), .A3(n_0_4_1217), 
      .A4(n_0_4_1218), .ZN(n_0_4_1219));
   NAND2_X1 i_0_4_1268 (.A1(n_0_64), .A2(\Memory[13] [48]), .ZN(n_0_4_1220));
   NAND2_X1 i_0_4_1269 (.A1(n_0_63), .A2(\Memory[12] [48]), .ZN(n_0_4_1221));
   NAND2_X1 i_0_4_1270 (.A1(n_0_62), .A2(\Memory[11] [48]), .ZN(n_0_4_1222));
   NAND3_X1 i_0_4_1271 (.A1(n_0_4_1220), .A2(n_0_4_1221), .A3(n_0_4_1222), 
      .ZN(n_0_4_1223));
   NOR2_X1 i_0_4_1272 (.A1(n_0_4_1219), .A2(n_0_4_1223), .ZN(n_0_4_1224));
   NAND3_X1 i_0_4_1273 (.A1(n_0_4_1205), .A2(n_0_4_1214), .A3(n_0_4_1224), 
      .ZN(dataOut2[48]));
   NAND2_X1 i_0_4_1274 (.A1(n_0_55), .A2(\Memory[4] [49]), .ZN(n_0_4_1225));
   NAND2_X1 i_0_4_1275 (.A1(n_0_58), .A2(\Memory[7] [49]), .ZN(n_0_4_1226));
   NAND2_X1 i_0_4_1276 (.A1(n_0_54), .A2(\Memory[3] [49]), .ZN(n_0_4_1227));
   NAND2_X1 i_0_4_1277 (.A1(n_0_53), .A2(\Memory[2] [49]), .ZN(n_0_4_1228));
   NAND4_X1 i_0_4_1278 (.A1(n_0_4_1225), .A2(n_0_4_1226), .A3(n_0_4_1227), 
      .A4(n_0_4_1228), .ZN(n_0_4_1229));
   INV_X1 i_0_4_1279 (.A(n_0_4_1229), .ZN(n_0_4_1230));
   NAND2_X1 i_0_4_1280 (.A1(n_0_67), .A2(\Memory[16] [49]), .ZN(n_0_4_1231));
   NAND2_X1 i_0_4_1281 (.A1(n_0_57), .A2(\Memory[6] [49]), .ZN(n_0_4_1232));
   NAND2_X1 i_0_4_1282 (.A1(n_0_56), .A2(\Memory[5] [49]), .ZN(n_0_4_1233));
   NAND3_X1 i_0_4_1283 (.A1(n_0_4_1231), .A2(n_0_4_1232), .A3(n_0_4_1233), 
      .ZN(n_0_4_1234));
   NAND2_X1 i_0_4_1284 (.A1(n_0_59), .A2(\Memory[8] [49]), .ZN(n_0_4_1235));
   NAND2_X1 i_0_4_1285 (.A1(n_0_52), .A2(\Memory[1] [49]), .ZN(n_0_4_1236));
   NAND2_X1 i_0_4_1286 (.A1(n_0_61), .A2(\Memory[10] [49]), .ZN(n_0_4_1237));
   NAND3_X1 i_0_4_1287 (.A1(n_0_4_1235), .A2(n_0_4_1236), .A3(n_0_4_1237), 
      .ZN(n_0_4_1238));
   NOR2_X1 i_0_4_1288 (.A1(n_0_4_1234), .A2(n_0_4_1238), .ZN(n_0_4_1239));
   NAND2_X1 i_0_4_1289 (.A1(n_0_65), .A2(\Memory[14] [49]), .ZN(n_0_4_1240));
   NAND2_X1 i_0_4_1290 (.A1(n_0_66), .A2(\Memory[15] [49]), .ZN(n_0_4_1241));
   NAND2_X1 i_0_4_1291 (.A1(n_0_51), .A2(\Memory[0] [49]), .ZN(n_0_4_1242));
   NAND2_X1 i_0_4_1292 (.A1(n_0_60), .A2(\Memory[9] [49]), .ZN(n_0_4_1243));
   NAND4_X1 i_0_4_1293 (.A1(n_0_4_1240), .A2(n_0_4_1241), .A3(n_0_4_1242), 
      .A4(n_0_4_1243), .ZN(n_0_4_1244));
   NAND2_X1 i_0_4_1294 (.A1(n_0_64), .A2(\Memory[13] [49]), .ZN(n_0_4_1245));
   NAND2_X1 i_0_4_1295 (.A1(n_0_63), .A2(\Memory[12] [49]), .ZN(n_0_4_1246));
   NAND2_X1 i_0_4_1296 (.A1(n_0_62), .A2(\Memory[11] [49]), .ZN(n_0_4_1247));
   NAND3_X1 i_0_4_1297 (.A1(n_0_4_1245), .A2(n_0_4_1246), .A3(n_0_4_1247), 
      .ZN(n_0_4_1248));
   NOR2_X1 i_0_4_1298 (.A1(n_0_4_1244), .A2(n_0_4_1248), .ZN(n_0_4_1249));
   NAND3_X1 i_0_4_1299 (.A1(n_0_4_1230), .A2(n_0_4_1239), .A3(n_0_4_1249), 
      .ZN(dataOut2[49]));
   NAND2_X1 i_0_4_1300 (.A1(n_0_55), .A2(\Memory[4] [50]), .ZN(n_0_4_1250));
   NAND2_X1 i_0_4_1301 (.A1(n_0_58), .A2(\Memory[7] [50]), .ZN(n_0_4_1251));
   NAND2_X1 i_0_4_1302 (.A1(n_0_54), .A2(\Memory[3] [50]), .ZN(n_0_4_1252));
   NAND2_X1 i_0_4_1303 (.A1(n_0_53), .A2(\Memory[2] [50]), .ZN(n_0_4_1253));
   NAND4_X1 i_0_4_1304 (.A1(n_0_4_1250), .A2(n_0_4_1251), .A3(n_0_4_1252), 
      .A4(n_0_4_1253), .ZN(n_0_4_1254));
   INV_X1 i_0_4_1305 (.A(n_0_4_1254), .ZN(n_0_4_1255));
   NAND2_X1 i_0_4_1306 (.A1(n_0_67), .A2(\Memory[16] [50]), .ZN(n_0_4_1256));
   NAND2_X1 i_0_4_1307 (.A1(n_0_57), .A2(\Memory[6] [50]), .ZN(n_0_4_1257));
   NAND2_X1 i_0_4_1308 (.A1(n_0_56), .A2(\Memory[5] [50]), .ZN(n_0_4_1258));
   NAND3_X1 i_0_4_1309 (.A1(n_0_4_1256), .A2(n_0_4_1257), .A3(n_0_4_1258), 
      .ZN(n_0_4_1259));
   NAND2_X1 i_0_4_1310 (.A1(n_0_59), .A2(\Memory[8] [50]), .ZN(n_0_4_1260));
   NAND2_X1 i_0_4_1311 (.A1(n_0_52), .A2(\Memory[1] [50]), .ZN(n_0_4_1261));
   NAND2_X1 i_0_4_1312 (.A1(n_0_61), .A2(\Memory[10] [50]), .ZN(n_0_4_1262));
   NAND3_X1 i_0_4_1313 (.A1(n_0_4_1260), .A2(n_0_4_1261), .A3(n_0_4_1262), 
      .ZN(n_0_4_1263));
   NOR2_X1 i_0_4_1314 (.A1(n_0_4_1259), .A2(n_0_4_1263), .ZN(n_0_4_1264));
   NAND2_X1 i_0_4_1315 (.A1(n_0_65), .A2(\Memory[14] [50]), .ZN(n_0_4_1265));
   NAND2_X1 i_0_4_1316 (.A1(n_0_66), .A2(\Memory[15] [50]), .ZN(n_0_4_1266));
   NAND2_X1 i_0_4_1317 (.A1(n_0_51), .A2(\Memory[0] [50]), .ZN(n_0_4_1267));
   NAND2_X1 i_0_4_1318 (.A1(n_0_60), .A2(\Memory[9] [50]), .ZN(n_0_4_1268));
   NAND4_X1 i_0_4_1319 (.A1(n_0_4_1265), .A2(n_0_4_1266), .A3(n_0_4_1267), 
      .A4(n_0_4_1268), .ZN(n_0_4_1269));
   NAND2_X1 i_0_4_1320 (.A1(n_0_64), .A2(\Memory[13] [50]), .ZN(n_0_4_1270));
   NAND2_X1 i_0_4_1321 (.A1(n_0_63), .A2(\Memory[12] [50]), .ZN(n_0_4_1271));
   NAND2_X1 i_0_4_1322 (.A1(n_0_62), .A2(\Memory[11] [50]), .ZN(n_0_4_1272));
   NAND3_X1 i_0_4_1323 (.A1(n_0_4_1270), .A2(n_0_4_1271), .A3(n_0_4_1272), 
      .ZN(n_0_4_1273));
   NOR2_X1 i_0_4_1324 (.A1(n_0_4_1269), .A2(n_0_4_1273), .ZN(n_0_4_1274));
   NAND3_X1 i_0_4_1325 (.A1(n_0_4_1255), .A2(n_0_4_1264), .A3(n_0_4_1274), 
      .ZN(dataOut2[50]));
   NAND2_X1 i_0_4_1326 (.A1(n_0_55), .A2(\Memory[4] [51]), .ZN(n_0_4_1275));
   NAND2_X1 i_0_4_1327 (.A1(n_0_58), .A2(\Memory[7] [51]), .ZN(n_0_4_1276));
   NAND2_X1 i_0_4_1328 (.A1(n_0_54), .A2(\Memory[3] [51]), .ZN(n_0_4_1277));
   NAND2_X1 i_0_4_1329 (.A1(n_0_53), .A2(\Memory[2] [51]), .ZN(n_0_4_1278));
   NAND4_X1 i_0_4_1330 (.A1(n_0_4_1275), .A2(n_0_4_1276), .A3(n_0_4_1277), 
      .A4(n_0_4_1278), .ZN(n_0_4_1279));
   INV_X1 i_0_4_1331 (.A(n_0_4_1279), .ZN(n_0_4_1280));
   NAND2_X1 i_0_4_1332 (.A1(n_0_67), .A2(\Memory[16] [51]), .ZN(n_0_4_1281));
   NAND2_X1 i_0_4_1333 (.A1(n_0_57), .A2(\Memory[6] [51]), .ZN(n_0_4_1282));
   NAND2_X1 i_0_4_1334 (.A1(n_0_56), .A2(\Memory[5] [51]), .ZN(n_0_4_1283));
   NAND3_X1 i_0_4_1335 (.A1(n_0_4_1281), .A2(n_0_4_1282), .A3(n_0_4_1283), 
      .ZN(n_0_4_1284));
   NAND2_X1 i_0_4_1336 (.A1(n_0_59), .A2(\Memory[8] [51]), .ZN(n_0_4_1285));
   NAND2_X1 i_0_4_1337 (.A1(n_0_52), .A2(\Memory[1] [51]), .ZN(n_0_4_1286));
   NAND2_X1 i_0_4_1338 (.A1(n_0_61), .A2(\Memory[10] [51]), .ZN(n_0_4_1287));
   NAND3_X1 i_0_4_1339 (.A1(n_0_4_1285), .A2(n_0_4_1286), .A3(n_0_4_1287), 
      .ZN(n_0_4_1288));
   NOR2_X1 i_0_4_1340 (.A1(n_0_4_1284), .A2(n_0_4_1288), .ZN(n_0_4_1289));
   NAND2_X1 i_0_4_1341 (.A1(n_0_65), .A2(\Memory[14] [51]), .ZN(n_0_4_1290));
   NAND2_X1 i_0_4_1342 (.A1(n_0_66), .A2(\Memory[15] [51]), .ZN(n_0_4_1291));
   NAND2_X1 i_0_4_1343 (.A1(n_0_51), .A2(\Memory[0] [51]), .ZN(n_0_4_1292));
   NAND2_X1 i_0_4_1344 (.A1(n_0_60), .A2(\Memory[9] [51]), .ZN(n_0_4_1293));
   NAND4_X1 i_0_4_1345 (.A1(n_0_4_1290), .A2(n_0_4_1291), .A3(n_0_4_1292), 
      .A4(n_0_4_1293), .ZN(n_0_4_1294));
   NAND2_X1 i_0_4_1346 (.A1(n_0_64), .A2(\Memory[13] [51]), .ZN(n_0_4_1295));
   NAND2_X1 i_0_4_1347 (.A1(n_0_63), .A2(\Memory[12] [51]), .ZN(n_0_4_1296));
   NAND2_X1 i_0_4_1348 (.A1(n_0_62), .A2(\Memory[11] [51]), .ZN(n_0_4_1297));
   NAND3_X1 i_0_4_1349 (.A1(n_0_4_1295), .A2(n_0_4_1296), .A3(n_0_4_1297), 
      .ZN(n_0_4_1298));
   NOR2_X1 i_0_4_1350 (.A1(n_0_4_1294), .A2(n_0_4_1298), .ZN(n_0_4_1299));
   NAND3_X1 i_0_4_1351 (.A1(n_0_4_1280), .A2(n_0_4_1289), .A3(n_0_4_1299), 
      .ZN(dataOut2[51]));
   NAND2_X1 i_0_4_1352 (.A1(n_0_55), .A2(\Memory[4] [52]), .ZN(n_0_4_1300));
   NAND2_X1 i_0_4_1353 (.A1(n_0_58), .A2(\Memory[7] [52]), .ZN(n_0_4_1301));
   NAND2_X1 i_0_4_1354 (.A1(n_0_54), .A2(\Memory[3] [52]), .ZN(n_0_4_1302));
   NAND2_X1 i_0_4_1355 (.A1(n_0_53), .A2(\Memory[2] [52]), .ZN(n_0_4_1303));
   NAND4_X1 i_0_4_1356 (.A1(n_0_4_1300), .A2(n_0_4_1301), .A3(n_0_4_1302), 
      .A4(n_0_4_1303), .ZN(n_0_4_1304));
   INV_X1 i_0_4_1357 (.A(n_0_4_1304), .ZN(n_0_4_1305));
   NAND2_X1 i_0_4_1358 (.A1(n_0_67), .A2(\Memory[16] [52]), .ZN(n_0_4_1306));
   NAND2_X1 i_0_4_1359 (.A1(n_0_57), .A2(\Memory[6] [52]), .ZN(n_0_4_1307));
   NAND2_X1 i_0_4_1360 (.A1(n_0_56), .A2(\Memory[5] [52]), .ZN(n_0_4_1308));
   NAND3_X1 i_0_4_1361 (.A1(n_0_4_1306), .A2(n_0_4_1307), .A3(n_0_4_1308), 
      .ZN(n_0_4_1309));
   NAND2_X1 i_0_4_1362 (.A1(n_0_59), .A2(\Memory[8] [52]), .ZN(n_0_4_1310));
   NAND2_X1 i_0_4_1363 (.A1(n_0_52), .A2(\Memory[1] [52]), .ZN(n_0_4_1311));
   NAND2_X1 i_0_4_1364 (.A1(n_0_61), .A2(\Memory[10] [52]), .ZN(n_0_4_1312));
   NAND3_X1 i_0_4_1365 (.A1(n_0_4_1310), .A2(n_0_4_1311), .A3(n_0_4_1312), 
      .ZN(n_0_4_1313));
   NOR2_X1 i_0_4_1366 (.A1(n_0_4_1309), .A2(n_0_4_1313), .ZN(n_0_4_1314));
   NAND2_X1 i_0_4_1367 (.A1(n_0_65), .A2(\Memory[14] [52]), .ZN(n_0_4_1315));
   NAND2_X1 i_0_4_1368 (.A1(n_0_66), .A2(\Memory[15] [52]), .ZN(n_0_4_1316));
   NAND2_X1 i_0_4_1369 (.A1(n_0_51), .A2(\Memory[0] [52]), .ZN(n_0_4_1317));
   NAND2_X1 i_0_4_1370 (.A1(n_0_60), .A2(\Memory[9] [52]), .ZN(n_0_4_1318));
   NAND4_X1 i_0_4_1371 (.A1(n_0_4_1315), .A2(n_0_4_1316), .A3(n_0_4_1317), 
      .A4(n_0_4_1318), .ZN(n_0_4_1319));
   NAND2_X1 i_0_4_1372 (.A1(n_0_64), .A2(\Memory[13] [52]), .ZN(n_0_4_1320));
   NAND2_X1 i_0_4_1373 (.A1(n_0_63), .A2(\Memory[12] [52]), .ZN(n_0_4_1321));
   NAND2_X1 i_0_4_1374 (.A1(n_0_62), .A2(\Memory[11] [52]), .ZN(n_0_4_1322));
   NAND3_X1 i_0_4_1375 (.A1(n_0_4_1320), .A2(n_0_4_1321), .A3(n_0_4_1322), 
      .ZN(n_0_4_1323));
   NOR2_X1 i_0_4_1376 (.A1(n_0_4_1319), .A2(n_0_4_1323), .ZN(n_0_4_1324));
   NAND3_X1 i_0_4_1377 (.A1(n_0_4_1305), .A2(n_0_4_1314), .A3(n_0_4_1324), 
      .ZN(dataOut2[52]));
   NAND2_X1 i_0_4_1378 (.A1(n_0_55), .A2(\Memory[4] [53]), .ZN(n_0_4_1325));
   NAND2_X1 i_0_4_1379 (.A1(n_0_58), .A2(\Memory[7] [53]), .ZN(n_0_4_1326));
   NAND2_X1 i_0_4_1380 (.A1(n_0_54), .A2(\Memory[3] [53]), .ZN(n_0_4_1327));
   NAND2_X1 i_0_4_1381 (.A1(n_0_53), .A2(\Memory[2] [53]), .ZN(n_0_4_1328));
   NAND4_X1 i_0_4_1382 (.A1(n_0_4_1325), .A2(n_0_4_1326), .A3(n_0_4_1327), 
      .A4(n_0_4_1328), .ZN(n_0_4_1329));
   INV_X1 i_0_4_1383 (.A(n_0_4_1329), .ZN(n_0_4_1330));
   NAND2_X1 i_0_4_1384 (.A1(n_0_67), .A2(\Memory[16] [53]), .ZN(n_0_4_1331));
   NAND2_X1 i_0_4_1385 (.A1(n_0_57), .A2(\Memory[6] [53]), .ZN(n_0_4_1332));
   NAND2_X1 i_0_4_1386 (.A1(n_0_56), .A2(\Memory[5] [53]), .ZN(n_0_4_1333));
   NAND3_X1 i_0_4_1387 (.A1(n_0_4_1331), .A2(n_0_4_1332), .A3(n_0_4_1333), 
      .ZN(n_0_4_1334));
   NAND2_X1 i_0_4_1388 (.A1(n_0_59), .A2(\Memory[8] [53]), .ZN(n_0_4_1335));
   NAND2_X1 i_0_4_1389 (.A1(n_0_52), .A2(\Memory[1] [53]), .ZN(n_0_4_1336));
   NAND2_X1 i_0_4_1390 (.A1(n_0_61), .A2(\Memory[10] [53]), .ZN(n_0_4_1337));
   NAND3_X1 i_0_4_1391 (.A1(n_0_4_1335), .A2(n_0_4_1336), .A3(n_0_4_1337), 
      .ZN(n_0_4_1338));
   NOR2_X1 i_0_4_1392 (.A1(n_0_4_1334), .A2(n_0_4_1338), .ZN(n_0_4_1339));
   NAND2_X1 i_0_4_1393 (.A1(n_0_65), .A2(\Memory[14] [53]), .ZN(n_0_4_1340));
   NAND2_X1 i_0_4_1394 (.A1(n_0_66), .A2(\Memory[15] [53]), .ZN(n_0_4_1341));
   NAND2_X1 i_0_4_1395 (.A1(n_0_51), .A2(\Memory[0] [53]), .ZN(n_0_4_1342));
   NAND2_X1 i_0_4_1396 (.A1(n_0_60), .A2(\Memory[9] [53]), .ZN(n_0_4_1343));
   NAND4_X1 i_0_4_1397 (.A1(n_0_4_1340), .A2(n_0_4_1341), .A3(n_0_4_1342), 
      .A4(n_0_4_1343), .ZN(n_0_4_1344));
   NAND2_X1 i_0_4_1398 (.A1(n_0_64), .A2(\Memory[13] [53]), .ZN(n_0_4_1345));
   NAND2_X1 i_0_4_1399 (.A1(n_0_63), .A2(\Memory[12] [53]), .ZN(n_0_4_1346));
   NAND2_X1 i_0_4_1400 (.A1(n_0_62), .A2(\Memory[11] [53]), .ZN(n_0_4_1347));
   NAND3_X1 i_0_4_1401 (.A1(n_0_4_1345), .A2(n_0_4_1346), .A3(n_0_4_1347), 
      .ZN(n_0_4_1348));
   NOR2_X1 i_0_4_1402 (.A1(n_0_4_1344), .A2(n_0_4_1348), .ZN(n_0_4_1349));
   NAND3_X1 i_0_4_1403 (.A1(n_0_4_1330), .A2(n_0_4_1339), .A3(n_0_4_1349), 
      .ZN(dataOut2[53]));
   NAND2_X1 i_0_4_1404 (.A1(n_0_55), .A2(\Memory[4] [54]), .ZN(n_0_4_1350));
   NAND2_X1 i_0_4_1405 (.A1(n_0_58), .A2(\Memory[7] [54]), .ZN(n_0_4_1351));
   NAND2_X1 i_0_4_1406 (.A1(n_0_54), .A2(\Memory[3] [54]), .ZN(n_0_4_1352));
   NAND2_X1 i_0_4_1407 (.A1(n_0_53), .A2(\Memory[2] [54]), .ZN(n_0_4_1353));
   NAND4_X1 i_0_4_1408 (.A1(n_0_4_1350), .A2(n_0_4_1351), .A3(n_0_4_1352), 
      .A4(n_0_4_1353), .ZN(n_0_4_1354));
   INV_X1 i_0_4_1409 (.A(n_0_4_1354), .ZN(n_0_4_1355));
   NAND2_X1 i_0_4_1410 (.A1(n_0_67), .A2(\Memory[16] [54]), .ZN(n_0_4_1356));
   NAND2_X1 i_0_4_1411 (.A1(n_0_57), .A2(\Memory[6] [54]), .ZN(n_0_4_1357));
   NAND2_X1 i_0_4_1412 (.A1(n_0_56), .A2(\Memory[5] [54]), .ZN(n_0_4_1358));
   NAND3_X1 i_0_4_1413 (.A1(n_0_4_1356), .A2(n_0_4_1357), .A3(n_0_4_1358), 
      .ZN(n_0_4_1359));
   NAND2_X1 i_0_4_1414 (.A1(n_0_59), .A2(\Memory[8] [54]), .ZN(n_0_4_1360));
   NAND2_X1 i_0_4_1415 (.A1(n_0_52), .A2(\Memory[1] [54]), .ZN(n_0_4_1361));
   NAND2_X1 i_0_4_1416 (.A1(n_0_61), .A2(\Memory[10] [54]), .ZN(n_0_4_1362));
   NAND3_X1 i_0_4_1417 (.A1(n_0_4_1360), .A2(n_0_4_1361), .A3(n_0_4_1362), 
      .ZN(n_0_4_1363));
   NOR2_X1 i_0_4_1418 (.A1(n_0_4_1359), .A2(n_0_4_1363), .ZN(n_0_4_1364));
   NAND2_X1 i_0_4_1419 (.A1(n_0_65), .A2(\Memory[14] [54]), .ZN(n_0_4_1365));
   NAND2_X1 i_0_4_1420 (.A1(n_0_66), .A2(\Memory[15] [54]), .ZN(n_0_4_1366));
   NAND2_X1 i_0_4_1421 (.A1(n_0_51), .A2(\Memory[0] [54]), .ZN(n_0_4_1367));
   NAND2_X1 i_0_4_1422 (.A1(n_0_60), .A2(\Memory[9] [54]), .ZN(n_0_4_1368));
   NAND4_X1 i_0_4_1423 (.A1(n_0_4_1365), .A2(n_0_4_1366), .A3(n_0_4_1367), 
      .A4(n_0_4_1368), .ZN(n_0_4_1369));
   NAND2_X1 i_0_4_1424 (.A1(n_0_64), .A2(\Memory[13] [54]), .ZN(n_0_4_1370));
   NAND2_X1 i_0_4_1425 (.A1(n_0_63), .A2(\Memory[12] [54]), .ZN(n_0_4_1371));
   NAND2_X1 i_0_4_1426 (.A1(n_0_62), .A2(\Memory[11] [54]), .ZN(n_0_4_1372));
   NAND3_X1 i_0_4_1427 (.A1(n_0_4_1370), .A2(n_0_4_1371), .A3(n_0_4_1372), 
      .ZN(n_0_4_1373));
   NOR2_X1 i_0_4_1428 (.A1(n_0_4_1369), .A2(n_0_4_1373), .ZN(n_0_4_1374));
   NAND3_X1 i_0_4_1429 (.A1(n_0_4_1355), .A2(n_0_4_1364), .A3(n_0_4_1374), 
      .ZN(dataOut2[54]));
   NAND2_X1 i_0_4_1430 (.A1(n_0_55), .A2(\Memory[4] [55]), .ZN(n_0_4_1375));
   NAND2_X1 i_0_4_1431 (.A1(n_0_58), .A2(\Memory[7] [55]), .ZN(n_0_4_1376));
   NAND2_X1 i_0_4_1432 (.A1(n_0_54), .A2(\Memory[3] [55]), .ZN(n_0_4_1377));
   NAND2_X1 i_0_4_1433 (.A1(n_0_53), .A2(\Memory[2] [55]), .ZN(n_0_4_1378));
   NAND4_X1 i_0_4_1434 (.A1(n_0_4_1375), .A2(n_0_4_1376), .A3(n_0_4_1377), 
      .A4(n_0_4_1378), .ZN(n_0_4_1379));
   INV_X1 i_0_4_1435 (.A(n_0_4_1379), .ZN(n_0_4_1380));
   NAND2_X1 i_0_4_1436 (.A1(n_0_67), .A2(\Memory[16] [55]), .ZN(n_0_4_1381));
   NAND2_X1 i_0_4_1437 (.A1(n_0_57), .A2(\Memory[6] [55]), .ZN(n_0_4_1382));
   NAND2_X1 i_0_4_1438 (.A1(n_0_56), .A2(\Memory[5] [55]), .ZN(n_0_4_1383));
   NAND3_X1 i_0_4_1439 (.A1(n_0_4_1381), .A2(n_0_4_1382), .A3(n_0_4_1383), 
      .ZN(n_0_4_1384));
   NAND2_X1 i_0_4_1440 (.A1(n_0_59), .A2(\Memory[8] [55]), .ZN(n_0_4_1385));
   NAND2_X1 i_0_4_1441 (.A1(n_0_52), .A2(\Memory[1] [55]), .ZN(n_0_4_1386));
   NAND2_X1 i_0_4_1442 (.A1(n_0_61), .A2(\Memory[10] [55]), .ZN(n_0_4_1387));
   NAND3_X1 i_0_4_1443 (.A1(n_0_4_1385), .A2(n_0_4_1386), .A3(n_0_4_1387), 
      .ZN(n_0_4_1388));
   NOR2_X1 i_0_4_1444 (.A1(n_0_4_1384), .A2(n_0_4_1388), .ZN(n_0_4_1389));
   NAND2_X1 i_0_4_1445 (.A1(n_0_65), .A2(\Memory[14] [55]), .ZN(n_0_4_1390));
   NAND2_X1 i_0_4_1446 (.A1(n_0_66), .A2(\Memory[15] [55]), .ZN(n_0_4_1391));
   NAND2_X1 i_0_4_1447 (.A1(n_0_51), .A2(\Memory[0] [55]), .ZN(n_0_4_1392));
   NAND2_X1 i_0_4_1448 (.A1(n_0_60), .A2(\Memory[9] [55]), .ZN(n_0_4_1393));
   NAND4_X1 i_0_4_1449 (.A1(n_0_4_1390), .A2(n_0_4_1391), .A3(n_0_4_1392), 
      .A4(n_0_4_1393), .ZN(n_0_4_1394));
   NAND2_X1 i_0_4_1450 (.A1(n_0_64), .A2(\Memory[13] [55]), .ZN(n_0_4_1395));
   NAND2_X1 i_0_4_1451 (.A1(n_0_63), .A2(\Memory[12] [55]), .ZN(n_0_4_1396));
   NAND2_X1 i_0_4_1452 (.A1(n_0_62), .A2(\Memory[11] [55]), .ZN(n_0_4_1397));
   NAND3_X1 i_0_4_1453 (.A1(n_0_4_1395), .A2(n_0_4_1396), .A3(n_0_4_1397), 
      .ZN(n_0_4_1398));
   NOR2_X1 i_0_4_1454 (.A1(n_0_4_1394), .A2(n_0_4_1398), .ZN(n_0_4_1399));
   NAND3_X1 i_0_4_1455 (.A1(n_0_4_1380), .A2(n_0_4_1389), .A3(n_0_4_1399), 
      .ZN(dataOut2[55]));
   NAND2_X1 i_0_4_1456 (.A1(n_0_55), .A2(\Memory[4] [56]), .ZN(n_0_4_1400));
   NAND2_X1 i_0_4_1457 (.A1(n_0_58), .A2(\Memory[7] [56]), .ZN(n_0_4_1401));
   NAND2_X1 i_0_4_1458 (.A1(n_0_54), .A2(\Memory[3] [56]), .ZN(n_0_4_1402));
   NAND2_X1 i_0_4_1459 (.A1(n_0_53), .A2(\Memory[2] [56]), .ZN(n_0_4_1403));
   NAND4_X1 i_0_4_1460 (.A1(n_0_4_1400), .A2(n_0_4_1401), .A3(n_0_4_1402), 
      .A4(n_0_4_1403), .ZN(n_0_4_1404));
   INV_X1 i_0_4_1461 (.A(n_0_4_1404), .ZN(n_0_4_1405));
   NAND2_X1 i_0_4_1462 (.A1(n_0_67), .A2(\Memory[16] [56]), .ZN(n_0_4_1406));
   NAND2_X1 i_0_4_1463 (.A1(n_0_57), .A2(\Memory[6] [56]), .ZN(n_0_4_1407));
   NAND2_X1 i_0_4_1464 (.A1(n_0_56), .A2(\Memory[5] [56]), .ZN(n_0_4_1408));
   NAND3_X1 i_0_4_1465 (.A1(n_0_4_1406), .A2(n_0_4_1407), .A3(n_0_4_1408), 
      .ZN(n_0_4_1409));
   NAND2_X1 i_0_4_1466 (.A1(n_0_59), .A2(\Memory[8] [56]), .ZN(n_0_4_1410));
   NAND2_X1 i_0_4_1467 (.A1(n_0_52), .A2(\Memory[1] [56]), .ZN(n_0_4_1411));
   NAND2_X1 i_0_4_1468 (.A1(n_0_61), .A2(\Memory[10] [56]), .ZN(n_0_4_1412));
   NAND3_X1 i_0_4_1469 (.A1(n_0_4_1410), .A2(n_0_4_1411), .A3(n_0_4_1412), 
      .ZN(n_0_4_1413));
   NOR2_X1 i_0_4_1470 (.A1(n_0_4_1409), .A2(n_0_4_1413), .ZN(n_0_4_1414));
   NAND2_X1 i_0_4_1471 (.A1(n_0_65), .A2(\Memory[14] [56]), .ZN(n_0_4_1415));
   NAND2_X1 i_0_4_1472 (.A1(n_0_66), .A2(\Memory[15] [56]), .ZN(n_0_4_1416));
   NAND2_X1 i_0_4_1473 (.A1(n_0_51), .A2(\Memory[0] [56]), .ZN(n_0_4_1417));
   NAND2_X1 i_0_4_1474 (.A1(n_0_60), .A2(\Memory[9] [56]), .ZN(n_0_4_1418));
   NAND4_X1 i_0_4_1475 (.A1(n_0_4_1415), .A2(n_0_4_1416), .A3(n_0_4_1417), 
      .A4(n_0_4_1418), .ZN(n_0_4_1419));
   NAND2_X1 i_0_4_1476 (.A1(n_0_64), .A2(\Memory[13] [56]), .ZN(n_0_4_1420));
   NAND2_X1 i_0_4_1477 (.A1(n_0_63), .A2(\Memory[12] [56]), .ZN(n_0_4_1421));
   NAND2_X1 i_0_4_1478 (.A1(n_0_62), .A2(\Memory[11] [56]), .ZN(n_0_4_1422));
   NAND3_X1 i_0_4_1479 (.A1(n_0_4_1420), .A2(n_0_4_1421), .A3(n_0_4_1422), 
      .ZN(n_0_4_1423));
   NOR2_X1 i_0_4_1480 (.A1(n_0_4_1419), .A2(n_0_4_1423), .ZN(n_0_4_1424));
   NAND3_X1 i_0_4_1481 (.A1(n_0_4_1405), .A2(n_0_4_1414), .A3(n_0_4_1424), 
      .ZN(dataOut2[56]));
   NAND2_X1 i_0_4_1482 (.A1(n_0_55), .A2(\Memory[4] [57]), .ZN(n_0_4_1425));
   NAND2_X1 i_0_4_1483 (.A1(n_0_58), .A2(\Memory[7] [57]), .ZN(n_0_4_1426));
   NAND2_X1 i_0_4_1484 (.A1(n_0_54), .A2(\Memory[3] [57]), .ZN(n_0_4_1427));
   NAND2_X1 i_0_4_1485 (.A1(n_0_53), .A2(\Memory[2] [57]), .ZN(n_0_4_1428));
   NAND4_X1 i_0_4_1486 (.A1(n_0_4_1425), .A2(n_0_4_1426), .A3(n_0_4_1427), 
      .A4(n_0_4_1428), .ZN(n_0_4_1429));
   INV_X1 i_0_4_1487 (.A(n_0_4_1429), .ZN(n_0_4_1430));
   NAND2_X1 i_0_4_1488 (.A1(n_0_67), .A2(\Memory[16] [57]), .ZN(n_0_4_1431));
   NAND2_X1 i_0_4_1489 (.A1(n_0_57), .A2(\Memory[6] [57]), .ZN(n_0_4_1432));
   NAND2_X1 i_0_4_1490 (.A1(n_0_56), .A2(\Memory[5] [57]), .ZN(n_0_4_1433));
   NAND3_X1 i_0_4_1491 (.A1(n_0_4_1431), .A2(n_0_4_1432), .A3(n_0_4_1433), 
      .ZN(n_0_4_1434));
   NAND2_X1 i_0_4_1492 (.A1(n_0_59), .A2(\Memory[8] [57]), .ZN(n_0_4_1435));
   NAND2_X1 i_0_4_1493 (.A1(n_0_52), .A2(\Memory[1] [57]), .ZN(n_0_4_1436));
   NAND2_X1 i_0_4_1494 (.A1(n_0_61), .A2(\Memory[10] [57]), .ZN(n_0_4_1437));
   NAND3_X1 i_0_4_1495 (.A1(n_0_4_1435), .A2(n_0_4_1436), .A3(n_0_4_1437), 
      .ZN(n_0_4_1438));
   NOR2_X1 i_0_4_1496 (.A1(n_0_4_1434), .A2(n_0_4_1438), .ZN(n_0_4_1439));
   NAND2_X1 i_0_4_1497 (.A1(n_0_65), .A2(\Memory[14] [57]), .ZN(n_0_4_1440));
   NAND2_X1 i_0_4_1498 (.A1(n_0_66), .A2(\Memory[15] [57]), .ZN(n_0_4_1441));
   NAND2_X1 i_0_4_1499 (.A1(n_0_51), .A2(\Memory[0] [57]), .ZN(n_0_4_1442));
   NAND2_X1 i_0_4_1500 (.A1(n_0_60), .A2(\Memory[9] [57]), .ZN(n_0_4_1443));
   NAND4_X1 i_0_4_1501 (.A1(n_0_4_1440), .A2(n_0_4_1441), .A3(n_0_4_1442), 
      .A4(n_0_4_1443), .ZN(n_0_4_1444));
   NAND2_X1 i_0_4_1502 (.A1(n_0_64), .A2(\Memory[13] [57]), .ZN(n_0_4_1445));
   NAND2_X1 i_0_4_1503 (.A1(n_0_63), .A2(\Memory[12] [57]), .ZN(n_0_4_1446));
   NAND2_X1 i_0_4_1504 (.A1(n_0_62), .A2(\Memory[11] [57]), .ZN(n_0_4_1447));
   NAND3_X1 i_0_4_1505 (.A1(n_0_4_1445), .A2(n_0_4_1446), .A3(n_0_4_1447), 
      .ZN(n_0_4_1448));
   NOR2_X1 i_0_4_1506 (.A1(n_0_4_1444), .A2(n_0_4_1448), .ZN(n_0_4_1449));
   NAND3_X1 i_0_4_1507 (.A1(n_0_4_1430), .A2(n_0_4_1439), .A3(n_0_4_1449), 
      .ZN(dataOut2[57]));
   NAND2_X1 i_0_4_1508 (.A1(n_0_55), .A2(\Memory[4] [58]), .ZN(n_0_4_1450));
   NAND2_X1 i_0_4_1509 (.A1(n_0_58), .A2(\Memory[7] [58]), .ZN(n_0_4_1451));
   NAND2_X1 i_0_4_1510 (.A1(n_0_54), .A2(\Memory[3] [58]), .ZN(n_0_4_1452));
   NAND2_X1 i_0_4_1511 (.A1(n_0_53), .A2(\Memory[2] [58]), .ZN(n_0_4_1453));
   NAND4_X1 i_0_4_1512 (.A1(n_0_4_1450), .A2(n_0_4_1451), .A3(n_0_4_1452), 
      .A4(n_0_4_1453), .ZN(n_0_4_1454));
   INV_X1 i_0_4_1513 (.A(n_0_4_1454), .ZN(n_0_4_1455));
   NAND2_X1 i_0_4_1514 (.A1(n_0_67), .A2(\Memory[16] [58]), .ZN(n_0_4_1456));
   NAND2_X1 i_0_4_1515 (.A1(n_0_57), .A2(\Memory[6] [58]), .ZN(n_0_4_1457));
   NAND2_X1 i_0_4_1516 (.A1(n_0_56), .A2(\Memory[5] [58]), .ZN(n_0_4_1458));
   NAND3_X1 i_0_4_1517 (.A1(n_0_4_1456), .A2(n_0_4_1457), .A3(n_0_4_1458), 
      .ZN(n_0_4_1459));
   NAND2_X1 i_0_4_1518 (.A1(n_0_59), .A2(\Memory[8] [58]), .ZN(n_0_4_1460));
   NAND2_X1 i_0_4_1519 (.A1(n_0_52), .A2(\Memory[1] [58]), .ZN(n_0_4_1461));
   NAND2_X1 i_0_4_1520 (.A1(n_0_61), .A2(\Memory[10] [58]), .ZN(n_0_4_1462));
   NAND3_X1 i_0_4_1521 (.A1(n_0_4_1460), .A2(n_0_4_1461), .A3(n_0_4_1462), 
      .ZN(n_0_4_1463));
   NOR2_X1 i_0_4_1522 (.A1(n_0_4_1459), .A2(n_0_4_1463), .ZN(n_0_4_1464));
   NAND2_X1 i_0_4_1523 (.A1(n_0_65), .A2(\Memory[14] [58]), .ZN(n_0_4_1465));
   NAND2_X1 i_0_4_1524 (.A1(n_0_66), .A2(\Memory[15] [58]), .ZN(n_0_4_1466));
   NAND2_X1 i_0_4_1525 (.A1(n_0_51), .A2(\Memory[0] [58]), .ZN(n_0_4_1467));
   NAND2_X1 i_0_4_1526 (.A1(n_0_60), .A2(\Memory[9] [58]), .ZN(n_0_4_1468));
   NAND4_X1 i_0_4_1527 (.A1(n_0_4_1465), .A2(n_0_4_1466), .A3(n_0_4_1467), 
      .A4(n_0_4_1468), .ZN(n_0_4_1469));
   NAND2_X1 i_0_4_1528 (.A1(n_0_64), .A2(\Memory[13] [58]), .ZN(n_0_4_1470));
   NAND2_X1 i_0_4_1529 (.A1(n_0_63), .A2(\Memory[12] [58]), .ZN(n_0_4_1471));
   NAND2_X1 i_0_4_1530 (.A1(n_0_62), .A2(\Memory[11] [58]), .ZN(n_0_4_1472));
   NAND3_X1 i_0_4_1531 (.A1(n_0_4_1470), .A2(n_0_4_1471), .A3(n_0_4_1472), 
      .ZN(n_0_4_1473));
   NOR2_X1 i_0_4_1532 (.A1(n_0_4_1469), .A2(n_0_4_1473), .ZN(n_0_4_1474));
   NAND3_X1 i_0_4_1533 (.A1(n_0_4_1455), .A2(n_0_4_1464), .A3(n_0_4_1474), 
      .ZN(dataOut2[58]));
   NAND2_X1 i_0_4_1534 (.A1(n_0_55), .A2(\Memory[4] [59]), .ZN(n_0_4_1475));
   NAND2_X1 i_0_4_1535 (.A1(n_0_58), .A2(\Memory[7] [59]), .ZN(n_0_4_1476));
   NAND2_X1 i_0_4_1536 (.A1(n_0_54), .A2(\Memory[3] [59]), .ZN(n_0_4_1477));
   NAND2_X1 i_0_4_1537 (.A1(n_0_53), .A2(\Memory[2] [59]), .ZN(n_0_4_1478));
   NAND4_X1 i_0_4_1538 (.A1(n_0_4_1475), .A2(n_0_4_1476), .A3(n_0_4_1477), 
      .A4(n_0_4_1478), .ZN(n_0_4_1479));
   INV_X1 i_0_4_1539 (.A(n_0_4_1479), .ZN(n_0_4_1480));
   NAND2_X1 i_0_4_1540 (.A1(n_0_67), .A2(\Memory[16] [59]), .ZN(n_0_4_1481));
   NAND2_X1 i_0_4_1541 (.A1(n_0_57), .A2(\Memory[6] [59]), .ZN(n_0_4_1482));
   NAND2_X1 i_0_4_1542 (.A1(n_0_56), .A2(\Memory[5] [59]), .ZN(n_0_4_1483));
   NAND3_X1 i_0_4_1543 (.A1(n_0_4_1481), .A2(n_0_4_1482), .A3(n_0_4_1483), 
      .ZN(n_0_4_1484));
   NAND2_X1 i_0_4_1544 (.A1(n_0_59), .A2(\Memory[8] [59]), .ZN(n_0_4_1485));
   NAND2_X1 i_0_4_1545 (.A1(n_0_52), .A2(\Memory[1] [59]), .ZN(n_0_4_1486));
   NAND2_X1 i_0_4_1546 (.A1(n_0_61), .A2(\Memory[10] [59]), .ZN(n_0_4_1487));
   NAND3_X1 i_0_4_1547 (.A1(n_0_4_1485), .A2(n_0_4_1486), .A3(n_0_4_1487), 
      .ZN(n_0_4_1488));
   NOR2_X1 i_0_4_1548 (.A1(n_0_4_1484), .A2(n_0_4_1488), .ZN(n_0_4_1489));
   NAND2_X1 i_0_4_1549 (.A1(n_0_65), .A2(\Memory[14] [59]), .ZN(n_0_4_1490));
   NAND2_X1 i_0_4_1550 (.A1(n_0_66), .A2(\Memory[15] [59]), .ZN(n_0_4_1491));
   NAND2_X1 i_0_4_1551 (.A1(n_0_51), .A2(\Memory[0] [59]), .ZN(n_0_4_1492));
   NAND2_X1 i_0_4_1552 (.A1(n_0_60), .A2(\Memory[9] [59]), .ZN(n_0_4_1493));
   NAND4_X1 i_0_4_1553 (.A1(n_0_4_1490), .A2(n_0_4_1491), .A3(n_0_4_1492), 
      .A4(n_0_4_1493), .ZN(n_0_4_1494));
   NAND2_X1 i_0_4_1554 (.A1(n_0_64), .A2(\Memory[13] [59]), .ZN(n_0_4_1495));
   NAND2_X1 i_0_4_1555 (.A1(n_0_63), .A2(\Memory[12] [59]), .ZN(n_0_4_1496));
   NAND2_X1 i_0_4_1556 (.A1(n_0_62), .A2(\Memory[11] [59]), .ZN(n_0_4_1497));
   NAND3_X1 i_0_4_1557 (.A1(n_0_4_1495), .A2(n_0_4_1496), .A3(n_0_4_1497), 
      .ZN(n_0_4_1498));
   NOR2_X1 i_0_4_1558 (.A1(n_0_4_1494), .A2(n_0_4_1498), .ZN(n_0_4_1499));
   NAND3_X1 i_0_4_1559 (.A1(n_0_4_1480), .A2(n_0_4_1489), .A3(n_0_4_1499), 
      .ZN(dataOut2[59]));
   NAND2_X1 i_0_4_1560 (.A1(n_0_55), .A2(\Memory[4] [60]), .ZN(n_0_4_1500));
   NAND2_X1 i_0_4_1561 (.A1(n_0_58), .A2(\Memory[7] [60]), .ZN(n_0_4_1501));
   NAND2_X1 i_0_4_1562 (.A1(n_0_54), .A2(\Memory[3] [60]), .ZN(n_0_4_1502));
   NAND2_X1 i_0_4_1563 (.A1(n_0_53), .A2(\Memory[2] [60]), .ZN(n_0_4_1503));
   NAND4_X1 i_0_4_1564 (.A1(n_0_4_1500), .A2(n_0_4_1501), .A3(n_0_4_1502), 
      .A4(n_0_4_1503), .ZN(n_0_4_1504));
   INV_X1 i_0_4_1565 (.A(n_0_4_1504), .ZN(n_0_4_1505));
   NAND2_X1 i_0_4_1566 (.A1(n_0_67), .A2(\Memory[16] [60]), .ZN(n_0_4_1506));
   NAND2_X1 i_0_4_1567 (.A1(n_0_57), .A2(\Memory[6] [60]), .ZN(n_0_4_1507));
   NAND2_X1 i_0_4_1568 (.A1(n_0_56), .A2(\Memory[5] [60]), .ZN(n_0_4_1508));
   NAND3_X1 i_0_4_1569 (.A1(n_0_4_1506), .A2(n_0_4_1507), .A3(n_0_4_1508), 
      .ZN(n_0_4_1509));
   NAND2_X1 i_0_4_1570 (.A1(n_0_59), .A2(\Memory[8] [60]), .ZN(n_0_4_1510));
   NAND2_X1 i_0_4_1571 (.A1(n_0_52), .A2(\Memory[1] [60]), .ZN(n_0_4_1511));
   NAND2_X1 i_0_4_1572 (.A1(n_0_61), .A2(\Memory[10] [60]), .ZN(n_0_4_1512));
   NAND3_X1 i_0_4_1573 (.A1(n_0_4_1510), .A2(n_0_4_1511), .A3(n_0_4_1512), 
      .ZN(n_0_4_1513));
   NOR2_X1 i_0_4_1574 (.A1(n_0_4_1509), .A2(n_0_4_1513), .ZN(n_0_4_1514));
   NAND2_X1 i_0_4_1575 (.A1(n_0_65), .A2(\Memory[14] [60]), .ZN(n_0_4_1515));
   NAND2_X1 i_0_4_1576 (.A1(n_0_66), .A2(\Memory[15] [60]), .ZN(n_0_4_1516));
   NAND2_X1 i_0_4_1577 (.A1(n_0_51), .A2(\Memory[0] [60]), .ZN(n_0_4_1517));
   NAND2_X1 i_0_4_1578 (.A1(n_0_60), .A2(\Memory[9] [60]), .ZN(n_0_4_1518));
   NAND4_X1 i_0_4_1579 (.A1(n_0_4_1515), .A2(n_0_4_1516), .A3(n_0_4_1517), 
      .A4(n_0_4_1518), .ZN(n_0_4_1519));
   NAND2_X1 i_0_4_1580 (.A1(n_0_64), .A2(\Memory[13] [60]), .ZN(n_0_4_1520));
   NAND2_X1 i_0_4_1581 (.A1(n_0_63), .A2(\Memory[12] [60]), .ZN(n_0_4_1521));
   NAND2_X1 i_0_4_1582 (.A1(n_0_62), .A2(\Memory[11] [60]), .ZN(n_0_4_1522));
   NAND3_X1 i_0_4_1583 (.A1(n_0_4_1520), .A2(n_0_4_1521), .A3(n_0_4_1522), 
      .ZN(n_0_4_1523));
   NOR2_X1 i_0_4_1584 (.A1(n_0_4_1519), .A2(n_0_4_1523), .ZN(n_0_4_1524));
   NAND3_X1 i_0_4_1585 (.A1(n_0_4_1505), .A2(n_0_4_1514), .A3(n_0_4_1524), 
      .ZN(dataOut2[60]));
   NAND2_X1 i_0_4_1586 (.A1(n_0_55), .A2(\Memory[4] [61]), .ZN(n_0_4_1525));
   NAND2_X1 i_0_4_1587 (.A1(n_0_58), .A2(\Memory[7] [61]), .ZN(n_0_4_1526));
   NAND2_X1 i_0_4_1588 (.A1(n_0_54), .A2(\Memory[3] [61]), .ZN(n_0_4_1527));
   NAND2_X1 i_0_4_1589 (.A1(n_0_53), .A2(\Memory[2] [61]), .ZN(n_0_4_1528));
   NAND4_X1 i_0_4_1590 (.A1(n_0_4_1525), .A2(n_0_4_1526), .A3(n_0_4_1527), 
      .A4(n_0_4_1528), .ZN(n_0_4_1529));
   INV_X1 i_0_4_1591 (.A(n_0_4_1529), .ZN(n_0_4_1530));
   NAND2_X1 i_0_4_1592 (.A1(n_0_67), .A2(\Memory[16] [61]), .ZN(n_0_4_1531));
   NAND2_X1 i_0_4_1593 (.A1(n_0_57), .A2(\Memory[6] [61]), .ZN(n_0_4_1532));
   NAND2_X1 i_0_4_1594 (.A1(n_0_56), .A2(\Memory[5] [61]), .ZN(n_0_4_1533));
   NAND3_X1 i_0_4_1595 (.A1(n_0_4_1531), .A2(n_0_4_1532), .A3(n_0_4_1533), 
      .ZN(n_0_4_1534));
   NAND2_X1 i_0_4_1596 (.A1(n_0_59), .A2(\Memory[8] [61]), .ZN(n_0_4_1535));
   NAND2_X1 i_0_4_1597 (.A1(n_0_52), .A2(\Memory[1] [61]), .ZN(n_0_4_1536));
   NAND2_X1 i_0_4_1598 (.A1(n_0_61), .A2(\Memory[10] [61]), .ZN(n_0_4_1537));
   NAND3_X1 i_0_4_1599 (.A1(n_0_4_1535), .A2(n_0_4_1536), .A3(n_0_4_1537), 
      .ZN(n_0_4_1538));
   NOR2_X1 i_0_4_1600 (.A1(n_0_4_1534), .A2(n_0_4_1538), .ZN(n_0_4_1539));
   NAND2_X1 i_0_4_1601 (.A1(n_0_65), .A2(\Memory[14] [61]), .ZN(n_0_4_1540));
   NAND2_X1 i_0_4_1602 (.A1(n_0_66), .A2(\Memory[15] [61]), .ZN(n_0_4_1541));
   NAND2_X1 i_0_4_1603 (.A1(n_0_51), .A2(\Memory[0] [61]), .ZN(n_0_4_1542));
   NAND2_X1 i_0_4_1604 (.A1(n_0_60), .A2(\Memory[9] [61]), .ZN(n_0_4_1543));
   NAND4_X1 i_0_4_1605 (.A1(n_0_4_1540), .A2(n_0_4_1541), .A3(n_0_4_1542), 
      .A4(n_0_4_1543), .ZN(n_0_4_1544));
   NAND2_X1 i_0_4_1606 (.A1(n_0_64), .A2(\Memory[13] [61]), .ZN(n_0_4_1545));
   NAND2_X1 i_0_4_1607 (.A1(n_0_63), .A2(\Memory[12] [61]), .ZN(n_0_4_1546));
   NAND2_X1 i_0_4_1608 (.A1(n_0_62), .A2(\Memory[11] [61]), .ZN(n_0_4_1547));
   NAND3_X1 i_0_4_1609 (.A1(n_0_4_1545), .A2(n_0_4_1546), .A3(n_0_4_1547), 
      .ZN(n_0_4_1548));
   NOR2_X1 i_0_4_1610 (.A1(n_0_4_1544), .A2(n_0_4_1548), .ZN(n_0_4_1549));
   NAND3_X1 i_0_4_1611 (.A1(n_0_4_1530), .A2(n_0_4_1539), .A3(n_0_4_1549), 
      .ZN(dataOut2[61]));
   NAND2_X1 i_0_4_1612 (.A1(n_0_55), .A2(\Memory[4] [62]), .ZN(n_0_4_1550));
   NAND2_X1 i_0_4_1613 (.A1(n_0_58), .A2(\Memory[7] [62]), .ZN(n_0_4_1551));
   NAND2_X1 i_0_4_1614 (.A1(n_0_54), .A2(\Memory[3] [62]), .ZN(n_0_4_1552));
   NAND2_X1 i_0_4_1615 (.A1(n_0_53), .A2(\Memory[2] [62]), .ZN(n_0_4_1553));
   NAND4_X1 i_0_4_1616 (.A1(n_0_4_1550), .A2(n_0_4_1551), .A3(n_0_4_1552), 
      .A4(n_0_4_1553), .ZN(n_0_4_1554));
   INV_X1 i_0_4_1617 (.A(n_0_4_1554), .ZN(n_0_4_1555));
   NAND2_X1 i_0_4_1618 (.A1(n_0_67), .A2(\Memory[16] [62]), .ZN(n_0_4_1556));
   NAND2_X1 i_0_4_1619 (.A1(n_0_57), .A2(\Memory[6] [62]), .ZN(n_0_4_1557));
   NAND2_X1 i_0_4_1620 (.A1(n_0_56), .A2(\Memory[5] [62]), .ZN(n_0_4_1558));
   NAND3_X1 i_0_4_1621 (.A1(n_0_4_1556), .A2(n_0_4_1557), .A3(n_0_4_1558), 
      .ZN(n_0_4_1559));
   NAND2_X1 i_0_4_1622 (.A1(n_0_59), .A2(\Memory[8] [62]), .ZN(n_0_4_1560));
   NAND2_X1 i_0_4_1623 (.A1(n_0_52), .A2(\Memory[1] [62]), .ZN(n_0_4_1561));
   NAND2_X1 i_0_4_1624 (.A1(n_0_61), .A2(\Memory[10] [62]), .ZN(n_0_4_1562));
   NAND3_X1 i_0_4_1625 (.A1(n_0_4_1560), .A2(n_0_4_1561), .A3(n_0_4_1562), 
      .ZN(n_0_4_1563));
   NOR2_X1 i_0_4_1626 (.A1(n_0_4_1559), .A2(n_0_4_1563), .ZN(n_0_4_1564));
   NAND2_X1 i_0_4_1627 (.A1(n_0_65), .A2(\Memory[14] [62]), .ZN(n_0_4_1565));
   NAND2_X1 i_0_4_1628 (.A1(n_0_66), .A2(\Memory[15] [62]), .ZN(n_0_4_1566));
   NAND2_X1 i_0_4_1629 (.A1(n_0_51), .A2(\Memory[0] [62]), .ZN(n_0_4_1567));
   NAND2_X1 i_0_4_1630 (.A1(n_0_60), .A2(\Memory[9] [62]), .ZN(n_0_4_1568));
   NAND4_X1 i_0_4_1631 (.A1(n_0_4_1565), .A2(n_0_4_1566), .A3(n_0_4_1567), 
      .A4(n_0_4_1568), .ZN(n_0_4_1569));
   NAND2_X1 i_0_4_1632 (.A1(n_0_64), .A2(\Memory[13] [62]), .ZN(n_0_4_1570));
   NAND2_X1 i_0_4_1633 (.A1(n_0_63), .A2(\Memory[12] [62]), .ZN(n_0_4_1571));
   NAND2_X1 i_0_4_1634 (.A1(n_0_62), .A2(\Memory[11] [62]), .ZN(n_0_4_1572));
   NAND3_X1 i_0_4_1635 (.A1(n_0_4_1570), .A2(n_0_4_1571), .A3(n_0_4_1572), 
      .ZN(n_0_4_1573));
   NOR2_X1 i_0_4_1636 (.A1(n_0_4_1569), .A2(n_0_4_1573), .ZN(n_0_4_1574));
   NAND3_X1 i_0_4_1637 (.A1(n_0_4_1555), .A2(n_0_4_1564), .A3(n_0_4_1574), 
      .ZN(dataOut2[62]));
   NAND2_X1 i_0_4_1638 (.A1(n_0_55), .A2(\Memory[4] [63]), .ZN(n_0_4_1575));
   NAND2_X1 i_0_4_1639 (.A1(n_0_58), .A2(\Memory[7] [63]), .ZN(n_0_4_1576));
   NAND2_X1 i_0_4_1640 (.A1(n_0_54), .A2(\Memory[3] [63]), .ZN(n_0_4_1577));
   NAND2_X1 i_0_4_1641 (.A1(n_0_53), .A2(\Memory[2] [63]), .ZN(n_0_4_1578));
   NAND4_X1 i_0_4_1642 (.A1(n_0_4_1575), .A2(n_0_4_1576), .A3(n_0_4_1577), 
      .A4(n_0_4_1578), .ZN(n_0_4_1579));
   INV_X1 i_0_4_1643 (.A(n_0_4_1579), .ZN(n_0_4_1580));
   NAND2_X1 i_0_4_1644 (.A1(n_0_67), .A2(\Memory[16] [63]), .ZN(n_0_4_1581));
   NAND2_X1 i_0_4_1645 (.A1(n_0_57), .A2(\Memory[6] [63]), .ZN(n_0_4_1582));
   NAND2_X1 i_0_4_1646 (.A1(n_0_56), .A2(\Memory[5] [63]), .ZN(n_0_4_1583));
   NAND3_X1 i_0_4_1647 (.A1(n_0_4_1581), .A2(n_0_4_1582), .A3(n_0_4_1583), 
      .ZN(n_0_4_1584));
   NAND2_X1 i_0_4_1648 (.A1(n_0_59), .A2(\Memory[8] [63]), .ZN(n_0_4_1585));
   NAND2_X1 i_0_4_1649 (.A1(n_0_52), .A2(\Memory[1] [63]), .ZN(n_0_4_1586));
   NAND2_X1 i_0_4_1650 (.A1(n_0_61), .A2(\Memory[10] [63]), .ZN(n_0_4_1587));
   NAND3_X1 i_0_4_1651 (.A1(n_0_4_1585), .A2(n_0_4_1586), .A3(n_0_4_1587), 
      .ZN(n_0_4_1588));
   NOR2_X1 i_0_4_1652 (.A1(n_0_4_1584), .A2(n_0_4_1588), .ZN(n_0_4_1589));
   NAND2_X1 i_0_4_1653 (.A1(n_0_65), .A2(\Memory[14] [63]), .ZN(n_0_4_1590));
   NAND2_X1 i_0_4_1654 (.A1(n_0_66), .A2(\Memory[15] [63]), .ZN(n_0_4_1591));
   NAND2_X1 i_0_4_1655 (.A1(n_0_51), .A2(\Memory[0] [63]), .ZN(n_0_4_1592));
   NAND2_X1 i_0_4_1656 (.A1(n_0_60), .A2(\Memory[9] [63]), .ZN(n_0_4_1593));
   NAND4_X1 i_0_4_1657 (.A1(n_0_4_1590), .A2(n_0_4_1591), .A3(n_0_4_1592), 
      .A4(n_0_4_1593), .ZN(n_0_4_1594));
   NAND2_X1 i_0_4_1658 (.A1(n_0_64), .A2(\Memory[13] [63]), .ZN(n_0_4_1595));
   NAND2_X1 i_0_4_1659 (.A1(n_0_63), .A2(\Memory[12] [63]), .ZN(n_0_4_1596));
   NAND2_X1 i_0_4_1660 (.A1(n_0_62), .A2(\Memory[11] [63]), .ZN(n_0_4_1597));
   NAND3_X1 i_0_4_1661 (.A1(n_0_4_1595), .A2(n_0_4_1596), .A3(n_0_4_1597), 
      .ZN(n_0_4_1598));
   NOR2_X1 i_0_4_1662 (.A1(n_0_4_1594), .A2(n_0_4_1598), .ZN(n_0_4_1599));
   NAND3_X1 i_0_4_1663 (.A1(n_0_4_1580), .A2(n_0_4_1589), .A3(n_0_4_1599), 
      .ZN(dataOut2[63]));
   AND2_X1 i_0_1_0 (.A1(n_0_1_21), .A2(dataIn[0]), .ZN(Memory[0]));
   AND2_X1 i_0_1_1 (.A1(n_0_1_21), .A2(dataIn[1]), .ZN(Memory[1]));
   AND2_X1 i_0_1_2 (.A1(n_0_1_21), .A2(dataIn[2]), .ZN(Memory[2]));
   AND2_X1 i_0_1_3 (.A1(n_0_1_21), .A2(dataIn[3]), .ZN(Memory[3]));
   AND2_X1 i_0_1_4 (.A1(n_0_1_21), .A2(dataIn[4]), .ZN(Memory[4]));
   AND2_X1 i_0_1_5 (.A1(n_0_1_21), .A2(dataIn[5]), .ZN(Memory[5]));
   AND2_X1 i_0_1_6 (.A1(n_0_1_21), .A2(dataIn[6]), .ZN(Memory[6]));
   AND2_X1 i_0_1_7 (.A1(n_0_1_21), .A2(dataIn[7]), .ZN(Memory[7]));
   AND2_X1 i_0_1_8 (.A1(n_0_1_21), .A2(dataIn[8]), .ZN(Memory[8]));
   AND2_X1 i_0_1_9 (.A1(n_0_1_21), .A2(dataIn[9]), .ZN(Memory[9]));
   AND2_X1 i_0_1_10 (.A1(n_0_1_21), .A2(dataIn[10]), .ZN(Memory[10]));
   AND2_X1 i_0_1_11 (.A1(n_0_1_21), .A2(dataIn[11]), .ZN(Memory[11]));
   AND2_X1 i_0_1_12 (.A1(n_0_1_21), .A2(dataIn[12]), .ZN(Memory[12]));
   AND2_X1 i_0_1_13 (.A1(n_0_1_21), .A2(dataIn[13]), .ZN(Memory[13]));
   AND2_X1 i_0_1_14 (.A1(n_0_1_21), .A2(dataIn[14]), .ZN(Memory[14]));
   AND2_X1 i_0_1_15 (.A1(n_0_1_21), .A2(dataIn[15]), .ZN(Memory[15]));
   AND2_X1 i_0_1_16 (.A1(n_0_1_21), .A2(dataIn[16]), .ZN(Memory[16]));
   AND2_X1 i_0_1_17 (.A1(n_0_1_21), .A2(dataIn[17]), .ZN(Memory[17]));
   AND2_X1 i_0_1_18 (.A1(n_0_1_21), .A2(dataIn[18]), .ZN(Memory[18]));
   AND2_X1 i_0_1_19 (.A1(n_0_1_21), .A2(dataIn[19]), .ZN(Memory[19]));
   AND2_X1 i_0_1_20 (.A1(n_0_1_21), .A2(dataIn[20]), .ZN(Memory[20]));
   AND2_X1 i_0_1_21 (.A1(n_0_1_21), .A2(dataIn[21]), .ZN(Memory[21]));
   AND2_X1 i_0_1_22 (.A1(n_0_1_21), .A2(dataIn[22]), .ZN(Memory[22]));
   AND2_X1 i_0_1_23 (.A1(n_0_1_21), .A2(dataIn[23]), .ZN(Memory[23]));
   AND2_X1 i_0_1_24 (.A1(n_0_1_21), .A2(dataIn[24]), .ZN(Memory[24]));
   AND2_X1 i_0_1_25 (.A1(n_0_1_21), .A2(dataIn[25]), .ZN(Memory[25]));
   AND2_X1 i_0_1_26 (.A1(n_0_1_21), .A2(dataIn[26]), .ZN(Memory[26]));
   AND2_X1 i_0_1_27 (.A1(n_0_1_21), .A2(dataIn[27]), .ZN(Memory[27]));
   AND2_X1 i_0_1_28 (.A1(n_0_1_21), .A2(dataIn[28]), .ZN(Memory[28]));
   AND2_X1 i_0_1_29 (.A1(n_0_1_21), .A2(dataIn[29]), .ZN(Memory[29]));
   AND2_X1 i_0_1_30 (.A1(n_0_1_21), .A2(dataIn[30]), .ZN(Memory[30]));
   AND2_X1 i_0_1_31 (.A1(n_0_1_21), .A2(dataIn[31]), .ZN(Memory[31]));
   AND2_X1 i_0_1_32 (.A1(n_0_1_21), .A2(dataIn[32]), .ZN(Memory[32]));
   AND2_X1 i_0_1_33 (.A1(n_0_1_21), .A2(dataIn[33]), .ZN(Memory[33]));
   AND2_X1 i_0_1_34 (.A1(n_0_1_21), .A2(dataIn[34]), .ZN(Memory[34]));
   AND2_X1 i_0_1_35 (.A1(n_0_1_21), .A2(dataIn[35]), .ZN(Memory[35]));
   AND2_X1 i_0_1_36 (.A1(n_0_1_21), .A2(dataIn[36]), .ZN(Memory[36]));
   AND2_X1 i_0_1_37 (.A1(n_0_1_21), .A2(dataIn[37]), .ZN(Memory[37]));
   AND2_X1 i_0_1_38 (.A1(n_0_1_21), .A2(dataIn[38]), .ZN(Memory[38]));
   AND2_X1 i_0_1_39 (.A1(n_0_1_21), .A2(dataIn[39]), .ZN(Memory[39]));
   AND2_X1 i_0_1_40 (.A1(n_0_1_21), .A2(dataIn[40]), .ZN(Memory[40]));
   AND2_X1 i_0_1_41 (.A1(n_0_1_21), .A2(dataIn[41]), .ZN(Memory[41]));
   AND2_X1 i_0_1_42 (.A1(n_0_1_21), .A2(dataIn[42]), .ZN(Memory[42]));
   AND2_X1 i_0_1_43 (.A1(n_0_1_21), .A2(dataIn[43]), .ZN(Memory[43]));
   AND2_X1 i_0_1_44 (.A1(n_0_1_21), .A2(dataIn[44]), .ZN(Memory[44]));
   AND2_X1 i_0_1_45 (.A1(n_0_1_21), .A2(dataIn[45]), .ZN(Memory[45]));
   AND2_X1 i_0_1_46 (.A1(n_0_1_21), .A2(dataIn[46]), .ZN(Memory[46]));
   AND2_X1 i_0_1_47 (.A1(n_0_1_21), .A2(dataIn[47]), .ZN(Memory[47]));
   AND2_X1 i_0_1_48 (.A1(n_0_1_21), .A2(dataIn[48]), .ZN(Memory[48]));
   AND2_X1 i_0_1_49 (.A1(n_0_1_21), .A2(dataIn[49]), .ZN(Memory[49]));
   AND2_X1 i_0_1_50 (.A1(n_0_1_21), .A2(dataIn[50]), .ZN(Memory[50]));
   AND2_X1 i_0_1_51 (.A1(n_0_1_21), .A2(dataIn[51]), .ZN(Memory[51]));
   AND2_X1 i_0_1_52 (.A1(n_0_1_21), .A2(dataIn[52]), .ZN(Memory[52]));
   AND2_X1 i_0_1_53 (.A1(n_0_1_21), .A2(dataIn[53]), .ZN(Memory[53]));
   AND2_X1 i_0_1_54 (.A1(n_0_1_21), .A2(dataIn[54]), .ZN(Memory[54]));
   AND2_X1 i_0_1_55 (.A1(n_0_1_21), .A2(dataIn[55]), .ZN(Memory[55]));
   AND2_X1 i_0_1_56 (.A1(n_0_1_21), .A2(dataIn[56]), .ZN(Memory[56]));
   AND2_X1 i_0_1_57 (.A1(n_0_1_21), .A2(dataIn[57]), .ZN(Memory[57]));
   AND2_X1 i_0_1_58 (.A1(n_0_1_21), .A2(dataIn[58]), .ZN(Memory[58]));
   AND2_X1 i_0_1_59 (.A1(n_0_1_21), .A2(dataIn[59]), .ZN(Memory[59]));
   AND2_X1 i_0_1_60 (.A1(n_0_1_21), .A2(dataIn[60]), .ZN(Memory[60]));
   AND2_X1 i_0_1_61 (.A1(n_0_1_21), .A2(dataIn[61]), .ZN(Memory[61]));
   AND2_X1 i_0_1_62 (.A1(n_0_1_21), .A2(dataIn[62]), .ZN(Memory[62]));
   AND2_X1 i_0_1_63 (.A1(n_0_1_21), .A2(dataIn[63]), .ZN(Memory[63]));
   OAI21_X1 i_0_1_64 (.A(n_0_1_21), .B1(n_0_1_13), .B2(n_0_1_3), .ZN(n_0_17));
   OAI21_X1 i_0_1_65 (.A(n_0_1_21), .B1(n_0_1_4), .B2(n_0_1_0), .ZN(n_0_18));
   OAI21_X1 i_0_1_66 (.A(n_0_1_21), .B1(n_0_1_5), .B2(n_0_1_0), .ZN(n_0_19));
   OAI21_X1 i_0_1_67 (.A(n_0_1_21), .B1(n_0_1_9), .B2(n_0_1_0), .ZN(n_0_20));
   OR2_X1 i_0_1_68 (.A1(n_0_1_14), .A2(n_0_1_3), .ZN(n_0_1_0));
   OAI21_X1 i_0_1_69 (.A(n_0_1_21), .B1(n_0_1_13), .B2(n_0_1_8), .ZN(n_0_21));
   OAI21_X1 i_0_1_70 (.A(n_0_1_21), .B1(n_0_1_4), .B2(n_0_1_1), .ZN(n_0_22));
   OAI21_X1 i_0_1_71 (.A(n_0_1_21), .B1(n_0_1_5), .B2(n_0_1_1), .ZN(n_0_23));
   OAI21_X1 i_0_1_72 (.A(n_0_1_21), .B1(n_0_1_9), .B2(n_0_1_1), .ZN(n_0_24));
   OR2_X1 i_0_1_73 (.A1(n_0_1_14), .A2(n_0_1_8), .ZN(n_0_1_1));
   OAI21_X1 i_0_1_74 (.A(n_0_1_21), .B1(n_0_1_17), .B2(n_0_1_2), .ZN(n_0_25));
   OAI21_X1 i_0_1_75 (.A(n_0_1_21), .B1(n_0_1_4), .B2(n_0_1_2), .ZN(n_0_26));
   OAI21_X1 i_0_1_76 (.A(n_0_1_21), .B1(n_0_1_5), .B2(n_0_1_2), .ZN(n_0_27));
   OAI21_X1 i_0_1_77 (.A(n_0_1_21), .B1(n_0_1_9), .B2(n_0_1_2), .ZN(n_0_28));
   OR2_X1 i_0_1_78 (.A1(n_0_1_7), .A2(n_0_1_3), .ZN(n_0_1_2));
   NAND2_X1 i_0_1_79 (.A1(n_0_1_11), .A2(n_0_1_20), .ZN(n_0_1_3));
   OAI21_X1 i_0_1_80 (.A(n_0_1_21), .B1(n_0_1_17), .B2(n_0_1_6), .ZN(n_0_29));
   OAI21_X1 i_0_1_81 (.A(n_0_1_21), .B1(n_0_1_6), .B2(n_0_1_4), .ZN(n_0_30));
   OR2_X1 i_0_1_82 (.A1(n_0_1_18), .A2(address_WR[1]), .ZN(n_0_1_4));
   OAI21_X1 i_0_1_83 (.A(n_0_1_21), .B1(n_0_1_6), .B2(n_0_1_5), .ZN(n_0_31));
   NAND2_X1 i_0_1_84 (.A1(n_0_1_18), .A2(address_WR[1]), .ZN(n_0_1_5));
   OAI21_X1 i_0_1_85 (.A(n_0_1_21), .B1(n_0_1_9), .B2(n_0_1_6), .ZN(n_0_32));
   OR2_X1 i_0_1_86 (.A1(n_0_1_8), .A2(n_0_1_7), .ZN(n_0_1_6));
   NAND4_X1 i_0_1_87 (.A1(WR_Enable), .A2(address_WR[3]), .A3(n_0_1_16), 
      .A4(n_0_1_15), .ZN(n_0_1_7));
   NAND3_X1 i_0_1_88 (.A1(n_0_1_12), .A2(n_0_1_20), .A3(address_WR[2]), .ZN(
      n_0_1_8));
   NAND2_X1 i_0_1_89 (.A1(address_WR[1]), .A2(address_WR[0]), .ZN(n_0_1_9));
   NOR2_X1 i_0_1_90 (.A1(n_0_1_13), .A2(n_0_1_10), .ZN(n_0_33));
   NAND3_X1 i_0_1_91 (.A1(n_0_1_11), .A2(n_0_1_21), .A3(address_WR[4]), .ZN(
      n_0_1_10));
   NOR3_X1 i_0_1_92 (.A1(address_WR[6]), .A2(address_WR[5]), .A3(address_WR[2]), 
      .ZN(n_0_1_11));
   NOR2_X1 i_0_1_93 (.A1(address_WR[6]), .A2(address_WR[5]), .ZN(n_0_1_12));
   OR2_X1 i_0_1_94 (.A1(n_0_1_17), .A2(n_0_1_14), .ZN(n_0_1_13));
   NAND4_X1 i_0_1_95 (.A1(WR_Enable), .A2(n_0_1_15), .A3(n_0_1_19), .A4(n_0_1_16), 
      .ZN(n_0_1_14));
   NOR4_X1 i_0_1_96 (.A1(address_WR[10]), .A2(address_WR[9]), .A3(address_WR[8]), 
      .A4(address_WR[7]), .ZN(n_0_1_15));
   NOR2_X1 i_0_1_97 (.A1(address_WR[12]), .A2(address_WR[11]), .ZN(n_0_1_16));
   OR2_X1 i_0_1_98 (.A1(address_WR[1]), .A2(address_WR[0]), .ZN(n_0_1_17));
   INV_X1 i_0_1_99 (.A(address_WR[0]), .ZN(n_0_1_18));
   INV_X1 i_0_1_100 (.A(address_WR[3]), .ZN(n_0_1_19));
   INV_X1 i_0_1_101 (.A(address_WR[4]), .ZN(n_0_1_20));
   INV_X1 i_0_1_102 (.A(RST), .ZN(n_0_1_21));
endmodule
