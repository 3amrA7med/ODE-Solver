/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Apr 24 21:42:34 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 4015801768 */

module add_sub_cla(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;

   INV_X1 i_0_0_0 (.A(n_0_0_0), .ZN(invalid));
   OAI21_X1 i_0_0_1 (.A(n_0_0_1), .B1(n_0_0_7), .B2(n_0_0_6), .ZN(n_0_0_0));
   OAI221_X1 i_0_0_2 (.A(n_0_0_2), .B1(n_0_0_23), .B2(n_0_0_4), .C1(n_0_0_21), 
      .C2(n_0_0_20), .ZN(n_0_0_1));
   NOR3_X1 i_0_0_3 (.A1(n_0_0_13), .A2(n_0_0_3), .A3(n_0_0_15), .ZN(n_0_0_2));
   OR4_X1 i_0_0_4 (.A1(out[12]), .A2(n_0_0_90), .A3(n_0_0_10), .A4(n_0_0_12), 
      .ZN(n_0_0_3));
   INV_X1 i_0_0_5 (.A(n_0_0_5), .ZN(n_0_0_4));
   OAI211_X1 i_0_0_6 (.A(n_0_0_27), .B(n_0_0_25), .C1(n_0_0_69), .C2(n_0_0_24), 
      .ZN(n_0_0_5));
   XNOR2_X1 i_0_0_7 (.A(n_0_0_90), .B(n_0_0_22), .ZN(n_0_0_6));
   OR3_X1 i_0_0_8 (.A1(n_0_0_16), .A2(n_0_0_8), .A3(n_0_0_20), .ZN(n_0_0_7));
   OAI211_X1 i_0_0_9 (.A(n_0_0_15), .B(n_0_0_9), .C1(n_0_0_19), .C2(n_0_0_18), 
      .ZN(n_0_0_8));
   AND4_X1 i_0_0_10 (.A1(out[12]), .A2(n_0_0_10), .A3(n_0_0_12), .A4(n_0_0_13), 
      .ZN(n_0_0_9));
   XNOR2_X1 i_0_0_11 (.A(n_0_0_33), .B(n_0_0_11), .ZN(n_0_0_10));
   AOI21_X1 i_0_0_12 (.A(n_0_0_32), .B1(n_0_0_37), .B2(n_0_0_35), .ZN(n_0_0_11));
   XOR2_X1 i_0_0_13 (.A(n_0_0_39), .B(n_0_0_31), .Z(n_0_0_12));
   XNOR2_X1 i_0_0_14 (.A(n_0_0_30), .B(n_0_0_14), .ZN(n_0_0_13));
   AOI21_X1 i_0_0_15 (.A(n_0_0_29), .B1(n_0_0_54), .B2(n_0_0_51), .ZN(n_0_0_14));
   XOR2_X1 i_0_0_16 (.A(n_0_0_57), .B(n_0_0_28), .Z(n_0_0_15));
   INV_X1 i_0_0_17 (.A(n_0_0_17), .ZN(n_0_0_16));
   OAI21_X1 i_0_0_18 (.A(n_0_0_19), .B1(n_0_0_79), .B2(n_0_0_18), .ZN(n_0_0_17));
   AOI22_X1 i_0_0_19 (.A1(n_0_0_80), .A2(n_0_0_70), .B1(n_0_0_84), .B2(n_0_0_26), 
      .ZN(n_0_0_18));
   OAI21_X1 i_0_0_20 (.A(n_0_0_70), .B1(n_0_0_84), .B2(n_0_0_26), .ZN(n_0_0_19));
   AND2_X1 i_0_0_21 (.A1(n_0_0_89), .A2(n_0_0_22), .ZN(n_0_0_20));
   OR2_X1 i_0_0_22 (.A1(n_0_0_90), .A2(n_0_0_21), .ZN(cout));
   NOR2_X1 i_0_0_23 (.A1(n_0_0_89), .A2(n_0_0_22), .ZN(n_0_0_21));
   NOR3_X1 i_0_0_24 (.A1(n_0_0_71), .A2(n_0_0_24), .A3(n_0_0_23), .ZN(n_0_0_22));
   NOR3_X1 i_0_0_25 (.A1(n_0_0_69), .A2(n_0_0_24), .A3(n_0_0_25), .ZN(n_0_0_23));
   AND2_X1 i_0_0_26 (.A1(n_0_0_84), .A2(n_0_0_80), .ZN(n_0_0_24));
   OAI22_X1 i_0_0_27 (.A1(n_0_0_84), .A2(n_0_0_80), .B1(n_0_0_69), .B2(n_0_0_26), 
      .ZN(n_0_0_25));
   INV_X1 i_0_0_28 (.A(n_0_0_27), .ZN(n_0_0_26));
   AOI21_X1 i_0_0_29 (.A(n_0_0_58), .B1(n_0_0_57), .B2(n_0_0_28), .ZN(n_0_0_27));
   OAI21_X1 i_0_0_30 (.A(n_0_0_50), .B1(n_0_0_30), .B2(n_0_0_29), .ZN(n_0_0_28));
   NOR2_X1 i_0_0_31 (.A1(n_0_0_54), .A2(n_0_0_51), .ZN(n_0_0_29));
   AOI21_X1 i_0_0_32 (.A(n_0_0_40), .B1(n_0_0_39), .B2(n_0_0_31), .ZN(n_0_0_30));
   OAI21_X1 i_0_0_33 (.A(n_0_0_34), .B1(n_0_0_33), .B2(n_0_0_32), .ZN(n_0_0_31));
   NOR2_X1 i_0_0_34 (.A1(n_0_0_37), .A2(n_0_0_35), .ZN(n_0_0_32));
   NOR2_X1 i_0_0_35 (.A1(n_0_0_97), .A2(n_0_0_94), .ZN(n_0_0_33));
   NAND2_X1 i_0_0_36 (.A1(n_0_0_37), .A2(n_0_0_35), .ZN(n_0_0_34));
   NAND2_X1 i_0_0_37 (.A1(n_0_0_102), .A2(n_0_0_36), .ZN(n_0_0_35));
   OAI221_X1 i_0_0_38 (.A(n_0_0_249), .B1(n_0_0_272), .B2(n_0_0_100), .C1(
      n_0_0_271), .C2(n_0_0_43), .ZN(n_0_0_36));
   XNOR2_X1 i_0_0_39 (.A(sub), .B(n_0_0_38), .ZN(n_0_0_37));
   AOI222_X1 i_0_0_40 (.A1(in2[12]), .A2(n_0_0_274), .B1(n_0_0_270), .B2(
      n_0_0_48), .C1(n_0_0_259), .C2(n_0_0_107), .ZN(n_0_0_38));
   AOI21_X1 i_0_0_41 (.A(n_0_0_40), .B1(n_0_0_45), .B2(n_0_0_41), .ZN(n_0_0_39));
   NOR2_X1 i_0_0_42 (.A1(n_0_0_45), .A2(n_0_0_41), .ZN(n_0_0_40));
   AND2_X1 i_0_0_43 (.A1(n_0_0_102), .A2(n_0_0_42), .ZN(n_0_0_41));
   OAI221_X1 i_0_0_44 (.A(n_0_0_249), .B1(n_0_0_272), .B2(n_0_0_43), .C1(
      n_0_0_271), .C2(n_0_0_53), .ZN(n_0_0_42));
   AOI22_X1 i_0_0_45 (.A1(n_0_0_247), .A2(n_0_0_229), .B1(n_0_0_248), .B2(
      n_0_0_44), .ZN(n_0_0_43));
   AOI22_X1 i_0_0_46 (.A1(in1[12]), .A2(n_0_0_246), .B1(in1[11]), .B2(n_0_0_245), 
      .ZN(n_0_0_44));
   XNOR2_X1 i_0_0_47 (.A(n_0_0_283), .B(n_0_0_46), .ZN(n_0_0_45));
   AOI21_X1 i_0_0_48 (.A(n_0_0_47), .B1(n_0_0_259), .B2(n_0_0_48), .ZN(n_0_0_46));
   OAI21_X1 i_0_0_49 (.A(n_0_0_106), .B1(n_0_0_269), .B2(n_0_0_56), .ZN(n_0_0_47));
   OAI21_X1 i_0_0_50 (.A(n_0_0_49), .B1(n_0_0_267), .B2(n_0_0_234), .ZN(n_0_0_48));
   OAI21_X1 i_0_0_51 (.A(n_0_0_109), .B1(in2[11]), .B2(n_0_0_264), .ZN(n_0_0_49));
   NAND2_X1 i_0_0_52 (.A1(n_0_0_54), .A2(n_0_0_51), .ZN(n_0_0_50));
   NAND2_X1 i_0_0_53 (.A1(n_0_0_102), .A2(n_0_0_52), .ZN(n_0_0_51));
   OAI221_X1 i_0_0_54 (.A(n_0_0_249), .B1(n_0_0_271), .B2(n_0_0_62), .C1(
      n_0_0_272), .C2(n_0_0_53), .ZN(n_0_0_52));
   OAI21_X1 i_0_0_55 (.A(n_0_0_64), .B1(n_0_0_248), .B2(n_0_0_241), .ZN(n_0_0_53));
   XNOR2_X1 i_0_0_56 (.A(n_0_0_283), .B(n_0_0_55), .ZN(n_0_0_54));
   OAI221_X1 i_0_0_57 (.A(n_0_0_106), .B1(n_0_0_269), .B2(n_0_0_67), .C1(
      n_0_0_258), .C2(n_0_0_56), .ZN(n_0_0_55));
   OAI22_X1 i_0_0_58 (.A1(in2[12]), .A2(n_0_0_266), .B1(n_0_0_267), .B2(
      n_0_0_256), .ZN(n_0_0_56));
   AOI21_X1 i_0_0_59 (.A(n_0_0_58), .B1(n_0_0_65), .B2(n_0_0_59), .ZN(n_0_0_57));
   NOR2_X1 i_0_0_60 (.A1(n_0_0_65), .A2(n_0_0_59), .ZN(n_0_0_58));
   AOI21_X1 i_0_0_61 (.A(n_0_0_103), .B1(n_0_0_63), .B2(n_0_0_60), .ZN(n_0_0_59));
   INV_X1 i_0_0_62 (.A(n_0_0_61), .ZN(n_0_0_60));
   OAI21_X1 i_0_0_63 (.A(n_0_0_249), .B1(n_0_0_272), .B2(n_0_0_62), .ZN(n_0_0_61));
   OAI21_X1 i_0_0_64 (.A(n_0_0_64), .B1(n_0_0_248), .B2(n_0_0_244), .ZN(n_0_0_62));
   OAI211_X1 i_0_0_65 (.A(n_0_0_272), .B(n_0_0_64), .C1(n_0_0_248), .C2(
      n_0_0_101), .ZN(n_0_0_63));
   NAND2_X1 i_0_0_66 (.A1(in1[12]), .A2(n_0_0_248), .ZN(n_0_0_64));
   XNOR2_X1 i_0_0_67 (.A(sub), .B(n_0_0_66), .ZN(n_0_0_65));
   OAI211_X1 i_0_0_68 (.A(n_0_0_106), .B(n_0_0_68), .C1(n_0_0_258), .C2(n_0_0_67), 
      .ZN(n_0_0_66));
   OAI22_X1 i_0_0_69 (.A1(in2[12]), .A2(n_0_0_266), .B1(n_0_0_267), .B2(
      n_0_0_262), .ZN(n_0_0_67));
   OAI221_X1 i_0_0_70 (.A(n_0_0_270), .B1(in2[12]), .B2(n_0_0_153), .C1(in2[10]), 
      .C2(n_0_0_152), .ZN(n_0_0_68));
   INV_X1 i_0_0_71 (.A(n_0_0_70), .ZN(n_0_0_69));
   AOI21_X1 i_0_0_72 (.A(n_0_0_71), .B1(n_0_0_76), .B2(n_0_0_72), .ZN(n_0_0_70));
   NOR2_X1 i_0_0_73 (.A1(n_0_0_76), .A2(n_0_0_72), .ZN(n_0_0_71));
   XOR2_X1 i_0_0_74 (.A(sub), .B(n_0_0_73), .Z(n_0_0_72));
   OAI22_X1 i_0_0_75 (.A1(in2[11]), .A2(n_0_0_74), .B1(in2[12]), .B2(n_0_0_75), 
      .ZN(n_0_0_73));
   INV_X1 i_0_0_76 (.A(n_0_0_75), .ZN(n_0_0_74));
   NOR2_X1 i_0_0_77 (.A1(n_0_0_258), .A2(n_0_0_152), .ZN(n_0_0_75));
   AOI22_X1 i_0_0_78 (.A1(in1[11]), .A2(n_0_0_78), .B1(in1[12]), .B2(n_0_0_77), 
      .ZN(n_0_0_76));
   INV_X1 i_0_0_79 (.A(n_0_0_78), .ZN(n_0_0_77));
   NOR2_X1 i_0_0_80 (.A1(n_0_0_272), .A2(n_0_0_82), .ZN(n_0_0_78));
   INV_X1 i_0_0_81 (.A(n_0_0_80), .ZN(n_0_0_79));
   OAI22_X1 i_0_0_82 (.A1(n_0_0_82), .A2(n_0_0_81), .B1(n_0_0_295), .B2(n_0_0_83), 
      .ZN(n_0_0_80));
   AOI22_X1 i_0_0_83 (.A1(in1[10]), .A2(n_0_0_271), .B1(in1[11]), .B2(n_0_0_272), 
      .ZN(n_0_0_81));
   INV_X1 i_0_0_84 (.A(n_0_0_83), .ZN(n_0_0_82));
   NOR3_X1 i_0_0_85 (.A1(n_0_0_275), .A2(n_0_0_246), .A3(n_0_0_248), .ZN(
      n_0_0_83));
   XOR2_X1 i_0_0_86 (.A(n_0_0_283), .B(n_0_0_85), .Z(n_0_0_84));
   AOI21_X1 i_0_0_87 (.A(n_0_0_86), .B1(in2[12]), .B2(n_0_0_88), .ZN(n_0_0_85));
   NOR2_X1 i_0_0_88 (.A1(n_0_0_88), .A2(n_0_0_87), .ZN(n_0_0_86));
   AOI22_X1 i_0_0_89 (.A1(in2[10]), .A2(n_0_0_271), .B1(in2[11]), .B2(n_0_0_272), 
      .ZN(n_0_0_87));
   NAND2_X1 i_0_0_90 (.A1(n_0_0_275), .A2(n_0_0_153), .ZN(n_0_0_88));
   NOR2_X1 i_0_0_91 (.A1(in1[12]), .A2(n_0_0_91), .ZN(n_0_0_89));
   AND2_X1 i_0_0_92 (.A1(in1[12]), .A2(n_0_0_91), .ZN(n_0_0_90));
   OAI22_X1 i_0_0_93 (.A1(n_0_0_286), .A2(sub), .B1(in2[12]), .B2(n_0_0_283), 
      .ZN(n_0_0_91));
   XOR2_X1 i_0_0_94 (.A(n_0_0_134), .B(n_0_0_133), .Z(out[0]));
   XOR2_X1 i_0_0_95 (.A(n_0_0_132), .B(n_0_0_131), .Z(out[1]));
   XNOR2_X1 i_0_0_96 (.A(n_0_0_129), .B(n_0_0_128), .ZN(out[2]));
   XNOR2_X1 i_0_0_97 (.A(n_0_0_127), .B(n_0_0_126), .ZN(out[3]));
   XOR2_X1 i_0_0_98 (.A(n_0_0_161), .B(n_0_0_124), .Z(out[4]));
   XOR2_X1 i_0_0_99 (.A(n_0_0_122), .B(n_0_0_121), .Z(out[5]));
   XOR2_X1 i_0_0_100 (.A(n_0_0_120), .B(n_0_0_119), .Z(out[6]));
   XNOR2_X1 i_0_0_101 (.A(n_0_0_118), .B(n_0_0_92), .ZN(out[7]));
   OAI21_X1 i_0_0_102 (.A(n_0_0_190), .B1(n_0_0_196), .B2(n_0_0_191), .ZN(
      n_0_0_92));
   XOR2_X1 i_0_0_103 (.A(n_0_0_200), .B(n_0_0_116), .Z(out[8]));
   XOR2_X1 i_0_0_104 (.A(n_0_0_115), .B(n_0_0_114), .Z(out[9]));
   XNOR2_X1 i_0_0_105 (.A(n_0_0_113), .B(n_0_0_93), .ZN(out[10]));
   OAI21_X1 i_0_0_106 (.A(n_0_0_223), .B1(n_0_0_230), .B2(n_0_0_224), .ZN(
      n_0_0_93));
   OAI22_X1 i_0_0_107 (.A1(n_0_0_235), .A2(n_0_0_111), .B1(n_0_0_236), .B2(
      n_0_0_112), .ZN(out[11]));
   AOI21_X1 i_0_0_108 (.A(n_0_0_94), .B1(n_0_0_110), .B2(n_0_0_95), .ZN(out[12]));
   NOR2_X1 i_0_0_109 (.A1(n_0_0_110), .A2(n_0_0_95), .ZN(n_0_0_94));
   INV_X1 i_0_0_110 (.A(n_0_0_96), .ZN(n_0_0_95));
   AOI21_X1 i_0_0_111 (.A(n_0_0_97), .B1(n_0_0_104), .B2(n_0_0_98), .ZN(n_0_0_96));
   NOR2_X1 i_0_0_112 (.A1(n_0_0_104), .A2(n_0_0_98), .ZN(n_0_0_97));
   AND2_X1 i_0_0_113 (.A1(n_0_0_102), .A2(n_0_0_99), .ZN(n_0_0_98));
   OAI221_X1 i_0_0_114 (.A(n_0_0_249), .B1(n_0_0_271), .B2(n_0_0_100), .C1(
      n_0_0_272), .C2(n_0_0_242), .ZN(n_0_0_99));
   OAI22_X1 i_0_0_115 (.A1(n_0_0_247), .A2(n_0_0_101), .B1(n_0_0_248), .B2(
      n_0_0_216), .ZN(n_0_0_100));
   AOI22_X1 i_0_0_116 (.A1(in1[10]), .A2(n_0_0_245), .B1(in1[12]), .B2(n_0_0_246), 
      .ZN(n_0_0_101));
   INV_X1 i_0_0_117 (.A(n_0_0_103), .ZN(n_0_0_102));
   NOR2_X1 i_0_0_118 (.A1(n_0_0_295), .A2(n_0_0_249), .ZN(n_0_0_103));
   XNOR2_X1 i_0_0_119 (.A(n_0_0_283), .B(n_0_0_105), .ZN(n_0_0_104));
   AOI222_X1 i_0_0_120 (.A1(n_0_0_260), .A2(n_0_0_259), .B1(in2[12]), .B2(
      n_0_0_274), .C1(n_0_0_270), .C2(n_0_0_107), .ZN(n_0_0_105));
   NAND2_X1 i_0_0_121 (.A1(in2[12]), .A2(n_0_0_274), .ZN(n_0_0_106));
   OAI21_X1 i_0_0_122 (.A(n_0_0_108), .B1(n_0_0_267), .B2(n_0_0_221), .ZN(
      n_0_0_107));
   OAI21_X1 i_0_0_123 (.A(n_0_0_109), .B1(in2[10]), .B2(n_0_0_264), .ZN(
      n_0_0_108));
   AOI21_X1 i_0_0_124 (.A(n_0_0_266), .B1(n_0_0_286), .B2(n_0_0_264), .ZN(
      n_0_0_109));
   OAI22_X1 i_0_0_125 (.A1(n_0_0_252), .A2(n_0_0_237), .B1(n_0_0_235), .B2(
      n_0_0_111), .ZN(n_0_0_110));
   INV_X1 i_0_0_126 (.A(n_0_0_112), .ZN(n_0_0_111));
   OAI21_X1 i_0_0_127 (.A(n_0_0_223), .B1(n_0_0_222), .B2(n_0_0_113), .ZN(
      n_0_0_112));
   OAI22_X1 i_0_0_128 (.A1(n_0_0_217), .A2(n_0_0_211), .B1(n_0_0_115), .B2(
      n_0_0_114), .ZN(n_0_0_113));
   XNOR2_X1 i_0_0_129 (.A(n_0_0_217), .B(n_0_0_211), .ZN(n_0_0_114));
   AOI21_X1 i_0_0_130 (.A(n_0_0_201), .B1(n_0_0_200), .B2(n_0_0_116), .ZN(
      n_0_0_115));
   INV_X1 i_0_0_131 (.A(n_0_0_117), .ZN(n_0_0_116));
   OAI21_X1 i_0_0_132 (.A(n_0_0_190), .B1(n_0_0_189), .B2(n_0_0_118), .ZN(
      n_0_0_117));
   OAI22_X1 i_0_0_133 (.A1(n_0_0_185), .A2(n_0_0_180), .B1(n_0_0_120), .B2(
      n_0_0_119), .ZN(n_0_0_118));
   XNOR2_X1 i_0_0_134 (.A(n_0_0_185), .B(n_0_0_180), .ZN(n_0_0_119));
   AOI21_X1 i_0_0_135 (.A(n_0_0_171), .B1(n_0_0_122), .B2(n_0_0_121), .ZN(
      n_0_0_120));
   AOI21_X1 i_0_0_136 (.A(n_0_0_171), .B1(n_0_0_176), .B2(n_0_0_172), .ZN(
      n_0_0_121));
   INV_X1 i_0_0_137 (.A(n_0_0_123), .ZN(n_0_0_122));
   AOI21_X1 i_0_0_138 (.A(n_0_0_162), .B1(n_0_0_161), .B2(n_0_0_124), .ZN(
      n_0_0_123));
   INV_X1 i_0_0_139 (.A(n_0_0_125), .ZN(n_0_0_124));
   OAI22_X1 i_0_0_140 (.A1(n_0_0_157), .A2(n_0_0_154), .B1(n_0_0_127), .B2(
      n_0_0_126), .ZN(n_0_0_125));
   XNOR2_X1 i_0_0_141 (.A(n_0_0_157), .B(n_0_0_154), .ZN(n_0_0_126));
   AOI21_X1 i_0_0_142 (.A(n_0_0_144), .B1(n_0_0_129), .B2(n_0_0_128), .ZN(
      n_0_0_127));
   AOI21_X1 i_0_0_143 (.A(n_0_0_144), .B1(n_0_0_149), .B2(n_0_0_145), .ZN(
      n_0_0_128));
   INV_X1 i_0_0_144 (.A(n_0_0_130), .ZN(n_0_0_129));
   OAI22_X1 i_0_0_145 (.A1(n_0_0_141), .A2(n_0_0_139), .B1(n_0_0_132), .B2(
      n_0_0_131), .ZN(n_0_0_130));
   XNOR2_X1 i_0_0_146 (.A(n_0_0_141), .B(n_0_0_139), .ZN(n_0_0_131));
   AOI21_X1 i_0_0_147 (.A(n_0_0_135), .B1(n_0_0_134), .B2(n_0_0_133), .ZN(
      n_0_0_132));
   AOI21_X1 i_0_0_148 (.A(n_0_0_135), .B1(n_0_0_137), .B2(n_0_0_136), .ZN(
      n_0_0_133));
   OR2_X1 i_0_0_149 (.A1(sub), .A2(cin), .ZN(n_0_0_134));
   NOR2_X1 i_0_0_150 (.A1(n_0_0_137), .A2(n_0_0_136), .ZN(n_0_0_135));
   NAND2_X1 i_0_0_151 (.A1(in1[0]), .A2(n_0_0_250), .ZN(n_0_0_136));
   XNOR2_X1 i_0_0_152 (.A(sub), .B(n_0_0_138), .ZN(n_0_0_137));
   NOR2_X1 i_0_0_153 (.A1(n_0_0_284), .A2(n_0_0_275), .ZN(n_0_0_138));
   AOI22_X1 i_0_0_154 (.A1(in1[1]), .A2(n_0_0_250), .B1(n_0_0_153), .B2(
      n_0_0_140), .ZN(n_0_0_139));
   NOR3_X1 i_0_0_155 (.A1(n_0_0_290), .A2(n_0_0_272), .A3(n_0_0_275), .ZN(
      n_0_0_140));
   XNOR2_X1 i_0_0_156 (.A(n_0_0_283), .B(n_0_0_142), .ZN(n_0_0_141));
   AOI22_X1 i_0_0_157 (.A1(in2[1]), .A2(n_0_0_274), .B1(n_0_0_259), .B2(
      n_0_0_143), .ZN(n_0_0_142));
   NOR2_X1 i_0_0_158 (.A1(n_0_0_284), .A2(n_0_0_251), .ZN(n_0_0_143));
   NOR2_X1 i_0_0_159 (.A1(n_0_0_149), .A2(n_0_0_145), .ZN(n_0_0_144));
   XNOR2_X1 i_0_0_160 (.A(sub), .B(n_0_0_146), .ZN(n_0_0_145));
   OAI21_X1 i_0_0_161 (.A(n_0_0_147), .B1(in2[2]), .B2(n_0_0_275), .ZN(n_0_0_146));
   OAI211_X1 i_0_0_162 (.A(n_0_0_275), .B(n_0_0_148), .C1(n_0_0_199), .C2(
      n_0_0_160), .ZN(n_0_0_147));
   NAND4_X1 i_0_0_163 (.A1(n_0_0_271), .A2(n_0_0_267), .A3(in2[1]), .A4(
      n_0_0_264), .ZN(n_0_0_148));
   OAI22_X1 i_0_0_164 (.A1(n_0_0_250), .A2(n_0_0_150), .B1(n_0_0_292), .B2(
      n_0_0_249), .ZN(n_0_0_149));
   AOI21_X1 i_0_0_165 (.A(n_0_0_151), .B1(n_0_0_272), .B2(n_0_0_156), .ZN(
      n_0_0_150));
   NOR3_X1 i_0_0_166 (.A1(n_0_0_291), .A2(n_0_0_272), .A3(n_0_0_152), .ZN(
      n_0_0_151));
   INV_X1 i_0_0_167 (.A(n_0_0_153), .ZN(n_0_0_152));
   NOR2_X1 i_0_0_168 (.A1(n_0_0_267), .A2(n_0_0_264), .ZN(n_0_0_153));
   AOI22_X1 i_0_0_169 (.A1(n_0_0_249), .A2(n_0_0_155), .B1(n_0_0_293), .B2(
      n_0_0_250), .ZN(n_0_0_154));
   OAI22_X1 i_0_0_170 (.A1(n_0_0_272), .A2(n_0_0_156), .B1(n_0_0_271), .B2(
      n_0_0_170), .ZN(n_0_0_155));
   NOR2_X1 i_0_0_171 (.A1(n_0_0_247), .A2(n_0_0_195), .ZN(n_0_0_156));
   XNOR2_X1 i_0_0_172 (.A(sub), .B(n_0_0_158), .ZN(n_0_0_157));
   OAI21_X1 i_0_0_173 (.A(n_0_0_159), .B1(in2[3]), .B2(n_0_0_275), .ZN(n_0_0_158));
   OAI221_X1 i_0_0_174 (.A(n_0_0_275), .B1(n_0_0_199), .B2(n_0_0_166), .C1(
      n_0_0_210), .C2(n_0_0_160), .ZN(n_0_0_159));
   NAND2_X1 i_0_0_175 (.A1(n_0_0_272), .A2(n_0_0_267), .ZN(n_0_0_160));
   AOI21_X1 i_0_0_176 (.A(n_0_0_162), .B1(n_0_0_167), .B2(n_0_0_163), .ZN(
      n_0_0_161));
   NOR2_X1 i_0_0_177 (.A1(n_0_0_167), .A2(n_0_0_163), .ZN(n_0_0_162));
   XOR2_X1 i_0_0_178 (.A(sub), .B(n_0_0_164), .Z(n_0_0_163));
   OAI21_X1 i_0_0_179 (.A(n_0_0_165), .B1(in2[4]), .B2(n_0_0_275), .ZN(n_0_0_164));
   OAI221_X1 i_0_0_180 (.A(n_0_0_275), .B1(n_0_0_210), .B2(n_0_0_166), .C1(
      n_0_0_271), .C2(n_0_0_178), .ZN(n_0_0_165));
   NAND2_X1 i_0_0_181 (.A1(n_0_0_271), .A2(n_0_0_267), .ZN(n_0_0_166));
   AOI22_X1 i_0_0_182 (.A1(n_0_0_249), .A2(n_0_0_168), .B1(in1[4]), .B2(
      n_0_0_250), .ZN(n_0_0_167));
   INV_X1 i_0_0_183 (.A(n_0_0_169), .ZN(n_0_0_168));
   AOI22_X1 i_0_0_184 (.A1(n_0_0_272), .A2(n_0_0_175), .B1(n_0_0_271), .B2(
      n_0_0_170), .ZN(n_0_0_169));
   NOR2_X1 i_0_0_185 (.A1(n_0_0_247), .A2(n_0_0_206), .ZN(n_0_0_170));
   NOR2_X1 i_0_0_186 (.A1(n_0_0_176), .A2(n_0_0_172), .ZN(n_0_0_171));
   AOI22_X1 i_0_0_187 (.A1(n_0_0_249), .A2(n_0_0_173), .B1(in1[5]), .B2(
      n_0_0_250), .ZN(n_0_0_172));
   INV_X1 i_0_0_188 (.A(n_0_0_174), .ZN(n_0_0_173));
   AOI22_X1 i_0_0_189 (.A1(n_0_0_271), .A2(n_0_0_175), .B1(n_0_0_272), .B2(
      n_0_0_183), .ZN(n_0_0_174));
   OAI22_X1 i_0_0_190 (.A1(n_0_0_247), .A2(n_0_0_215), .B1(n_0_0_290), .B2(
      n_0_0_184), .ZN(n_0_0_175));
   XNOR2_X1 i_0_0_191 (.A(n_0_0_283), .B(n_0_0_177), .ZN(n_0_0_176));
   AOI222_X1 i_0_0_192 (.A1(n_0_0_259), .A2(n_0_0_179), .B1(in2[5]), .B2(
      n_0_0_274), .C1(n_0_0_270), .C2(n_0_0_187), .ZN(n_0_0_177));
   INV_X1 i_0_0_193 (.A(n_0_0_179), .ZN(n_0_0_178));
   OAI22_X1 i_0_0_194 (.A1(n_0_0_284), .A2(n_0_0_188), .B1(n_0_0_266), .B2(
      n_0_0_220), .ZN(n_0_0_179));
   OAI22_X1 i_0_0_195 (.A1(n_0_0_250), .A2(n_0_0_181), .B1(in1[6]), .B2(
      n_0_0_249), .ZN(n_0_0_180));
   INV_X1 i_0_0_196 (.A(n_0_0_182), .ZN(n_0_0_181));
   OAI22_X1 i_0_0_197 (.A1(n_0_0_272), .A2(n_0_0_183), .B1(n_0_0_271), .B2(
      n_0_0_194), .ZN(n_0_0_182));
   OAI22_X1 i_0_0_198 (.A1(n_0_0_247), .A2(n_0_0_228), .B1(n_0_0_291), .B2(
      n_0_0_184), .ZN(n_0_0_183));
   NAND2_X1 i_0_0_199 (.A1(n_0_0_247), .A2(n_0_0_246), .ZN(n_0_0_184));
   XNOR2_X1 i_0_0_200 (.A(n_0_0_283), .B(n_0_0_186), .ZN(n_0_0_185));
   AOI222_X1 i_0_0_201 (.A1(n_0_0_270), .A2(n_0_0_198), .B1(in2[6]), .B2(
      n_0_0_274), .C1(n_0_0_259), .C2(n_0_0_187), .ZN(n_0_0_186));
   OAI22_X1 i_0_0_202 (.A1(n_0_0_266), .A2(n_0_0_233), .B1(n_0_0_285), .B2(
      n_0_0_188), .ZN(n_0_0_187));
   NAND2_X1 i_0_0_203 (.A1(n_0_0_266), .A2(n_0_0_264), .ZN(n_0_0_188));
   NOR2_X1 i_0_0_204 (.A1(n_0_0_196), .A2(n_0_0_191), .ZN(n_0_0_189));
   NAND2_X1 i_0_0_205 (.A1(n_0_0_196), .A2(n_0_0_191), .ZN(n_0_0_190));
   OAI22_X1 i_0_0_206 (.A1(n_0_0_250), .A2(n_0_0_192), .B1(in1[7]), .B2(
      n_0_0_249), .ZN(n_0_0_191));
   INV_X1 i_0_0_207 (.A(n_0_0_193), .ZN(n_0_0_192));
   OAI22_X1 i_0_0_208 (.A1(n_0_0_271), .A2(n_0_0_205), .B1(n_0_0_272), .B2(
      n_0_0_194), .ZN(n_0_0_193));
   OAI22_X1 i_0_0_209 (.A1(n_0_0_248), .A2(n_0_0_195), .B1(n_0_0_247), .B2(
      n_0_0_240), .ZN(n_0_0_194));
   AOI22_X1 i_0_0_210 (.A1(in1[0]), .A2(n_0_0_245), .B1(in1[2]), .B2(n_0_0_246), 
      .ZN(n_0_0_195));
   XNOR2_X1 i_0_0_211 (.A(n_0_0_283), .B(n_0_0_197), .ZN(n_0_0_196));
   OAI222_X1 i_0_0_212 (.A1(n_0_0_269), .A2(n_0_0_209), .B1(in2[7]), .B2(
      n_0_0_275), .C1(n_0_0_258), .C2(n_0_0_198), .ZN(n_0_0_197));
   OAI22_X1 i_0_0_213 (.A1(n_0_0_266), .A2(n_0_0_255), .B1(n_0_0_267), .B2(
      n_0_0_199), .ZN(n_0_0_198));
   AOI22_X1 i_0_0_214 (.A1(in2[2]), .A2(n_0_0_264), .B1(in2[0]), .B2(n_0_0_265), 
      .ZN(n_0_0_199));
   AOI21_X1 i_0_0_215 (.A(n_0_0_201), .B1(n_0_0_207), .B2(n_0_0_202), .ZN(
      n_0_0_200));
   NOR2_X1 i_0_0_216 (.A1(n_0_0_207), .A2(n_0_0_202), .ZN(n_0_0_201));
   OAI22_X1 i_0_0_217 (.A1(n_0_0_250), .A2(n_0_0_203), .B1(in1[8]), .B2(
      n_0_0_249), .ZN(n_0_0_202));
   INV_X1 i_0_0_218 (.A(n_0_0_204), .ZN(n_0_0_203));
   OAI22_X1 i_0_0_219 (.A1(n_0_0_271), .A2(n_0_0_214), .B1(n_0_0_272), .B2(
      n_0_0_205), .ZN(n_0_0_204));
   OAI22_X1 i_0_0_220 (.A1(n_0_0_248), .A2(n_0_0_206), .B1(n_0_0_247), .B2(
      n_0_0_243), .ZN(n_0_0_205));
   AOI22_X1 i_0_0_221 (.A1(in1[1]), .A2(n_0_0_245), .B1(in1[3]), .B2(n_0_0_246), 
      .ZN(n_0_0_206));
   XNOR2_X1 i_0_0_222 (.A(n_0_0_283), .B(n_0_0_208), .ZN(n_0_0_207));
   OAI222_X1 i_0_0_223 (.A1(n_0_0_269), .A2(n_0_0_219), .B1(in2[8]), .B2(
      n_0_0_275), .C1(n_0_0_258), .C2(n_0_0_209), .ZN(n_0_0_208));
   OAI22_X1 i_0_0_224 (.A1(n_0_0_266), .A2(n_0_0_261), .B1(n_0_0_267), .B2(
      n_0_0_210), .ZN(n_0_0_209));
   AOI22_X1 i_0_0_225 (.A1(in2[3]), .A2(n_0_0_264), .B1(in2[1]), .B2(n_0_0_265), 
      .ZN(n_0_0_210));
   OAI22_X1 i_0_0_226 (.A1(n_0_0_250), .A2(n_0_0_212), .B1(in1[9]), .B2(
      n_0_0_249), .ZN(n_0_0_211));
   INV_X1 i_0_0_227 (.A(n_0_0_213), .ZN(n_0_0_212));
   OAI22_X1 i_0_0_228 (.A1(n_0_0_271), .A2(n_0_0_227), .B1(n_0_0_272), .B2(
      n_0_0_214), .ZN(n_0_0_213));
   OAI22_X1 i_0_0_229 (.A1(n_0_0_247), .A2(n_0_0_216), .B1(n_0_0_248), .B2(
      n_0_0_215), .ZN(n_0_0_214));
   AOI22_X1 i_0_0_230 (.A1(in1[2]), .A2(n_0_0_245), .B1(in1[4]), .B2(n_0_0_246), 
      .ZN(n_0_0_215));
   AOI22_X1 i_0_0_231 (.A1(in1[6]), .A2(n_0_0_245), .B1(in1[8]), .B2(n_0_0_246), 
      .ZN(n_0_0_216));
   XNOR2_X1 i_0_0_232 (.A(n_0_0_283), .B(n_0_0_218), .ZN(n_0_0_217));
   OAI222_X1 i_0_0_233 (.A1(n_0_0_269), .A2(n_0_0_232), .B1(in2[9]), .B2(
      n_0_0_275), .C1(n_0_0_258), .C2(n_0_0_219), .ZN(n_0_0_218));
   OAI22_X1 i_0_0_234 (.A1(n_0_0_266), .A2(n_0_0_221), .B1(n_0_0_267), .B2(
      n_0_0_220), .ZN(n_0_0_219));
   AOI22_X1 i_0_0_235 (.A1(in2[4]), .A2(n_0_0_264), .B1(in2[2]), .B2(n_0_0_265), 
      .ZN(n_0_0_220));
   AOI22_X1 i_0_0_236 (.A1(in2[8]), .A2(n_0_0_264), .B1(in2[6]), .B2(n_0_0_265), 
      .ZN(n_0_0_221));
   NOR2_X1 i_0_0_237 (.A1(n_0_0_230), .A2(n_0_0_224), .ZN(n_0_0_222));
   NAND2_X1 i_0_0_238 (.A1(n_0_0_230), .A2(n_0_0_224), .ZN(n_0_0_223));
   OAI22_X1 i_0_0_239 (.A1(n_0_0_250), .A2(n_0_0_225), .B1(in1[10]), .B2(
      n_0_0_249), .ZN(n_0_0_224));
   INV_X1 i_0_0_240 (.A(n_0_0_226), .ZN(n_0_0_225));
   OAI22_X1 i_0_0_241 (.A1(n_0_0_271), .A2(n_0_0_239), .B1(n_0_0_272), .B2(
      n_0_0_227), .ZN(n_0_0_226));
   OAI22_X1 i_0_0_242 (.A1(n_0_0_247), .A2(n_0_0_229), .B1(n_0_0_248), .B2(
      n_0_0_228), .ZN(n_0_0_227));
   AOI22_X1 i_0_0_243 (.A1(in1[3]), .A2(n_0_0_245), .B1(in1[5]), .B2(n_0_0_246), 
      .ZN(n_0_0_228));
   AOI22_X1 i_0_0_244 (.A1(in1[7]), .A2(n_0_0_245), .B1(in1[9]), .B2(n_0_0_246), 
      .ZN(n_0_0_229));
   XOR2_X1 i_0_0_245 (.A(sub), .B(n_0_0_231), .Z(n_0_0_230));
   OAI222_X1 i_0_0_246 (.A1(n_0_0_258), .A2(n_0_0_232), .B1(in2[10]), .B2(
      n_0_0_275), .C1(n_0_0_269), .C2(n_0_0_254), .ZN(n_0_0_231));
   OAI22_X1 i_0_0_247 (.A1(n_0_0_266), .A2(n_0_0_234), .B1(n_0_0_267), .B2(
      n_0_0_233), .ZN(n_0_0_232));
   AOI22_X1 i_0_0_248 (.A1(in2[5]), .A2(n_0_0_264), .B1(in2[3]), .B2(n_0_0_265), 
      .ZN(n_0_0_233));
   AOI22_X1 i_0_0_249 (.A1(in2[9]), .A2(n_0_0_264), .B1(in2[7]), .B2(n_0_0_265), 
      .ZN(n_0_0_234));
   INV_X1 i_0_0_250 (.A(n_0_0_236), .ZN(n_0_0_235));
   XOR2_X1 i_0_0_251 (.A(n_0_0_252), .B(n_0_0_237), .Z(n_0_0_236));
   OAI22_X1 i_0_0_252 (.A1(n_0_0_250), .A2(n_0_0_238), .B1(n_0_0_294), .B2(
      n_0_0_249), .ZN(n_0_0_237));
   AOI22_X1 i_0_0_253 (.A1(n_0_0_272), .A2(n_0_0_242), .B1(n_0_0_271), .B2(
      n_0_0_239), .ZN(n_0_0_238));
   OAI22_X1 i_0_0_254 (.A1(n_0_0_247), .A2(n_0_0_241), .B1(n_0_0_248), .B2(
      n_0_0_240), .ZN(n_0_0_239));
   AOI22_X1 i_0_0_255 (.A1(in1[4]), .A2(n_0_0_245), .B1(in1[6]), .B2(n_0_0_246), 
      .ZN(n_0_0_240));
   AOI22_X1 i_0_0_256 (.A1(in1[8]), .A2(n_0_0_245), .B1(in1[10]), .B2(n_0_0_246), 
      .ZN(n_0_0_241));
   OAI22_X1 i_0_0_257 (.A1(n_0_0_247), .A2(n_0_0_244), .B1(n_0_0_248), .B2(
      n_0_0_243), .ZN(n_0_0_242));
   AOI22_X1 i_0_0_258 (.A1(in1[5]), .A2(n_0_0_245), .B1(in1[7]), .B2(n_0_0_246), 
      .ZN(n_0_0_243));
   AOI22_X1 i_0_0_259 (.A1(in1[9]), .A2(n_0_0_245), .B1(in1[11]), .B2(n_0_0_246), 
      .ZN(n_0_0_244));
   INV_X1 i_0_0_260 (.A(n_0_0_246), .ZN(n_0_0_245));
   XOR2_X1 i_0_0_261 (.A(n_0_0_281), .B(n_0_0_278), .Z(n_0_0_246));
   INV_X1 i_0_0_262 (.A(n_0_0_248), .ZN(n_0_0_247));
   XOR2_X1 i_0_0_263 (.A(n_0_0_277), .B(n_0_0_276), .Z(n_0_0_248));
   INV_X1 i_0_0_264 (.A(n_0_0_250), .ZN(n_0_0_249));
   OAI21_X1 i_0_0_265 (.A(n_0_0_274), .B1(n_0_0_271), .B2(n_0_0_251), .ZN(
      n_0_0_250));
   NAND2_X1 i_0_0_266 (.A1(n_0_0_267), .A2(n_0_0_264), .ZN(n_0_0_251));
   XNOR2_X1 i_0_0_267 (.A(sub), .B(n_0_0_253), .ZN(n_0_0_252));
   OAI222_X1 i_0_0_268 (.A1(n_0_0_258), .A2(n_0_0_254), .B1(in2[11]), .B2(
      n_0_0_275), .C1(n_0_0_269), .C2(n_0_0_260), .ZN(n_0_0_253));
   OAI22_X1 i_0_0_269 (.A1(n_0_0_266), .A2(n_0_0_257), .B1(n_0_0_267), .B2(
      n_0_0_255), .ZN(n_0_0_254));
   AOI22_X1 i_0_0_270 (.A1(in2[6]), .A2(n_0_0_264), .B1(in2[4]), .B2(n_0_0_265), 
      .ZN(n_0_0_255));
   INV_X1 i_0_0_271 (.A(n_0_0_257), .ZN(n_0_0_256));
   AOI22_X1 i_0_0_272 (.A1(in2[10]), .A2(n_0_0_264), .B1(in2[8]), .B2(n_0_0_265), 
      .ZN(n_0_0_257));
   INV_X1 i_0_0_273 (.A(n_0_0_259), .ZN(n_0_0_258));
   NOR2_X1 i_0_0_274 (.A1(n_0_0_274), .A2(n_0_0_272), .ZN(n_0_0_259));
   OAI22_X1 i_0_0_275 (.A1(n_0_0_266), .A2(n_0_0_263), .B1(n_0_0_267), .B2(
      n_0_0_261), .ZN(n_0_0_260));
   AOI22_X1 i_0_0_276 (.A1(in2[7]), .A2(n_0_0_264), .B1(in2[5]), .B2(n_0_0_265), 
      .ZN(n_0_0_261));
   INV_X1 i_0_0_277 (.A(n_0_0_263), .ZN(n_0_0_262));
   AOI22_X1 i_0_0_278 (.A1(in2[11]), .A2(n_0_0_264), .B1(in2[9]), .B2(n_0_0_265), 
      .ZN(n_0_0_263));
   INV_X1 i_0_0_279 (.A(n_0_0_265), .ZN(n_0_0_264));
   XOR2_X1 i_0_0_280 (.A(n_0_0_279), .B(n_0_0_273), .Z(n_0_0_265));
   INV_X1 i_0_0_281 (.A(n_0_0_267), .ZN(n_0_0_266));
   XOR2_X1 i_0_0_282 (.A(n_0_0_276), .B(n_0_0_268), .Z(n_0_0_267));
   OAI21_X1 i_0_0_283 (.A(n_0_0_282), .B1(n_0_0_280), .B2(n_0_0_273), .ZN(
      n_0_0_268));
   INV_X1 i_0_0_284 (.A(n_0_0_270), .ZN(n_0_0_269));
   NOR2_X1 i_0_0_285 (.A1(n_0_0_274), .A2(n_0_0_271), .ZN(n_0_0_270));
   INV_X1 i_0_0_286 (.A(n_0_0_272), .ZN(n_0_0_271));
   NOR2_X1 i_0_0_287 (.A1(n_0_0_281), .A2(n_0_0_273), .ZN(n_0_0_272));
   NOR2_X1 i_0_0_288 (.A1(in1[13]), .A2(n_0_0_287), .ZN(n_0_0_273));
   OAI22_X1 i_0_0_289 (.A1(n_0_0_296), .A2(n_0_0_274), .B1(n_0_0_287), .B2(
      n_0_0_275), .ZN(out[13]));
   OAI22_X1 i_0_0_290 (.A1(n_0_0_297), .A2(n_0_0_274), .B1(n_0_0_288), .B2(
      n_0_0_275), .ZN(out[14]));
   INV_X1 i_0_0_291 (.A(n_0_0_275), .ZN(n_0_0_274));
   OAI22_X1 i_0_0_292 (.A1(n_0_0_298), .A2(in2[15]), .B1(n_0_0_277), .B2(
      n_0_0_276), .ZN(n_0_0_275));
   OAI22_X1 i_0_0_293 (.A1(n_0_0_298), .A2(in2[15]), .B1(in1[15]), .B2(n_0_0_289), 
      .ZN(n_0_0_276));
   AOI22_X1 i_0_0_294 (.A1(in1[14]), .A2(n_0_0_288), .B1(n_0_0_281), .B2(
      n_0_0_278), .ZN(n_0_0_277));
   INV_X1 i_0_0_295 (.A(n_0_0_279), .ZN(n_0_0_278));
   OAI21_X1 i_0_0_296 (.A(n_0_0_282), .B1(in1[14]), .B2(n_0_0_288), .ZN(
      n_0_0_279));
   NOR2_X1 i_0_0_297 (.A1(in1[14]), .A2(n_0_0_288), .ZN(n_0_0_280));
   NOR2_X1 i_0_0_298 (.A1(n_0_0_296), .A2(in2[13]), .ZN(n_0_0_281));
   NAND2_X1 i_0_0_299 (.A1(in1[14]), .A2(n_0_0_288), .ZN(n_0_0_282));
   NAND2_X1 i_0_0_300 (.A1(n_0_0_298), .A2(n_0_0_289), .ZN(out[15]));
   INV_X1 i_0_0_301 (.A(sub), .ZN(n_0_0_283));
   INV_X1 i_0_0_302 (.A(in2[0]), .ZN(n_0_0_284));
   INV_X1 i_0_0_303 (.A(in2[1]), .ZN(n_0_0_285));
   INV_X1 i_0_0_304 (.A(in2[12]), .ZN(n_0_0_286));
   INV_X1 i_0_0_305 (.A(in2[13]), .ZN(n_0_0_287));
   INV_X1 i_0_0_306 (.A(in2[14]), .ZN(n_0_0_288));
   INV_X1 i_0_0_307 (.A(in2[15]), .ZN(n_0_0_289));
   INV_X1 i_0_0_308 (.A(in1[0]), .ZN(n_0_0_290));
   INV_X1 i_0_0_309 (.A(in1[1]), .ZN(n_0_0_291));
   INV_X1 i_0_0_310 (.A(in1[2]), .ZN(n_0_0_292));
   INV_X1 i_0_0_311 (.A(in1[3]), .ZN(n_0_0_293));
   INV_X1 i_0_0_312 (.A(in1[11]), .ZN(n_0_0_294));
   INV_X1 i_0_0_313 (.A(in1[12]), .ZN(n_0_0_295));
   INV_X1 i_0_0_314 (.A(in1[13]), .ZN(n_0_0_296));
   INV_X1 i_0_0_315 (.A(in1[14]), .ZN(n_0_0_297));
   INV_X1 i_0_0_316 (.A(in1[15]), .ZN(n_0_0_298));
endmodule
