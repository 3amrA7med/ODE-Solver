/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Apr 24 00:10:33 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2590224225 */

module datapath(num_of_X, p_0);
   input [63:0]num_of_X;
   output [63:0]p_0;

   NAND2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0[1]));
   NAND2_X1 i_1 (.A1(num_of_X[1]), .A2(num_of_X[0]), .ZN(n_0));
   NAND2_X1 i_2 (.A1(n_1), .A2(n_4), .ZN(p_0[2]));
   NAND2_X1 i_3 (.A1(n_2), .A2(num_of_X[2]), .ZN(n_1));
   NAND2_X1 i_4 (.A1(n_230), .A2(n_237), .ZN(n_2));
   NAND2_X1 i_5 (.A1(n_3), .A2(n_229), .ZN(p_0[3]));
   NAND2_X1 i_6 (.A1(n_4), .A2(num_of_X[3]), .ZN(n_3));
   NAND3_X1 i_7 (.A1(n_230), .A2(n_237), .A3(n_231), .ZN(n_4));
   NAND2_X1 i_8 (.A1(n_12), .A2(n_5), .ZN(p_0[4]));
   NAND2_X1 i_9 (.A1(n_229), .A2(num_of_X[4]), .ZN(n_5));
   NAND2_X1 i_10 (.A1(n_8), .A2(n_6), .ZN(p_0[5]));
   NAND2_X1 i_11 (.A1(n_12), .A2(num_of_X[5]), .ZN(n_6));
   NAND2_X1 i_32 (.A1(n_26), .A2(n_21), .ZN(p_0[12]));
   NAND2_X1 i_33 (.A1(n_58), .A2(num_of_X[12]), .ZN(n_21));
   XNOR2_X1 i_34 (.A(n_26), .B(num_of_X[13]), .ZN(p_0[13]));
   NAND2_X1 i_35 (.A1(n_22), .A2(n_24), .ZN(p_0[14]));
   OAI21_X1 i_36 (.A(num_of_X[14]), .B1(n_26), .B2(num_of_X[13]), .ZN(n_22));
   OAI21_X1 i_37 (.A(n_209), .B1(n_23), .B2(n_215), .ZN(p_0[15]));
   INV_X1 i_38 (.A(n_24), .ZN(n_23));
   NAND3_X1 i_39 (.A1(n_25), .A2(n_214), .A3(n_213), .ZN(n_24));
   INV_X1 i_40 (.A(n_26), .ZN(n_25));
   NAND2_X1 i_41 (.A1(n_57), .A2(n_212), .ZN(n_26));
   XNOR2_X1 i_42 (.A(n_209), .B(num_of_X[16]), .ZN(p_0[16]));
   NAND2_X1 i_43 (.A1(n_27), .A2(n_29), .ZN(p_0[17]));
   OAI21_X1 i_44 (.A(num_of_X[17]), .B1(n_209), .B2(num_of_X[16]), .ZN(n_27));
   OAI21_X1 i_45 (.A(n_39), .B1(n_28), .B2(n_206), .ZN(p_0[18]));
   INV_X1 i_46 (.A(n_29), .ZN(n_28));
   NAND3_X1 i_47 (.A1(n_208), .A2(n_205), .A3(n_204), .ZN(n_29));
   XNOR2_X1 i_48 (.A(n_39), .B(num_of_X[19]), .ZN(p_0[19]));
   NAND2_X1 i_49 (.A1(n_30), .A2(n_32), .ZN(p_0[20]));
   OAI21_X1 i_50 (.A(num_of_X[20]), .B1(n_39), .B2(num_of_X[19]), .ZN(n_30));
   OAI21_X1 i_51 (.A(n_34), .B1(n_31), .B2(n_201), .ZN(p_0[21]));
   INV_X1 i_52 (.A(n_32), .ZN(n_31));
   NAND3_X1 i_53 (.A1(n_38), .A2(n_200), .A3(n_207), .ZN(n_32));
   NAND2_X1 i_54 (.A1(n_33), .A2(n_37), .ZN(p_0[22]));
   NAND2_X1 i_55 (.A1(n_34), .A2(num_of_X[22]), .ZN(n_33));
   NAND3_X1 i_56 (.A1(n_38), .A2(n_207), .A3(n_198), .ZN(n_34));
   OAI21_X1 i_57 (.A(n_35), .B1(n_36), .B2(n_197), .ZN(p_0[23]));
   NAND4_X1 i_58 (.A1(n_38), .A2(n_207), .A3(n_198), .A4(n_194), .ZN(n_35));
   INV_X1 i_59 (.A(n_37), .ZN(n_36));
   NAND4_X1 i_60 (.A1(n_38), .A2(n_196), .A3(n_207), .A4(n_198), .ZN(n_37));
   INV_X1 i_61 (.A(n_39), .ZN(n_38));
   NAND2_X1 i_62 (.A1(n_208), .A2(n_202), .ZN(n_39));
   XNOR2_X1 i_63 (.A(n_50), .B(num_of_X[24]), .ZN(p_0[24]));
   NAND2_X1 i_64 (.A1(n_40), .A2(n_42), .ZN(p_0[25]));
   OAI21_X1 i_65 (.A(num_of_X[25]), .B1(n_50), .B2(num_of_X[24]), .ZN(n_40));
   OAI21_X1 i_66 (.A(n_56), .B1(n_41), .B2(n_186), .ZN(p_0[26]));
   INV_X1 i_67 (.A(n_42), .ZN(n_41));
   NAND3_X1 i_68 (.A1(n_49), .A2(n_185), .A3(n_184), .ZN(n_42));
   NAND2_X1 i_69 (.A1(n_43), .A2(n_61), .ZN(p_0[27]));
   NAND2_X1 i_70 (.A1(n_56), .A2(num_of_X[27]), .ZN(n_43));
   NAND2_X1 i_71 (.A1(n_46), .A2(n_44), .ZN(p_0[28]));
   NAND2_X1 i_72 (.A1(n_61), .A2(num_of_X[28]), .ZN(n_44));
   OAI21_X1 i_73 (.A(n_48), .B1(n_45), .B2(n_190), .ZN(p_0[29]));
   INV_X1 i_74 (.A(n_46), .ZN(n_45));
   NAND4_X1 i_75 (.A1(n_49), .A2(n_189), .A3(n_180), .A4(n_182), .ZN(n_46));
   OAI22_X1 i_76 (.A1(n_47), .A2(n_191), .B1(n_188), .B2(n_61), .ZN(p_0[30]));
   INV_X1 i_77 (.A(n_48), .ZN(n_47));
   NAND4_X1 i_78 (.A1(n_49), .A2(n_180), .A3(n_51), .A4(n_182), .ZN(n_48));
   INV_X1 i_79 (.A(n_50), .ZN(n_49));
   NAND2_X1 i_80 (.A1(n_208), .A2(n_192), .ZN(n_50));
   INV_X1 i_81 (.A(n_52), .ZN(n_51));
   NAND2_X1 i_82 (.A1(n_190), .A2(n_189), .ZN(n_52));
   NOR2_X1 i_83 (.A1(n_59), .A2(n_53), .ZN(p_0[31]));
   INV_X1 i_84 (.A(n_54), .ZN(n_53));
   NAND4_X1 i_85 (.A1(n_55), .A2(num_of_X[31]), .A3(n_180), .A4(n_187), .ZN(n_54));
   INV_X1 i_86 (.A(n_56), .ZN(n_55));
   NAND4_X1 i_87 (.A1(n_57), .A2(n_210), .A3(n_248), .A4(n_182), .ZN(n_56));
   INV_X1 i_88 (.A(n_58), .ZN(n_57));
   AOI21_X1 i_90 (.A(num_of_X[31]), .B1(n_60), .B2(n_187), .ZN(n_59));
   INV_X1 i_91 (.A(n_61), .ZN(n_60));
   NAND4_X1 i_92 (.A1(n_208), .A2(n_180), .A3(n_248), .A4(n_182), .ZN(n_61));
   XNOR2_X1 i_93 (.A(n_91), .B(n_166), .ZN(p_0[32]));
   NAND2_X1 i_94 (.A1(n_62), .A2(n_65), .ZN(p_0[33]));
   NAND2_X1 i_95 (.A1(n_63), .A2(num_of_X[33]), .ZN(n_62));
   NAND2_X1 i_96 (.A1(n_91), .A2(n_166), .ZN(n_63));
   OAI21_X1 i_97 (.A(n_67), .B1(n_64), .B2(n_168), .ZN(p_0[34]));
   INV_X1 i_98 (.A(n_65), .ZN(n_64));
   NAND3_X1 i_99 (.A1(n_91), .A2(n_167), .A3(n_166), .ZN(n_65));
   NAND2_X1 i_100 (.A1(n_66), .A2(n_72), .ZN(p_0[35]));
   NAND2_X1 i_101 (.A1(n_67), .A2(num_of_X[35]), .ZN(n_66));
   NAND2_X1 i_102 (.A1(n_91), .A2(n_164), .ZN(n_67));
   XNOR2_X1 i_103 (.A(n_72), .B(num_of_X[36]), .ZN(p_0[36]));
   OAI22_X1 i_104 (.A1(n_68), .A2(n_172), .B1(n_70), .B2(n_72), .ZN(p_0[37]));
   NOR2_X1 i_105 (.A1(n_72), .A2(num_of_X[36]), .ZN(n_68));
   OAI22_X1 i_106 (.A1(n_69), .A2(n_173), .B1(n_170), .B2(n_72), .ZN(p_0[38]));
   NOR2_X1 i_107 (.A1(n_72), .A2(n_70), .ZN(n_69));
   NAND2_X1 i_108 (.A1(n_172), .A2(n_171), .ZN(n_70));
   OAI21_X1 i_109 (.A(n_74), .B1(n_71), .B2(n_163), .ZN(p_0[39]));
   NOR2_X1 i_110 (.A1(n_72), .A2(n_170), .ZN(n_71));
   NAND4_X1 i_111 (.A1(n_208), .A2(n_162), .A3(n_174), .A4(n_164), .ZN(n_72));
   NAND2_X1 i_112 (.A1(n_73), .A2(n_76), .ZN(p_0[40]));
   NAND2_X1 i_113 (.A1(n_74), .A2(num_of_X[40]), .ZN(n_73));
   NAND2_X1 i_114 (.A1(n_91), .A2(n_86), .ZN(n_74));
   OAI21_X1 i_115 (.A(n_78), .B1(n_75), .B2(n_152), .ZN(p_0[41]));
   INV_X1 i_116 (.A(n_76), .ZN(n_75));
   NAND3_X1 i_117 (.A1(n_91), .A2(n_151), .A3(n_86), .ZN(n_76));
   XNOR2_X1 i_118 (.A(n_78), .B(num_of_X[42]), .ZN(p_0[42]));
   OAI21_X1 i_119 (.A(n_83), .B1(n_77), .B2(n_148), .ZN(p_0[43]));
   NOR2_X1 i_120 (.A1(n_78), .A2(num_of_X[42]), .ZN(n_77));
   NAND4_X1 i_121 (.A1(n_208), .A2(n_174), .A3(n_86), .A4(n_149), .ZN(n_78));
   XNOR2_X1 i_122 (.A(n_83), .B(num_of_X[44]), .ZN(p_0[44]));
   OAI22_X1 i_123 (.A1(n_79), .A2(n_156), .B1(n_81), .B2(n_83), .ZN(p_0[45]));
   NOR2_X1 i_124 (.A1(n_83), .A2(num_of_X[44]), .ZN(n_79));
   OAI22_X1 i_125 (.A1(n_80), .A2(n_157), .B1(n_154), .B2(n_83), .ZN(p_0[46]));
   NOR2_X1 i_126 (.A1(n_83), .A2(n_81), .ZN(n_80));
   NAND2_X1 i_127 (.A1(n_156), .A2(n_155), .ZN(n_81));
   OAI21_X1 i_128 (.A(n_88), .B1(n_82), .B2(n_158), .ZN(p_0[47]));
   NOR2_X1 i_129 (.A1(n_83), .A2(n_154), .ZN(n_82));
   NAND4_X1 i_130 (.A1(n_208), .A2(n_174), .A3(n_86), .A4(n_84), .ZN(n_83));
   INV_X1 i_131 (.A(n_85), .ZN(n_84));
   NAND2_X1 i_132 (.A1(n_149), .A2(n_145), .ZN(n_85));
   INV_X1 i_133 (.A(n_159), .ZN(n_86));
   NAND2_X1 i_134 (.A1(n_87), .A2(n_90), .ZN(p_0[48]));
   NAND2_X1 i_135 (.A1(n_88), .A2(num_of_X[48]), .ZN(n_87));
   NAND2_X1 i_136 (.A1(n_91), .A2(n_143), .ZN(n_88));
   OAI21_X1 i_137 (.A(n_93), .B1(n_89), .B2(n_134), .ZN(p_0[49]));
   INV_X1 i_138 (.A(n_90), .ZN(n_89));
   NAND3_X1 i_139 (.A1(n_91), .A2(n_133), .A3(n_143), .ZN(n_90));
   NOR2_X1 i_140 (.A1(n_209), .A2(n_175), .ZN(n_91));
   XNOR2_X1 i_141 (.A(n_93), .B(num_of_X[50]), .ZN(p_0[50]));
   OAI21_X1 i_142 (.A(n_98), .B1(n_92), .B2(n_136), .ZN(p_0[51]));
   NOR2_X1 i_143 (.A1(n_93), .A2(num_of_X[50]), .ZN(n_92));
   NAND4_X1 i_144 (.A1(n_208), .A2(n_174), .A3(n_143), .A4(n_131), .ZN(n_93));
   XNOR2_X1 i_145 (.A(n_98), .B(num_of_X[52]), .ZN(p_0[52]));
   OAI22_X1 i_146 (.A1(n_94), .A2(n_140), .B1(n_96), .B2(n_98), .ZN(p_0[53]));
   NOR2_X1 i_147 (.A1(n_98), .A2(num_of_X[52]), .ZN(n_94));
   OAI22_X1 i_148 (.A1(n_95), .A2(n_141), .B1(n_138), .B2(n_98), .ZN(p_0[54]));
   NOR2_X1 i_149 (.A1(n_98), .A2(n_96), .ZN(n_95));
   NAND2_X1 i_150 (.A1(n_140), .A2(n_139), .ZN(n_96));
   OAI21_X1 i_151 (.A(n_103), .B1(n_97), .B2(n_142), .ZN(p_0[55]));
   NOR2_X1 i_152 (.A1(n_98), .A2(n_138), .ZN(n_97));
   NAND4_X1 i_153 (.A1(n_208), .A2(n_174), .A3(n_143), .A4(n_129), .ZN(n_98));
   XNOR2_X1 i_154 (.A(n_103), .B(num_of_X[56]), .ZN(p_0[56]));
   OAI22_X1 i_155 (.A1(n_99), .A2(n_126), .B1(n_101), .B2(n_103), .ZN(p_0[57]));
   NOR2_X1 i_156 (.A1(n_103), .A2(num_of_X[56]), .ZN(n_99));
   OAI22_X1 i_157 (.A1(n_100), .A2(n_127), .B1(n_106), .B2(n_103), .ZN(p_0[58]));
   NOR2_X1 i_158 (.A1(n_103), .A2(n_101), .ZN(n_100));
   NAND2_X1 i_159 (.A1(n_126), .A2(n_125), .ZN(n_101));
   OAI21_X1 i_160 (.A(n_120), .B1(n_102), .B2(n_128), .ZN(p_0[59]));
   NOR2_X1 i_161 (.A1(n_103), .A2(n_106), .ZN(n_102));
   NAND4_X1 i_162 (.A1(n_208), .A2(n_174), .A3(n_143), .A4(n_104), .ZN(n_103));
   INV_X1 i_163 (.A(n_105), .ZN(n_104));
   NAND3_X1 i_164 (.A1(n_129), .A2(n_142), .A3(n_137), .ZN(n_105));
   NAND3_X1 i_165 (.A1(n_127), .A2(n_126), .A3(n_125), .ZN(n_106));
   INV_X1 i_177 (.A(n_115), .ZN(n_114));
   INV_X1 i_179 (.A(num_of_X[60]), .ZN(n_116));
   NAND2_X1 i_13 (.A1(n_228), .A2(n_233), .ZN(n_12));
   OAI21_X1 i_14 (.A(n_10), .B1(n_7), .B2(n_235), .ZN(p_0[6]));
   INV_X1 i_15 (.A(n_8), .ZN(n_7));
   NAND3_X1 i_16 (.A1(n_228), .A2(n_234), .A3(n_233), .ZN(n_8));
   OAI21_X1 i_17 (.A(n_15), .B1(n_9), .B2(n_236), .ZN(p_0[7]));
   INV_X1 i_18 (.A(n_10), .ZN(n_9));
   NAND3_X1 i_19 (.A1(n_228), .A2(n_233), .A3(n_11), .ZN(n_10));
   INV_X1 i_20 (.A(n_13), .ZN(n_11));
   NAND2_X1 i_21 (.A1(n_235), .A2(n_234), .ZN(n_13));
   NAND2_X1 i_22 (.A1(n_14), .A2(n_17), .ZN(p_0[8]));
   NAND2_X1 i_23 (.A1(n_15), .A2(num_of_X[8]), .ZN(n_14));
   INV_X1 i_24 (.A(n_226), .ZN(n_15));
   NAND2_X1 i_25 (.A1(n_16), .A2(n_19), .ZN(p_0[9]));
   NAND2_X1 i_26 (.A1(n_17), .A2(num_of_X[9]), .ZN(n_16));
   NAND3_X1 i_27 (.A1(n_228), .A2(n_218), .A3(n_222), .ZN(n_17));
   OAI21_X1 i_28 (.A(n_223), .B1(n_18), .B2(n_220), .ZN(p_0[10]));
   INV_X1 i_29 (.A(n_19), .ZN(n_18));
   NAND4_X1 i_30 (.A1(n_228), .A2(n_222), .A3(n_219), .A4(n_218), .ZN(n_19));
   NAND2_X1 i_31 (.A1(n_20), .A2(n_58), .ZN(p_0[11]));
   NAND2_X1 i_89 (.A1(n_223), .A2(num_of_X[11]), .ZN(n_20));
   NAND4_X1 i_281 (.A1(n_228), .A2(n_222), .A3(n_218), .A4(n_224), .ZN(n_223));
   INV_X1 i_282 (.A(n_225), .ZN(n_224));
   NAND2_X1 i_283 (.A1(n_219), .A2(n_220), .ZN(n_225));
   NAND2_X1 i_289 (.A1(n_216), .A2(n_226), .ZN(n_58));
   NOR2_X1 i_290 (.A1(n_229), .A2(n_232), .ZN(n_226));
   INV_X1 i_12 (.A(n_107), .ZN(n_129));
   NAND2_X1 i_166 (.A1(n_165), .A2(n_131), .ZN(n_107));
   INV_X1 i_167 (.A(num_of_X[51]), .ZN(n_136));
   INV_X1 i_168 (.A(num_of_X[48]), .ZN(n_133));
   INV_X1 i_169 (.A(num_of_X[49]), .ZN(n_134));
   NOR2_X1 i_170 (.A1(num_of_X[40]), .A2(num_of_X[41]), .ZN(n_149));
   INV_X1 i_171 (.A(num_of_X[43]), .ZN(n_148));
   INV_X1 i_172 (.A(num_of_X[35]), .ZN(n_162));
   INV_X1 i_173 (.A(num_of_X[39]), .ZN(n_163));
   INV_X1 i_174 (.A(num_of_X[22]), .ZN(n_196));
   INV_X1 i_175 (.A(num_of_X[23]), .ZN(n_197));
   INV_X1 i_176 (.A(num_of_X[20]), .ZN(n_200));
   INV_X1 i_178 (.A(num_of_X[21]), .ZN(n_201));
   NAND2_X1 i_180 (.A1(n_108), .A2(n_110), .ZN(p_0[60]));
   NAND2_X1 i_181 (.A1(n_120), .A2(num_of_X[60]), .ZN(n_108));
   NAND2_X1 i_182 (.A1(n_121), .A2(n_208), .ZN(n_120));
   OAI21_X1 i_183 (.A(n_113), .B1(n_109), .B2(n_118), .ZN(p_0[61]));
   INV_X1 i_184 (.A(n_110), .ZN(n_109));
   NAND4_X1 i_185 (.A1(n_208), .A2(n_150), .A3(n_111), .A4(n_143), .ZN(n_110));
   INV_X1 i_186 (.A(num_of_X[60]), .ZN(n_111));
   OAI21_X1 i_187 (.A(n_135), .B1(n_112), .B2(n_147), .ZN(p_0[62]));
   INV_X1 i_188 (.A(n_113), .ZN(n_112));
   NAND4_X1 i_189 (.A1(n_208), .A2(n_150), .A3(n_143), .A4(n_117), .ZN(n_113));
   INV_X1 i_190 (.A(n_115), .ZN(n_117));
   NAND2_X1 i_191 (.A1(n_116), .A2(n_118), .ZN(n_115));
   INV_X1 i_192 (.A(num_of_X[61]), .ZN(n_118));
   NAND2_X1 i_193 (.A1(n_132), .A2(n_119), .ZN(p_0[63]));
   NAND4_X1 i_194 (.A1(n_121), .A2(n_130), .A3(n_208), .A4(n_144), .ZN(n_119));
   INV_X1 i_195 (.A(n_122), .ZN(n_121));
   NAND3_X1 i_196 (.A1(n_174), .A2(n_143), .A3(n_123), .ZN(n_122));
   INV_X1 i_197 (.A(n_124), .ZN(n_123));
   NAND2_X1 i_198 (.A1(n_160), .A2(n_169), .ZN(n_124));
   INV_X1 i_199 (.A(n_175), .ZN(n_174));
   NAND2_X1 i_200 (.A1(n_192), .A2(n_178), .ZN(n_175));
   INV_X1 i_201 (.A(num_of_X[63]), .ZN(n_130));
   NAND2_X1 i_202 (.A1(n_135), .A2(num_of_X[63]), .ZN(n_132));
   NAND4_X1 i_203 (.A1(n_208), .A2(n_150), .A3(n_143), .A4(n_144), .ZN(n_135));
   INV_X1 i_204 (.A(n_146), .ZN(n_144));
   NAND2_X1 i_205 (.A1(n_114), .A2(n_147), .ZN(n_146));
   INV_X1 i_206 (.A(num_of_X[62]), .ZN(n_147));
   INV_X1 i_207 (.A(n_153), .ZN(n_150));
   NAND4_X1 i_208 (.A1(n_192), .A2(n_178), .A3(n_160), .A4(n_169), .ZN(n_153));
   INV_X1 i_209 (.A(n_161), .ZN(n_160));
   NAND3_X1 i_210 (.A1(n_137), .A2(n_131), .A3(n_165), .ZN(n_161));
   NOR2_X1 i_211 (.A1(num_of_X[50]), .A2(num_of_X[51]), .ZN(n_165));
   NOR2_X1 i_212 (.A1(num_of_X[48]), .A2(num_of_X[49]), .ZN(n_131));
   INV_X1 i_213 (.A(n_138), .ZN(n_137));
   NAND3_X1 i_214 (.A1(n_139), .A2(n_141), .A3(n_140), .ZN(n_138));
   INV_X1 i_215 (.A(num_of_X[52]), .ZN(n_139));
   INV_X1 i_216 (.A(num_of_X[53]), .ZN(n_140));
   INV_X1 i_217 (.A(num_of_X[54]), .ZN(n_141));
   NOR2_X1 i_218 (.A1(n_176), .A2(n_177), .ZN(n_169));
   NAND3_X1 i_219 (.A1(n_125), .A2(n_126), .A3(n_142), .ZN(n_176));
   INV_X1 i_220 (.A(num_of_X[55]), .ZN(n_142));
   INV_X1 i_221 (.A(num_of_X[56]), .ZN(n_125));
   INV_X1 i_222 (.A(num_of_X[57]), .ZN(n_126));
   NAND2_X1 i_223 (.A1(n_128), .A2(n_127), .ZN(n_177));
   INV_X1 i_224 (.A(num_of_X[58]), .ZN(n_127));
   INV_X1 i_225 (.A(num_of_X[59]), .ZN(n_128));
   INV_X1 i_226 (.A(n_179), .ZN(n_178));
   NAND3_X1 i_227 (.A1(n_182), .A2(n_187), .A3(n_181), .ZN(n_179));
   INV_X1 i_228 (.A(n_183), .ZN(n_181));
   NAND2_X1 i_229 (.A1(n_193), .A2(n_180), .ZN(n_183));
   INV_X1 i_230 (.A(num_of_X[27]), .ZN(n_180));
   INV_X1 i_231 (.A(num_of_X[31]), .ZN(n_193));
   INV_X1 i_232 (.A(n_195), .ZN(n_182));
   NAND3_X1 i_233 (.A1(n_184), .A2(n_185), .A3(n_186), .ZN(n_195));
   INV_X1 i_234 (.A(num_of_X[24]), .ZN(n_184));
   INV_X1 i_235 (.A(num_of_X[25]), .ZN(n_185));
   INV_X1 i_236 (.A(num_of_X[26]), .ZN(n_186));
   INV_X1 i_237 (.A(n_188), .ZN(n_187));
   NAND3_X1 i_238 (.A1(n_189), .A2(n_191), .A3(n_190), .ZN(n_188));
   INV_X1 i_239 (.A(num_of_X[28]), .ZN(n_189));
   INV_X1 i_240 (.A(num_of_X[29]), .ZN(n_190));
   INV_X1 i_241 (.A(num_of_X[30]), .ZN(n_191));
   INV_X1 i_242 (.A(n_199), .ZN(n_192));
   NAND4_X1 i_243 (.A1(n_202), .A2(n_207), .A3(n_194), .A4(n_198), .ZN(n_199));
   NOR2_X1 i_244 (.A1(num_of_X[20]), .A2(num_of_X[21]), .ZN(n_198));
   NOR2_X1 i_245 (.A1(num_of_X[22]), .A2(num_of_X[23]), .ZN(n_194));
   INV_X1 i_246 (.A(n_203), .ZN(n_202));
   NAND3_X1 i_247 (.A1(n_204), .A2(n_205), .A3(n_206), .ZN(n_203));
   INV_X1 i_248 (.A(num_of_X[16]), .ZN(n_204));
   INV_X1 i_249 (.A(num_of_X[17]), .ZN(n_205));
   INV_X1 i_250 (.A(num_of_X[18]), .ZN(n_206));
   INV_X1 i_251 (.A(num_of_X[19]), .ZN(n_207));
   INV_X1 i_252 (.A(n_211), .ZN(n_143));
   NAND2_X1 i_253 (.A1(n_240), .A2(n_217), .ZN(n_211));
   INV_X1 i_254 (.A(n_221), .ZN(n_217));
   NAND3_X1 i_255 (.A1(n_239), .A2(n_227), .A3(n_145), .ZN(n_221));
   INV_X1 i_256 (.A(n_238), .ZN(n_227));
   NAND3_X1 i_257 (.A1(n_151), .A2(n_158), .A3(n_152), .ZN(n_238));
   INV_X1 i_258 (.A(num_of_X[40]), .ZN(n_151));
   INV_X1 i_259 (.A(num_of_X[41]), .ZN(n_152));
   INV_X1 i_260 (.A(num_of_X[47]), .ZN(n_158));
   NOR2_X1 i_261 (.A1(num_of_X[42]), .A2(num_of_X[43]), .ZN(n_145));
   INV_X1 i_262 (.A(n_154), .ZN(n_239));
   NAND3_X1 i_263 (.A1(n_155), .A2(n_157), .A3(n_156), .ZN(n_154));
   INV_X1 i_264 (.A(num_of_X[44]), .ZN(n_155));
   INV_X1 i_265 (.A(num_of_X[45]), .ZN(n_156));
   INV_X1 i_266 (.A(num_of_X[46]), .ZN(n_157));
   INV_X1 i_267 (.A(n_159), .ZN(n_240));
   NAND3_X1 i_268 (.A1(n_243), .A2(n_164), .A3(n_241), .ZN(n_159));
   NOR2_X1 i_269 (.A1(num_of_X[35]), .A2(num_of_X[39]), .ZN(n_241));
   INV_X1 i_270 (.A(n_242), .ZN(n_164));
   NAND3_X1 i_271 (.A1(n_167), .A2(n_168), .A3(n_166), .ZN(n_242));
   INV_X1 i_272 (.A(num_of_X[32]), .ZN(n_166));
   INV_X1 i_273 (.A(num_of_X[33]), .ZN(n_167));
   INV_X1 i_274 (.A(num_of_X[34]), .ZN(n_168));
   INV_X1 i_275 (.A(n_170), .ZN(n_243));
   NAND3_X1 i_276 (.A1(n_171), .A2(n_173), .A3(n_172), .ZN(n_170));
   INV_X1 i_277 (.A(num_of_X[36]), .ZN(n_171));
   INV_X1 i_278 (.A(num_of_X[37]), .ZN(n_172));
   INV_X1 i_279 (.A(num_of_X[38]), .ZN(n_173));
   INV_X1 i_280 (.A(n_209), .ZN(n_208));
   NAND4_X1 i_284 (.A1(n_222), .A2(n_228), .A3(n_216), .A4(n_210), .ZN(n_209));
   INV_X1 i_285 (.A(n_244), .ZN(n_210));
   NAND4_X1 i_286 (.A1(n_213), .A2(n_212), .A3(n_214), .A4(n_215), .ZN(n_244));
   INV_X1 i_287 (.A(num_of_X[12]), .ZN(n_212));
   INV_X1 i_288 (.A(num_of_X[13]), .ZN(n_213));
   INV_X1 i_291 (.A(num_of_X[14]), .ZN(n_214));
   INV_X1 i_292 (.A(num_of_X[15]), .ZN(n_215));
   INV_X1 i_293 (.A(n_232), .ZN(n_222));
   NAND4_X1 i_294 (.A1(n_234), .A2(n_233), .A3(n_235), .A4(n_236), .ZN(n_232));
   INV_X1 i_295 (.A(num_of_X[4]), .ZN(n_233));
   INV_X1 i_296 (.A(num_of_X[5]), .ZN(n_234));
   INV_X1 i_297 (.A(num_of_X[6]), .ZN(n_235));
   INV_X1 i_298 (.A(num_of_X[7]), .ZN(n_236));
   INV_X1 i_299 (.A(n_245), .ZN(n_216));
   NAND4_X1 i_300 (.A1(n_219), .A2(n_218), .A3(n_220), .A4(n_246), .ZN(n_245));
   INV_X1 i_301 (.A(num_of_X[8]), .ZN(n_218));
   INV_X1 i_302 (.A(num_of_X[9]), .ZN(n_219));
   INV_X1 i_303 (.A(num_of_X[10]), .ZN(n_220));
   INV_X1 i_304 (.A(num_of_X[11]), .ZN(n_246));
   INV_X1 i_305 (.A(n_229), .ZN(n_228));
   NAND4_X1 i_306 (.A1(n_237), .A2(n_230), .A3(n_231), .A4(n_247), .ZN(n_229));
   INV_X1 i_307 (.A(num_of_X[0]), .ZN(n_237));
   INV_X1 i_308 (.A(num_of_X[1]), .ZN(n_230));
   INV_X1 i_309 (.A(num_of_X[2]), .ZN(n_231));
   INV_X1 i_310 (.A(num_of_X[3]), .ZN(n_247));
   BUF_X1 rt_shieldBuf__1 (.A(n_192), .Z(n_248));
endmodule

module datapath__0_19(num_of_T, p_0);
   input [63:0]num_of_T;
   output [63:0]p_0;

   NAND2_X1 i_5 (.A1(n_3), .A2(n_259), .ZN(p_0[3]));
   NAND2_X1 i_6 (.A1(n_4), .A2(num_of_T[3]), .ZN(n_3));
   NAND2_X1 i_10 (.A1(n_8), .A2(n_6), .ZN(p_0[5]));
   NAND2_X1 i_11 (.A1(n_251), .A2(num_of_T[5]), .ZN(n_6));
   XNOR2_X1 i_17 (.A(n_14), .B(num_of_T[9]), .ZN(p_0[9]));
   NAND2_X1 i_18 (.A1(n_10), .A2(n_12), .ZN(p_0[10]));
   OAI21_X1 i_19 (.A(num_of_T[10]), .B1(n_14), .B2(num_of_T[9]), .ZN(n_10));
   OAI21_X1 i_20 (.A(n_22), .B1(n_11), .B2(n_223), .ZN(p_0[11]));
   INV_X1 i_21 (.A(n_12), .ZN(n_11));
   NAND3_X1 i_22 (.A1(n_13), .A2(n_222), .A3(n_221), .ZN(n_12));
   INV_X1 i_23 (.A(n_14), .ZN(n_13));
   NAND2_X1 i_25 (.A1(n_20), .A2(n_15), .ZN(p_0[12]));
   NAND2_X1 i_26 (.A1(n_22), .A2(num_of_T[12]), .ZN(n_15));
   XNOR2_X1 i_27 (.A(n_20), .B(num_of_T[13]), .ZN(p_0[13]));
   NAND2_X1 i_28 (.A1(n_16), .A2(n_18), .ZN(p_0[14]));
   OAI21_X1 i_29 (.A(num_of_T[14]), .B1(n_20), .B2(num_of_T[13]), .ZN(n_16));
   OAI21_X1 i_30 (.A(n_305), .B1(n_17), .B2(n_217), .ZN(p_0[15]));
   INV_X1 i_31 (.A(n_18), .ZN(n_17));
   NAND3_X1 i_32 (.A1(n_19), .A2(n_216), .A3(n_215), .ZN(n_18));
   INV_X1 i_33 (.A(n_20), .ZN(n_19));
   NAND2_X1 i_34 (.A1(n_21), .A2(n_214), .ZN(n_20));
   INV_X1 i_35 (.A(n_22), .ZN(n_21));
   NAND2_X1 i_36 (.A1(n_23), .A2(n_218), .ZN(n_22));
   NAND2_X1 i_39 (.A1(n_24), .A2(n_26), .ZN(p_0[17]));
   OAI21_X1 i_40 (.A(num_of_T[17]), .B1(n_305), .B2(num_of_T[16]), .ZN(n_24));
   OAI21_X1 i_41 (.A(n_38), .B1(n_25), .B2(n_209), .ZN(p_0[18]));
   INV_X1 i_42 (.A(n_26), .ZN(n_25));
   NAND3_X1 i_43 (.A1(n_210), .A2(n_208), .A3(n_207), .ZN(n_26));
   NAND2_X1 i_44 (.A1(n_36), .A2(n_27), .ZN(p_0[19]));
   NAND2_X1 i_45 (.A1(n_38), .A2(num_of_T[19]), .ZN(n_27));
   NAND2_X1 i_46 (.A1(n_30), .A2(n_28), .ZN(p_0[20]));
   NAND2_X1 i_47 (.A1(n_36), .A2(num_of_T[20]), .ZN(n_28));
   NAND2_X1 i_51 (.A1(n_31), .A2(n_33), .ZN(p_0[22]));
   NAND2_X1 i_52 (.A1(n_34), .A2(num_of_T[22]), .ZN(n_31));
   OAI21_X1 i_53 (.A(n_32), .B1(n_34), .B2(n_39), .ZN(p_0[23]));
   NAND2_X1 i_54 (.A1(n_33), .A2(num_of_T[23]), .ZN(n_32));
   NAND4_X1 i_55 (.A1(n_37), .A2(n_199), .A3(n_198), .A4(n_201), .ZN(n_33));
   NAND2_X1 i_61 (.A1(n_200), .A2(n_199), .ZN(n_39));
   XNOR2_X1 i_62 (.A(n_44), .B(num_of_T[24]), .ZN(p_0[24]));
   NAND2_X1 i_63 (.A1(n_40), .A2(n_42), .ZN(p_0[25]));
   OAI21_X1 i_64 (.A(num_of_T[25]), .B1(n_44), .B2(num_of_T[24]), .ZN(n_40));
   OAI21_X1 i_65 (.A(n_57), .B1(n_41), .B2(n_304), .ZN(p_0[26]));
   INV_X1 i_66 (.A(n_42), .ZN(n_41));
   NAND3_X1 i_67 (.A1(n_43), .A2(n_302), .A3(n_186), .ZN(n_42));
   INV_X1 i_68 (.A(n_44), .ZN(n_43));
   NAND2_X1 i_69 (.A1(n_210), .A2(n_194), .ZN(n_44));
   NAND2_X1 i_70 (.A1(n_55), .A2(n_45), .ZN(p_0[27]));
   NAND2_X1 i_71 (.A1(n_57), .A2(num_of_T[27]), .ZN(n_45));
   NAND2_X1 i_72 (.A1(n_46), .A2(n_48), .ZN(p_0[28]));
   NAND2_X1 i_73 (.A1(n_55), .A2(num_of_T[28]), .ZN(n_46));
   OAI21_X1 i_74 (.A(n_50), .B1(n_192), .B2(n_47), .ZN(p_0[29]));
   INV_X1 i_75 (.A(n_48), .ZN(n_47));
   NAND3_X1 i_76 (.A1(n_56), .A2(n_191), .A3(n_296), .ZN(n_48));
   OAI22_X1 i_77 (.A1(n_49), .A2(n_193), .B1(n_55), .B2(n_190), .ZN(p_0[30]));
   INV_X1 i_78 (.A(n_50), .ZN(n_49));
   NAND4_X1 i_79 (.A1(n_56), .A2(n_192), .A3(n_191), .A4(n_296), .ZN(n_50));
   NOR2_X1 i_80 (.A1(n_53), .A2(n_51), .ZN(p_0[31]));
   INV_X1 i_81 (.A(n_52), .ZN(n_51));
   NAND4_X1 i_82 (.A1(n_56), .A2(num_of_T[31]), .A3(n_296), .A4(n_189), .ZN(n_52));
   AOI21_X1 i_83 (.A(num_of_T[31]), .B1(n_54), .B2(n_189), .ZN(n_53));
   INV_X1 i_84 (.A(n_55), .ZN(n_54));
   NAND2_X1 i_85 (.A1(n_56), .A2(n_296), .ZN(n_55));
   INV_X1 i_86 (.A(n_57), .ZN(n_56));
   NAND3_X1 i_87 (.A1(n_210), .A2(n_194), .A3(n_184), .ZN(n_57));
   XNOR2_X1 i_88 (.A(n_94), .B(num_of_T[32]), .ZN(p_0[32]));
   NAND2_X1 i_89 (.A1(n_58), .A2(n_60), .ZN(p_0[33]));
   OAI21_X1 i_90 (.A(num_of_T[33]), .B1(n_94), .B2(num_of_T[32]), .ZN(n_58));
   OAI21_X1 i_91 (.A(n_62), .B1(n_59), .B2(n_170), .ZN(p_0[34]));
   INV_X1 i_92 (.A(n_60), .ZN(n_59));
   NAND3_X1 i_93 (.A1(n_93), .A2(n_169), .A3(n_168), .ZN(n_60));
   XNOR2_X1 i_94 (.A(n_62), .B(num_of_T[35]), .ZN(p_0[35]));
   OAI21_X1 i_98 (.A(n_66), .B1(n_63), .B2(n_174), .ZN(p_0[37]));
   INV_X1 i_99 (.A(n_64), .ZN(n_63));
   OAI21_X1 i_101 (.A(n_70), .B1(n_65), .B2(n_175), .ZN(p_0[38]));
   INV_X1 i_102 (.A(n_66), .ZN(n_65));
   NAND4_X1 i_103 (.A1(n_93), .A2(n_164), .A3(n_67), .A4(n_166), .ZN(n_66));
   INV_X1 i_104 (.A(n_68), .ZN(n_67));
   NAND2_X1 i_105 (.A1(n_174), .A2(n_173), .ZN(n_68));
   NAND2_X1 i_109 (.A1(n_73), .A2(n_71), .ZN(p_0[40]));
   NAND2_X1 i_110 (.A1(n_81), .A2(num_of_T[40]), .ZN(n_71));
   NAND2_X1 i_114 (.A1(n_74), .A2(n_77), .ZN(p_0[42]));
   NAND2_X1 i_115 (.A1(n_75), .A2(num_of_T[42]), .ZN(n_74));
   OAI21_X1 i_117 (.A(n_79), .B1(n_150), .B2(n_76), .ZN(p_0[43]));
   INV_X1 i_118 (.A(n_77), .ZN(n_76));
   NAND4_X1 i_119 (.A1(n_93), .A2(n_149), .A3(n_92), .A4(n_151), .ZN(n_77));
   OAI21_X1 i_125 (.A(n_85), .B1(n_82), .B2(n_158), .ZN(p_0[45]));
   INV_X1 i_126 (.A(n_83), .ZN(n_82));
   OAI21_X1 i_128 (.A(n_89), .B1(n_84), .B2(n_159), .ZN(p_0[46]));
   INV_X1 i_129 (.A(n_85), .ZN(n_84));
   NAND4_X1 i_130 (.A1(n_93), .A2(n_92), .A3(n_86), .A4(n_90), .ZN(n_85));
   INV_X1 i_131 (.A(n_87), .ZN(n_86));
   NAND2_X1 i_132 (.A1(n_158), .A2(n_157), .ZN(n_87));
   OAI21_X1 i_133 (.A(n_144), .B1(n_88), .B2(n_160), .ZN(p_0[47]));
   INV_X1 i_134 (.A(n_89), .ZN(n_88));
   NAND4_X1 i_135 (.A1(n_93), .A2(n_92), .A3(n_155), .A4(n_90), .ZN(n_89));
   NAND2_X1 i_137 (.A1(n_151), .A2(n_147), .ZN(n_91));
   NAND2_X1 i_141 (.A1(n_97), .A2(n_95), .ZN(p_0[48]));
   NAND2_X1 i_142 (.A1(n_144), .A2(num_of_T[48]), .ZN(n_95));
   OAI21_X1 i_143 (.A(n_99), .B1(n_96), .B2(n_244), .ZN(p_0[49]));
   INV_X1 i_144 (.A(n_97), .ZN(n_96));
   NAND2_X1 i_145 (.A1(n_143), .A2(n_243), .ZN(n_97));
   NAND2_X1 i_146 (.A1(n_98), .A2(n_101), .ZN(p_0[50]));
   NAND2_X1 i_147 (.A1(n_99), .A2(num_of_T[50]), .ZN(n_98));
   NAND3_X1 i_148 (.A1(n_143), .A2(n_244), .A3(n_243), .ZN(n_99));
   OAI21_X1 i_149 (.A(n_103), .B1(n_100), .B2(n_242), .ZN(p_0[51]));
   INV_X1 i_150 (.A(n_101), .ZN(n_100));
   NAND4_X1 i_151 (.A1(n_143), .A2(n_241), .A3(n_244), .A4(n_243), .ZN(n_101));
   NAND2_X1 i_152 (.A1(n_102), .A2(n_105), .ZN(p_0[52]));
   NAND2_X1 i_153 (.A1(n_103), .A2(num_of_T[52]), .ZN(n_102));
   NAND2_X1 i_154 (.A1(n_143), .A2(n_106), .ZN(n_103));
   OAI21_X1 i_155 (.A(n_109), .B1(n_104), .B2(n_238), .ZN(p_0[53]));
   INV_X1 i_156 (.A(n_105), .ZN(n_104));
   NAND3_X1 i_157 (.A1(n_143), .A2(n_237), .A3(n_106), .ZN(n_105));
   INV_X1 i_158 (.A(n_107), .ZN(n_106));
   NAND3_X1 i_159 (.A1(n_243), .A2(n_244), .A3(n_239), .ZN(n_107));
   OAI21_X1 i_160 (.A(n_111), .B1(n_108), .B2(n_245), .ZN(p_0[54]));
   INV_X1 i_161 (.A(n_109), .ZN(n_108));
   NAND2_X1 i_162 (.A1(n_143), .A2(n_233), .ZN(n_109));
   OAI21_X1 i_163 (.A(n_113), .B1(n_110), .B2(n_246), .ZN(p_0[55]));
   INV_X1 i_164 (.A(n_111), .ZN(n_110));
   NAND2_X1 i_165 (.A1(n_143), .A2(n_120), .ZN(n_111));
   NAND2_X1 i_166 (.A1(n_112), .A2(n_115), .ZN(p_0[56]));
   NAND2_X1 i_167 (.A1(n_113), .A2(num_of_T[56]), .ZN(n_112));
   NAND2_X1 i_168 (.A1(n_143), .A2(n_118), .ZN(n_113));
   OAI21_X1 i_169 (.A(n_117), .B1(n_114), .B2(n_231), .ZN(p_0[57]));
   INV_X1 i_170 (.A(n_115), .ZN(n_114));
   NAND3_X1 i_171 (.A1(n_143), .A2(n_230), .A3(n_118), .ZN(n_115));
   OAI21_X1 i_172 (.A(n_123), .B1(n_116), .B2(n_232), .ZN(p_0[58]));
   INV_X1 i_173 (.A(n_117), .ZN(n_116));
   NAND4_X1 i_174 (.A1(n_143), .A2(n_231), .A3(n_118), .A4(n_230), .ZN(n_117));
   INV_X1 i_175 (.A(n_119), .ZN(n_118));
   NAND2_X1 i_176 (.A1(n_120), .A2(n_246), .ZN(n_119));
   INV_X1 i_177 (.A(n_121), .ZN(n_120));
   NAND2_X1 i_178 (.A1(n_233), .A2(n_245), .ZN(n_121));
   OAI21_X1 i_179 (.A(n_125), .B1(n_122), .B2(n_247), .ZN(p_0[59]));
   INV_X1 i_180 (.A(n_123), .ZN(n_122));
   NAND2_X1 i_181 (.A1(n_143), .A2(n_226), .ZN(n_123));
   NAND2_X1 i_199 (.A1(n_138), .A2(n_142), .ZN(n_137));
   NAND2_X1 i_201 (.A1(n_141), .A2(n_140), .ZN(n_139));
   INV_X1 i_209 (.A(n_148), .ZN(n_147));
   NAND2_X1 i_210 (.A1(n_150), .A2(n_149), .ZN(n_148));
   INV_X1 i_211 (.A(num_of_T[42]), .ZN(n_149));
   INV_X1 i_212 (.A(num_of_T[43]), .ZN(n_150));
   INV_X1 i_213 (.A(n_152), .ZN(n_151));
   NAND2_X1 i_214 (.A1(n_154), .A2(n_153), .ZN(n_152));
   NAND3_X1 i_218 (.A1(n_159), .A2(n_158), .A3(n_157), .ZN(n_156));
   INV_X1 i_219 (.A(num_of_T[44]), .ZN(n_157));
   INV_X1 i_220 (.A(num_of_T[45]), .ZN(n_158));
   INV_X1 i_221 (.A(num_of_T[46]), .ZN(n_159));
   INV_X1 i_222 (.A(num_of_T[47]), .ZN(n_160));
   NAND3_X1 i_291 (.A1(n_231), .A2(n_230), .A3(n_232), .ZN(n_229));
   INV_X1 i_292 (.A(num_of_T[56]), .ZN(n_230));
   INV_X1 i_293 (.A(num_of_T[57]), .ZN(n_231));
   INV_X1 i_294 (.A(num_of_T[58]), .ZN(n_232));
   INV_X1 i_310 (.A(num_of_T[63]), .ZN(n_248));
   NAND2_X1 i_314 (.A1(n_257), .A2(n_252), .ZN(p_0[7]));
   NAND2_X1 i_315 (.A1(n_253), .A2(num_of_T[7]), .ZN(n_252));
   NAND2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0[1]));
   NAND2_X1 i_1 (.A1(num_of_T[0]), .A2(num_of_T[1]), .ZN(n_0));
   OAI21_X1 i_2 (.A(n_4), .B1(n_1), .B2(n_269), .ZN(p_0[2]));
   INV_X1 i_3 (.A(n_2), .ZN(n_1));
   NAND2_X1 i_4 (.A1(n_272), .A2(n_266), .ZN(n_2));
   NAND3_X1 i_7 (.A1(n_269), .A2(n_272), .A3(n_266), .ZN(n_4));
   OAI21_X1 i_8 (.A(n_253), .B1(n_5), .B2(n_258), .ZN(p_0[6]));
   NAND4_X1 i_9 (.A1(n_262), .A2(n_258), .A3(n_256), .A4(n_271), .ZN(n_253));
   INV_X1 i_12 (.A(n_8), .ZN(n_5));
   NAND3_X1 i_13 (.A1(n_262), .A2(n_256), .A3(n_271), .ZN(n_8));
   NAND2_X1 i_14 (.A1(n_14), .A2(n_7), .ZN(p_0[8]));
   NAND2_X1 i_15 (.A1(n_257), .A2(num_of_T[8]), .ZN(n_7));
   NAND2_X1 i_16 (.A1(n_23), .A2(n_250), .ZN(n_14));
   INV_X1 i_24 (.A(n_257), .ZN(n_23));
   NAND2_X1 i_37 (.A1(n_262), .A2(n_254), .ZN(n_257));
   INV_X1 i_38 (.A(n_9), .ZN(p_0[16]));
   NAND2_X1 i_273 (.A1(n_213), .A2(n_212), .ZN(n_9));
   NAND4_X1 i_274 (.A1(n_262), .A2(n_219), .A3(num_of_T[16]), .A4(n_254), 
      .ZN(n_212));
   NAND2_X1 i_275 (.A1(n_305), .A2(n_261), .ZN(n_213));
   INV_X1 i_321 (.A(num_of_T[16]), .ZN(n_261));
   NAND2_X1 i_323 (.A1(n_263), .A2(n_251), .ZN(p_0[4]));
   NAND2_X1 i_324 (.A1(n_259), .A2(num_of_T[4]), .ZN(n_263));
   NAND3_X1 i_326 (.A1(n_264), .A2(n_267), .A3(n_271), .ZN(n_251));
   INV_X1 i_327 (.A(n_265), .ZN(n_264));
   NAND2_X1 i_328 (.A1(n_272), .A2(n_266), .ZN(n_265));
   INV_X1 i_331 (.A(n_268), .ZN(n_267));
   NAND2_X1 i_332 (.A1(n_269), .A2(n_270), .ZN(n_268));
   INV_X1 i_111 (.A(n_72), .ZN(n_219));
   NAND2_X1 i_112 (.A1(n_218), .A2(n_273), .ZN(n_72));
   INV_X1 i_113 (.A(n_124), .ZN(n_226));
   NAND3_X1 i_116 (.A1(n_233), .A2(n_178), .A3(n_162), .ZN(n_124));
   INV_X1 i_138 (.A(n_228), .ZN(n_194));
   NAND2_X1 i_140 (.A1(n_240), .A2(n_207), .ZN(n_126));
   OAI21_X1 i_182 (.A(n_75), .B1(n_154), .B2(n_127), .ZN(p_0[41]));
   INV_X1 i_183 (.A(n_73), .ZN(n_127));
   NAND3_X1 i_184 (.A1(n_93), .A2(n_153), .A3(n_92), .ZN(n_73));
   INV_X1 i_185 (.A(num_of_T[40]), .ZN(n_153));
   NAND2_X1 i_186 (.A1(n_80), .A2(n_151), .ZN(n_75));
   INV_X1 i_189 (.A(num_of_T[41]), .ZN(n_154));
   NAND2_X1 i_228 (.A1(n_246), .A2(n_245), .ZN(n_163));
   INV_X1 i_229 (.A(num_of_T[54]), .ZN(n_245));
   INV_X1 i_230 (.A(num_of_T[55]), .ZN(n_246));
   INV_X1 i_245 (.A(n_144), .ZN(n_143));
   NAND4_X1 i_246 (.A1(n_202), .A2(n_210), .A3(n_179), .A4(n_196), .ZN(n_144));
   INV_X1 i_247 (.A(n_180), .ZN(n_179));
   INV_X1 i_262 (.A(n_197), .ZN(n_196));
   INV_X1 i_340 (.A(num_of_T[63]), .ZN(n_277));
   NAND2_X1 i_48 (.A1(n_92), .A2(n_155), .ZN(n_180));
   INV_X1 i_49 (.A(n_29), .ZN(n_240));
   NAND2_X1 i_50 (.A1(n_209), .A2(n_208), .ZN(n_29));
   NAND2_X1 i_56 (.A1(n_285), .A2(n_281), .ZN(n_228));
   INV_X1 i_57 (.A(n_35), .ZN(n_233));
   NAND2_X1 i_58 (.A1(n_292), .A2(n_239), .ZN(n_35));
   INV_X1 i_59 (.A(n_81), .ZN(n_80));
   INV_X1 i_127 (.A(n_78), .ZN(n_184));
   NAND3_X1 i_136 (.A1(n_304), .A2(n_302), .A3(n_186), .ZN(n_78));
   NAND2_X1 i_139 (.A1(n_37), .A2(n_198), .ZN(n_36));
   INV_X1 i_187 (.A(n_38), .ZN(n_37));
   NAND2_X1 i_188 (.A1(n_210), .A2(n_130), .ZN(n_38));
   OAI21_X1 i_190 (.A(n_34), .B1(n_128), .B2(n_284), .ZN(p_0[21]));
   INV_X1 i_191 (.A(n_30), .ZN(n_128));
   NAND4_X1 i_192 (.A1(n_210), .A2(n_283), .A3(n_198), .A4(n_130), .ZN(n_30));
   NAND4_X1 i_193 (.A1(n_210), .A2(n_198), .A3(n_130), .A4(n_201), .ZN(n_34));
   INV_X1 i_194 (.A(n_129), .ZN(n_201));
   NAND2_X1 i_195 (.A1(n_284), .A2(n_283), .ZN(n_129));
   INV_X1 i_196 (.A(n_126), .ZN(n_130));
   OAI21_X1 i_197 (.A(n_83), .B1(n_133), .B2(n_135), .ZN(p_0[44]));
   NAND4_X1 i_198 (.A1(n_210), .A2(n_202), .A3(n_92), .A4(n_131), .ZN(n_83));
   INV_X1 i_200 (.A(n_132), .ZN(n_131));
   NAND2_X1 i_202 (.A1(n_90), .A2(n_157), .ZN(n_132));
   INV_X1 i_203 (.A(n_79), .ZN(n_133));
   NAND4_X1 i_204 (.A1(n_210), .A2(n_202), .A3(n_90), .A4(n_92), .ZN(n_79));
   INV_X1 i_205 (.A(n_134), .ZN(n_92));
   NAND2_X1 i_206 (.A1(n_206), .A2(n_166), .ZN(n_134));
   INV_X1 i_207 (.A(n_91), .ZN(n_90));
   INV_X1 i_208 (.A(num_of_T[44]), .ZN(n_135));
   OAI21_X1 i_215 (.A(n_146), .B1(n_136), .B2(n_140), .ZN(p_0[60]));
   INV_X1 i_216 (.A(n_125), .ZN(n_136));
   NAND4_X1 i_217 (.A1(n_306), .A2(n_204), .A3(n_202), .A4(n_288), .ZN(n_125));
   OAI21_X1 i_223 (.A(n_176), .B1(n_145), .B2(n_141), .ZN(p_0[61]));
   INV_X1 i_224 (.A(n_146), .ZN(n_145));
   NAND4_X1 i_225 (.A1(n_306), .A2(n_204), .A3(n_202), .A4(n_161), .ZN(n_146));
   INV_X1 i_226 (.A(n_167), .ZN(n_161));
   NAND4_X1 i_227 (.A1(n_292), .A2(n_140), .A3(n_239), .A4(n_290), .ZN(n_167));
   INV_X1 i_231 (.A(num_of_T[60]), .ZN(n_140));
   INV_X1 i_232 (.A(num_of_T[61]), .ZN(n_141));
   OAI21_X1 i_233 (.A(n_185), .B1(n_172), .B2(n_142), .ZN(p_0[62]));
   INV_X1 i_234 (.A(n_176), .ZN(n_172));
   NAND4_X1 i_235 (.A1(n_210), .A2(n_204), .A3(n_202), .A4(n_177), .ZN(n_176));
   INV_X1 i_236 (.A(n_181), .ZN(n_177));
   NAND4_X1 i_237 (.A1(n_292), .A2(n_138), .A3(n_239), .A4(n_290), .ZN(n_181));
   INV_X1 i_238 (.A(n_139), .ZN(n_138));
   INV_X1 i_239 (.A(num_of_T[62]), .ZN(n_142));
   OAI21_X1 i_240 (.A(n_287), .B1(n_183), .B2(n_248), .ZN(p_0[63]));
   INV_X1 i_241 (.A(n_185), .ZN(n_183));
   NAND4_X1 i_242 (.A1(n_210), .A2(n_204), .A3(n_202), .A4(n_195), .ZN(n_185));
   INV_X1 i_243 (.A(n_203), .ZN(n_195));
   NAND4_X1 i_244 (.A1(n_292), .A2(n_295), .A3(n_239), .A4(n_290), .ZN(n_203));
   INV_X1 i_248 (.A(n_205), .ZN(n_204));
   NAND4_X1 i_249 (.A1(n_206), .A2(n_155), .A3(n_249), .A4(n_166), .ZN(n_205));
   NOR2_X1 i_250 (.A1(n_235), .A2(n_220), .ZN(n_206));
   NAND2_X1 i_251 (.A1(n_234), .A2(n_227), .ZN(n_220));
   INV_X1 i_252 (.A(num_of_T[35]), .ZN(n_227));
   INV_X1 i_253 (.A(num_of_T[39]), .ZN(n_234));
   NAND3_X1 i_254 (.A1(n_175), .A2(n_174), .A3(n_173), .ZN(n_235));
   INV_X1 i_255 (.A(num_of_T[36]), .ZN(n_173));
   INV_X1 i_256 (.A(num_of_T[37]), .ZN(n_174));
   INV_X1 i_257 (.A(num_of_T[38]), .ZN(n_175));
   NAND3_X1 i_259 (.A1(n_170), .A2(n_169), .A3(n_168), .ZN(n_236));
   INV_X1 i_260 (.A(num_of_T[32]), .ZN(n_168));
   INV_X1 i_261 (.A(num_of_T[33]), .ZN(n_169));
   INV_X1 i_263 (.A(num_of_T[34]), .ZN(n_170));
   INV_X1 i_264 (.A(n_197), .ZN(n_249));
   NAND3_X1 i_265 (.A1(n_151), .A2(n_160), .A3(n_147), .ZN(n_197));
   INV_X1 i_266 (.A(n_156), .ZN(n_155));
   NAND4_X1 i_271 (.A1(n_262), .A2(n_273), .A3(n_254), .A4(n_218), .ZN(n_211));
   INV_X1 i_272 (.A(n_255), .ZN(n_218));
   NAND4_X1 i_276 (.A1(n_223), .A2(n_222), .A3(n_221), .A4(n_250), .ZN(n_255));
   INV_X1 i_277 (.A(num_of_T[8]), .ZN(n_250));
   INV_X1 i_278 (.A(num_of_T[9]), .ZN(n_221));
   INV_X1 i_279 (.A(num_of_T[10]), .ZN(n_222));
   INV_X1 i_280 (.A(num_of_T[11]), .ZN(n_223));
   INV_X1 i_281 (.A(n_260), .ZN(n_254));
   NAND4_X1 i_282 (.A1(n_274), .A2(n_258), .A3(n_256), .A4(n_271), .ZN(n_260));
   INV_X1 i_283 (.A(num_of_T[4]), .ZN(n_271));
   INV_X1 i_284 (.A(num_of_T[5]), .ZN(n_256));
   INV_X1 i_285 (.A(num_of_T[6]), .ZN(n_258));
   INV_X1 i_286 (.A(num_of_T[7]), .ZN(n_274));
   INV_X1 i_287 (.A(n_275), .ZN(n_273));
   NAND4_X1 i_288 (.A1(n_217), .A2(n_216), .A3(n_215), .A4(n_214), .ZN(n_275));
   INV_X1 i_289 (.A(num_of_T[12]), .ZN(n_214));
   INV_X1 i_290 (.A(num_of_T[13]), .ZN(n_215));
   INV_X1 i_295 (.A(num_of_T[14]), .ZN(n_216));
   INV_X1 i_296 (.A(num_of_T[15]), .ZN(n_217));
   INV_X1 i_297 (.A(n_259), .ZN(n_262));
   NAND4_X1 i_298 (.A1(n_270), .A2(n_269), .A3(n_266), .A4(n_272), .ZN(n_259));
   INV_X1 i_299 (.A(num_of_T[0]), .ZN(n_272));
   INV_X1 i_300 (.A(num_of_T[1]), .ZN(n_266));
   INV_X1 i_301 (.A(num_of_T[2]), .ZN(n_269));
   INV_X1 i_302 (.A(num_of_T[3]), .ZN(n_270));
   NAND3_X1 i_313 (.A1(n_193), .A2(n_192), .A3(n_191), .ZN(n_190));
   INV_X1 i_316 (.A(num_of_T[28]), .ZN(n_191));
   INV_X1 i_317 (.A(num_of_T[29]), .ZN(n_192));
   INV_X1 i_318 (.A(num_of_T[30]), .ZN(n_193));
   NAND4_X1 i_320 (.A1(n_284), .A2(n_283), .A3(n_209), .A4(n_208), .ZN(n_282));
   INV_X1 i_322 (.A(num_of_T[17]), .ZN(n_208));
   INV_X1 i_325 (.A(num_of_T[18]), .ZN(n_209));
   INV_X1 i_329 (.A(num_of_T[20]), .ZN(n_283));
   INV_X1 i_330 (.A(num_of_T[21]), .ZN(n_284));
   NAND4_X1 i_334 (.A1(n_200), .A2(n_199), .A3(n_198), .A4(n_207), .ZN(n_286));
   INV_X1 i_335 (.A(num_of_T[16]), .ZN(n_207));
   INV_X1 i_336 (.A(num_of_T[19]), .ZN(n_198));
   INV_X1 i_337 (.A(num_of_T[22]), .ZN(n_199));
   INV_X1 i_338 (.A(num_of_T[23]), .ZN(n_200));
   NAND4_X1 i_339 (.A1(n_288), .A2(n_143), .A3(n_295), .A4(n_277), .ZN(n_287));
   INV_X1 i_341 (.A(n_289), .ZN(n_288));
   NAND3_X1 i_342 (.A1(n_292), .A2(n_239), .A3(n_290), .ZN(n_289));
   INV_X1 i_343 (.A(n_291), .ZN(n_290));
   NAND3_X1 i_344 (.A1(n_247), .A2(n_178), .A3(n_162), .ZN(n_291));
   INV_X1 i_345 (.A(n_163), .ZN(n_162));
   INV_X1 i_346 (.A(n_229), .ZN(n_178));
   INV_X1 i_347 (.A(num_of_T[59]), .ZN(n_247));
   INV_X1 i_348 (.A(n_293), .ZN(n_292));
   NAND4_X1 i_349 (.A1(n_238), .A2(n_237), .A3(n_244), .A4(n_243), .ZN(n_293));
   INV_X1 i_350 (.A(num_of_T[48]), .ZN(n_243));
   INV_X1 i_351 (.A(num_of_T[49]), .ZN(n_244));
   INV_X1 i_352 (.A(num_of_T[52]), .ZN(n_237));
   INV_X1 i_353 (.A(num_of_T[53]), .ZN(n_238));
   INV_X1 i_354 (.A(n_294), .ZN(n_239));
   NAND2_X1 i_355 (.A1(n_242), .A2(n_241), .ZN(n_294));
   INV_X1 i_356 (.A(num_of_T[50]), .ZN(n_241));
   INV_X1 i_357 (.A(num_of_T[51]), .ZN(n_242));
   INV_X1 i_358 (.A(n_137), .ZN(n_295));
   BUF_X1 rt_shieldBuf__1 (.A(n_182), .Z(n_296));
   NAND3_X1 i_60 (.A1(n_306), .A2(n_303), .A3(n_276), .ZN(n_70));
   NAND2_X1 i_95 (.A1(n_93), .A2(n_166), .ZN(n_62));
   INV_X1 i_96 (.A(n_93), .ZN(n_94));
   NOR2_X1 i_97 (.A1(n_211), .A2(n_280), .ZN(n_93));
   NAND2_X1 i_100 (.A1(n_64), .A2(n_165), .ZN(p_0[36]));
   NAND4_X1 i_106 (.A1(n_210), .A2(n_166), .A3(n_202), .A4(n_61), .ZN(n_64));
   INV_X1 i_107 (.A(n_69), .ZN(n_61));
   NAND2_X1 i_108 (.A1(n_164), .A2(n_173), .ZN(n_69));
   OAI21_X1 i_120 (.A(num_of_T[36]), .B1(n_211), .B2(n_171), .ZN(n_165));
   NAND4_X1 i_121 (.A1(n_297), .A2(n_164), .A3(n_166), .A4(n_285), .ZN(n_171));
   NAND2_X1 i_122 (.A1(n_224), .A2(n_81), .ZN(p_0[39]));
   OAI21_X1 i_123 (.A(num_of_T[39]), .B1(n_305), .B2(n_225), .ZN(n_224));
   NAND2_X1 i_124 (.A1(n_276), .A2(n_303), .ZN(n_225));
   INV_X1 i_258 (.A(n_278), .ZN(n_276));
   NAND4_X1 i_267 (.A1(n_285), .A2(n_164), .A3(n_279), .A4(n_166), .ZN(n_278));
   INV_X1 i_268 (.A(n_236), .ZN(n_166));
   INV_X1 i_269 (.A(n_235), .ZN(n_279));
   INV_X1 i_270 (.A(num_of_T[35]), .ZN(n_164));
   NAND3_X1 i_303 (.A1(n_210), .A2(n_92), .A3(n_202), .ZN(n_81));
   INV_X1 i_304 (.A(n_280), .ZN(n_202));
   NAND2_X1 i_305 (.A1(n_297), .A2(n_285), .ZN(n_280));
   INV_X1 i_306 (.A(n_298), .ZN(n_297));
   NAND4_X1 i_307 (.A1(n_281), .A2(n_186), .A3(n_189), .A4(n_299), .ZN(n_298));
   INV_X1 i_308 (.A(n_300), .ZN(n_299));
   NAND4_X1 i_309 (.A1(n_301), .A2(n_182), .A3(n_187), .A4(n_188), .ZN(n_300));
   INV_X1 i_311 (.A(num_of_T[25]), .ZN(n_187));
   INV_X1 i_312 (.A(num_of_T[26]), .ZN(n_188));
   INV_X1 i_319 (.A(num_of_T[27]), .ZN(n_182));
   INV_X1 i_333 (.A(num_of_T[31]), .ZN(n_301));
   INV_X1 i_359 (.A(n_282), .ZN(n_281));
   INV_X1 i_360 (.A(n_190), .ZN(n_189));
   INV_X1 i_361 (.A(num_of_T[24]), .ZN(n_186));
   INV_X1 i_362 (.A(n_286), .ZN(n_285));
   INV_X1 i_363 (.A(n_211), .ZN(n_210));
   BUF_X1 rt_shieldBuf__1__1__0 (.A(n_187), .Z(n_302));
   BUF_X1 rt_shieldBuf__1__1__1 (.A(n_297), .Z(n_303));
   BUF_X1 rt_shieldBuf__1__1__2 (.A(n_188), .Z(n_304));
   BUF_X1 rt_shieldBuf__1__1__3 (.A(n_211), .Z(n_305));
   BUF_X1 rt_shieldBuf__1__1__4 (.A(n_210), .Z(n_306));
endmodule

module datapath__1_253(X_Count, p_0, T_Count, num_of_X);
   input [7:0]X_Count;
   output [12:0]p_0;
   input [7:0]T_Count;
   input [12:0]num_of_X;

   INV_X1 i_0 (.A(n_0), .ZN(p_0[0]));
   XOR2_X1 i_1 (.A(X_Count[0]), .B(n_1), .Z(n_0));
   NAND2_X1 i_2 (.A1(T_Count[0]), .A2(n_657), .ZN(n_1));
   XNOR2_X1 i_3 (.A(n_2), .B(n_322), .ZN(p_0[1]));
   NAND2_X1 i_4 (.A1(n_3), .A2(n_325), .ZN(n_2));
   INV_X1 i_5 (.A(n_324), .ZN(n_3));
   XOR2_X1 i_6 (.A(n_321), .B(n_4), .Z(p_0[2]));
   XNOR2_X1 i_7 (.A(n_329), .B(n_333), .ZN(n_4));
   XOR2_X1 i_8 (.A(n_319), .B(n_5), .Z(p_0[3]));
   NAND2_X1 i_9 (.A1(n_338), .A2(n_336), .ZN(n_5));
   XOR2_X1 i_10 (.A(n_7), .B(n_6), .Z(p_0[4]));
   NAND2_X1 i_11 (.A1(n_346), .A2(n_349), .ZN(n_6));
   NAND2_X1 i_12 (.A1(n_338), .A2(n_318), .ZN(n_7));
   INV_X1 i_13 (.A(n_8), .ZN(p_0[5]));
   XOR2_X1 i_14 (.A(n_316), .B(n_9), .Z(n_8));
   NAND2_X1 i_15 (.A1(n_359), .A2(n_362), .ZN(n_9));
   INV_X1 i_16 (.A(n_10), .ZN(p_0[6]));
   XNOR2_X1 i_17 (.A(n_11), .B(n_315), .ZN(n_10));
   NAND2_X1 i_18 (.A1(n_373), .A2(n_371), .ZN(n_11));
   AOI22_X1 i_49 (.A1(n_317), .A2(n_349), .B1(n_368), .B2(n_360), .ZN(n_37));
   NAND2_X1 i_71 (.A1(n_209), .A2(n_197), .ZN(n_58));
   XOR2_X1 i_85 (.A(n_74), .B(n_73), .Z(n_72));
   NAND2_X1 i_86 (.A1(T_Count[4]), .A2(num_of_X[8]), .ZN(n_73));
   NAND2_X1 i_87 (.A1(n_255), .A2(num_of_X[9]), .ZN(n_74));
   INV_X1 i_90 (.A(n_178), .ZN(n_77));
   XOR2_X1 i_98 (.A(n_87), .B(n_86), .Z(n_85));
   NAND2_X1 i_99 (.A1(T_Count[2]), .A2(num_of_X[10]), .ZN(n_86));
   NAND2_X1 i_100 (.A1(T_Count[0]), .A2(num_of_X[12]), .ZN(n_87));
   NAND2_X1 i_101 (.A1(T_Count[1]), .A2(num_of_X[11]), .ZN(n_88));
   XNOR2_X1 i_104 (.A(n_92), .B(n_95), .ZN(n_91));
   XOR2_X1 i_105 (.A(n_94), .B(n_93), .Z(n_92));
   OAI21_X1 i_106 (.A(n_203), .B1(n_200), .B2(n_205), .ZN(n_93));
   NAND2_X1 i_107 (.A1(T_Count[6]), .A2(num_of_X[6]), .ZN(n_94));
   XNOR2_X1 i_108 (.A(n_188), .B(n_96), .ZN(n_95));
   NAND2_X1 i_109 (.A1(T_Count[5]), .A2(num_of_X[7]), .ZN(n_96));
   INV_X1 i_110 (.A(n_98), .ZN(n_97));
   OAI21_X1 i_111 (.A(n_187), .B1(n_99), .B2(n_184), .ZN(n_98));
   INV_X1 i_112 (.A(n_190), .ZN(n_99));
   NAND2_X1 i_192 (.A1(T_Count[5]), .A2(num_of_X[6]), .ZN(n_179));
   NAND2_X1 i_197 (.A1(n_255), .A2(num_of_X[8]), .ZN(n_184));
   NAND2_X1 i_199 (.A1(n_190), .A2(n_187), .ZN(n_186));
   NAND3_X1 i_200 (.A1(n_188), .A2(T_Count[6]), .A3(num_of_X[4]), .ZN(n_187));
   INV_X1 i_201 (.A(n_189), .ZN(n_188));
   NAND2_X1 i_202 (.A1(T_Count[7]), .A2(num_of_X[5]), .ZN(n_189));
   OAI22_X1 i_203 (.A1(n_306), .A2(n_431), .B1(n_417), .B2(n_298), .ZN(n_190));
   INV_X1 i_213 (.A(n_201), .ZN(n_200));
   NAND4_X1 i_214 (.A1(T_Count[1]), .A2(T_Count[0]), .A3(num_of_X[11]), .A4(
      num_of_X[10]), .ZN(n_201));
   INV_X1 i_215 (.A(n_203), .ZN(n_202));
   OAI21_X1 i_216 (.A(n_204), .B1(n_491), .B2(n_277), .ZN(n_203));
   NAND2_X1 i_217 (.A1(T_Count[0]), .A2(num_of_X[11]), .ZN(n_204));
   INV_X1 i_218 (.A(n_206), .ZN(n_205));
   NAND2_X1 i_219 (.A1(T_Count[2]), .A2(num_of_X[9]), .ZN(n_206));
   NAND2_X1 i_279 (.A1(n_283), .A2(n_296), .ZN(n_266));
   NAND3_X1 i_336 (.A1(X_Count[0]), .A2(T_Count[0]), .A3(n_657), .ZN(n_323));
   NAND3_X1 i_344 (.A1(n_539), .A2(n_538), .A3(n_537), .ZN(n_331));
   AOI21_X1 i_345 (.A(n_538), .B1(n_539), .B2(n_537), .ZN(n_332));
   NAND3_X1 i_347 (.A1(n_335), .A2(n_525), .A3(n_526), .ZN(n_334));
   NAND2_X1 i_348 (.A1(T_Count[2]), .A2(n_657), .ZN(n_335));
   NAND2_X1 i_350 (.A1(n_344), .A2(n_343), .ZN(n_337));
   NOR2_X1 i_352 (.A1(n_341), .A2(n_340), .ZN(n_339));
   AOI21_X1 i_353 (.A(n_523), .B1(n_527), .B2(n_528), .ZN(n_340));
   INV_X1 i_354 (.A(n_342), .ZN(n_341));
   NAND3_X1 i_355 (.A1(n_528), .A2(n_527), .A3(n_523), .ZN(n_342));
   NAND3_X1 i_356 (.A1(n_517), .A2(n_513), .A3(n_516), .ZN(n_343));
   NAND2_X1 i_357 (.A1(n_345), .A2(n_515), .ZN(n_344));
   NAND2_X1 i_358 (.A1(n_513), .A2(n_517), .ZN(n_345));
   INV_X1 i_360 (.A(n_350), .ZN(n_347));
   NAND2_X1 i_361 (.A1(n_356), .A2(n_521), .ZN(n_348));
   NAND2_X1 i_363 (.A1(n_353), .A2(n_351), .ZN(n_350));
   OAI21_X1 i_364 (.A(n_506), .B1(n_352), .B2(n_511), .ZN(n_351));
   INV_X1 i_365 (.A(n_512), .ZN(n_352));
   NAND4_X1 i_366 (.A1(n_354), .A2(n_512), .A3(n_508), .A4(n_507), .ZN(n_353));
   NAND2_X1 i_367 (.A1(n_355), .A2(n_532), .ZN(n_354));
   NAND2_X1 i_368 (.A1(n_514), .A2(n_513), .ZN(n_355));
   NAND2_X1 i_369 (.A1(n_357), .A2(n_358), .ZN(n_356));
   NAND2_X1 i_370 (.A1(n_522), .A2(n_528), .ZN(n_357));
   INV_X1 i_371 (.A(n_542), .ZN(n_358));
   INV_X1 i_373 (.A(n_363), .ZN(n_360));
   NAND3_X1 i_377 (.A1(n_552), .A2(n_580), .A3(n_577), .ZN(n_364));
   NAND3_X1 i_378 (.A1(n_366), .A2(n_557), .A3(n_553), .ZN(n_365));
   NAND2_X1 i_379 (.A1(n_577), .A2(n_580), .ZN(n_366));
   NAND2_X1 i_396 (.A1(n_449), .A2(n_448), .ZN(n_383));
   INV_X1 i_409 (.A(n_646), .ZN(n_396));
   NAND2_X1 i_416 (.A1(n_407), .A2(n_405), .ZN(n_403));
   OR2_X1 i_417 (.A1(n_407), .A2(n_405), .ZN(n_404));
   NAND2_X1 i_419 (.A1(n_464), .A2(n_460), .ZN(n_406));
   NAND2_X1 i_420 (.A1(n_409), .A2(n_408), .ZN(n_407));
   NAND2_X1 i_423 (.A1(n_412), .A2(n_411), .ZN(n_410));
   NAND2_X1 i_426 (.A1(n_414), .A2(n_415), .ZN(n_413));
   NAND2_X1 i_433 (.A1(n_423), .A2(n_421), .ZN(n_420));
   NAND2_X1 i_636 (.A1(n_625), .A2(n_624), .ZN(n_623));
   BUF_X1 rt_shieldBuf__1 (.A(num_of_X[0]), .Z(n_657));
   NAND2_X1 i_19 (.A1(n_292), .A2(n_304), .ZN(n_449));
   INV_X1 i_20 (.A(T_Count[7]), .ZN(n_306));
   INV_X1 i_21 (.A(n_136), .ZN(n_315));
   NAND2_X1 i_22 (.A1(n_319), .A2(n_336), .ZN(n_318));
   INV_X1 i_23 (.A(n_138), .ZN(n_319));
   NAND2_X1 i_24 (.A1(n_523), .A2(n_334), .ZN(n_333));
   INV_X1 i_25 (.A(n_143), .ZN(n_329));
   INV_X1 i_26 (.A(n_12), .ZN(p_0[7]));
   XOR2_X1 i_27 (.A(n_134), .B(n_13), .Z(n_12));
   NAND2_X1 i_28 (.A1(n_131), .A2(n_161), .ZN(n_13));
   INV_X1 i_29 (.A(n_14), .ZN(p_0[8]));
   XNOR2_X1 i_30 (.A(n_130), .B(n_15), .ZN(n_14));
   NAND2_X1 i_31 (.A1(n_127), .A2(n_169), .ZN(n_15));
   INV_X1 i_32 (.A(n_16), .ZN(p_0[9]));
   XNOR2_X1 i_33 (.A(n_125), .B(n_17), .ZN(n_16));
   AND2_X1 i_34 (.A1(n_83), .A2(n_54), .ZN(n_17));
   NAND2_X1 i_35 (.A1(n_20), .A2(n_18), .ZN(p_0[10]));
   NAND3_X1 i_36 (.A1(n_27), .A2(n_83), .A3(n_19), .ZN(n_18));
   NAND2_X1 i_37 (.A1(n_40), .A2(n_64), .ZN(n_19));
   NAND3_X1 i_38 (.A1(n_21), .A2(n_64), .A3(n_40), .ZN(n_20));
   NAND2_X1 i_39 (.A1(n_27), .A2(n_83), .ZN(n_21));
   INV_X1 i_40 (.A(n_22), .ZN(p_0[11]));
   OAI21_X1 i_41 (.A(n_23), .B1(n_28), .B2(n_42), .ZN(n_22));
   NAND2_X1 i_42 (.A1(n_26), .A2(n_24), .ZN(n_23));
   INV_X1 i_43 (.A(n_25), .ZN(n_24));
   NAND2_X1 i_44 (.A1(n_42), .A2(n_40), .ZN(n_25));
   NAND2_X1 i_45 (.A1(n_27), .A2(n_36), .ZN(n_26));
   OAI21_X1 i_46 (.A(n_30), .B1(n_130), .B2(n_126), .ZN(n_27));
   AOI21_X1 i_47 (.A(n_39), .B1(n_29), .B2(n_36), .ZN(n_28));
   OAI21_X1 i_48 (.A(n_30), .B1(n_32), .B2(n_126), .ZN(n_29));
   INV_X1 i_50 (.A(n_31), .ZN(n_30));
   NAND2_X1 i_51 (.A1(n_54), .A2(n_169), .ZN(n_31));
   AOI21_X1 i_52 (.A(n_160), .B1(n_33), .B2(n_131), .ZN(n_32));
   NAND2_X1 i_53 (.A1(n_34), .A2(n_373), .ZN(n_33));
   OAI21_X1 i_54 (.A(n_371), .B1(n_37), .B2(n_35), .ZN(n_34));
   INV_X1 i_55 (.A(n_362), .ZN(n_35));
   INV_X1 i_56 (.A(n_38), .ZN(n_36));
   NAND2_X1 i_57 (.A1(n_64), .A2(n_83), .ZN(n_38));
   INV_X1 i_58 (.A(n_40), .ZN(n_39));
   NAND3_X1 i_59 (.A1(n_51), .A2(n_41), .A3(n_67), .ZN(n_40));
   INV_X1 i_60 (.A(n_670), .ZN(n_41));
   NAND2_X1 i_61 (.A1(n_59), .A2(n_43), .ZN(n_42));
   NAND3_X1 i_62 (.A1(n_61), .A2(n_66), .A3(n_442), .ZN(n_43));
   NAND2_X1 i_63 (.A1(n_45), .A2(n_44), .ZN(p_0[12]));
   NAND4_X1 i_64 (.A1(n_55), .A2(n_47), .A3(n_398), .A4(n_394), .ZN(n_44));
   NAND2_X1 i_65 (.A1(n_46), .A2(n_393), .ZN(n_45));
   NAND2_X1 i_66 (.A1(n_55), .A2(n_47), .ZN(n_46));
   INV_X1 i_67 (.A(n_48), .ZN(n_47));
   NAND2_X1 i_68 (.A1(n_52), .A2(n_49), .ZN(n_48));
   NAND4_X1 i_69 (.A1(n_50), .A2(n_51), .A3(n_442), .A4(n_61), .ZN(n_49));
   NAND2_X1 i_70 (.A1(n_670), .A2(n_67), .ZN(n_50));
   INV_X1 i_72 (.A(n_65), .ZN(n_51));
   NAND3_X1 i_73 (.A1(n_59), .A2(n_64), .A3(n_53), .ZN(n_52));
   INV_X1 i_74 (.A(n_54), .ZN(n_53));
   NAND3_X1 i_75 (.A1(n_89), .A2(n_670), .A3(n_128), .ZN(n_54));
   NAND2_X1 i_76 (.A1(n_125), .A2(n_56), .ZN(n_55));
   INV_X1 i_77 (.A(n_57), .ZN(n_56));
   NAND3_X1 i_78 (.A1(n_59), .A2(n_83), .A3(n_64), .ZN(n_57));
   NAND2_X1 i_79 (.A1(n_60), .A2(n_67), .ZN(n_59));
   NAND2_X1 i_80 (.A1(n_61), .A2(n_442), .ZN(n_60));
   OAI21_X1 i_81 (.A(n_495), .B1(n_63), .B2(n_62), .ZN(n_61));
   AOI21_X1 i_82 (.A(n_472), .B1(n_455), .B2(n_452), .ZN(n_62));
   INV_X1 i_83 (.A(n_451), .ZN(n_63));
   OAI21_X1 i_84 (.A(n_670), .B1(n_66), .B2(n_65), .ZN(n_64));
   AOI21_X1 i_88 (.A(n_68), .B1(n_71), .B2(n_70), .ZN(n_65));
   INV_X1 i_89 (.A(n_67), .ZN(n_66));
   NAND3_X1 i_91 (.A1(n_71), .A2(n_68), .A3(n_70), .ZN(n_67));
   NAND2_X1 i_92 (.A1(n_69), .A2(n_102), .ZN(n_68));
   NAND2_X1 i_93 (.A1(n_105), .A2(n_103), .ZN(n_69));
   NAND3_X1 i_94 (.A1(n_82), .A2(n_76), .A3(n_585), .ZN(n_70));
   NAND2_X1 i_95 (.A1(n_75), .A2(n_81), .ZN(n_71));
   NAND2_X1 i_96 (.A1(n_76), .A2(n_585), .ZN(n_75));
   NAND2_X1 i_97 (.A1(n_80), .A2(n_78), .ZN(n_76));
   OAI21_X1 i_102 (.A(n_120), .B1(n_79), .B2(n_118), .ZN(n_78));
   INV_X1 i_103 (.A(n_588), .ZN(n_79));
   INV_X1 i_113 (.A(n_622), .ZN(n_80));
   INV_X1 i_114 (.A(n_82), .ZN(n_81));
   NAND2_X1 i_115 (.A1(n_499), .A2(n_497), .ZN(n_82));
   NAND2_X1 i_116 (.A1(n_84), .A2(n_227), .ZN(n_83));
   NAND2_X1 i_117 (.A1(n_89), .A2(n_670), .ZN(n_84));
   NAND2_X1 i_118 (.A1(n_90), .A2(n_100), .ZN(n_89));
   NAND2_X1 i_119 (.A1(n_282), .A2(n_313), .ZN(n_90));
   INV_X1 i_120 (.A(n_281), .ZN(n_100));
   NAND2_X1 i_124 (.A1(n_102), .A2(n_103), .ZN(n_101));
   NAND2_X1 i_125 (.A1(n_106), .A2(n_107), .ZN(n_102));
   NAND2_X1 i_126 (.A1(n_112), .A2(n_111), .ZN(n_106));
   NAND2_X1 i_127 (.A1(n_109), .A2(n_409), .ZN(n_107));
   NAND4_X1 i_128 (.A1(n_112), .A2(n_109), .A3(n_111), .A4(n_409), .ZN(n_103));
   NAND2_X1 i_129 (.A1(n_408), .A2(n_405), .ZN(n_109));
   NAND4_X1 i_130 (.A1(n_423), .A2(n_421), .A3(n_411), .A4(n_412), .ZN(n_408));
   NAND2_X1 i_131 (.A1(n_581), .A2(n_413), .ZN(n_412));
   NAND3_X1 i_132 (.A1(n_414), .A2(n_415), .A3(n_582), .ZN(n_411));
   NAND3_X1 i_133 (.A1(n_110), .A2(n_567), .A3(n_564), .ZN(n_423));
   NAND2_X1 i_134 (.A1(n_573), .A2(n_548), .ZN(n_110));
   NAND3_X1 i_135 (.A1(n_549), .A2(n_573), .A3(n_548), .ZN(n_421));
   NAND2_X1 i_136 (.A1(n_263), .A2(n_406), .ZN(n_405));
   NAND2_X1 i_137 (.A1(n_420), .A2(n_410), .ZN(n_409));
   NAND3_X1 i_138 (.A1(n_562), .A2(n_550), .A3(n_546), .ZN(n_111));
   NAND2_X1 i_139 (.A1(n_113), .A2(n_114), .ZN(n_112));
   NAND2_X1 i_140 (.A1(n_562), .A2(n_546), .ZN(n_113));
   INV_X1 i_141 (.A(n_550), .ZN(n_114));
   INV_X1 i_142 (.A(n_105), .ZN(n_104));
   NAND2_X1 i_143 (.A1(n_117), .A2(n_119), .ZN(n_105));
   OAI21_X1 i_144 (.A(n_588), .B1(n_118), .B2(n_613), .ZN(n_117));
   INV_X1 i_145 (.A(n_587), .ZN(n_118));
   NAND4_X1 i_146 (.A1(n_120), .A2(n_595), .A3(n_589), .A4(n_587), .ZN(n_119));
   NAND2_X1 i_147 (.A1(n_122), .A2(n_121), .ZN(n_120));
   NAND2_X1 i_148 (.A1(n_614), .A2(n_616), .ZN(n_121));
   NAND2_X1 i_149 (.A1(n_619), .A2(n_617), .ZN(n_122));
   OAI21_X1 i_151 (.A(n_115), .B1(n_232), .B2(n_231), .ZN(n_108));
   OAI21_X1 i_152 (.A(n_169), .B1(n_130), .B2(n_126), .ZN(n_125));
   INV_X1 i_121 (.A(n_127), .ZN(n_126));
   OAI21_X1 i_122 (.A(n_171), .B1(n_128), .B2(n_129), .ZN(n_127));
   INV_X1 i_123 (.A(n_227), .ZN(n_128));
   AOI21_X1 i_150 (.A(n_392), .B1(n_276), .B2(n_230), .ZN(n_129));
   AOI21_X1 i_153 (.A(n_160), .B1(n_134), .B2(n_131), .ZN(n_130));
   NAND2_X1 i_158 (.A1(n_132), .A2(n_133), .ZN(n_131));
   NAND2_X1 i_159 (.A1(n_165), .A2(n_171), .ZN(n_132));
   NAND2_X1 i_160 (.A1(n_163), .A2(n_162), .ZN(n_133));
   NAND2_X1 i_161 (.A1(n_135), .A2(n_373), .ZN(n_134));
   NAND2_X1 i_162 (.A1(n_371), .A2(n_136), .ZN(n_135));
   NAND2_X1 i_163 (.A1(n_137), .A2(n_362), .ZN(n_136));
   NAND2_X1 i_164 (.A1(n_359), .A2(n_316), .ZN(n_137));
   NAND2_X1 i_165 (.A1(n_368), .A2(n_360), .ZN(n_359));
   NAND2_X1 i_166 (.A1(n_207), .A2(n_147), .ZN(n_368));
   NAND2_X1 i_167 (.A1(n_317), .A2(n_349), .ZN(n_316));
   NAND3_X1 i_168 (.A1(n_521), .A2(n_350), .A3(n_356), .ZN(n_349));
   OAI211_X1 i_183 (.A(n_338), .B(n_346), .C1(n_138), .C2(n_146), .ZN(n_317));
   NAND2_X1 i_170 (.A1(n_348), .A2(n_347), .ZN(n_346));
   NAND3_X1 i_171 (.A1(n_344), .A2(n_343), .A3(n_339), .ZN(n_338));
   AOI21_X1 i_172 (.A(n_142), .B1(n_321), .B2(n_139), .ZN(n_138));
   NAND3_X1 i_173 (.A1(n_523), .A2(n_334), .A3(n_143), .ZN(n_139));
   OAI21_X1 i_174 (.A(n_325), .B1(n_324), .B2(n_322), .ZN(n_321));
   AOI21_X1 i_175 (.A(n_140), .B1(n_226), .B2(n_141), .ZN(n_324));
   NAND3_X1 i_176 (.A1(n_226), .A2(n_141), .A3(n_140), .ZN(n_325));
   NAND2_X1 i_177 (.A1(T_Count[1]), .A2(n_657), .ZN(n_140));
   NAND3_X1 i_178 (.A1(X_Count[1]), .A2(T_Count[0]), .A3(num_of_X[1]), .ZN(n_141));
   INV_X1 i_179 (.A(n_323), .ZN(n_322));
   AOI21_X1 i_180 (.A(n_143), .B1(n_523), .B2(n_334), .ZN(n_142));
   NAND2_X1 i_181 (.A1(n_331), .A2(n_144), .ZN(n_143));
   INV_X1 i_182 (.A(n_332), .ZN(n_144));
   INV_X1 i_184 (.A(n_336), .ZN(n_146));
   OAI21_X1 i_185 (.A(n_337), .B1(n_341), .B2(n_340), .ZN(n_336));
   NAND3_X1 i_186 (.A1(n_207), .A2(n_147), .A3(n_363), .ZN(n_362));
   NAND2_X1 i_187 (.A1(n_365), .A2(n_364), .ZN(n_363));
   NAND2_X1 i_188 (.A1(n_210), .A2(n_521), .ZN(n_147));
   NAND3_X1 i_189 (.A1(n_151), .A2(n_148), .A3(n_150), .ZN(n_371));
   INV_X1 i_190 (.A(n_159), .ZN(n_148));
   NAND2_X1 i_191 (.A1(n_149), .A2(n_159), .ZN(n_373));
   NAND2_X1 i_193 (.A1(n_151), .A2(n_150), .ZN(n_149));
   NAND3_X1 i_194 (.A1(n_173), .A2(n_207), .A3(n_153), .ZN(n_150));
   NAND2_X1 i_195 (.A1(n_152), .A2(n_158), .ZN(n_151));
   OAI21_X1 i_196 (.A(n_153), .B1(n_196), .B2(n_156), .ZN(n_152));
   NAND2_X1 i_198 (.A1(n_154), .A2(n_177), .ZN(n_153));
   INV_X1 i_204 (.A(n_155), .ZN(n_154));
   NAND3_X1 i_205 (.A1(n_314), .A2(n_199), .A3(n_580), .ZN(n_155));
   AOI21_X1 i_206 (.A(n_157), .B1(n_552), .B2(n_577), .ZN(n_156));
   INV_X1 i_207 (.A(n_580), .ZN(n_157));
   NOR2_X1 i_208 (.A1(n_521), .A2(n_210), .ZN(n_158));
   XNOR2_X1 i_209 (.A(n_272), .B(n_383), .ZN(n_159));
   INV_X1 i_210 (.A(n_161), .ZN(n_160));
   NAND4_X1 i_211 (.A1(n_165), .A2(n_171), .A3(n_163), .A4(n_162), .ZN(n_161));
   NAND3_X1 i_212 (.A1(n_256), .A2(n_254), .A3(n_124), .ZN(n_162));
   OAI21_X1 i_220 (.A(n_314), .B1(n_164), .B2(n_231), .ZN(n_163));
   INV_X1 i_221 (.A(n_124), .ZN(n_164));
   OAI21_X1 i_222 (.A(n_166), .B1(n_168), .B2(n_167), .ZN(n_165));
   XNOR2_X1 i_223 (.A(n_623), .B(n_396), .ZN(n_166));
   INV_X1 i_224 (.A(n_173), .ZN(n_167));
   INV_X1 i_225 (.A(n_175), .ZN(n_168));
   OAI211_X1 i_226 (.A(n_227), .B(n_170), .C1(n_228), .C2(n_392), .ZN(n_169));
   INV_X1 i_227 (.A(n_171), .ZN(n_170));
   NAND3_X1 i_154 (.A1(n_175), .A2(n_173), .A3(n_172), .ZN(n_171));
   XNOR2_X1 i_229 (.A(n_646), .B(n_623), .ZN(n_172));
   NAND2_X1 i_230 (.A1(n_174), .A2(n_198), .ZN(n_173));
   NAND2_X1 i_231 (.A1(n_177), .A2(n_580), .ZN(n_174));
   NAND2_X1 i_232 (.A1(n_176), .A2(n_207), .ZN(n_175));
   NAND3_X1 i_233 (.A1(n_177), .A2(n_196), .A3(n_580), .ZN(n_176));
   NAND2_X1 i_234 (.A1(n_552), .A2(n_577), .ZN(n_177));
   NAND2_X1 i_235 (.A1(n_553), .A2(n_557), .ZN(n_552));
   NAND3_X1 i_236 (.A1(n_180), .A2(n_671), .A3(n_284), .ZN(n_557));
   INV_X1 i_237 (.A(n_273), .ZN(n_180));
   OAI21_X1 i_238 (.A(n_675), .B1(n_181), .B2(n_273), .ZN(n_553));
   INV_X1 i_239 (.A(n_284), .ZN(n_181));
   NAND2_X1 i_240 (.A1(n_183), .A2(n_182), .ZN(n_577));
   NAND2_X1 i_241 (.A1(n_185), .A2(n_195), .ZN(n_182));
   NAND2_X1 i_242 (.A1(n_192), .A2(n_194), .ZN(n_183));
   NAND4_X1 i_243 (.A1(n_192), .A2(n_185), .A3(n_195), .A4(n_194), .ZN(n_580));
   NAND3_X1 i_244 (.A1(n_191), .A2(T_Count[1]), .A3(num_of_X[4]), .ZN(n_185));
   NAND2_X1 i_245 (.A1(n_389), .A2(n_388), .ZN(n_191));
   NAND2_X1 i_246 (.A1(n_193), .A2(n_310), .ZN(n_192));
   NAND2_X1 i_247 (.A1(n_307), .A2(n_312), .ZN(n_193));
   NAND3_X1 i_248 (.A1(n_307), .A2(n_312), .A3(n_311), .ZN(n_194));
   NAND3_X1 i_249 (.A1(n_389), .A2(n_388), .A3(n_387), .ZN(n_195));
   INV_X1 i_250 (.A(n_198), .ZN(n_196));
   NAND2_X1 i_251 (.A1(n_314), .A2(n_199), .ZN(n_198));
   NAND4_X1 i_252 (.A1(n_376), .A2(n_379), .A3(n_361), .A4(n_326), .ZN(n_199));
   NAND2_X1 i_253 (.A1(n_208), .A2(n_215), .ZN(n_207));
   INV_X1 i_254 (.A(n_210), .ZN(n_208));
   OAI21_X1 i_255 (.A(n_512), .B1(n_506), .B2(n_511), .ZN(n_210));
   AOI21_X1 i_256 (.A(n_214), .B1(n_514), .B2(n_513), .ZN(n_511));
   NAND2_X1 i_257 (.A1(n_508), .A2(n_507), .ZN(n_506));
   NAND3_X1 i_258 (.A1(n_287), .A2(n_291), .A3(n_290), .ZN(n_507));
   NAND2_X1 i_259 (.A1(n_211), .A2(n_212), .ZN(n_508));
   NAND2_X1 i_260 (.A1(n_287), .A2(n_290), .ZN(n_211));
   INV_X1 i_261 (.A(n_291), .ZN(n_212));
   NAND3_X1 i_262 (.A1(n_513), .A2(n_214), .A3(n_514), .ZN(n_512));
   OR2_X1 i_263 (.A1(n_280), .A2(n_538), .ZN(n_513));
   NAND2_X1 i_264 (.A1(n_517), .A2(n_515), .ZN(n_514));
   INV_X1 i_265 (.A(n_516), .ZN(n_515));
   NAND2_X1 i_266 (.A1(T_Count[3]), .A2(num_of_X[0]), .ZN(n_516));
   OAI21_X1 i_267 (.A(n_213), .B1(n_491), .B2(n_584), .ZN(n_517));
   NAND2_X1 i_268 (.A1(T_Count[2]), .A2(num_of_X[1]), .ZN(n_213));
   INV_X1 i_269 (.A(T_Count[1]), .ZN(n_491));
   INV_X1 i_270 (.A(n_532), .ZN(n_214));
   INV_X1 i_271 (.A(n_521), .ZN(n_215));
   NAND3_X1 i_272 (.A1(n_542), .A2(n_522), .A3(n_528), .ZN(n_521));
   NAND2_X1 i_273 (.A1(n_217), .A2(n_216), .ZN(n_542));
   NAND3_X1 i_274 (.A1(n_278), .A2(n_235), .A3(n_236), .ZN(n_216));
   NAND3_X1 i_275 (.A1(n_218), .A2(T_Count[4]), .A3(num_of_X[0]), .ZN(n_217));
   NAND2_X1 i_276 (.A1(n_235), .A2(n_278), .ZN(n_218));
   NAND3_X1 i_277 (.A1(n_219), .A2(n_532), .A3(n_223), .ZN(n_528));
   NAND2_X1 i_278 (.A1(n_539), .A2(n_220), .ZN(n_219));
   NAND2_X1 i_280 (.A1(n_527), .A2(n_523), .ZN(n_522));
   NAND3_X1 i_281 (.A1(n_222), .A2(n_220), .A3(n_539), .ZN(n_527));
   NAND2_X1 i_282 (.A1(n_537), .A2(n_538), .ZN(n_220));
   NAND2_X1 i_283 (.A1(T_Count[1]), .A2(num_of_X[1]), .ZN(n_538));
   NAND3_X1 i_284 (.A1(X_Count[2]), .A2(T_Count[0]), .A3(num_of_X[2]), .ZN(n_537));
   OAI21_X1 i_285 (.A(n_221), .B1(n_665), .B2(n_584), .ZN(n_539));
   INV_X1 i_286 (.A(X_Count[2]), .ZN(n_221));
   NAND2_X1 i_287 (.A1(n_532), .A2(n_223), .ZN(n_222));
   NAND3_X1 i_288 (.A1(X_Count[3]), .A2(T_Count[0]), .A3(num_of_X[3]), .ZN(n_223));
   NAND2_X1 i_289 (.A1(n_224), .A2(n_225), .ZN(n_532));
   NAND2_X1 i_290 (.A1(T_Count[0]), .A2(num_of_X[3]), .ZN(n_224));
   INV_X1 i_291 (.A(X_Count[3]), .ZN(n_225));
   NAND3_X1 i_292 (.A1(n_226), .A2(T_Count[2]), .A3(num_of_X[0]), .ZN(n_523));
   NAND2_X1 i_293 (.A1(n_525), .A2(n_526), .ZN(n_226));
   NAND2_X1 i_294 (.A1(T_Count[0]), .A2(num_of_X[1]), .ZN(n_525));
   INV_X1 i_295 (.A(X_Count[1]), .ZN(n_526));
   NAND3_X1 i_155 (.A1(n_230), .A2(n_276), .A3(n_392), .ZN(n_227));
   INV_X1 i_297 (.A(n_229), .ZN(n_228));
   NAND2_X1 i_298 (.A1(n_230), .A2(n_276), .ZN(n_229));
   OAI211_X1 i_156 (.A(n_116), .B(n_115), .C1(n_232), .C2(n_231), .ZN(n_230));
   NOR2_X1 i_157 (.A1(n_258), .A2(n_271), .ZN(n_231));
   AOI21_X1 i_169 (.A(n_314), .B1(n_258), .B2(n_271), .ZN(n_232));
   NAND4_X1 i_228 (.A1(n_239), .A2(n_244), .A3(n_238), .A4(n_625), .ZN(n_115));
   NAND2_X1 i_296 (.A1(n_237), .A2(n_241), .ZN(n_116));
   NAND2_X1 i_306 (.A1(n_239), .A2(n_238), .ZN(n_237));
   NAND4_X1 i_307 (.A1(n_595), .A2(n_594), .A3(n_592), .A4(n_591), .ZN(n_238));
   NAND2_X1 i_308 (.A1(n_240), .A2(n_590), .ZN(n_239));
   NAND2_X1 i_309 (.A1(n_594), .A2(n_595), .ZN(n_240));
   NAND2_X1 i_310 (.A1(n_244), .A2(n_625), .ZN(n_241));
   NAND2_X1 i_311 (.A1(n_243), .A2(n_242), .ZN(n_625));
   NAND2_X1 i_312 (.A1(n_247), .A2(n_249), .ZN(n_242));
   NAND2_X1 i_313 (.A1(n_245), .A2(n_250), .ZN(n_243));
   NAND2_X1 i_314 (.A1(n_624), .A2(n_646), .ZN(n_244));
   NAND4_X1 i_315 (.A1(n_245), .A2(n_247), .A3(n_250), .A4(n_249), .ZN(n_624));
   NAND2_X1 i_316 (.A1(n_246), .A2(n_608), .ZN(n_245));
   NAND2_X1 i_317 (.A1(n_610), .A2(n_607), .ZN(n_246));
   NAND3_X1 i_318 (.A1(n_248), .A2(T_Count[1]), .A3(num_of_X[6]), .ZN(n_247));
   NAND2_X1 i_319 (.A1(n_567), .A2(n_566), .ZN(n_248));
   NAND3_X1 i_320 (.A1(n_567), .A2(n_566), .A3(n_565), .ZN(n_249));
   NAND3_X1 i_321 (.A1(n_610), .A2(n_609), .A3(n_607), .ZN(n_250));
   OAI21_X1 i_322 (.A(n_251), .B1(n_252), .B2(n_602), .ZN(n_646));
   NAND3_X1 i_323 (.A1(n_603), .A2(n_602), .A3(n_598), .ZN(n_251));
   INV_X1 i_324 (.A(n_253), .ZN(n_252));
   NAND2_X1 i_325 (.A1(n_603), .A2(n_598), .ZN(n_253));
   INV_X1 i_327 (.A(n_271), .ZN(n_123));
   NAND2_X1 i_329 (.A1(n_271), .A2(n_258), .ZN(n_124));
   NAND2_X1 i_299 (.A1(n_145), .A2(n_233), .ZN(n_258));
   NAND2_X1 i_331 (.A1(n_260), .A2(n_261), .ZN(n_145));
   NAND2_X1 i_332 (.A1(n_263), .A2(n_464), .ZN(n_260));
   INV_X1 i_333 (.A(n_460), .ZN(n_261));
   NAND3_X1 i_334 (.A1(n_263), .A2(n_460), .A3(n_464), .ZN(n_233));
   NAND2_X1 i_335 (.A1(n_264), .A2(n_265), .ZN(n_263));
   NAND2_X1 i_337 (.A1(n_267), .A2(n_372), .ZN(n_264));
   INV_X1 i_338 (.A(n_268), .ZN(n_265));
   NAND3_X1 i_339 (.A1(n_268), .A2(n_372), .A3(n_267), .ZN(n_464));
   NAND2_X1 i_340 (.A1(n_367), .A2(n_328), .ZN(n_267));
   NAND2_X1 i_341 (.A1(n_269), .A2(n_301), .ZN(n_268));
   NAND2_X1 i_342 (.A1(n_300), .A2(n_299), .ZN(n_269));
   NAND2_X1 i_346 (.A1(n_270), .A2(n_385), .ZN(n_460));
   NAND3_X1 i_349 (.A1(n_386), .A2(n_389), .A3(n_381), .ZN(n_270));
   AOI22_X1 i_300 (.A1(n_272), .A2(n_448), .B1(n_304), .B2(n_292), .ZN(n_271));
   NAND4_X1 i_301 (.A1(n_293), .A2(n_312), .A3(n_305), .A4(n_297), .ZN(n_448));
   OAI21_X1 i_304 (.A(n_284), .B1(n_675), .B2(n_273), .ZN(n_272));
   AOI21_X1 i_305 (.A(n_285), .B1(n_289), .B2(n_287), .ZN(n_273));
   INV_X1 i_376 (.A(n_278), .ZN(n_234));
   NAND2_X1 i_380 (.A1(n_280), .A2(n_279), .ZN(n_278));
   NAND2_X1 i_381 (.A1(T_Count[3]), .A2(num_of_X[1]), .ZN(n_279));
   NAND2_X1 i_382 (.A1(T_Count[2]), .A2(num_of_X[2]), .ZN(n_280));
   NAND4_X1 i_383 (.A1(T_Count[3]), .A2(T_Count[2]), .A3(num_of_X[2]), .A4(
      num_of_X[1]), .ZN(n_235));
   NAND2_X1 i_384 (.A1(T_Count[4]), .A2(num_of_X[0]), .ZN(n_236));
   NAND3_X1 i_359 (.A1(n_289), .A2(n_287), .A3(n_285), .ZN(n_284));
   INV_X1 i_386 (.A(n_286), .ZN(n_285));
   NAND2_X1 i_387 (.A1(T_Count[5]), .A2(num_of_X[0]), .ZN(n_286));
   OAI21_X1 i_388 (.A(n_288), .B1(n_665), .B2(n_431), .ZN(n_287));
   INV_X1 i_389 (.A(X_Count[4]), .ZN(n_288));
   NAND2_X1 i_390 (.A1(n_290), .A2(n_291), .ZN(n_289));
   NAND3_X1 i_391 (.A1(X_Count[4]), .A2(T_Count[0]), .A3(num_of_X[4]), .ZN(n_290));
   NAND2_X1 i_392 (.A1(T_Count[1]), .A2(num_of_X[3]), .ZN(n_291));
   NAND2_X1 i_362 (.A1(n_293), .A2(n_297), .ZN(n_292));
   NAND2_X1 i_394 (.A1(n_294), .A2(n_295), .ZN(n_293));
   NAND2_X1 i_395 (.A1(n_301), .A2(n_300), .ZN(n_294));
   INV_X1 i_397 (.A(n_299), .ZN(n_295));
   NAND3_X1 i_398 (.A1(n_301), .A2(n_300), .A3(n_299), .ZN(n_297));
   NAND2_X1 i_399 (.A1(T_Count[1]), .A2(num_of_X[5]), .ZN(n_299));
   NAND3_X1 i_400 (.A1(X_Count[6]), .A2(T_Count[0]), .A3(num_of_X[6]), .ZN(n_300));
   NAND2_X1 i_401 (.A1(n_302), .A2(n_303), .ZN(n_301));
   NAND2_X1 i_402 (.A1(T_Count[0]), .A2(num_of_X[6]), .ZN(n_302));
   INV_X1 i_403 (.A(X_Count[6]), .ZN(n_303));
   NAND2_X1 i_372 (.A1(n_305), .A2(n_312), .ZN(n_304));
   NAND2_X1 i_405 (.A1(n_307), .A2(n_310), .ZN(n_305));
   OAI21_X1 i_406 (.A(n_308), .B1(n_309), .B2(n_584), .ZN(n_307));
   NAND2_X1 i_407 (.A1(T_Count[2]), .A2(num_of_X[3]), .ZN(n_308));
   INV_X1 i_408 (.A(T_Count[3]), .ZN(n_309));
   INV_X1 i_410 (.A(n_311), .ZN(n_310));
   NAND2_X1 i_411 (.A1(T_Count[4]), .A2(num_of_X[1]), .ZN(n_311));
   NAND4_X1 i_412 (.A1(T_Count[3]), .A2(T_Count[2]), .A3(num_of_X[3]), .A4(
      num_of_X[2]), .ZN(n_312));
   INV_X1 i_413 (.A(n_314), .ZN(n_254));
   NAND2_X1 i_414 (.A1(n_375), .A2(n_320), .ZN(n_314));
   NAND2_X1 i_415 (.A1(n_326), .A2(n_361), .ZN(n_320));
   NAND2_X1 i_418 (.A1(n_327), .A2(n_328), .ZN(n_326));
   NAND2_X1 i_421 (.A1(n_372), .A2(n_367), .ZN(n_327));
   INV_X1 i_422 (.A(n_374), .ZN(n_328));
   NAND3_X1 i_424 (.A1(n_367), .A2(n_372), .A3(n_374), .ZN(n_361));
   NAND2_X1 i_425 (.A1(n_370), .A2(n_369), .ZN(n_367));
   NAND2_X1 i_427 (.A1(T_Count[3]), .A2(num_of_X[3]), .ZN(n_369));
   NAND2_X1 i_428 (.A1(T_Count[2]), .A2(num_of_X[4]), .ZN(n_370));
   NAND4_X1 i_429 (.A1(T_Count[3]), .A2(T_Count[2]), .A3(num_of_X[4]), .A4(
      num_of_X[3]), .ZN(n_372));
   NAND2_X1 i_430 (.A1(T_Count[5]), .A2(num_of_X[1]), .ZN(n_374));
   NAND2_X1 i_431 (.A1(n_379), .A2(n_376), .ZN(n_375));
   NAND2_X1 i_432 (.A1(n_377), .A2(n_378), .ZN(n_376));
   INV_X1 i_434 (.A(n_380), .ZN(n_377));
   NAND2_X1 i_435 (.A1(n_386), .A2(n_389), .ZN(n_378));
   NAND3_X1 i_436 (.A1(n_380), .A2(n_389), .A3(n_386), .ZN(n_379));
   NAND2_X1 i_437 (.A1(n_385), .A2(n_381), .ZN(n_380));
   NAND2_X1 i_438 (.A1(n_384), .A2(n_382), .ZN(n_381));
   NAND2_X1 i_439 (.A1(T_Count[6]), .A2(num_of_X[0]), .ZN(n_382));
   NAND2_X1 i_440 (.A1(T_Count[4]), .A2(num_of_X[2]), .ZN(n_384));
   NAND4_X1 i_441 (.A1(T_Count[6]), .A2(T_Count[4]), .A3(num_of_X[2]), .A4(
      num_of_X[0]), .ZN(n_385));
   NAND2_X1 i_442 (.A1(n_388), .A2(n_387), .ZN(n_386));
   NAND2_X1 i_443 (.A1(T_Count[1]), .A2(num_of_X[4]), .ZN(n_387));
   NAND3_X1 i_444 (.A1(X_Count[5]), .A2(T_Count[0]), .A3(num_of_X[5]), .ZN(n_388));
   NAND2_X1 i_445 (.A1(n_390), .A2(n_391), .ZN(n_389));
   NAND2_X1 i_446 (.A1(T_Count[0]), .A2(num_of_X[5]), .ZN(n_390));
   INV_X1 i_447 (.A(X_Count[5]), .ZN(n_391));
   NAND2_X1 i_374 (.A1(n_404), .A2(n_403), .ZN(n_392));
   NAND2_X1 i_449 (.A1(n_394), .A2(n_398), .ZN(n_393));
   OAI21_X1 i_450 (.A(n_395), .B1(n_397), .B2(n_440), .ZN(n_394));
   INV_X1 i_451 (.A(n_399), .ZN(n_395));
   INV_X1 i_452 (.A(n_438), .ZN(n_397));
   NAND3_X1 i_453 (.A1(n_439), .A2(n_438), .A3(n_399), .ZN(n_398));
   NAND2_X1 i_454 (.A1(n_401), .A2(n_400), .ZN(n_399));
   NAND3_X1 i_455 (.A1(n_416), .A2(n_426), .A3(n_419), .ZN(n_400));
   NAND2_X1 i_456 (.A1(n_402), .A2(n_425), .ZN(n_401));
   NAND2_X1 i_457 (.A1(n_416), .A2(n_419), .ZN(n_402));
   NAND3_X1 i_458 (.A1(n_418), .A2(n_58), .A3(n_467), .ZN(n_416));
   NAND2_X1 i_459 (.A1(n_424), .A2(n_452), .ZN(n_418));
   NAND3_X1 i_460 (.A1(n_424), .A2(n_452), .A3(n_422), .ZN(n_419));
   NAND2_X1 i_461 (.A1(n_467), .A2(n_58), .ZN(n_422));
   NAND2_X1 i_462 (.A1(n_455), .A2(n_472), .ZN(n_424));
   INV_X1 i_463 (.A(n_426), .ZN(n_425));
   NAND2_X1 i_464 (.A1(n_429), .A2(n_427), .ZN(n_426));
   NAND3_X1 i_465 (.A1(n_432), .A2(n_428), .A3(n_434), .ZN(n_427));
   INV_X1 i_466 (.A(n_437), .ZN(n_428));
   NAND2_X1 i_467 (.A1(n_430), .A2(n_437), .ZN(n_429));
   NAND2_X1 i_468 (.A1(n_432), .A2(n_434), .ZN(n_430));
   NAND2_X1 i_469 (.A1(n_433), .A2(n_72), .ZN(n_432));
   NAND2_X1 i_470 (.A1(n_435), .A2(n_479), .ZN(n_433));
   NAND3_X1 i_471 (.A1(n_435), .A2(n_436), .A3(n_479), .ZN(n_434));
   NAND2_X1 i_472 (.A1(n_493), .A2(n_476), .ZN(n_435));
   INV_X1 i_473 (.A(n_72), .ZN(n_436));
   AOI21_X1 i_474 (.A(n_77), .B1(n_484), .B2(n_489), .ZN(n_437));
   NAND3_X1 i_475 (.A1(n_441), .A2(n_666), .A3(n_443), .ZN(n_438));
   INV_X1 i_476 (.A(n_440), .ZN(n_439));
   AOI21_X1 i_477 (.A(n_666), .B1(n_441), .B2(n_443), .ZN(n_440));
   NAND2_X1 i_478 (.A1(n_442), .A2(n_445), .ZN(n_441));
   NAND3_X1 i_479 (.A1(n_494), .A2(n_446), .A3(n_451), .ZN(n_442));
   NAND4_X1 i_480 (.A1(n_494), .A2(n_446), .A3(n_451), .A4(n_444), .ZN(n_443));
   INV_X1 i_481 (.A(n_445), .ZN(n_444));
   XNOR2_X1 i_482 (.A(n_85), .B(n_88), .ZN(n_445));
   NAND2_X1 i_483 (.A1(n_447), .A2(n_450), .ZN(n_446));
   NAND2_X1 i_484 (.A1(n_452), .A2(n_455), .ZN(n_447));
   INV_X1 i_485 (.A(n_472), .ZN(n_450));
   NAND3_X1 i_486 (.A1(n_452), .A2(n_455), .A3(n_472), .ZN(n_451));
   NAND3_X1 i_487 (.A1(n_453), .A2(n_454), .A3(n_458), .ZN(n_452));
   NAND2_X1 i_488 (.A1(n_456), .A2(n_502), .ZN(n_453));
   INV_X1 i_489 (.A(n_459), .ZN(n_454));
   OAI211_X1 i_490 (.A(n_502), .B(n_456), .C1(n_457), .C2(n_459), .ZN(n_455));
   NAND3_X1 i_491 (.A1(n_545), .A2(n_501), .A3(n_562), .ZN(n_456));
   INV_X1 i_492 (.A(n_458), .ZN(n_457));
   NAND3_X1 i_493 (.A1(n_209), .A2(n_467), .A3(n_197), .ZN(n_458));
   AOI21_X1 i_494 (.A(n_197), .B1(n_467), .B2(n_209), .ZN(n_459));
   NAND2_X1 i_495 (.A1(n_461), .A2(n_462), .ZN(n_197));
   OAI21_X1 i_496 (.A(n_205), .B1(n_200), .B2(n_202), .ZN(n_461));
   NAND3_X1 i_497 (.A1(n_203), .A2(n_206), .A3(n_201), .ZN(n_462));
   OAI21_X1 i_498 (.A(n_465), .B1(n_463), .B2(n_466), .ZN(n_209));
   AOI21_X1 i_499 (.A(n_470), .B1(n_544), .B2(n_559), .ZN(n_463));
   INV_X1 i_500 (.A(n_468), .ZN(n_465));
   INV_X1 i_501 (.A(n_536), .ZN(n_466));
   OAI211_X1 i_502 (.A(n_468), .B(n_536), .C1(n_471), .C2(n_470), .ZN(n_467));
   NAND2_X1 i_503 (.A1(n_469), .A2(n_519), .ZN(n_468));
   NAND2_X1 i_504 (.A1(n_510), .A2(n_520), .ZN(n_469));
   INV_X1 i_505 (.A(n_535), .ZN(n_470));
   INV_X1 i_506 (.A(n_543), .ZN(n_471));
   NAND2_X1 i_507 (.A1(n_474), .A2(n_473), .ZN(n_472));
   NAND3_X1 i_508 (.A1(n_493), .A2(n_479), .A3(n_476), .ZN(n_473));
   NAND2_X1 i_509 (.A1(n_492), .A2(n_475), .ZN(n_474));
   NAND2_X1 i_510 (.A1(n_476), .A2(n_479), .ZN(n_475));
   NAND2_X1 i_511 (.A1(n_477), .A2(n_478), .ZN(n_476));
   NAND2_X1 i_512 (.A1(n_482), .A2(n_486), .ZN(n_477));
   NAND2_X1 i_513 (.A1(n_481), .A2(n_480), .ZN(n_478));
   NAND4_X1 i_514 (.A1(n_482), .A2(n_486), .A3(n_481), .A4(n_480), .ZN(n_479));
   NAND3_X1 i_515 (.A1(n_255), .A2(num_of_X[8]), .A3(n_186), .ZN(n_480));
   NAND3_X1 i_516 (.A1(n_187), .A2(n_184), .A3(n_190), .ZN(n_481));
   NAND2_X1 i_517 (.A1(n_483), .A2(n_484), .ZN(n_482));
   INV_X1 i_518 (.A(n_487), .ZN(n_483));
   OAI21_X1 i_519 (.A(n_663), .B1(n_485), .B2(n_659), .ZN(n_484));
   INV_X1 i_520 (.A(n_662), .ZN(n_485));
   NAND3_X1 i_521 (.A1(n_487), .A2(n_490), .A3(n_663), .ZN(n_486));
   NAND2_X1 i_522 (.A1(n_489), .A2(n_178), .ZN(n_487));
   OAI21_X1 i_523 (.A(n_179), .B1(n_575), .B2(n_488), .ZN(n_178));
   INV_X1 i_524 (.A(num_of_X[7]), .ZN(n_488));
   NAND3_X1 i_525 (.A1(n_641), .A2(num_of_X[7]), .A3(num_of_X[6]), .ZN(n_489));
   NAND2_X1 i_526 (.A1(n_662), .A2(n_661), .ZN(n_490));
   INV_X1 i_527 (.A(n_493), .ZN(n_492));
   OAI21_X1 i_528 (.A(n_631), .B1(n_629), .B2(n_655), .ZN(n_493));
   INV_X1 i_529 (.A(n_495), .ZN(n_494));
   NAND2_X1 i_530 (.A1(n_496), .A2(n_585), .ZN(n_495));
   OAI211_X1 i_531 (.A(n_497), .B(n_499), .C1(n_622), .C2(n_586), .ZN(n_496));
   NAND3_X1 i_532 (.A1(n_498), .A2(n_502), .A3(n_501), .ZN(n_497));
   NAND2_X1 i_533 (.A1(n_545), .A2(n_562), .ZN(n_498));
   NAND3_X1 i_534 (.A1(n_500), .A2(n_562), .A3(n_545), .ZN(n_499));
   NAND2_X1 i_535 (.A1(n_502), .A2(n_501), .ZN(n_500));
   NAND4_X1 i_536 (.A1(n_531), .A2(n_530), .A3(n_505), .A4(n_504), .ZN(n_501));
   NAND2_X1 i_537 (.A1(n_529), .A2(n_503), .ZN(n_502));
   NAND2_X1 i_538 (.A1(n_505), .A2(n_504), .ZN(n_503));
   NAND3_X1 i_539 (.A1(n_510), .A2(n_524), .A3(n_519), .ZN(n_504));
   NAND2_X1 i_540 (.A1(n_509), .A2(n_520), .ZN(n_505));
   NAND2_X1 i_541 (.A1(n_510), .A2(n_519), .ZN(n_509));
   OAI21_X1 i_542 (.A(n_518), .B1(n_417), .B2(n_431), .ZN(n_510));
   NAND2_X1 i_543 (.A1(T_Count[7]), .A2(num_of_X[3]), .ZN(n_518));
   NAND4_X1 i_544 (.A1(T_Count[7]), .A2(T_Count[6]), .A3(num_of_X[4]), .A4(
      num_of_X[3]), .ZN(n_519));
   INV_X1 i_545 (.A(n_524), .ZN(n_520));
   NAND2_X1 i_546 (.A1(T_Count[3]), .A2(num_of_X[7]), .ZN(n_524));
   NAND2_X1 i_547 (.A1(n_531), .A2(n_530), .ZN(n_529));
   NAND3_X1 i_548 (.A1(n_534), .A2(n_559), .A3(n_544), .ZN(n_530));
   NAND2_X1 i_549 (.A1(n_543), .A2(n_533), .ZN(n_531));
   INV_X1 i_550 (.A(n_534), .ZN(n_533));
   NAND2_X1 i_551 (.A1(n_536), .A2(n_535), .ZN(n_534));
   NAND4_X1 i_552 (.A1(T_Count[5]), .A2(T_Count[4]), .A3(num_of_X[6]), .A4(
      num_of_X[5]), .ZN(n_535));
   OAI21_X1 i_553 (.A(n_540), .B1(n_575), .B2(n_541), .ZN(n_536));
   NAND2_X1 i_554 (.A1(T_Count[5]), .A2(num_of_X[5]), .ZN(n_540));
   INV_X1 i_555 (.A(num_of_X[6]), .ZN(n_541));
   NAND2_X1 i_556 (.A1(n_544), .A2(n_559), .ZN(n_543));
   NAND2_X1 i_557 (.A1(n_556), .A2(n_558), .ZN(n_544));
   NAND2_X1 i_558 (.A1(n_546), .A2(n_550), .ZN(n_545));
   NAND3_X1 i_559 (.A1(n_578), .A2(n_547), .A3(n_573), .ZN(n_546));
   NAND2_X1 i_560 (.A1(n_549), .A2(n_548), .ZN(n_547));
   NAND2_X1 i_561 (.A1(n_571), .A2(n_570), .ZN(n_548));
   NAND2_X1 i_562 (.A1(n_564), .A2(n_567), .ZN(n_549));
   NOR2_X1 i_563 (.A1(n_554), .A2(n_551), .ZN(n_550));
   AOI21_X1 i_564 (.A(n_558), .B1(n_556), .B2(n_559), .ZN(n_551));
   INV_X1 i_565 (.A(n_555), .ZN(n_554));
   NAND3_X1 i_566 (.A1(n_559), .A2(n_558), .A3(n_556), .ZN(n_555));
   NAND4_X1 i_567 (.A1(T_Count[1]), .A2(T_Count[0]), .A3(num_of_X[9]), .A4(
      num_of_X[8]), .ZN(n_556));
   NAND2_X1 i_568 (.A1(T_Count[2]), .A2(num_of_X[7]), .ZN(n_558));
   OAI21_X1 i_569 (.A(n_560), .B1(n_665), .B2(n_561), .ZN(n_559));
   NAND2_X1 i_570 (.A1(T_Count[1]), .A2(num_of_X[8]), .ZN(n_560));
   INV_X1 i_571 (.A(num_of_X[9]), .ZN(n_561));
   OAI21_X1 i_572 (.A(n_576), .B1(n_572), .B2(n_563), .ZN(n_562));
   AOI22_X1 i_573 (.A1(n_564), .A2(n_567), .B1(n_571), .B2(n_570), .ZN(n_563));
   NAND2_X1 i_574 (.A1(n_566), .A2(n_565), .ZN(n_564));
   NAND2_X1 i_575 (.A1(T_Count[1]), .A2(num_of_X[6]), .ZN(n_565));
   NAND3_X1 i_576 (.A1(X_Count[7]), .A2(T_Count[0]), .A3(num_of_X[7]), .ZN(n_566));
   NAND2_X1 i_577 (.A1(n_568), .A2(n_569), .ZN(n_567));
   NAND2_X1 i_578 (.A1(T_Count[0]), .A2(num_of_X[7]), .ZN(n_568));
   INV_X1 i_579 (.A(X_Count[7]), .ZN(n_569));
   INV_X1 i_580 (.A(n_600), .ZN(n_570));
   INV_X1 i_581 (.A(n_645), .ZN(n_571));
   INV_X1 i_582 (.A(n_573), .ZN(n_572));
   OAI21_X1 i_583 (.A(n_574), .B1(n_575), .B2(n_431), .ZN(n_573));
   NAND2_X1 i_584 (.A1(T_Count[5]), .A2(num_of_X[3]), .ZN(n_574));
   INV_X1 i_585 (.A(num_of_X[4]), .ZN(n_431));
   INV_X1 i_586 (.A(T_Count[4]), .ZN(n_575));
   INV_X1 i_587 (.A(n_578), .ZN(n_576));
   NAND2_X1 i_588 (.A1(n_579), .A2(n_414), .ZN(n_578));
   NAND3_X1 i_589 (.A1(n_601), .A2(T_Count[7]), .A3(num_of_X[2]), .ZN(n_414));
   NAND2_X1 i_590 (.A1(n_415), .A2(n_581), .ZN(n_579));
   INV_X1 i_591 (.A(n_582), .ZN(n_581));
   NAND2_X1 i_592 (.A1(T_Count[3]), .A2(num_of_X[5]), .ZN(n_582));
   OAI21_X1 i_593 (.A(n_583), .B1(n_417), .B2(n_584), .ZN(n_415));
   NAND2_X1 i_594 (.A1(T_Count[7]), .A2(num_of_X[1]), .ZN(n_583));
   INV_X1 i_595 (.A(num_of_X[2]), .ZN(n_584));
   INV_X1 i_596 (.A(T_Count[6]), .ZN(n_417));
   NAND2_X1 i_597 (.A1(n_586), .A2(n_622), .ZN(n_585));
   AOI21_X1 i_598 (.A(n_613), .B1(n_588), .B2(n_587), .ZN(n_586));
   NAND4_X1 i_599 (.A1(n_619), .A2(n_617), .A3(n_616), .A4(n_614), .ZN(n_587));
   NAND2_X1 i_600 (.A1(n_589), .A2(n_595), .ZN(n_588));
   NAND2_X1 i_601 (.A1(n_594), .A2(n_590), .ZN(n_589));
   NAND2_X1 i_602 (.A1(n_592), .A2(n_591), .ZN(n_590));
   NAND3_X1 i_603 (.A1(n_651), .A2(n_650), .A3(n_648), .ZN(n_591));
   OAI21_X1 i_604 (.A(n_647), .B1(n_593), .B2(n_649), .ZN(n_592));
   INV_X1 i_605 (.A(n_651), .ZN(n_593));
   NAND3_X1 i_606 (.A1(n_605), .A2(n_603), .A3(n_597), .ZN(n_594));
   NAND2_X1 i_607 (.A1(n_604), .A2(n_596), .ZN(n_595));
   NAND2_X1 i_608 (.A1(n_597), .A2(n_603), .ZN(n_596));
   NAND2_X1 i_609 (.A1(n_598), .A2(n_601), .ZN(n_597));
   NAND2_X1 i_610 (.A1(n_600), .A2(n_599), .ZN(n_598));
   NAND2_X1 i_611 (.A1(T_Count[5]), .A2(num_of_X[2]), .ZN(n_599));
   NAND2_X1 i_612 (.A1(T_Count[4]), .A2(num_of_X[3]), .ZN(n_600));
   INV_X1 i_613 (.A(n_602), .ZN(n_601));
   NAND2_X1 i_614 (.A1(T_Count[6]), .A2(num_of_X[1]), .ZN(n_602));
   NAND3_X1 i_615 (.A1(n_641), .A2(num_of_X[3]), .A3(num_of_X[2]), .ZN(n_603));
   INV_X1 i_616 (.A(n_605), .ZN(n_604));
   OAI21_X1 i_617 (.A(n_610), .B1(n_606), .B2(n_608), .ZN(n_605));
   INV_X1 i_618 (.A(n_607), .ZN(n_606));
   NAND4_X1 i_619 (.A1(T_Count[7]), .A2(T_Count[2]), .A3(num_of_X[5]), .A4(
      num_of_X[0]), .ZN(n_607));
   INV_X1 i_620 (.A(n_609), .ZN(n_608));
   NAND2_X1 i_621 (.A1(T_Count[3]), .A2(num_of_X[4]), .ZN(n_609));
   OAI21_X1 i_622 (.A(n_611), .B1(n_612), .B2(n_298), .ZN(n_610));
   NAND2_X1 i_623 (.A1(T_Count[7]), .A2(num_of_X[0]), .ZN(n_611));
   INV_X1 i_624 (.A(num_of_X[5]), .ZN(n_298));
   INV_X1 i_625 (.A(T_Count[2]), .ZN(n_612));
   AOI22_X1 i_626 (.A1(n_619), .A2(n_617), .B1(n_614), .B2(n_616), .ZN(n_613));
   NAND2_X1 i_627 (.A1(n_615), .A2(n_636), .ZN(n_614));
   NAND2_X1 i_628 (.A1(n_634), .A2(n_638), .ZN(n_615));
   NAND3_X1 i_629 (.A1(n_638), .A2(n_634), .A3(n_637), .ZN(n_616));
   NAND3_X1 i_630 (.A1(n_618), .A2(n_651), .A3(n_621), .ZN(n_617));
   NAND2_X1 i_631 (.A1(n_296), .A2(n_643), .ZN(n_618));
   NAND3_X1 i_632 (.A1(n_620), .A2(n_643), .A3(n_296), .ZN(n_619));
   NAND2_X1 i_633 (.A1(n_621), .A2(n_651), .ZN(n_620));
   NAND2_X1 i_634 (.A1(n_650), .A2(n_648), .ZN(n_621));
   NAND2_X1 i_635 (.A1(n_628), .A2(n_626), .ZN(n_622));
   NAND3_X1 i_637 (.A1(n_631), .A2(n_655), .A3(n_627), .ZN(n_626));
   NAND2_X1 i_638 (.A1(n_633), .A2(n_266), .ZN(n_627));
   OAI21_X1 i_639 (.A(n_654), .B1(n_630), .B2(n_629), .ZN(n_628));
   AOI22_X1 i_640 (.A1(n_283), .A2(n_296), .B1(n_635), .B2(n_634), .ZN(n_629));
   INV_X1 i_641 (.A(n_631), .ZN(n_630));
   NAND3_X1 i_642 (.A1(n_632), .A2(n_283), .A3(n_296), .ZN(n_631));
   INV_X1 i_643 (.A(n_633), .ZN(n_632));
   NAND2_X1 i_644 (.A1(n_635), .A2(n_634), .ZN(n_633));
   NAND4_X1 i_645 (.A1(T_Count[7]), .A2(T_Count[6]), .A3(num_of_X[3]), .A4(
      num_of_X[2]), .ZN(n_634));
   NAND2_X1 i_646 (.A1(n_638), .A2(n_636), .ZN(n_635));
   INV_X1 i_647 (.A(n_637), .ZN(n_636));
   NAND2_X1 i_648 (.A1(T_Count[3]), .A2(num_of_X[6]), .ZN(n_637));
   NAND2_X1 i_649 (.A1(n_640), .A2(n_639), .ZN(n_638));
   NAND2_X1 i_650 (.A1(T_Count[7]), .A2(num_of_X[2]), .ZN(n_639));
   NAND2_X1 i_651 (.A1(T_Count[6]), .A2(num_of_X[3]), .ZN(n_640));
   NAND3_X1 i_652 (.A1(n_641), .A2(num_of_X[5]), .A3(num_of_X[4]), .ZN(n_296));
   INV_X1 i_653 (.A(n_642), .ZN(n_641));
   NAND2_X1 i_654 (.A1(T_Count[5]), .A2(T_Count[4]), .ZN(n_642));
   OAI211_X1 i_655 (.A(n_651), .B(n_643), .C1(n_649), .C2(n_647), .ZN(n_283));
   NAND2_X1 i_656 (.A1(n_645), .A2(n_644), .ZN(n_643));
   NAND2_X1 i_657 (.A1(T_Count[4]), .A2(num_of_X[5]), .ZN(n_644));
   NAND2_X1 i_658 (.A1(T_Count[5]), .A2(num_of_X[4]), .ZN(n_645));
   INV_X1 i_659 (.A(n_648), .ZN(n_647));
   NAND2_X1 i_660 (.A1(T_Count[2]), .A2(num_of_X[6]), .ZN(n_648));
   INV_X1 i_661 (.A(n_650), .ZN(n_649));
   NAND4_X1 i_662 (.A1(T_Count[1]), .A2(T_Count[0]), .A3(num_of_X[8]), .A4(
      num_of_X[7]), .ZN(n_650));
   NAND2_X1 i_663 (.A1(n_653), .A2(n_652), .ZN(n_651));
   NAND2_X1 i_664 (.A1(T_Count[1]), .A2(num_of_X[7]), .ZN(n_652));
   NAND2_X1 i_665 (.A1(T_Count[0]), .A2(num_of_X[8]), .ZN(n_653));
   INV_X1 i_666 (.A(n_655), .ZN(n_654));
   NAND2_X1 i_667 (.A1(n_656), .A2(n_660), .ZN(n_655));
   NAND2_X1 i_668 (.A1(n_658), .A2(n_659), .ZN(n_656));
   NAND2_X1 i_669 (.A1(n_663), .A2(n_662), .ZN(n_658));
   INV_X1 i_670 (.A(n_661), .ZN(n_659));
   NAND3_X1 i_671 (.A1(n_663), .A2(n_662), .A3(n_661), .ZN(n_660));
   NAND2_X1 i_672 (.A1(T_Count[2]), .A2(num_of_X[8]), .ZN(n_661));
   NAND4_X1 i_673 (.A1(T_Count[1]), .A2(T_Count[0]), .A3(num_of_X[10]), .A4(
      num_of_X[9]), .ZN(n_662));
   OAI21_X1 i_674 (.A(n_664), .B1(n_665), .B2(n_277), .ZN(n_663));
   NAND2_X1 i_675 (.A1(T_Count[1]), .A2(num_of_X[9]), .ZN(n_664));
   INV_X1 i_676 (.A(num_of_X[10]), .ZN(n_277));
   INV_X1 i_677 (.A(T_Count[0]), .ZN(n_665));
   INV_X1 i_678 (.A(n_667), .ZN(n_666));
   XNOR2_X1 i_679 (.A(n_91), .B(n_97), .ZN(n_667));
   BUF_X1 rt_shieldBuf__1__1__0 (.A(T_Count[3]), .Z(n_255));
   NAND3_X1 i_302 (.A1(n_123), .A2(n_233), .A3(n_145), .ZN(n_256));
   NAND2_X1 i_303 (.A1(n_124), .A2(n_254), .ZN(n_257));
   NAND2_X1 i_326 (.A1(n_116), .A2(n_115), .ZN(n_259));
   NAND2_X1 i_328 (.A1(n_145), .A2(n_233), .ZN(n_262));
   INV_X1 i_351 (.A(n_262), .ZN(n_274));
   NAND2_X1 i_448 (.A1(n_123), .A2(n_274), .ZN(n_275));
   NAND3_X1 i_375 (.A1(n_257), .A2(n_259), .A3(n_275), .ZN(n_276));
   NAND2_X1 i_385 (.A1(n_108), .A2(n_116), .ZN(n_281));
   NAND2_X1 i_393 (.A1(n_101), .A2(n_104), .ZN(n_282));
   NAND3_X1 i_404 (.A1(n_105), .A2(n_102), .A3(n_103), .ZN(n_313));
   NAND2_X1 i_680 (.A1(n_101), .A2(n_104), .ZN(n_330));
   NAND2_X1 i_681 (.A1(n_108), .A2(n_116), .ZN(n_668));
   NAND2_X1 i_684 (.A1(n_105), .A2(n_677), .ZN(n_669));
   NAND3_X1 i_685 (.A1(n_330), .A2(n_668), .A3(n_669), .ZN(n_670));
   OAI21_X1 i_682 (.A(n_235), .B1(n_234), .B2(n_236), .ZN(n_671));
   INV_X1 i_683 (.A(n_235), .ZN(n_672));
   INV_X1 i_686 (.A(n_234), .ZN(n_673));
   INV_X1 i_687 (.A(n_236), .ZN(n_674));
   AOI21_X1 i_688 (.A(n_672), .B1(n_673), .B2(n_674), .ZN(n_675));
   NAND2_X1 i_330 (.A1(n_103), .A2(n_102), .ZN(n_676));
   INV_X1 i_343 (.A(n_676), .ZN(n_677));
endmodule

module datapath__1_501(p_0, X_Count, p_1);
   input [63:0]p_0;
   input [7:0]X_Count;
   output p_1;

   XNOR2_X1 i_0 (.A(X_Count[0]), .B(p_0[0]), .ZN(n_0));
   INV_X1 i_1 (.A(n_0), .ZN(n_1));
   XNOR2_X1 i_2 (.A(X_Count[1]), .B(p_0[1]), .ZN(n_2));
   INV_X1 i_3 (.A(n_2), .ZN(n_3));
   XNOR2_X1 i_4 (.A(X_Count[2]), .B(p_0[2]), .ZN(n_4));
   INV_X1 i_5 (.A(n_4), .ZN(n_5));
   XNOR2_X1 i_6 (.A(X_Count[3]), .B(p_0[3]), .ZN(n_6));
   INV_X1 i_7 (.A(n_6), .ZN(n_7));
   XNOR2_X1 i_8 (.A(X_Count[4]), .B(p_0[4]), .ZN(n_8));
   INV_X1 i_9 (.A(n_8), .ZN(n_9));
   XNOR2_X1 i_10 (.A(X_Count[5]), .B(p_0[5]), .ZN(n_10));
   INV_X1 i_11 (.A(n_10), .ZN(n_11));
   XNOR2_X1 i_12 (.A(X_Count[6]), .B(p_0[6]), .ZN(n_12));
   INV_X1 i_13 (.A(n_12), .ZN(n_13));
   XNOR2_X1 i_14 (.A(X_Count[7]), .B(p_0[7]), .ZN(n_14));
   INV_X1 i_15 (.A(n_14), .ZN(n_15));
   NOR2_X1 i_16 (.A1(p_0[63]), .A2(p_0[62]), .ZN(n_16));
   NOR2_X1 i_17 (.A1(p_0[61]), .A2(p_0[60]), .ZN(n_17));
   NOR2_X1 i_18 (.A1(p_0[59]), .A2(p_0[58]), .ZN(n_18));
   NOR2_X1 i_19 (.A1(p_0[57]), .A2(p_0[56]), .ZN(n_19));
   NOR2_X1 i_20 (.A1(p_0[55]), .A2(p_0[54]), .ZN(n_20));
   NOR2_X1 i_21 (.A1(p_0[53]), .A2(p_0[52]), .ZN(n_21));
   NOR2_X1 i_22 (.A1(p_0[51]), .A2(p_0[50]), .ZN(n_22));
   NOR2_X1 i_23 (.A1(p_0[49]), .A2(p_0[48]), .ZN(n_23));
   NOR2_X1 i_24 (.A1(p_0[47]), .A2(p_0[46]), .ZN(n_24));
   NOR2_X1 i_25 (.A1(p_0[45]), .A2(p_0[44]), .ZN(n_25));
   NOR2_X1 i_26 (.A1(p_0[43]), .A2(p_0[42]), .ZN(n_26));
   NOR2_X1 i_27 (.A1(p_0[41]), .A2(p_0[40]), .ZN(n_27));
   NOR2_X1 i_28 (.A1(p_0[39]), .A2(p_0[38]), .ZN(n_28));
   NOR2_X1 i_29 (.A1(p_0[37]), .A2(p_0[36]), .ZN(n_29));
   NOR2_X1 i_30 (.A1(p_0[35]), .A2(p_0[34]), .ZN(n_30));
   NOR2_X1 i_31 (.A1(p_0[33]), .A2(p_0[32]), .ZN(n_31));
   NOR2_X1 i_32 (.A1(p_0[31]), .A2(p_0[30]), .ZN(n_32));
   NOR2_X1 i_33 (.A1(p_0[29]), .A2(p_0[28]), .ZN(n_33));
   NOR2_X1 i_34 (.A1(p_0[27]), .A2(p_0[26]), .ZN(n_34));
   NOR2_X1 i_35 (.A1(p_0[25]), .A2(p_0[24]), .ZN(n_35));
   NOR2_X1 i_36 (.A1(p_0[23]), .A2(p_0[22]), .ZN(n_36));
   NOR2_X1 i_37 (.A1(p_0[21]), .A2(p_0[20]), .ZN(n_37));
   NOR2_X1 i_38 (.A1(p_0[19]), .A2(p_0[18]), .ZN(n_38));
   NOR2_X1 i_39 (.A1(p_0[17]), .A2(p_0[16]), .ZN(n_39));
   NOR2_X1 i_40 (.A1(p_0[15]), .A2(p_0[14]), .ZN(n_40));
   NOR2_X1 i_41 (.A1(p_0[13]), .A2(p_0[12]), .ZN(n_41));
   NOR2_X1 i_42 (.A1(p_0[11]), .A2(p_0[10]), .ZN(n_42));
   NOR2_X1 i_43 (.A1(p_0[9]), .A2(p_0[8]), .ZN(n_43));
   NOR2_X1 i_44 (.A1(n_15), .A2(n_13), .ZN(n_44));
   NOR2_X1 i_45 (.A1(n_11), .A2(n_9), .ZN(n_45));
   NOR2_X1 i_46 (.A1(n_7), .A2(n_5), .ZN(n_46));
   NOR2_X1 i_47 (.A1(n_3), .A2(n_1), .ZN(n_47));
   NAND4_X1 i_48 (.A1(n_16), .A2(n_17), .A3(n_18), .A4(n_19), .ZN(n_48));
   NAND4_X1 i_49 (.A1(n_20), .A2(n_21), .A3(n_22), .A4(n_23), .ZN(n_49));
   NAND4_X1 i_50 (.A1(n_24), .A2(n_25), .A3(n_26), .A4(n_27), .ZN(n_50));
   NAND4_X1 i_51 (.A1(n_28), .A2(n_29), .A3(n_30), .A4(n_31), .ZN(n_51));
   NAND4_X1 i_52 (.A1(n_32), .A2(n_33), .A3(n_34), .A4(n_35), .ZN(n_52));
   NAND4_X1 i_53 (.A1(n_36), .A2(n_37), .A3(n_38), .A4(n_39), .ZN(n_53));
   NAND4_X1 i_54 (.A1(n_40), .A2(n_41), .A3(n_42), .A4(n_43), .ZN(n_54));
   NAND4_X1 i_55 (.A1(n_44), .A2(n_45), .A3(n_46), .A4(n_47), .ZN(n_55));
   NOR2_X1 i_56 (.A1(n_48), .A2(n_49), .ZN(n_56));
   NOR2_X1 i_57 (.A1(n_50), .A2(n_51), .ZN(n_57));
   NOR2_X1 i_58 (.A1(n_52), .A2(n_53), .ZN(n_58));
   NOR2_X1 i_59 (.A1(n_54), .A2(n_55), .ZN(n_59));
   NAND4_X1 i_60 (.A1(n_56), .A2(n_57), .A3(n_58), .A4(n_59), .ZN(n_60));
   INV_X1 i_61 (.A(n_60), .ZN(p_1));
endmodule

module datapath__1_506(p_0, T_Count, p_1);
   input [63:0]p_0;
   input [7:0]T_Count;
   output p_1;

   XNOR2_X1 i_0 (.A(T_Count[0]), .B(p_0[0]), .ZN(n_0));
   INV_X1 i_1 (.A(n_0), .ZN(n_1));
   XNOR2_X1 i_2 (.A(T_Count[1]), .B(p_0[1]), .ZN(n_2));
   INV_X1 i_3 (.A(n_2), .ZN(n_3));
   XNOR2_X1 i_4 (.A(T_Count[2]), .B(p_0[2]), .ZN(n_4));
   INV_X1 i_5 (.A(n_4), .ZN(n_5));
   XNOR2_X1 i_6 (.A(T_Count[3]), .B(p_0[3]), .ZN(n_6));
   INV_X1 i_7 (.A(n_6), .ZN(n_7));
   XNOR2_X1 i_8 (.A(T_Count[4]), .B(p_0[4]), .ZN(n_8));
   INV_X1 i_9 (.A(n_8), .ZN(n_9));
   XNOR2_X1 i_10 (.A(T_Count[5]), .B(p_0[5]), .ZN(n_10));
   INV_X1 i_11 (.A(n_10), .ZN(n_11));
   XNOR2_X1 i_12 (.A(T_Count[6]), .B(p_0[6]), .ZN(n_12));
   INV_X1 i_13 (.A(n_12), .ZN(n_13));
   XNOR2_X1 i_14 (.A(T_Count[7]), .B(p_0[7]), .ZN(n_14));
   INV_X1 i_15 (.A(n_14), .ZN(n_15));
   NOR2_X1 i_16 (.A1(p_0[63]), .A2(p_0[62]), .ZN(n_16));
   NOR2_X1 i_17 (.A1(p_0[61]), .A2(p_0[60]), .ZN(n_17));
   NOR2_X1 i_18 (.A1(p_0[59]), .A2(p_0[58]), .ZN(n_18));
   NOR2_X1 i_19 (.A1(p_0[57]), .A2(p_0[56]), .ZN(n_19));
   NOR2_X1 i_20 (.A1(p_0[55]), .A2(p_0[54]), .ZN(n_20));
   NOR2_X1 i_21 (.A1(p_0[53]), .A2(p_0[52]), .ZN(n_21));
   NOR2_X1 i_22 (.A1(p_0[51]), .A2(p_0[50]), .ZN(n_22));
   NOR2_X1 i_23 (.A1(p_0[49]), .A2(p_0[48]), .ZN(n_23));
   NOR2_X1 i_24 (.A1(p_0[47]), .A2(p_0[46]), .ZN(n_24));
   NOR2_X1 i_25 (.A1(p_0[45]), .A2(p_0[44]), .ZN(n_25));
   NOR2_X1 i_26 (.A1(p_0[43]), .A2(p_0[42]), .ZN(n_26));
   NOR2_X1 i_27 (.A1(p_0[41]), .A2(p_0[40]), .ZN(n_27));
   NOR2_X1 i_28 (.A1(p_0[39]), .A2(p_0[38]), .ZN(n_28));
   NOR2_X1 i_29 (.A1(p_0[37]), .A2(p_0[36]), .ZN(n_29));
   NOR2_X1 i_30 (.A1(p_0[35]), .A2(p_0[34]), .ZN(n_30));
   NOR2_X1 i_31 (.A1(p_0[33]), .A2(p_0[32]), .ZN(n_31));
   NOR2_X1 i_32 (.A1(p_0[31]), .A2(p_0[30]), .ZN(n_32));
   NOR2_X1 i_33 (.A1(p_0[29]), .A2(p_0[28]), .ZN(n_33));
   NOR2_X1 i_34 (.A1(p_0[27]), .A2(p_0[26]), .ZN(n_34));
   NOR2_X1 i_35 (.A1(p_0[25]), .A2(p_0[24]), .ZN(n_35));
   NOR2_X1 i_36 (.A1(p_0[23]), .A2(p_0[22]), .ZN(n_36));
   NOR2_X1 i_37 (.A1(p_0[21]), .A2(p_0[20]), .ZN(n_37));
   NOR2_X1 i_38 (.A1(p_0[19]), .A2(p_0[18]), .ZN(n_38));
   NOR2_X1 i_39 (.A1(p_0[17]), .A2(p_0[16]), .ZN(n_39));
   NOR2_X1 i_40 (.A1(p_0[15]), .A2(p_0[14]), .ZN(n_40));
   NOR2_X1 i_41 (.A1(p_0[13]), .A2(p_0[12]), .ZN(n_41));
   NOR2_X1 i_42 (.A1(p_0[11]), .A2(p_0[10]), .ZN(n_42));
   NOR2_X1 i_43 (.A1(p_0[9]), .A2(p_0[8]), .ZN(n_43));
   NOR2_X1 i_44 (.A1(n_15), .A2(n_13), .ZN(n_44));
   NOR2_X1 i_45 (.A1(n_11), .A2(n_9), .ZN(n_45));
   NOR2_X1 i_46 (.A1(n_7), .A2(n_5), .ZN(n_46));
   NOR2_X1 i_47 (.A1(n_3), .A2(n_1), .ZN(n_47));
   NAND4_X1 i_48 (.A1(n_16), .A2(n_17), .A3(n_18), .A4(n_19), .ZN(n_48));
   NAND4_X1 i_49 (.A1(n_20), .A2(n_21), .A3(n_22), .A4(n_23), .ZN(n_49));
   NAND4_X1 i_50 (.A1(n_24), .A2(n_25), .A3(n_26), .A4(n_27), .ZN(n_50));
   NAND4_X1 i_51 (.A1(n_28), .A2(n_29), .A3(n_30), .A4(n_31), .ZN(n_51));
   NAND4_X1 i_52 (.A1(n_32), .A2(n_33), .A3(n_34), .A4(n_35), .ZN(n_52));
   NAND4_X1 i_53 (.A1(n_36), .A2(n_37), .A3(n_38), .A4(n_39), .ZN(n_53));
   NAND4_X1 i_54 (.A1(n_40), .A2(n_41), .A3(n_42), .A4(n_43), .ZN(n_54));
   NAND4_X1 i_55 (.A1(n_44), .A2(n_45), .A3(n_46), .A4(n_47), .ZN(n_55));
   NOR2_X1 i_56 (.A1(n_48), .A2(n_49), .ZN(n_56));
   NOR2_X1 i_57 (.A1(n_50), .A2(n_51), .ZN(n_57));
   NOR2_X1 i_58 (.A1(n_52), .A2(n_53), .ZN(n_58));
   NOR2_X1 i_59 (.A1(n_54), .A2(n_55), .ZN(n_59));
   NAND4_X1 i_60 (.A1(n_56), .A2(n_57), .A3(n_58), .A4(n_59), .ZN(n_60));
   INV_X1 i_61 (.A(n_60), .ZN(p_1));
endmodule

module Results_Sender(RST, CLK, Sending_Enable, CPU_Bus, Done_Sending, 
      RAM_Data_A, RAM_Data_B, RAM_Address_A, RAM_Address_B);
   input RST;
   input CLK;
   input Sending_Enable;
   output [31:0]CPU_Bus;
   output Done_Sending;
   input [63:0]RAM_Data_A;
   input [63:0]RAM_Data_B;
   output [12:0]RAM_Address_A;
   output [12:0]RAM_Address_B;

   wire [1:0]Partial_Data_Count;
   wire [1:0]T_OR_X;
   wire [7:0]X_Count;
   wire [7:0]T_Count;
   wire [1:0]Init_Count;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire [63:0]num_of_T;
   wire [63:0]num_of_X;
   wire n_0_0;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_183;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_22_0;
   wire Init_Counter_genblk1_1_counterBits_n_4;
   wire Init_Counter_genblk1_1_counterBits_n_2;
   wire Init_Counter_firstBit_n_4;
   wire Init_Counter_firstBit_n_2;
   wire T_Counter_genblk1_7_counterBits_n_4;
   wire T_Counter_genblk1_7_counterBits_n_2;
   wire T_Counter_genblk1_6_counterBits_n_4;
   wire T_Counter_genblk1_6_counterBits_n_2;
   wire n_0_22_1;
   wire T_Counter_genblk1_5_counterBits_n_4;
   wire T_Counter_genblk1_5_counterBits_n_2;
   wire T_Counter_genblk1_4_counterBits_n_4;
   wire T_Counter_genblk1_4_counterBits_n_2;
   wire n_0_22_2;
   wire n_0_22_3;
   wire T_Counter_genblk1_3_counterBits_n_4;
   wire T_Counter_genblk1_3_counterBits_n_2;
   wire n_0_22_4;
   wire T_Counter_genblk1_2_counterBits_n_4;
   wire T_Counter_genblk1_2_counterBits_n_2;
   wire n_0_22_5;
   wire T_Counter_genblk1_1_counterBits_n_4;
   wire T_Counter_genblk1_1_counterBits_n_2;
   wire T_Counter_firstBit_n_4;
   wire T_Counter_firstBit_n_2;
   wire n_0_22_6;
   wire n_0_22_7;
   wire X_Counter_genblk1_7_counterBits_n_4;
   wire X_Counter_genblk1_7_counterBits_n_2;
   wire X_Counter_genblk1_6_counterBits_n_4;
   wire X_Counter_genblk1_6_counterBits_n_2;
   wire n_0_22_8;
   wire X_Counter_genblk1_5_counterBits_n_4;
   wire X_Counter_genblk1_5_counterBits_n_2;
   wire X_Counter_genblk1_4_counterBits_n_4;
   wire X_Counter_genblk1_4_counterBits_n_2;
   wire n_0_22_9;
   wire n_0_22_10;
   wire X_Counter_genblk1_3_counterBits_n_4;
   wire X_Counter_genblk1_3_counterBits_n_2;
   wire n_0_22_11;
   wire X_Counter_genblk1_2_counterBits_n_4;
   wire X_Counter_genblk1_2_counterBits_n_2;
   wire n_0_22_12;
   wire X_Counter_genblk1_1_counterBits_n_4;
   wire X_Counter_genblk1_1_counterBits_n_2;
   wire X_Counter_firstBit_n_4;
   wire X_Counter_firstBit_n_2;
   wire n_0_22_13;
   wire n_0_22_14;
   wire T_OR_X_COUNTER_firstBit_n_4;
   wire T_OR_X_COUNTER_firstBit_n_2;
   wire _64data_Counter_firstBit_n_4;
   wire _64data_Counter_firstBit_n_2;
   wire n_0_341;
   wire n_0_342;
   wire n_0_22_15;
   wire n_0_22_16;
   wire n_0_22_17;
   wire n_0_22_18;
   wire n_0_22_19;
   wire n_0_22_20;
   wire n_0_22_21;
   wire n_0_22_22;
   wire n_0_22_23;
   wire n_0_22_24;
   wire n_0_22_25;
   wire n_0_22_26;
   wire n_0_22_27;
   wire n_0_22_28;
   wire n_0_22_29;
   wire n_0_22_30;
   wire n_0_22_31;
   wire n_0_22_32;
   wire n_0_22_33;
   wire n_0_22_34;
   wire n_0_22_35;
   wire n_0_22_36;
   wire n_0_22_37;
   wire n_0_22_38;
   wire n_0_22_39;
   wire n_0_22_40;
   wire n_0_22_41;
   wire n_0_22_42;
   wire n_0_22_43;
   wire n_0_22_44;
   wire n_0_22_45;
   wire n_0_22_46;
   wire n_0_22_47;
   wire n_0_22_48;
   wire n_0_22_49;
   wire n_0_22_50;
   wire n_0_22_51;
   wire n_0_22_52;
   wire n_0_22_53;
   wire n_0_22_54;
   wire n_0_22_55;
   wire n_0_22_56;
   wire n_0_22_57;
   wire n_0_22_58;
   wire n_0_22_59;
   wire n_0_22_60;
   wire n_0_22_61;
   wire n_0_22_62;
   wire n_0_22_63;
   wire n_0_22_64;
   wire n_0_22_65;
   wire n_0_22_66;
   wire n_0_22_67;
   wire n_0_22_68;
   wire n_0_22_69;
   wire n_0_22_70;
   wire n_0_22_71;
   wire n_0_22_72;
   wire n_0_22_73;
   wire n_0_22_74;
   wire n_0_22_75;
   wire n_0_22_76;
   wire n_0_22_77;
   wire n_0_22_78;
   wire n_0_22_79;
   wire n_0_22_80;
   wire n_0_140;
   wire n_0_22_81;
   wire n_0_22_82;
   wire n_0_22_83;
   wire n_0_22_84;
   wire n_0_139;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_159;
   wire n_0_25_0;
   wire n_0_160;
   wire n_0_25_1;
   wire n_0_161;
   wire n_0_25_2;
   wire n_0_162;
   wire n_0_25_3;
   wire n_0_163;
   wire n_0_25_4;
   wire n_0_164;
   wire n_0_165;
   wire n_0_360;
   wire n_0_25_5;
   wire n_0_361;
   wire n_0_25_6;
   wire n_0_362;
   wire n_0_25_7;
   wire n_0_25_8;
   wire n_0_25_9;
   wire n_0_158;
   wire n_0_363;
   wire n_0_25_10;
   wire n_0_25_11;
   wire n_0_25_12;
   wire n_0_25_13;
   wire n_0_25_14;
   wire n_0_25_15;
   wire n_0_25_16;
   wire n_0_25_17;
   wire n_0_25_18;
   wire n_0_25_19;
   wire n_0_25_20;
   wire n_0_25_21;
   wire n_0_25_22;
   wire n_0_25_23;
   wire n_0_25_24;
   wire n_0_25_25;
   wire n_0_25_26;
   wire n_0_25_27;
   wire n_0_25_28;
   wire n_0_25_29;
   wire n_0_25_30;
   wire n_0_25_31;
   wire n_0_25_32;
   wire n_0_25_33;
   wire n_0_25_34;
   wire n_0_25_35;
   wire n_0_25_36;
   wire n_0_25_37;
   wire n_0_25_38;
   wire n_0_109;
   wire n_0_340;
   wire n_0_25_39;
   wire n_0_343;
   wire n_0_137;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire X_Counter_firstBit_Q_reg_enable_mux_n_0;
   wire X_Counter_firstBit_Q_reg_enable_mux_n_1;
   wire n_0_114;
   wire X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_n_0;
   wire X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_n_1;
   wire X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_n_2;
   wire n_0_115;
   wire X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_n_0;
   wire X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_n_1;
   wire X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_n_2;
   wire n_0_134;
   wire X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_n_0;
   wire X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_n_1;
   wire X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_n_2;
   wire n_0_135;
   wire X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_n_0;
   wire X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_n_1;
   wire X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_n_2;
   wire n_0_180;
   wire X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_n_0;
   wire X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_n_1;
   wire X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_n_2;
   wire n_0_181;
   wire X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_n_0;
   wire X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_n_1;
   wire X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_n_2;
   wire n_0_182;
   wire X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_n_0;
   wire X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_n_1;
   wire X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_n_2;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_242;
   wire n_0_243;
   wire n_0_308;
   wire n_0_136;
   wire n_0_30_0;
   wire n_0_138;
   wire n_0_30_1;
   wire n_0_30_2;
   wire n_0_30_3;
   wire n_0_30_4;
   wire n_0_344;
   wire n_0_157;
   wire n_0_4_0;
   wire n_0_4_1;
   wire n_0_5_0;
   wire n_0_5_1;
   wire n_0_5_2;
   wire n_0_5_3;
   wire n_0_5_4;
   wire n_0_5_5;
   wire n_0_5_6;
   wire n_0_5_7;
   wire n_0_5_8;
   wire n_0_5_9;
   wire n_0_5_10;
   wire n_0_5_11;
   wire n_0_5_12;
   wire n_0_5_13;
   wire n_0_5_14;
   wire n_0_345;
   wire n_0_6_0;
   wire n_0_6_1;
   wire n_0_6_2;
   wire n_0_6_3;
   wire n_0_6_4;
   wire n_0_6_5;
   wire n_0_6_6;
   wire n_0_6_7;
   wire n_0_6_8;
   wire n_0_346;
   wire n_0_347;
   wire n_0_7_0;
   wire n_0_7_1;
   wire n_0_7_2;
   wire n_0_7_3;
   wire n_0_7_4;
   wire n_0_7_5;
   wire n_0_7_6;
   wire n_0_7_7;
   wire n_0_8_0;
   wire n_0_8_1;
   wire n_0_8_2;
   wire n_0_8_3;
   wire n_0_8_4;
   wire n_0_8_5;
   wire n_0_8_6;
   wire n_0_8_7;
   wire n_0_8_8;
   wire n_0_8_9;
   wire n_0_348;
   wire n_0_349;
   wire n_0_9_0;
   wire n_0_9_1;
   wire n_0_9_2;
   wire n_0_9_3;
   wire n_0_9_4;
   wire n_0_9_5;
   wire n_0_9_6;
   wire n_0_9_7;
   wire n_0_350;
   wire n_0_10_0;
   wire n_0_10_1;
   wire n_0_10_2;
   wire n_0_10_3;
   wire n_0_10_4;
   wire n_0_10_5;
   wire n_0_10_6;
   wire n_0_10_7;
   wire n_0_11_0;
   wire n_0_11_1;
   wire n_0_11_2;
   wire n_0_11_3;
   wire n_0_11_4;
   wire n_0_11_5;
   wire n_0_11_6;
   wire n_0_11_7;
   wire n_0_11_8;
   wire n_0_11_9;
   wire n_0_11_10;
   wire n_0_351;
   wire n_0_12_0;
   wire n_0_12_1;
   wire n_0_12_2;
   wire n_0_12_3;
   wire n_0_12_4;
   wire n_0_12_5;
   wire n_0_12_6;
   wire n_0_12_7;
   wire n_0_12_8;
   wire n_0_12_9;
   wire n_0_12_10;
   wire n_0_352;
   wire n_0_13_0;
   wire n_0_13_1;
   wire n_0_13_2;
   wire n_0_13_3;
   wire n_0_13_4;
   wire n_0_13_5;
   wire n_0_13_6;
   wire n_0_13_7;
   wire n_0_13_8;
   wire n_0_13_9;
   wire n_0_13_10;
   wire n_0_353;
   wire n_0_14_0;
   wire n_0_14_1;
   wire n_0_14_2;
   wire n_0_14_3;
   wire n_0_14_4;
   wire n_0_14_5;
   wire n_0_14_6;
   wire n_0_14_7;
   wire n_0_14_8;
   wire n_0_14_9;
   wire n_0_14_10;
   wire n_0_354;
   wire n_0_15_0;
   wire n_0_15_1;
   wire n_0_15_2;
   wire n_0_15_3;
   wire n_0_15_4;
   wire n_0_15_5;
   wire n_0_15_6;
   wire n_0_15_7;
   wire n_0_15_8;
   wire n_0_15_9;
   wire n_0_15_10;
   wire n_0_355;
   wire n_0_16_0;
   wire n_0_16_1;
   wire n_0_16_2;
   wire n_0_16_3;
   wire n_0_16_4;
   wire n_0_16_5;
   wire n_0_16_6;
   wire n_0_16_7;
   wire n_0_16_8;
   wire n_0_16_9;
   wire n_0_16_10;
   wire n_0_356;
   wire n_0_17_0;
   wire n_0_17_1;
   wire n_0_17_2;
   wire n_0_17_3;
   wire n_0_17_4;
   wire n_0_17_5;
   wire n_0_17_6;
   wire n_0_17_7;
   wire n_0_17_8;
   wire n_0_17_9;
   wire n_0_17_10;
   wire n_0_357;
   wire n_0_19_0;
   wire n_0_19_1;
   wire n_0_19_2;
   wire n_0_19_3;
   wire n_0_19_4;
   wire n_0_19_5;
   wire n_0_19_6;
   wire n_0_19_7;
   wire n_0_19_8;
   wire n_0_19_9;
   wire n_0_19_10;
   wire n_0_358;
   wire n_0_21_0;
   wire n_0_21_1;
   wire n_0_21_2;
   wire n_0_21_3;
   wire n_0_21_4;
   wire n_0_359;
   wire n_0_26_2;
   wire n_0_26_3;
   wire n_0_26_5;
   wire n_0_26_6;
   wire n_0_26_7;
   wire n_0_26_8;
   wire n_0_26_9;
   wire n_0_26_10;
   wire n_0_26_0;
   wire n_0_26_1;
   wire n_0_26_4;
   wire n_0_364;
   wire n_0_18_1;
   wire n_0_18_0;
   wire n_0_18_3;
   wire n_0_18_4;
   wire n_0_18_5;
   wire n_0_18_2;
   wire n_0_365;
   wire n_0_18_6;
   wire n_0_18_7;
   wire n_0_18_8;
   wire n_0_18_9;
   wire T_OR_X_Enable;
   wire _64data_Enable;
   wire T_Count_Enable;
   wire X_Count_Enable;
   wire Init_Count_Enable;

   assign RAM_Address_B[12] = 1'b0;
   assign RAM_Address_B[11] = 1'b0;
   assign RAM_Address_B[10] = 1'b0;
   assign RAM_Address_B[9] = 1'b0;
   assign RAM_Address_B[8] = 1'b0;
   assign RAM_Address_B[7] = 1'b0;
   assign RAM_Address_B[6] = 1'b0;
   assign RAM_Address_B[5] = 1'b0;
   assign RAM_Address_B[4] = 1'b0;
   assign RAM_Address_B[3] = 1'b0;
   assign RAM_Address_B[2] = 1'b0;
   assign RAM_Address_B[1] = 1'b1;
   assign RAM_Address_B[0] = 1'b0;

   DFF_X1 _64data_Counter_firstBit_Q_reg (.D(n_0_111), .CK(CLK), .Q(
      Partial_Data_Count[0]), .QN());
   DFF_X1 T_OR_X_COUNTER_firstBit_Q_reg (.D(n_0_112), .CK(CLK), .Q(T_OR_X[0]), 
      .QN());
   DFF_X1 X_Counter_firstBit_Q_reg (.D(n_0_113), .CK(CLK), .Q(X_Count[0]), .QN());
   DFF_X1 X_Counter_genblk1_1_counterBits_Q_reg (.D(n_0_114), .CK(CLK), .Q(
      X_Count[1]), .QN());
   DFF_X1 X_Counter_genblk1_2_counterBits_Q_reg (.D(n_0_115), .CK(CLK), .Q(
      X_Count[2]), .QN());
   DFF_X1 X_Counter_genblk1_3_counterBits_Q_reg (.D(n_0_134), .CK(CLK), .Q(
      X_Count[3]), .QN());
   DFF_X1 X_Counter_genblk1_4_counterBits_Q_reg (.D(n_0_135), .CK(CLK), .Q(
      X_Count[4]), .QN());
   DFF_X1 X_Counter_genblk1_5_counterBits_Q_reg (.D(n_0_180), .CK(CLK), .Q(
      X_Count[5]), .QN());
   DFF_X1 X_Counter_genblk1_6_counterBits_Q_reg (.D(n_0_181), .CK(CLK), .Q(
      X_Count[6]), .QN());
   DFF_X1 X_Counter_genblk1_7_counterBits_Q_reg (.D(n_0_182), .CK(CLK), .Q(
      X_Count[7]), .QN());
   DFF_X2 T_Counter_firstBit_Q_reg (.D(n_0_184), .CK(CLK), .Q(T_Count[0]), .QN());
   DFF_X2 T_Counter_genblk1_1_counterBits_Q_reg (.D(n_0_185), .CK(CLK), .Q(
      T_Count[1]), .QN());
   DFF_X1 T_Counter_genblk1_2_counterBits_Q_reg (.D(n_0_186), .CK(CLK), .Q(
      T_Count[2]), .QN());
   DFF_X1 T_Counter_genblk1_3_counterBits_Q_reg (.D(n_0_187), .CK(CLK), .Q(
      T_Count[3]), .QN());
   DFF_X1 T_Counter_genblk1_4_counterBits_Q_reg (.D(n_0_188), .CK(CLK), .Q(
      T_Count[4]), .QN());
   DFF_X1 T_Counter_genblk1_5_counterBits_Q_reg (.D(n_0_189), .CK(CLK), .Q(
      T_Count[5]), .QN());
   DFF_X1 T_Counter_genblk1_6_counterBits_Q_reg (.D(n_0_190), .CK(CLK), .Q(
      T_Count[6]), .QN());
   DFF_X1 T_Counter_genblk1_7_counterBits_Q_reg (.D(n_0_242), .CK(CLK), .Q(
      T_Count[7]), .QN());
   DFF_X1 Init_Counter_firstBit_Q_reg (.D(n_0_243), .CK(CLK), .Q(Init_Count[0]), 
      .QN());
   DFF_X1 Init_Counter_genblk1_1_counterBits_Q_reg (.D(n_0_308), .CK(CLK), 
      .Q(Init_Count[1]), .QN());
   datapath i_0_2 (.num_of_X(num_of_X), .p_0({n_0_63, n_0_62, n_0_61, n_0_60, 
      n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, 
      n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, 
      n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, 
      n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, 
      n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, 
      n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, 
      n_0_4, n_0_3, n_0_2, n_0_1, uc_0}));
   datapath__0_19 i_0_0 (.num_of_T(num_of_T), .p_0({n_0_133, n_0_132, n_0_131, 
      n_0_130, n_0_129, n_0_128, n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, 
      n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_108, 
      n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, 
      n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, 
      n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, 
      n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, 
      n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, 
      uc_1}));
   DFF_X1 \CPU_Bus_reg[31]  (.D(n_0_339), .CK(CLK), .Q(CPU_Bus[31]), .QN());
   DFF_X1 \CPU_Bus_reg[30]  (.D(n_0_338), .CK(CLK), .Q(CPU_Bus[30]), .QN());
   DFF_X1 \CPU_Bus_reg[29]  (.D(n_0_337), .CK(CLK), .Q(CPU_Bus[29]), .QN());
   DFF_X1 \CPU_Bus_reg[28]  (.D(n_0_336), .CK(CLK), .Q(CPU_Bus[28]), .QN());
   DFF_X1 \CPU_Bus_reg[27]  (.D(n_0_335), .CK(CLK), .Q(CPU_Bus[27]), .QN());
   DFF_X1 \CPU_Bus_reg[26]  (.D(n_0_334), .CK(CLK), .Q(CPU_Bus[26]), .QN());
   DFF_X1 \CPU_Bus_reg[25]  (.D(n_0_333), .CK(CLK), .Q(CPU_Bus[25]), .QN());
   DFF_X1 \CPU_Bus_reg[24]  (.D(n_0_332), .CK(CLK), .Q(CPU_Bus[24]), .QN());
   DFF_X1 \CPU_Bus_reg[23]  (.D(n_0_331), .CK(CLK), .Q(CPU_Bus[23]), .QN());
   DFF_X1 \CPU_Bus_reg[22]  (.D(n_0_330), .CK(CLK), .Q(CPU_Bus[22]), .QN());
   DFF_X1 \CPU_Bus_reg[21]  (.D(n_0_329), .CK(CLK), .Q(CPU_Bus[21]), .QN());
   DFF_X1 \CPU_Bus_reg[20]  (.D(n_0_328), .CK(CLK), .Q(CPU_Bus[20]), .QN());
   DFF_X1 \CPU_Bus_reg[19]  (.D(n_0_327), .CK(CLK), .Q(CPU_Bus[19]), .QN());
   DFF_X1 \CPU_Bus_reg[18]  (.D(n_0_326), .CK(CLK), .Q(CPU_Bus[18]), .QN());
   DFF_X1 \CPU_Bus_reg[17]  (.D(n_0_325), .CK(CLK), .Q(CPU_Bus[17]), .QN());
   DFF_X1 \CPU_Bus_reg[16]  (.D(n_0_324), .CK(CLK), .Q(CPU_Bus[16]), .QN());
   DFF_X1 \CPU_Bus_reg[15]  (.D(n_0_323), .CK(CLK), .Q(CPU_Bus[15]), .QN());
   DFF_X1 \CPU_Bus_reg[14]  (.D(n_0_322), .CK(CLK), .Q(CPU_Bus[14]), .QN());
   DFF_X1 \CPU_Bus_reg[13]  (.D(n_0_321), .CK(CLK), .Q(CPU_Bus[13]), .QN());
   DFF_X1 \CPU_Bus_reg[12]  (.D(n_0_320), .CK(CLK), .Q(CPU_Bus[12]), .QN());
   DFF_X1 \CPU_Bus_reg[11]  (.D(n_0_319), .CK(CLK), .Q(CPU_Bus[11]), .QN());
   DFF_X1 \CPU_Bus_reg[10]  (.D(n_0_318), .CK(CLK), .Q(CPU_Bus[10]), .QN());
   DFF_X1 \CPU_Bus_reg[9]  (.D(n_0_317), .CK(CLK), .Q(CPU_Bus[9]), .QN());
   DFF_X1 \CPU_Bus_reg[8]  (.D(n_0_316), .CK(CLK), .Q(CPU_Bus[8]), .QN());
   DFF_X1 \CPU_Bus_reg[7]  (.D(n_0_315), .CK(CLK), .Q(CPU_Bus[7]), .QN());
   DFF_X1 \CPU_Bus_reg[6]  (.D(n_0_314), .CK(CLK), .Q(CPU_Bus[6]), .QN());
   DFF_X1 \CPU_Bus_reg[5]  (.D(n_0_313), .CK(CLK), .Q(CPU_Bus[5]), .QN());
   DFF_X1 \CPU_Bus_reg[4]  (.D(n_0_312), .CK(CLK), .Q(CPU_Bus[4]), .QN());
   DFF_X1 \CPU_Bus_reg[3]  (.D(n_0_311), .CK(CLK), .Q(CPU_Bus[3]), .QN());
   DFF_X1 \CPU_Bus_reg[2]  (.D(n_0_310), .CK(CLK), .Q(CPU_Bus[2]), .QN());
   DFF_X1 \CPU_Bus_reg[1]  (.D(n_0_309), .CK(CLK), .Q(CPU_Bus[1]), .QN());
   DFF_X1 \CPU_Bus_reg[0]  (.D(n_0_307), .CK(CLK), .Q(CPU_Bus[0]), .QN());
   DFF_X1 \num_of_T_reg[63]  (.D(n_0_306), .CK(n_0_0), .Q(num_of_T[63]), .QN());
   DFF_X1 \num_of_T_reg[62]  (.D(n_0_305), .CK(n_0_0), .Q(num_of_T[62]), .QN());
   DFF_X1 \num_of_T_reg[61]  (.D(n_0_304), .CK(n_0_0), .Q(num_of_T[61]), .QN());
   DFF_X1 \num_of_T_reg[60]  (.D(n_0_303), .CK(n_0_0), .Q(num_of_T[60]), .QN());
   DFF_X1 \num_of_T_reg[59]  (.D(n_0_302), .CK(n_0_0), .Q(num_of_T[59]), .QN());
   DFF_X1 \num_of_T_reg[58]  (.D(n_0_301), .CK(n_0_0), .Q(num_of_T[58]), .QN());
   DFF_X1 \num_of_T_reg[57]  (.D(n_0_300), .CK(n_0_0), .Q(num_of_T[57]), .QN());
   DFF_X1 \num_of_T_reg[56]  (.D(n_0_299), .CK(n_0_0), .Q(num_of_T[56]), .QN());
   DFF_X1 \num_of_T_reg[55]  (.D(n_0_298), .CK(n_0_0), .Q(num_of_T[55]), .QN());
   DFF_X1 \num_of_T_reg[54]  (.D(n_0_297), .CK(n_0_0), .Q(num_of_T[54]), .QN());
   DFF_X1 \num_of_T_reg[53]  (.D(n_0_296), .CK(n_0_0), .Q(num_of_T[53]), .QN());
   DFF_X1 \num_of_T_reg[52]  (.D(n_0_295), .CK(n_0_0), .Q(num_of_T[52]), .QN());
   DFF_X1 \num_of_T_reg[51]  (.D(n_0_294), .CK(n_0_0), .Q(num_of_T[51]), .QN());
   DFF_X1 \num_of_T_reg[50]  (.D(n_0_293), .CK(n_0_0), .Q(num_of_T[50]), .QN());
   DFF_X1 \num_of_T_reg[49]  (.D(n_0_292), .CK(n_0_0), .Q(num_of_T[49]), .QN());
   DFF_X1 \num_of_T_reg[48]  (.D(n_0_291), .CK(n_0_0), .Q(num_of_T[48]), .QN());
   DFF_X1 \num_of_T_reg[47]  (.D(n_0_290), .CK(n_0_0), .Q(num_of_T[47]), .QN());
   DFF_X1 \num_of_T_reg[46]  (.D(n_0_289), .CK(n_0_0), .Q(num_of_T[46]), .QN());
   DFF_X1 \num_of_T_reg[45]  (.D(n_0_288), .CK(n_0_0), .Q(num_of_T[45]), .QN());
   DFF_X1 \num_of_T_reg[44]  (.D(n_0_287), .CK(n_0_0), .Q(num_of_T[44]), .QN());
   DFF_X1 \num_of_T_reg[43]  (.D(n_0_286), .CK(n_0_0), .Q(num_of_T[43]), .QN());
   DFF_X1 \num_of_T_reg[42]  (.D(n_0_285), .CK(n_0_0), .Q(num_of_T[42]), .QN());
   DFF_X1 \num_of_T_reg[41]  (.D(n_0_284), .CK(n_0_0), .Q(num_of_T[41]), .QN());
   DFF_X1 \num_of_T_reg[40]  (.D(n_0_283), .CK(n_0_0), .Q(num_of_T[40]), .QN());
   DFF_X1 \num_of_T_reg[39]  (.D(n_0_282), .CK(n_0_0), .Q(num_of_T[39]), .QN());
   DFF_X1 \num_of_T_reg[38]  (.D(n_0_281), .CK(n_0_0), .Q(num_of_T[38]), .QN());
   DFF_X1 \num_of_T_reg[37]  (.D(n_0_280), .CK(n_0_0), .Q(num_of_T[37]), .QN());
   DFF_X1 \num_of_T_reg[36]  (.D(n_0_279), .CK(n_0_0), .Q(num_of_T[36]), .QN());
   DFF_X1 \num_of_T_reg[35]  (.D(n_0_278), .CK(n_0_0), .Q(num_of_T[35]), .QN());
   DFF_X1 \num_of_T_reg[34]  (.D(n_0_277), .CK(n_0_0), .Q(num_of_T[34]), .QN());
   DFF_X1 \num_of_T_reg[33]  (.D(n_0_276), .CK(n_0_0), .Q(num_of_T[33]), .QN());
   DFF_X1 \num_of_T_reg[32]  (.D(n_0_275), .CK(n_0_0), .Q(num_of_T[32]), .QN());
   DFF_X1 \num_of_T_reg[31]  (.D(n_0_274), .CK(n_0_0), .Q(num_of_T[31]), .QN());
   DFF_X1 \num_of_T_reg[30]  (.D(n_0_273), .CK(n_0_0), .Q(num_of_T[30]), .QN());
   DFF_X1 \num_of_T_reg[29]  (.D(n_0_272), .CK(n_0_0), .Q(num_of_T[29]), .QN());
   DFF_X1 \num_of_T_reg[28]  (.D(n_0_271), .CK(n_0_0), .Q(num_of_T[28]), .QN());
   DFF_X1 \num_of_T_reg[27]  (.D(n_0_270), .CK(n_0_0), .Q(num_of_T[27]), .QN());
   DFF_X1 \num_of_T_reg[26]  (.D(n_0_269), .CK(n_0_0), .Q(num_of_T[26]), .QN());
   DFF_X1 \num_of_T_reg[25]  (.D(n_0_268), .CK(n_0_0), .Q(num_of_T[25]), .QN());
   DFF_X1 \num_of_T_reg[24]  (.D(n_0_267), .CK(n_0_0), .Q(num_of_T[24]), .QN());
   DFF_X1 \num_of_T_reg[23]  (.D(n_0_266), .CK(n_0_0), .Q(num_of_T[23]), .QN());
   DFF_X1 \num_of_T_reg[22]  (.D(n_0_265), .CK(n_0_0), .Q(num_of_T[22]), .QN());
   DFF_X1 \num_of_T_reg[21]  (.D(n_0_264), .CK(n_0_0), .Q(num_of_T[21]), .QN());
   DFF_X1 \num_of_T_reg[20]  (.D(n_0_263), .CK(n_0_0), .Q(num_of_T[20]), .QN());
   DFF_X1 \num_of_T_reg[19]  (.D(n_0_262), .CK(n_0_0), .Q(num_of_T[19]), .QN());
   DFF_X1 \num_of_T_reg[18]  (.D(n_0_261), .CK(n_0_0), .Q(num_of_T[18]), .QN());
   DFF_X1 \num_of_T_reg[17]  (.D(n_0_260), .CK(n_0_0), .Q(num_of_T[17]), .QN());
   DFF_X1 \num_of_T_reg[16]  (.D(n_0_259), .CK(n_0_0), .Q(num_of_T[16]), .QN());
   DFF_X1 \num_of_T_reg[15]  (.D(n_0_258), .CK(n_0_0), .Q(num_of_T[15]), .QN());
   DFF_X1 \num_of_T_reg[14]  (.D(n_0_257), .CK(n_0_0), .Q(num_of_T[14]), .QN());
   DFF_X1 \num_of_T_reg[13]  (.D(n_0_256), .CK(n_0_0), .Q(num_of_T[13]), .QN());
   DFF_X1 \num_of_T_reg[12]  (.D(n_0_255), .CK(n_0_0), .Q(num_of_T[12]), .QN());
   DFF_X1 \num_of_T_reg[11]  (.D(n_0_254), .CK(n_0_0), .Q(num_of_T[11]), .QN());
   DFF_X1 \num_of_T_reg[10]  (.D(n_0_253), .CK(n_0_0), .Q(num_of_T[10]), .QN());
   DFF_X1 \num_of_T_reg[9]  (.D(n_0_252), .CK(n_0_0), .Q(num_of_T[9]), .QN());
   DFF_X1 \num_of_T_reg[8]  (.D(n_0_251), .CK(n_0_0), .Q(num_of_T[8]), .QN());
   DFF_X1 \num_of_T_reg[7]  (.D(n_0_250), .CK(n_0_0), .Q(num_of_T[7]), .QN());
   DFF_X1 \num_of_T_reg[6]  (.D(n_0_249), .CK(n_0_0), .Q(num_of_T[6]), .QN());
   DFF_X1 \num_of_T_reg[5]  (.D(n_0_248), .CK(n_0_0), .Q(num_of_T[5]), .QN());
   DFF_X1 \num_of_T_reg[4]  (.D(n_0_247), .CK(n_0_0), .Q(num_of_T[4]), .QN());
   DFF_X1 \num_of_T_reg[3]  (.D(n_0_246), .CK(n_0_0), .Q(num_of_T[3]), .QN());
   DFF_X1 \num_of_T_reg[2]  (.D(n_0_245), .CK(n_0_0), .Q(num_of_T[2]), .QN());
   DFF_X1 \num_of_T_reg[1]  (.D(n_0_244), .CK(n_0_0), .Q(num_of_T[1]), .QN());
   DFF_X1 \num_of_T_reg[0]  (.D(n_0_241), .CK(n_0_0), .Q(num_of_T[0]), .QN());
   DFF_X1 \num_of_X_reg[63]  (.D(n_0_239), .CK(n_0_0), .Q(num_of_X[63]), .QN());
   DFF_X1 \num_of_X_reg[62]  (.D(n_0_238), .CK(n_0_0), .Q(num_of_X[62]), .QN());
   DFF_X1 \num_of_X_reg[61]  (.D(n_0_237), .CK(n_0_0), .Q(num_of_X[61]), .QN());
   DFF_X1 \num_of_X_reg[60]  (.D(n_0_236), .CK(n_0_0), .Q(num_of_X[60]), .QN());
   DFF_X1 \num_of_X_reg[59]  (.D(n_0_235), .CK(n_0_0), .Q(num_of_X[59]), .QN());
   DFF_X1 \num_of_X_reg[58]  (.D(n_0_234), .CK(n_0_0), .Q(num_of_X[58]), .QN());
   DFF_X1 \num_of_X_reg[57]  (.D(n_0_233), .CK(n_0_0), .Q(num_of_X[57]), .QN());
   DFF_X1 \num_of_X_reg[56]  (.D(n_0_232), .CK(n_0_0), .Q(num_of_X[56]), .QN());
   DFF_X1 \num_of_X_reg[55]  (.D(n_0_231), .CK(n_0_0), .Q(num_of_X[55]), .QN());
   DFF_X1 \num_of_X_reg[54]  (.D(n_0_230), .CK(n_0_0), .Q(num_of_X[54]), .QN());
   DFF_X1 \num_of_X_reg[53]  (.D(n_0_229), .CK(n_0_0), .Q(num_of_X[53]), .QN());
   DFF_X1 \num_of_X_reg[52]  (.D(n_0_228), .CK(n_0_0), .Q(num_of_X[52]), .QN());
   DFF_X1 \num_of_X_reg[51]  (.D(n_0_227), .CK(n_0_0), .Q(num_of_X[51]), .QN());
   DFF_X1 \num_of_X_reg[50]  (.D(n_0_226), .CK(n_0_0), .Q(num_of_X[50]), .QN());
   DFF_X1 \num_of_X_reg[49]  (.D(n_0_225), .CK(n_0_0), .Q(num_of_X[49]), .QN());
   DFF_X1 \num_of_X_reg[48]  (.D(n_0_224), .CK(n_0_0), .Q(num_of_X[48]), .QN());
   DFF_X1 \num_of_X_reg[47]  (.D(n_0_223), .CK(n_0_0), .Q(num_of_X[47]), .QN());
   DFF_X1 \num_of_X_reg[46]  (.D(n_0_222), .CK(n_0_0), .Q(num_of_X[46]), .QN());
   DFF_X1 \num_of_X_reg[45]  (.D(n_0_221), .CK(n_0_0), .Q(num_of_X[45]), .QN());
   DFF_X1 \num_of_X_reg[44]  (.D(n_0_220), .CK(n_0_0), .Q(num_of_X[44]), .QN());
   DFF_X1 \num_of_X_reg[43]  (.D(n_0_219), .CK(n_0_0), .Q(num_of_X[43]), .QN());
   DFF_X1 \num_of_X_reg[42]  (.D(n_0_218), .CK(n_0_0), .Q(num_of_X[42]), .QN());
   DFF_X1 \num_of_X_reg[41]  (.D(n_0_217), .CK(n_0_0), .Q(num_of_X[41]), .QN());
   DFF_X1 \num_of_X_reg[40]  (.D(n_0_216), .CK(n_0_0), .Q(num_of_X[40]), .QN());
   DFF_X1 \num_of_X_reg[39]  (.D(n_0_215), .CK(n_0_0), .Q(num_of_X[39]), .QN());
   DFF_X1 \num_of_X_reg[38]  (.D(n_0_214), .CK(n_0_0), .Q(num_of_X[38]), .QN());
   DFF_X1 \num_of_X_reg[37]  (.D(n_0_213), .CK(n_0_0), .Q(num_of_X[37]), .QN());
   DFF_X1 \num_of_X_reg[36]  (.D(n_0_212), .CK(n_0_0), .Q(num_of_X[36]), .QN());
   DFF_X1 \num_of_X_reg[35]  (.D(n_0_211), .CK(n_0_0), .Q(num_of_X[35]), .QN());
   DFF_X1 \num_of_X_reg[34]  (.D(n_0_210), .CK(n_0_0), .Q(num_of_X[34]), .QN());
   DFF_X1 \num_of_X_reg[33]  (.D(n_0_209), .CK(n_0_0), .Q(num_of_X[33]), .QN());
   DFF_X1 \num_of_X_reg[32]  (.D(n_0_208), .CK(n_0_0), .Q(num_of_X[32]), .QN());
   DFF_X1 \num_of_X_reg[31]  (.D(n_0_207), .CK(n_0_0), .Q(num_of_X[31]), .QN());
   DFF_X1 \num_of_X_reg[30]  (.D(n_0_206), .CK(n_0_0), .Q(num_of_X[30]), .QN());
   DFF_X1 \num_of_X_reg[29]  (.D(n_0_205), .CK(n_0_0), .Q(num_of_X[29]), .QN());
   DFF_X1 \num_of_X_reg[28]  (.D(n_0_204), .CK(n_0_0), .Q(num_of_X[28]), .QN());
   DFF_X1 \num_of_X_reg[27]  (.D(n_0_203), .CK(n_0_0), .Q(num_of_X[27]), .QN());
   DFF_X1 \num_of_X_reg[26]  (.D(n_0_202), .CK(n_0_0), .Q(num_of_X[26]), .QN());
   DFF_X1 \num_of_X_reg[25]  (.D(n_0_201), .CK(n_0_0), .Q(num_of_X[25]), .QN());
   DFF_X1 \num_of_X_reg[24]  (.D(n_0_200), .CK(n_0_0), .Q(num_of_X[24]), .QN());
   DFF_X1 \num_of_X_reg[23]  (.D(n_0_199), .CK(n_0_0), .Q(num_of_X[23]), .QN());
   DFF_X1 \num_of_X_reg[22]  (.D(n_0_198), .CK(n_0_0), .Q(num_of_X[22]), .QN());
   DFF_X1 \num_of_X_reg[21]  (.D(n_0_197), .CK(n_0_0), .Q(num_of_X[21]), .QN());
   DFF_X1 \num_of_X_reg[20]  (.D(n_0_196), .CK(n_0_0), .Q(num_of_X[20]), .QN());
   DFF_X1 \num_of_X_reg[19]  (.D(n_0_195), .CK(n_0_0), .Q(num_of_X[19]), .QN());
   DFF_X1 \num_of_X_reg[18]  (.D(n_0_194), .CK(n_0_0), .Q(num_of_X[18]), .QN());
   DFF_X1 \num_of_X_reg[17]  (.D(n_0_193), .CK(n_0_0), .Q(num_of_X[17]), .QN());
   DFF_X1 \num_of_X_reg[16]  (.D(n_0_192), .CK(n_0_0), .Q(num_of_X[16]), .QN());
   DFF_X1 \num_of_X_reg[15]  (.D(n_0_191), .CK(n_0_0), .Q(num_of_X[15]), .QN());
   DFF_X1 \num_of_X_reg[14]  (.D(n_0_183), .CK(n_0_0), .Q(num_of_X[14]), .QN());
   DFF_X1 \num_of_X_reg[13]  (.D(n_0_179), .CK(n_0_0), .Q(num_of_X[13]), .QN());
   DFF_X1 \num_of_X_reg[12]  (.D(n_0_178), .CK(n_0_0), .Q(num_of_X[12]), .QN());
   DFF_X1 \num_of_X_reg[11]  (.D(n_0_177), .CK(n_0_0), .Q(num_of_X[11]), .QN());
   DFF_X1 \num_of_X_reg[10]  (.D(n_0_176), .CK(n_0_0), .Q(num_of_X[10]), .QN());
   DFF_X1 \num_of_X_reg[9]  (.D(n_0_175), .CK(n_0_0), .Q(num_of_X[9]), .QN());
   DFF_X1 \num_of_X_reg[8]  (.D(n_0_174), .CK(n_0_0), .Q(num_of_X[8]), .QN());
   DFF_X1 \num_of_X_reg[7]  (.D(n_0_173), .CK(n_0_0), .Q(num_of_X[7]), .QN());
   DFF_X1 \num_of_X_reg[6]  (.D(n_0_172), .CK(n_0_0), .Q(num_of_X[6]), .QN());
   DFF_X1 \num_of_X_reg[5]  (.D(n_0_171), .CK(n_0_0), .Q(num_of_X[5]), .QN());
   DFF_X1 \num_of_X_reg[4]  (.D(n_0_170), .CK(n_0_0), .Q(num_of_X[4]), .QN());
   DFF_X2 \num_of_X_reg[2]  (.D(n_0_168), .CK(n_0_0), .Q(num_of_X[2]), .QN());
   DFF_X1 \num_of_X_reg[1]  (.D(n_0_167), .CK(n_0_0), .Q(num_of_X[1]), .QN());
   DFF_X1 \num_of_X_reg[0]  (.D(n_0_166), .CK(n_0_0), .Q(num_of_X[0]), .QN());
   CLKGATETST_X1 clk_gate_num_of_T_reg (.CK(CLK), .E(n_0_240), .SE(1'b0), 
      .GCK(n_0_0));
   AND2_X1 i_0_22_0 (.A1(n_0_139), .A2(RAM_Data_B[0]), .ZN(n_0_166));
   AND2_X1 i_0_22_1 (.A1(n_0_139), .A2(RAM_Data_B[1]), .ZN(n_0_167));
   AND2_X1 i_0_22_2 (.A1(n_0_139), .A2(RAM_Data_B[2]), .ZN(n_0_168));
   AND2_X1 i_0_22_3 (.A1(n_0_139), .A2(RAM_Data_B[3]), .ZN(n_0_169));
   AND2_X1 i_0_22_4 (.A1(n_0_139), .A2(RAM_Data_B[4]), .ZN(n_0_170));
   AND2_X1 i_0_22_5 (.A1(n_0_139), .A2(RAM_Data_B[5]), .ZN(n_0_171));
   AND2_X1 i_0_22_6 (.A1(n_0_139), .A2(RAM_Data_B[6]), .ZN(n_0_172));
   AND2_X1 i_0_22_7 (.A1(n_0_139), .A2(RAM_Data_B[7]), .ZN(n_0_173));
   AND2_X1 i_0_22_8 (.A1(n_0_139), .A2(RAM_Data_B[8]), .ZN(n_0_174));
   AND2_X1 i_0_22_9 (.A1(n_0_139), .A2(RAM_Data_B[9]), .ZN(n_0_175));
   AND2_X1 i_0_22_10 (.A1(n_0_139), .A2(RAM_Data_B[10]), .ZN(n_0_176));
   AND2_X1 i_0_22_11 (.A1(n_0_139), .A2(RAM_Data_B[11]), .ZN(n_0_177));
   AND2_X1 i_0_22_12 (.A1(n_0_139), .A2(RAM_Data_B[12]), .ZN(n_0_178));
   AND2_X1 i_0_22_13 (.A1(n_0_139), .A2(RAM_Data_B[13]), .ZN(n_0_179));
   AND2_X1 i_0_22_14 (.A1(n_0_139), .A2(RAM_Data_B[14]), .ZN(n_0_183));
   AND2_X1 i_0_22_15 (.A1(n_0_139), .A2(RAM_Data_B[15]), .ZN(n_0_191));
   AND2_X1 i_0_22_16 (.A1(n_0_139), .A2(RAM_Data_B[16]), .ZN(n_0_192));
   AND2_X1 i_0_22_17 (.A1(n_0_139), .A2(RAM_Data_B[17]), .ZN(n_0_193));
   AND2_X1 i_0_22_18 (.A1(n_0_139), .A2(RAM_Data_B[18]), .ZN(n_0_194));
   AND2_X1 i_0_22_19 (.A1(n_0_139), .A2(RAM_Data_B[19]), .ZN(n_0_195));
   AND2_X1 i_0_22_20 (.A1(n_0_139), .A2(RAM_Data_B[20]), .ZN(n_0_196));
   AND2_X1 i_0_22_21 (.A1(n_0_139), .A2(RAM_Data_B[21]), .ZN(n_0_197));
   AND2_X1 i_0_22_22 (.A1(n_0_139), .A2(RAM_Data_B[22]), .ZN(n_0_198));
   AND2_X1 i_0_22_23 (.A1(n_0_139), .A2(RAM_Data_B[23]), .ZN(n_0_199));
   AND2_X1 i_0_22_24 (.A1(n_0_139), .A2(RAM_Data_B[24]), .ZN(n_0_200));
   AND2_X1 i_0_22_25 (.A1(n_0_139), .A2(RAM_Data_B[25]), .ZN(n_0_201));
   AND2_X1 i_0_22_26 (.A1(n_0_139), .A2(RAM_Data_B[26]), .ZN(n_0_202));
   AND2_X1 i_0_22_27 (.A1(n_0_139), .A2(RAM_Data_B[27]), .ZN(n_0_203));
   AND2_X1 i_0_22_28 (.A1(n_0_139), .A2(RAM_Data_B[28]), .ZN(n_0_204));
   AND2_X1 i_0_22_29 (.A1(n_0_139), .A2(RAM_Data_B[29]), .ZN(n_0_205));
   AND2_X1 i_0_22_30 (.A1(n_0_139), .A2(RAM_Data_B[30]), .ZN(n_0_206));
   AND2_X1 i_0_22_31 (.A1(n_0_139), .A2(RAM_Data_B[31]), .ZN(n_0_207));
   AND2_X1 i_0_22_32 (.A1(n_0_139), .A2(RAM_Data_B[32]), .ZN(n_0_208));
   AND2_X1 i_0_22_33 (.A1(n_0_139), .A2(RAM_Data_B[33]), .ZN(n_0_209));
   AND2_X1 i_0_22_34 (.A1(n_0_139), .A2(RAM_Data_B[34]), .ZN(n_0_210));
   AND2_X1 i_0_22_35 (.A1(n_0_139), .A2(RAM_Data_B[35]), .ZN(n_0_211));
   AND2_X1 i_0_22_36 (.A1(n_0_139), .A2(RAM_Data_B[36]), .ZN(n_0_212));
   AND2_X1 i_0_22_37 (.A1(n_0_139), .A2(RAM_Data_B[37]), .ZN(n_0_213));
   AND2_X1 i_0_22_38 (.A1(n_0_139), .A2(RAM_Data_B[38]), .ZN(n_0_214));
   AND2_X1 i_0_22_39 (.A1(n_0_139), .A2(RAM_Data_B[39]), .ZN(n_0_215));
   AND2_X1 i_0_22_40 (.A1(n_0_139), .A2(RAM_Data_B[40]), .ZN(n_0_216));
   AND2_X1 i_0_22_41 (.A1(n_0_139), .A2(RAM_Data_B[41]), .ZN(n_0_217));
   AND2_X1 i_0_22_42 (.A1(n_0_139), .A2(RAM_Data_B[42]), .ZN(n_0_218));
   AND2_X1 i_0_22_43 (.A1(n_0_139), .A2(RAM_Data_B[43]), .ZN(n_0_219));
   AND2_X1 i_0_22_44 (.A1(n_0_139), .A2(RAM_Data_B[44]), .ZN(n_0_220));
   AND2_X1 i_0_22_45 (.A1(n_0_139), .A2(RAM_Data_B[45]), .ZN(n_0_221));
   AND2_X1 i_0_22_46 (.A1(n_0_139), .A2(RAM_Data_B[46]), .ZN(n_0_222));
   AND2_X1 i_0_22_47 (.A1(n_0_139), .A2(RAM_Data_B[47]), .ZN(n_0_223));
   AND2_X1 i_0_22_48 (.A1(n_0_139), .A2(RAM_Data_B[48]), .ZN(n_0_224));
   AND2_X1 i_0_22_49 (.A1(n_0_139), .A2(RAM_Data_B[49]), .ZN(n_0_225));
   AND2_X1 i_0_22_50 (.A1(n_0_139), .A2(RAM_Data_B[50]), .ZN(n_0_226));
   AND2_X1 i_0_22_51 (.A1(n_0_139), .A2(RAM_Data_B[51]), .ZN(n_0_227));
   AND2_X1 i_0_22_52 (.A1(n_0_139), .A2(RAM_Data_B[52]), .ZN(n_0_228));
   AND2_X1 i_0_22_53 (.A1(n_0_139), .A2(RAM_Data_B[53]), .ZN(n_0_229));
   AND2_X1 i_0_22_54 (.A1(n_0_139), .A2(RAM_Data_B[54]), .ZN(n_0_230));
   AND2_X1 i_0_22_55 (.A1(n_0_139), .A2(RAM_Data_B[55]), .ZN(n_0_231));
   AND2_X1 i_0_22_56 (.A1(n_0_139), .A2(RAM_Data_B[56]), .ZN(n_0_232));
   AND2_X1 i_0_22_57 (.A1(n_0_139), .A2(RAM_Data_B[57]), .ZN(n_0_233));
   AND2_X1 i_0_22_58 (.A1(n_0_139), .A2(RAM_Data_B[58]), .ZN(n_0_234));
   AND2_X1 i_0_22_59 (.A1(n_0_139), .A2(RAM_Data_B[59]), .ZN(n_0_235));
   AND2_X1 i_0_22_60 (.A1(n_0_139), .A2(RAM_Data_B[60]), .ZN(n_0_236));
   AND2_X1 i_0_22_61 (.A1(n_0_139), .A2(RAM_Data_B[61]), .ZN(n_0_237));
   AND2_X1 i_0_22_62 (.A1(n_0_139), .A2(RAM_Data_B[62]), .ZN(n_0_238));
   AND2_X1 i_0_22_63 (.A1(n_0_139), .A2(RAM_Data_B[63]), .ZN(n_0_239));
   OR2_X1 i_0_22_64 (.A1(RST), .A2(n_0_344), .ZN(n_0_240));
   NOR2_X1 i_0_22_65 (.A1(RST), .A2(n_0_22_16), .ZN(n_0_241));
   NOR2_X1 i_0_22_66 (.A1(RST), .A2(n_0_22_17), .ZN(n_0_244));
   NOR2_X1 i_0_22_67 (.A1(RST), .A2(n_0_22_18), .ZN(n_0_245));
   NOR2_X1 i_0_22_68 (.A1(RST), .A2(n_0_22_19), .ZN(n_0_246));
   NOR2_X1 i_0_22_69 (.A1(RST), .A2(n_0_22_20), .ZN(n_0_247));
   NOR2_X1 i_0_22_70 (.A1(RST), .A2(n_0_22_21), .ZN(n_0_248));
   NOR2_X1 i_0_22_71 (.A1(RST), .A2(n_0_22_22), .ZN(n_0_249));
   NOR2_X1 i_0_22_72 (.A1(RST), .A2(n_0_22_23), .ZN(n_0_250));
   NOR2_X1 i_0_22_73 (.A1(RST), .A2(n_0_22_24), .ZN(n_0_251));
   NOR2_X1 i_0_22_74 (.A1(RST), .A2(n_0_22_25), .ZN(n_0_252));
   NOR2_X1 i_0_22_75 (.A1(RST), .A2(n_0_22_26), .ZN(n_0_253));
   NOR2_X1 i_0_22_76 (.A1(RST), .A2(n_0_22_27), .ZN(n_0_254));
   NOR2_X1 i_0_22_77 (.A1(RST), .A2(n_0_22_28), .ZN(n_0_255));
   NOR2_X1 i_0_22_78 (.A1(RST), .A2(n_0_22_29), .ZN(n_0_256));
   NOR2_X1 i_0_22_79 (.A1(RST), .A2(n_0_22_30), .ZN(n_0_257));
   NOR2_X1 i_0_22_80 (.A1(RST), .A2(n_0_22_31), .ZN(n_0_258));
   NOR2_X1 i_0_22_81 (.A1(RST), .A2(n_0_22_32), .ZN(n_0_259));
   NOR2_X1 i_0_22_82 (.A1(RST), .A2(n_0_22_33), .ZN(n_0_260));
   NOR2_X1 i_0_22_83 (.A1(RST), .A2(n_0_22_34), .ZN(n_0_261));
   NOR2_X1 i_0_22_84 (.A1(RST), .A2(n_0_22_35), .ZN(n_0_262));
   NOR2_X1 i_0_22_85 (.A1(RST), .A2(n_0_22_36), .ZN(n_0_263));
   NOR2_X1 i_0_22_86 (.A1(RST), .A2(n_0_22_37), .ZN(n_0_264));
   NOR2_X1 i_0_22_87 (.A1(RST), .A2(n_0_22_38), .ZN(n_0_265));
   NOR2_X1 i_0_22_88 (.A1(RST), .A2(n_0_22_39), .ZN(n_0_266));
   NOR2_X1 i_0_22_89 (.A1(RST), .A2(n_0_22_40), .ZN(n_0_267));
   NOR2_X1 i_0_22_90 (.A1(RST), .A2(n_0_22_41), .ZN(n_0_268));
   NOR2_X1 i_0_22_91 (.A1(RST), .A2(n_0_22_42), .ZN(n_0_269));
   NOR2_X1 i_0_22_92 (.A1(RST), .A2(n_0_22_43), .ZN(n_0_270));
   NOR2_X1 i_0_22_93 (.A1(RST), .A2(n_0_22_44), .ZN(n_0_271));
   NOR2_X1 i_0_22_94 (.A1(RST), .A2(n_0_22_45), .ZN(n_0_272));
   NOR2_X1 i_0_22_95 (.A1(RST), .A2(n_0_22_46), .ZN(n_0_273));
   NOR2_X1 i_0_22_96 (.A1(RST), .A2(n_0_22_47), .ZN(n_0_274));
   NOR2_X1 i_0_22_97 (.A1(RST), .A2(n_0_22_48), .ZN(n_0_275));
   NOR2_X1 i_0_22_98 (.A1(RST), .A2(n_0_22_49), .ZN(n_0_276));
   NOR2_X1 i_0_22_99 (.A1(RST), .A2(n_0_22_50), .ZN(n_0_277));
   NOR2_X1 i_0_22_100 (.A1(RST), .A2(n_0_22_51), .ZN(n_0_278));
   NOR2_X1 i_0_22_101 (.A1(RST), .A2(n_0_22_52), .ZN(n_0_279));
   NOR2_X1 i_0_22_102 (.A1(RST), .A2(n_0_22_53), .ZN(n_0_280));
   NOR2_X1 i_0_22_103 (.A1(RST), .A2(n_0_22_54), .ZN(n_0_281));
   NOR2_X1 i_0_22_104 (.A1(RST), .A2(n_0_22_55), .ZN(n_0_282));
   NOR2_X1 i_0_22_105 (.A1(RST), .A2(n_0_22_56), .ZN(n_0_283));
   NOR2_X1 i_0_22_106 (.A1(RST), .A2(n_0_22_57), .ZN(n_0_284));
   NOR2_X1 i_0_22_107 (.A1(RST), .A2(n_0_22_58), .ZN(n_0_285));
   NOR2_X1 i_0_22_108 (.A1(RST), .A2(n_0_22_59), .ZN(n_0_286));
   NOR2_X1 i_0_22_109 (.A1(RST), .A2(n_0_22_60), .ZN(n_0_287));
   NOR2_X1 i_0_22_110 (.A1(RST), .A2(n_0_22_61), .ZN(n_0_288));
   NOR2_X1 i_0_22_111 (.A1(RST), .A2(n_0_22_62), .ZN(n_0_289));
   NOR2_X1 i_0_22_112 (.A1(RST), .A2(n_0_22_63), .ZN(n_0_290));
   NOR2_X1 i_0_22_113 (.A1(RST), .A2(n_0_22_64), .ZN(n_0_291));
   NOR2_X1 i_0_22_114 (.A1(RST), .A2(n_0_22_65), .ZN(n_0_292));
   NOR2_X1 i_0_22_115 (.A1(RST), .A2(n_0_22_66), .ZN(n_0_293));
   NOR2_X1 i_0_22_116 (.A1(RST), .A2(n_0_22_67), .ZN(n_0_294));
   NOR2_X1 i_0_22_117 (.A1(RST), .A2(n_0_22_68), .ZN(n_0_295));
   NOR2_X1 i_0_22_118 (.A1(RST), .A2(n_0_22_69), .ZN(n_0_296));
   NOR2_X1 i_0_22_119 (.A1(RST), .A2(n_0_22_70), .ZN(n_0_297));
   NOR2_X1 i_0_22_120 (.A1(RST), .A2(n_0_22_71), .ZN(n_0_298));
   NOR2_X1 i_0_22_121 (.A1(RST), .A2(n_0_22_72), .ZN(n_0_299));
   NOR2_X1 i_0_22_122 (.A1(RST), .A2(n_0_22_73), .ZN(n_0_300));
   NOR2_X1 i_0_22_123 (.A1(RST), .A2(n_0_22_74), .ZN(n_0_301));
   NOR2_X1 i_0_22_124 (.A1(RST), .A2(n_0_22_75), .ZN(n_0_302));
   NOR2_X1 i_0_22_125 (.A1(RST), .A2(n_0_22_76), .ZN(n_0_303));
   NOR2_X1 i_0_22_126 (.A1(RST), .A2(n_0_22_77), .ZN(n_0_304));
   NOR2_X1 i_0_22_127 (.A1(RST), .A2(n_0_22_78), .ZN(n_0_305));
   NOR2_X1 i_0_22_128 (.A1(RST), .A2(n_0_22_79), .ZN(n_0_306));
   OAI22_X1 i_0_22_129 (.A1(n_0_22_16), .A2(n_0_22_0), .B1(n_0_22_48), .B2(
      n_0_22_15), .ZN(n_0_307));
   OAI22_X1 i_0_22_130 (.A1(n_0_22_17), .A2(n_0_22_0), .B1(n_0_22_49), .B2(
      n_0_22_15), .ZN(n_0_309));
   OAI22_X1 i_0_22_131 (.A1(n_0_22_18), .A2(n_0_22_0), .B1(n_0_22_50), .B2(
      n_0_22_15), .ZN(n_0_310));
   OAI22_X1 i_0_22_132 (.A1(n_0_22_19), .A2(n_0_22_0), .B1(n_0_22_51), .B2(
      n_0_22_15), .ZN(n_0_311));
   OAI22_X1 i_0_22_133 (.A1(n_0_22_20), .A2(n_0_22_0), .B1(n_0_22_52), .B2(
      n_0_22_15), .ZN(n_0_312));
   OAI22_X1 i_0_22_134 (.A1(n_0_22_21), .A2(n_0_22_0), .B1(n_0_22_53), .B2(
      n_0_22_15), .ZN(n_0_313));
   OAI22_X1 i_0_22_135 (.A1(n_0_22_22), .A2(n_0_22_0), .B1(n_0_22_54), .B2(
      n_0_22_15), .ZN(n_0_314));
   OAI22_X1 i_0_22_136 (.A1(n_0_22_23), .A2(n_0_22_0), .B1(n_0_22_55), .B2(
      n_0_22_15), .ZN(n_0_315));
   OAI22_X1 i_0_22_137 (.A1(n_0_22_24), .A2(n_0_22_0), .B1(n_0_22_56), .B2(
      n_0_22_15), .ZN(n_0_316));
   OAI22_X1 i_0_22_138 (.A1(n_0_22_25), .A2(n_0_22_0), .B1(n_0_22_57), .B2(
      n_0_22_15), .ZN(n_0_317));
   OAI22_X1 i_0_22_139 (.A1(n_0_22_26), .A2(n_0_22_0), .B1(n_0_22_58), .B2(
      n_0_22_15), .ZN(n_0_318));
   OAI22_X1 i_0_22_140 (.A1(n_0_22_27), .A2(n_0_22_0), .B1(n_0_22_59), .B2(
      n_0_22_15), .ZN(n_0_319));
   OAI22_X1 i_0_22_141 (.A1(n_0_22_28), .A2(n_0_22_0), .B1(n_0_22_60), .B2(
      n_0_22_15), .ZN(n_0_320));
   OAI22_X1 i_0_22_142 (.A1(n_0_22_29), .A2(n_0_22_0), .B1(n_0_22_61), .B2(
      n_0_22_15), .ZN(n_0_321));
   OAI22_X1 i_0_22_143 (.A1(n_0_22_30), .A2(n_0_22_0), .B1(n_0_22_62), .B2(
      n_0_22_15), .ZN(n_0_322));
   OAI22_X1 i_0_22_144 (.A1(n_0_22_31), .A2(n_0_22_0), .B1(n_0_22_63), .B2(
      n_0_22_15), .ZN(n_0_323));
   OAI22_X1 i_0_22_145 (.A1(n_0_22_32), .A2(n_0_22_0), .B1(n_0_22_64), .B2(
      n_0_22_15), .ZN(n_0_324));
   OAI22_X1 i_0_22_146 (.A1(n_0_22_33), .A2(n_0_22_0), .B1(n_0_22_65), .B2(
      n_0_22_15), .ZN(n_0_325));
   OAI22_X1 i_0_22_147 (.A1(n_0_22_34), .A2(n_0_22_0), .B1(n_0_22_66), .B2(
      n_0_22_15), .ZN(n_0_326));
   OAI22_X1 i_0_22_148 (.A1(n_0_22_35), .A2(n_0_22_0), .B1(n_0_22_67), .B2(
      n_0_22_15), .ZN(n_0_327));
   OAI22_X1 i_0_22_149 (.A1(n_0_22_36), .A2(n_0_22_0), .B1(n_0_22_68), .B2(
      n_0_22_15), .ZN(n_0_328));
   OAI22_X1 i_0_22_150 (.A1(n_0_22_37), .A2(n_0_22_0), .B1(n_0_22_69), .B2(
      n_0_22_15), .ZN(n_0_329));
   OAI22_X1 i_0_22_151 (.A1(n_0_22_38), .A2(n_0_22_0), .B1(n_0_22_70), .B2(
      n_0_22_15), .ZN(n_0_330));
   OAI22_X1 i_0_22_152 (.A1(n_0_22_39), .A2(n_0_22_0), .B1(n_0_22_71), .B2(
      n_0_22_15), .ZN(n_0_331));
   OAI22_X1 i_0_22_153 (.A1(n_0_22_40), .A2(n_0_22_0), .B1(n_0_22_72), .B2(
      n_0_22_15), .ZN(n_0_332));
   OAI22_X1 i_0_22_154 (.A1(n_0_22_41), .A2(n_0_22_0), .B1(n_0_22_73), .B2(
      n_0_22_15), .ZN(n_0_333));
   OAI22_X1 i_0_22_155 (.A1(n_0_22_42), .A2(n_0_22_0), .B1(n_0_22_74), .B2(
      n_0_22_15), .ZN(n_0_334));
   OAI22_X1 i_0_22_156 (.A1(n_0_22_43), .A2(n_0_22_0), .B1(n_0_22_75), .B2(
      n_0_22_15), .ZN(n_0_335));
   OAI22_X1 i_0_22_157 (.A1(n_0_22_44), .A2(n_0_22_0), .B1(n_0_22_76), .B2(
      n_0_22_15), .ZN(n_0_336));
   OAI22_X1 i_0_22_158 (.A1(n_0_22_45), .A2(n_0_22_0), .B1(n_0_22_77), .B2(
      n_0_22_15), .ZN(n_0_337));
   OAI22_X1 i_0_22_159 (.A1(n_0_22_46), .A2(n_0_22_0), .B1(n_0_22_78), .B2(
      n_0_22_15), .ZN(n_0_338));
   OAI22_X1 i_0_22_160 (.A1(n_0_22_47), .A2(n_0_22_0), .B1(n_0_22_79), .B2(
      n_0_22_15), .ZN(n_0_339));
   NOR2_X1 i_0_22_161 (.A1(n_0_361), .A2(n_0_360), .ZN(n_0_22_0));
   NOR2_X1 i_0_22_162 (.A1(RST), .A2(Init_Count[1]), .ZN(
      Init_Counter_genblk1_1_counterBits_n_4));
   AOI21_X1 i_0_22_163 (.A(Init_Counter_firstBit_n_4), .B1(n_0_139), .B2(
      n_0_22_80), .ZN(Init_Counter_genblk1_1_counterBits_n_2));
   NOR2_X1 i_0_22_164 (.A1(RST), .A2(Init_Count[0]), .ZN(
      Init_Counter_firstBit_n_4));
   NAND2_X1 i_0_22_165 (.A1(n_0_139), .A2(n_0_22_80), .ZN(
      Init_Counter_firstBit_n_2));
   NOR2_X1 i_0_22_166 (.A1(T_Count[7]), .A2(n_0_22_6), .ZN(
      T_Counter_genblk1_7_counterBits_n_4));
   AOI21_X1 i_0_22_167 (.A(T_Counter_genblk1_6_counterBits_n_4), .B1(n_0_22_7), 
      .B2(n_0_22_1), .ZN(T_Counter_genblk1_7_counterBits_n_2));
   NOR2_X1 i_0_22_168 (.A1(T_Count[6]), .A2(n_0_22_6), .ZN(
      T_Counter_genblk1_6_counterBits_n_4));
   NAND2_X1 i_0_22_169 (.A1(n_0_22_7), .A2(n_0_22_1), .ZN(
      T_Counter_genblk1_6_counterBits_n_2));
   NAND3_X1 i_0_22_170 (.A1(T_Count[4]), .A2(n_0_22_3), .A3(T_Count[5]), 
      .ZN(n_0_22_1));
   NOR2_X1 i_0_22_171 (.A1(T_Count[5]), .A2(n_0_22_6), .ZN(
      T_Counter_genblk1_5_counterBits_n_4));
   NOR2_X1 i_0_22_172 (.A1(n_0_22_2), .A2(T_Counter_genblk1_4_counterBits_n_4), 
      .ZN(T_Counter_genblk1_5_counterBits_n_2));
   NOR2_X1 i_0_22_173 (.A1(T_Count[4]), .A2(n_0_22_6), .ZN(
      T_Counter_genblk1_4_counterBits_n_4));
   INV_X1 i_0_22_174 (.A(n_0_22_2), .ZN(T_Counter_genblk1_4_counterBits_n_2));
   NOR2_X1 i_0_22_175 (.A1(n_0_22_6), .A2(n_0_22_3), .ZN(n_0_22_2));
   NOR2_X1 i_0_22_176 (.A1(n_0_22_81), .A2(n_0_22_4), .ZN(n_0_22_3));
   NOR2_X1 i_0_22_177 (.A1(T_Count[3]), .A2(n_0_22_6), .ZN(
      T_Counter_genblk1_3_counterBits_n_4));
   NAND2_X1 i_0_22_178 (.A1(n_0_22_7), .A2(n_0_22_4), .ZN(
      T_Counter_genblk1_3_counterBits_n_2));
   NAND4_X1 i_0_22_179 (.A1(T_Count_Enable), .A2(T_Count[1]), .A3(T_Count[0]), 
      .A4(T_Count[2]), .ZN(n_0_22_4));
   NOR2_X1 i_0_22_180 (.A1(T_Count[2]), .A2(n_0_22_6), .ZN(
      T_Counter_genblk1_2_counterBits_n_4));
   NAND2_X1 i_0_22_181 (.A1(n_0_22_7), .A2(n_0_22_5), .ZN(
      T_Counter_genblk1_2_counterBits_n_2));
   NAND3_X1 i_0_22_182 (.A1(T_Count_Enable), .A2(T_Count[0]), .A3(T_Count[1]), 
      .ZN(n_0_22_5));
   NOR2_X1 i_0_22_183 (.A1(T_Count[1]), .A2(n_0_22_6), .ZN(
      T_Counter_genblk1_1_counterBits_n_4));
   OAI21_X1 i_0_22_184 (.A(n_0_22_7), .B1(n_0_22_82), .B2(n_0_140), .ZN(
      T_Counter_genblk1_1_counterBits_n_2));
   NOR2_X1 i_0_22_185 (.A1(T_Count[0]), .A2(n_0_22_6), .ZN(
      T_Counter_firstBit_n_4));
   NAND2_X1 i_0_22_186 (.A1(n_0_22_82), .A2(n_0_22_7), .ZN(
      T_Counter_firstBit_n_2));
   INV_X1 i_0_22_187 (.A(n_0_22_7), .ZN(n_0_22_6));
   AOI21_X1 i_0_22_188 (.A(RST), .B1(T_Count_Enable), .B2(n_0_109), .ZN(n_0_22_7));
   NOR2_X1 i_0_22_189 (.A1(X_Count[7]), .A2(n_0_22_13), .ZN(
      X_Counter_genblk1_7_counterBits_n_4));
   AOI21_X1 i_0_22_190 (.A(X_Counter_genblk1_6_counterBits_n_4), .B1(n_0_22_14), 
      .B2(n_0_22_8), .ZN(X_Counter_genblk1_7_counterBits_n_2));
   NOR2_X1 i_0_22_191 (.A1(X_Count[6]), .A2(n_0_22_13), .ZN(
      X_Counter_genblk1_6_counterBits_n_4));
   NAND2_X1 i_0_22_192 (.A1(n_0_22_14), .A2(n_0_22_8), .ZN(
      X_Counter_genblk1_6_counterBits_n_2));
   NAND3_X1 i_0_22_193 (.A1(X_Count[4]), .A2(n_0_22_10), .A3(X_Count[5]), 
      .ZN(n_0_22_8));
   NOR2_X1 i_0_22_194 (.A1(X_Count[5]), .A2(n_0_22_13), .ZN(
      X_Counter_genblk1_5_counterBits_n_4));
   NOR2_X1 i_0_22_195 (.A1(n_0_22_9), .A2(X_Counter_genblk1_4_counterBits_n_4), 
      .ZN(X_Counter_genblk1_5_counterBits_n_2));
   NOR2_X1 i_0_22_196 (.A1(X_Count[4]), .A2(n_0_22_13), .ZN(
      X_Counter_genblk1_4_counterBits_n_4));
   INV_X1 i_0_22_197 (.A(n_0_22_9), .ZN(X_Counter_genblk1_4_counterBits_n_2));
   NOR2_X1 i_0_22_198 (.A1(n_0_22_13), .A2(n_0_22_10), .ZN(n_0_22_9));
   NOR2_X1 i_0_22_199 (.A1(n_0_22_83), .A2(n_0_22_11), .ZN(n_0_22_10));
   NOR2_X1 i_0_22_200 (.A1(X_Count[3]), .A2(n_0_22_13), .ZN(
      X_Counter_genblk1_3_counterBits_n_4));
   NAND2_X1 i_0_22_201 (.A1(n_0_22_14), .A2(n_0_22_11), .ZN(
      X_Counter_genblk1_3_counterBits_n_2));
   NAND4_X1 i_0_22_202 (.A1(X_Count_Enable), .A2(X_Count[1]), .A3(X_Count[0]), 
      .A4(X_Count[2]), .ZN(n_0_22_11));
   NOR2_X1 i_0_22_203 (.A1(X_Count[2]), .A2(n_0_22_13), .ZN(
      X_Counter_genblk1_2_counterBits_n_4));
   NAND2_X1 i_0_22_204 (.A1(n_0_22_14), .A2(n_0_22_12), .ZN(
      X_Counter_genblk1_2_counterBits_n_2));
   NAND3_X1 i_0_22_205 (.A1(X_Count_Enable), .A2(X_Count[0]), .A3(X_Count[1]), 
      .ZN(n_0_22_12));
   NOR2_X1 i_0_22_206 (.A1(X_Count[1]), .A2(n_0_22_13), .ZN(
      X_Counter_genblk1_1_counterBits_n_4));
   AOI21_X1 i_0_22_207 (.A(X_Counter_firstBit_n_4), .B1(n_0_22_84), .B2(
      n_0_22_14), .ZN(X_Counter_genblk1_1_counterBits_n_2));
   NOR2_X1 i_0_22_208 (.A1(X_Count[0]), .A2(n_0_22_13), .ZN(
      X_Counter_firstBit_n_4));
   NAND2_X1 i_0_22_209 (.A1(n_0_22_84), .A2(n_0_22_14), .ZN(
      X_Counter_firstBit_n_2));
   INV_X1 i_0_22_210 (.A(n_0_22_14), .ZN(n_0_22_13));
   AOI21_X1 i_0_22_211 (.A(RST), .B1(X_Count_Enable), .B2(n_0_155), .ZN(
      n_0_22_14));
   NOR2_X1 i_0_22_212 (.A1(RST), .A2(T_OR_X[0]), .ZN(T_OR_X_COUNTER_firstBit_n_4));
   OR2_X1 i_0_22_213 (.A1(RST), .A2(T_OR_X_Enable), .ZN(
      T_OR_X_COUNTER_firstBit_n_2));
   NOR2_X1 i_0_22_214 (.A1(Partial_Data_Count[0]), .A2(RST), .ZN(
      _64data_Counter_firstBit_n_4));
   OR2_X1 i_0_22_215 (.A1(_64data_Enable), .A2(RST), .ZN(
      _64data_Counter_firstBit_n_2));
   OR2_X1 i_0_22_216 (.A1(n_0_141), .A2(n_0_136), .ZN(n_0_341));
   NOR2_X1 i_0_22_217 (.A1(_64data_Enable), .A2(n_0_136), .ZN(n_0_342));
   INV_X1 i_0_22_218 (.A(n_0_362), .ZN(n_0_22_15));
   INV_X1 i_0_22_219 (.A(RAM_Data_A[0]), .ZN(n_0_22_16));
   INV_X1 i_0_22_220 (.A(RAM_Data_A[1]), .ZN(n_0_22_17));
   INV_X1 i_0_22_221 (.A(RAM_Data_A[2]), .ZN(n_0_22_18));
   INV_X1 i_0_22_222 (.A(RAM_Data_A[3]), .ZN(n_0_22_19));
   INV_X1 i_0_22_223 (.A(RAM_Data_A[4]), .ZN(n_0_22_20));
   INV_X1 i_0_22_224 (.A(RAM_Data_A[5]), .ZN(n_0_22_21));
   INV_X1 i_0_22_225 (.A(RAM_Data_A[6]), .ZN(n_0_22_22));
   INV_X1 i_0_22_226 (.A(RAM_Data_A[7]), .ZN(n_0_22_23));
   INV_X1 i_0_22_227 (.A(RAM_Data_A[8]), .ZN(n_0_22_24));
   INV_X1 i_0_22_228 (.A(RAM_Data_A[9]), .ZN(n_0_22_25));
   INV_X1 i_0_22_229 (.A(RAM_Data_A[10]), .ZN(n_0_22_26));
   INV_X1 i_0_22_230 (.A(RAM_Data_A[11]), .ZN(n_0_22_27));
   INV_X1 i_0_22_231 (.A(RAM_Data_A[12]), .ZN(n_0_22_28));
   INV_X1 i_0_22_232 (.A(RAM_Data_A[13]), .ZN(n_0_22_29));
   INV_X1 i_0_22_233 (.A(RAM_Data_A[14]), .ZN(n_0_22_30));
   INV_X1 i_0_22_234 (.A(RAM_Data_A[15]), .ZN(n_0_22_31));
   INV_X1 i_0_22_235 (.A(RAM_Data_A[16]), .ZN(n_0_22_32));
   INV_X1 i_0_22_236 (.A(RAM_Data_A[17]), .ZN(n_0_22_33));
   INV_X1 i_0_22_237 (.A(RAM_Data_A[18]), .ZN(n_0_22_34));
   INV_X1 i_0_22_238 (.A(RAM_Data_A[19]), .ZN(n_0_22_35));
   INV_X1 i_0_22_239 (.A(RAM_Data_A[20]), .ZN(n_0_22_36));
   INV_X1 i_0_22_240 (.A(RAM_Data_A[21]), .ZN(n_0_22_37));
   INV_X1 i_0_22_241 (.A(RAM_Data_A[22]), .ZN(n_0_22_38));
   INV_X1 i_0_22_242 (.A(RAM_Data_A[23]), .ZN(n_0_22_39));
   INV_X1 i_0_22_243 (.A(RAM_Data_A[24]), .ZN(n_0_22_40));
   INV_X1 i_0_22_244 (.A(RAM_Data_A[25]), .ZN(n_0_22_41));
   INV_X1 i_0_22_245 (.A(RAM_Data_A[26]), .ZN(n_0_22_42));
   INV_X1 i_0_22_246 (.A(RAM_Data_A[27]), .ZN(n_0_22_43));
   INV_X1 i_0_22_247 (.A(RAM_Data_A[28]), .ZN(n_0_22_44));
   INV_X1 i_0_22_248 (.A(RAM_Data_A[29]), .ZN(n_0_22_45));
   INV_X1 i_0_22_249 (.A(RAM_Data_A[30]), .ZN(n_0_22_46));
   INV_X1 i_0_22_250 (.A(RAM_Data_A[31]), .ZN(n_0_22_47));
   INV_X1 i_0_22_251 (.A(RAM_Data_A[32]), .ZN(n_0_22_48));
   INV_X1 i_0_22_252 (.A(RAM_Data_A[33]), .ZN(n_0_22_49));
   INV_X1 i_0_22_253 (.A(RAM_Data_A[34]), .ZN(n_0_22_50));
   INV_X1 i_0_22_254 (.A(RAM_Data_A[35]), .ZN(n_0_22_51));
   INV_X1 i_0_22_255 (.A(RAM_Data_A[36]), .ZN(n_0_22_52));
   INV_X1 i_0_22_256 (.A(RAM_Data_A[37]), .ZN(n_0_22_53));
   INV_X1 i_0_22_257 (.A(RAM_Data_A[38]), .ZN(n_0_22_54));
   INV_X1 i_0_22_258 (.A(RAM_Data_A[39]), .ZN(n_0_22_55));
   INV_X1 i_0_22_259 (.A(RAM_Data_A[40]), .ZN(n_0_22_56));
   INV_X1 i_0_22_260 (.A(RAM_Data_A[41]), .ZN(n_0_22_57));
   INV_X1 i_0_22_261 (.A(RAM_Data_A[42]), .ZN(n_0_22_58));
   INV_X1 i_0_22_262 (.A(RAM_Data_A[43]), .ZN(n_0_22_59));
   INV_X1 i_0_22_263 (.A(RAM_Data_A[44]), .ZN(n_0_22_60));
   INV_X1 i_0_22_264 (.A(RAM_Data_A[45]), .ZN(n_0_22_61));
   INV_X1 i_0_22_265 (.A(RAM_Data_A[46]), .ZN(n_0_22_62));
   INV_X1 i_0_22_266 (.A(RAM_Data_A[47]), .ZN(n_0_22_63));
   INV_X1 i_0_22_267 (.A(RAM_Data_A[48]), .ZN(n_0_22_64));
   INV_X1 i_0_22_268 (.A(RAM_Data_A[49]), .ZN(n_0_22_65));
   INV_X1 i_0_22_269 (.A(RAM_Data_A[50]), .ZN(n_0_22_66));
   INV_X1 i_0_22_270 (.A(RAM_Data_A[51]), .ZN(n_0_22_67));
   INV_X1 i_0_22_271 (.A(RAM_Data_A[52]), .ZN(n_0_22_68));
   INV_X1 i_0_22_272 (.A(RAM_Data_A[53]), .ZN(n_0_22_69));
   INV_X1 i_0_22_273 (.A(RAM_Data_A[54]), .ZN(n_0_22_70));
   INV_X1 i_0_22_274 (.A(RAM_Data_A[55]), .ZN(n_0_22_71));
   INV_X1 i_0_22_275 (.A(RAM_Data_A[56]), .ZN(n_0_22_72));
   INV_X1 i_0_22_276 (.A(RAM_Data_A[57]), .ZN(n_0_22_73));
   INV_X1 i_0_22_277 (.A(RAM_Data_A[58]), .ZN(n_0_22_74));
   INV_X1 i_0_22_278 (.A(RAM_Data_A[59]), .ZN(n_0_22_75));
   INV_X1 i_0_22_279 (.A(RAM_Data_A[60]), .ZN(n_0_22_76));
   INV_X1 i_0_22_280 (.A(RAM_Data_A[61]), .ZN(n_0_22_77));
   INV_X1 i_0_22_281 (.A(RAM_Data_A[62]), .ZN(n_0_22_78));
   INV_X1 i_0_22_282 (.A(RAM_Data_A[63]), .ZN(n_0_22_79));
   INV_X1 i_0_22_283 (.A(Init_Count_Enable), .ZN(n_0_22_80));
   INV_X1 i_0_22_284 (.A(T_Count[0]), .ZN(n_0_140));
   INV_X1 i_0_22_285 (.A(T_Count[3]), .ZN(n_0_22_81));
   INV_X1 i_0_22_286 (.A(T_Count_Enable), .ZN(n_0_22_82));
   INV_X1 i_0_22_287 (.A(X_Count[3]), .ZN(n_0_22_83));
   INV_X1 i_0_22_288 (.A(X_Count_Enable), .ZN(n_0_22_84));
   INV_X1 i_0_22_289 (.A(RST), .ZN(n_0_139));
   INV_X1 i_0_22_290 (.A(Partial_Data_Count[0]), .ZN(n_0_141));
   datapath__1_253 i_0_1 (.X_Count(X_Count), .p_0({n_0_154, n_0_153, n_0_152, 
      n_0_151, n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, 
      n_0_143, n_0_142}), .T_Count(T_Count), .num_of_X({num_of_X[12], 
      num_of_X[11], num_of_X[10], num_of_X[9], num_of_X[8], num_of_X[7], 
      num_of_X[6], num_of_X[5], num_of_X[4], num_of_X[3], num_of_X[2], 
      num_of_X[1], num_of_X[0]}));
   datapath__1_501 i_0_23 (.p_0({n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, 
      n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, 
      n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, 
      n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, 
      n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, 
      n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, 
      n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, 
      n_0_2, n_0_1, n_0_110}), .X_Count(X_Count), .p_1(n_0_155));
   datapath__1_506 i_0_24 (.p_0({n_0_133, n_0_132, n_0_131, n_0_130, n_0_129, 
      n_0_128, n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, 
      n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_108, n_0_107, n_0_106, 
      n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, 
      n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, 
      n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, 
      n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, 
      n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_363}), 
      .T_Count(T_Count), .p_1(n_0_156));
   HA_X1 i_0_25_0 (.A(T_Count[2]), .B(n_0_25_9), .CO(n_0_25_0), .S(n_0_159));
   HA_X1 i_0_25_1 (.A(T_Count[3]), .B(n_0_25_0), .CO(n_0_25_1), .S(n_0_160));
   HA_X1 i_0_25_2 (.A(T_Count[4]), .B(n_0_25_1), .CO(n_0_25_2), .S(n_0_161));
   HA_X1 i_0_25_3 (.A(T_Count[5]), .B(n_0_25_2), .CO(n_0_25_3), .S(n_0_162));
   HA_X1 i_0_25_4 (.A(T_Count[6]), .B(n_0_25_3), .CO(n_0_25_4), .S(n_0_163));
   HA_X1 i_0_25_5 (.A(T_Count[7]), .B(n_0_25_4), .CO(n_0_165), .S(n_0_164));
   NOR3_X1 i_0_25_6 (.A1(n_0_341), .A2(RST), .A3(n_0_342), .ZN(n_0_360));
   INV_X1 i_0_25_7 (.A(n_0_342), .ZN(n_0_25_5));
   NOR2_X1 i_0_25_8 (.A1(n_0_25_5), .A2(RST), .ZN(n_0_361));
   INV_X1 i_0_25_9 (.A(n_0_341), .ZN(n_0_25_6));
   NOR3_X1 i_0_25_10 (.A1(n_0_25_6), .A2(RST), .A3(n_0_342), .ZN(n_0_362));
   INV_X1 i_0_25_11 (.A(T_Count[1]), .ZN(n_0_25_7));
   INV_X1 i_0_25_12 (.A(T_Count[0]), .ZN(n_0_25_8));
   NAND2_X1 i_0_25_13 (.A1(n_0_25_7), .A2(n_0_25_8), .ZN(n_0_25_9));
   OAI21_X1 i_0_25_14 (.A(n_0_25_9), .B1(n_0_25_7), .B2(n_0_25_8), .ZN(n_0_158));
   INV_X1 i_0_25_15 (.A(num_of_T[0]), .ZN(n_0_363));
   NOR4_X1 i_0_25_16 (.A1(num_of_T[19]), .A2(num_of_T[16]), .A3(num_of_T[22]), 
      .A4(num_of_T[21]), .ZN(n_0_25_10));
   NOR4_X1 i_0_25_17 (.A1(num_of_T[10]), .A2(num_of_T[9]), .A3(num_of_T[15]), 
      .A4(num_of_T[12]), .ZN(n_0_25_11));
   NOR4_X1 i_0_25_18 (.A1(num_of_T[34]), .A2(num_of_T[33]), .A3(num_of_T[39]), 
      .A4(num_of_T[36]), .ZN(n_0_25_12));
   NOR4_X1 i_0_25_19 (.A1(num_of_T[27]), .A2(num_of_T[24]), .A3(num_of_T[30]), 
      .A4(num_of_T[29]), .ZN(n_0_25_13));
   NAND4_X1 i_0_25_20 (.A1(n_0_25_10), .A2(n_0_25_11), .A3(n_0_25_12), .A4(
      n_0_25_13), .ZN(n_0_25_14));
   XNOR2_X1 i_0_25_21 (.A(num_of_T[1]), .B(T_Count[1]), .ZN(n_0_25_15));
   OAI221_X1 i_0_25_22 (.A(n_0_25_15), .B1(n_0_363), .B2(T_Count[0]), .C1(
      n_0_25_8), .C2(num_of_T[0]), .ZN(n_0_25_16));
   XOR2_X1 i_0_25_23 (.A(num_of_T[4]), .B(T_Count[4]), .Z(n_0_25_17));
   XOR2_X1 i_0_25_24 (.A(num_of_T[5]), .B(T_Count[5]), .Z(n_0_25_18));
   NOR4_X1 i_0_25_25 (.A1(n_0_25_14), .A2(n_0_25_16), .A3(n_0_25_17), .A4(
      n_0_25_18), .ZN(n_0_25_19));
   NOR4_X1 i_0_25_26 (.A1(num_of_T[50]), .A2(num_of_T[49]), .A3(num_of_T[55]), 
      .A4(num_of_T[52]), .ZN(n_0_25_20));
   NOR4_X1 i_0_25_27 (.A1(num_of_T[43]), .A2(num_of_T[40]), .A3(num_of_T[46]), 
      .A4(num_of_T[45]), .ZN(n_0_25_21));
   NOR4_X1 i_0_25_28 (.A1(num_of_T[59]), .A2(num_of_T[56]), .A3(num_of_T[62]), 
      .A4(num_of_T[61]), .ZN(n_0_25_22));
   NOR4_X1 i_0_25_29 (.A1(num_of_T[58]), .A2(num_of_T[57]), .A3(num_of_T[63]), 
      .A4(num_of_T[60]), .ZN(n_0_25_23));
   NOR4_X1 i_0_25_30 (.A1(num_of_T[51]), .A2(num_of_T[48]), .A3(num_of_T[54]), 
      .A4(num_of_T[53]), .ZN(n_0_25_24));
   NOR4_X1 i_0_25_31 (.A1(num_of_T[42]), .A2(num_of_T[41]), .A3(num_of_T[47]), 
      .A4(num_of_T[44]), .ZN(n_0_25_25));
   AND4_X1 i_0_25_32 (.A1(n_0_25_22), .A2(n_0_25_23), .A3(n_0_25_24), .A4(
      n_0_25_25), .ZN(n_0_25_26));
   NAND4_X1 i_0_25_33 (.A1(n_0_25_19), .A2(n_0_25_20), .A3(n_0_25_21), .A4(
      n_0_25_26), .ZN(n_0_25_27));
   XNOR2_X1 i_0_25_34 (.A(num_of_T[3]), .B(T_Count[3]), .ZN(n_0_25_28));
   XNOR2_X1 i_0_25_35 (.A(num_of_T[2]), .B(T_Count[2]), .ZN(n_0_25_29));
   NAND2_X1 i_0_25_36 (.A1(n_0_25_28), .A2(n_0_25_29), .ZN(n_0_25_30));
   XNOR2_X1 i_0_25_37 (.A(num_of_T[7]), .B(T_Count[7]), .ZN(n_0_25_31));
   XNOR2_X1 i_0_25_38 (.A(num_of_T[6]), .B(T_Count[6]), .ZN(n_0_25_32));
   NAND2_X1 i_0_25_39 (.A1(n_0_25_31), .A2(n_0_25_32), .ZN(n_0_25_33));
   NOR4_X1 i_0_25_40 (.A1(num_of_T[18]), .A2(num_of_T[17]), .A3(num_of_T[23]), 
      .A4(num_of_T[20]), .ZN(n_0_25_34));
   NOR4_X1 i_0_25_41 (.A1(num_of_T[11]), .A2(num_of_T[8]), .A3(num_of_T[14]), 
      .A4(num_of_T[13]), .ZN(n_0_25_35));
   NOR4_X1 i_0_25_42 (.A1(num_of_T[35]), .A2(num_of_T[32]), .A3(num_of_T[38]), 
      .A4(num_of_T[37]), .ZN(n_0_25_36));
   NOR4_X1 i_0_25_43 (.A1(num_of_T[26]), .A2(num_of_T[25]), .A3(num_of_T[31]), 
      .A4(num_of_T[28]), .ZN(n_0_25_37));
   NAND4_X1 i_0_25_44 (.A1(n_0_25_34), .A2(n_0_25_35), .A3(n_0_25_36), .A4(
      n_0_25_37), .ZN(n_0_25_38));
   NOR4_X1 i_0_25_45 (.A1(n_0_25_27), .A2(n_0_25_30), .A3(n_0_25_33), .A4(
      n_0_25_38), .ZN(n_0_109));
   NOR2_X1 i_0_25_46 (.A1(Init_Count[1]), .A2(Init_Count[0]), .ZN(n_0_340));
   INV_X1 i_0_25_47 (.A(Init_Count[1]), .ZN(n_0_25_39));
   NOR2_X1 i_0_25_48 (.A1(n_0_25_39), .A2(Init_Count[0]), .ZN(n_0_343));
   INV_X1 i_0_25_49 (.A(CLK), .ZN(n_0_137));
   INV_X1 i_0_25_50 (.A(num_of_X[0]), .ZN(n_0_110));
   MUX2_X1 _64data_Counter_firstBit_Q_reg_enable_mux_0 (.A(Partial_Data_Count[0]), 
      .B(_64data_Counter_firstBit_n_4), .S(_64data_Counter_firstBit_n_2), 
      .Z(n_0_111));
   MUX2_X1 T_OR_X_COUNTER_firstBit_Q_reg_enable_mux_0 (.A(T_OR_X[0]), .B(
      T_OR_X_COUNTER_firstBit_n_4), .S(T_OR_X_COUNTER_firstBit_n_2), .Z(n_0_112));
   AOI21_X1 X_Counter_firstBit_Q_reg_enable_mux_0 (.A(
      X_Counter_firstBit_Q_reg_enable_mux_n_0), .B1(
      X_Counter_firstBit_Q_reg_enable_mux_n_1), .B2(X_Counter_firstBit_n_2), 
      .ZN(n_0_113));
   NOR2_X1 X_Counter_firstBit_Q_reg_enable_mux_1 (.A1(X_Counter_firstBit_n_2), 
      .A2(X_Count[0]), .ZN(X_Counter_firstBit_Q_reg_enable_mux_n_0));
   INV_X1 X_Counter_firstBit_Q_reg_enable_mux_2 (.A(X_Counter_firstBit_n_4), 
      .ZN(X_Counter_firstBit_Q_reg_enable_mux_n_1));
   NAND2_X1 X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_0 (.A1(
      X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_n_1), .A2(
      X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_n_0), .ZN(n_0_114));
   NAND2_X1 X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_1 (.A1(
      X_Counter_genblk1_1_counterBits_n_2), .A2(
      X_Counter_genblk1_1_counterBits_n_4), .ZN(
      X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_n_0));
   NAND2_X1 X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_2 (.A1(
      X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_n_2), .A2(X_Count[1]), 
      .ZN(X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_n_1));
   INV_X1 X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_3 (.A(
      X_Counter_genblk1_1_counterBits_n_2), .ZN(
      X_Counter_genblk1_1_counterBits_Q_reg_enable_mux_n_2));
   NAND2_X1 X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_0 (.A1(
      X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_n_1), .A2(
      X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_n_0), .ZN(n_0_115));
   NAND2_X1 X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_1 (.A1(
      X_Counter_genblk1_2_counterBits_n_2), .A2(
      X_Counter_genblk1_2_counterBits_n_4), .ZN(
      X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_n_0));
   NAND2_X1 X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_2 (.A1(
      X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_n_2), .A2(X_Count[2]), 
      .ZN(X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_n_1));
   INV_X1 X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_3 (.A(
      X_Counter_genblk1_2_counterBits_n_2), .ZN(
      X_Counter_genblk1_2_counterBits_Q_reg_enable_mux_n_2));
   NAND2_X1 X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_0 (.A1(
      X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_n_1), .A2(
      X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_n_0), .ZN(n_0_134));
   NAND2_X1 X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_1 (.A1(
      X_Counter_genblk1_3_counterBits_n_2), .A2(
      X_Counter_genblk1_3_counterBits_n_4), .ZN(
      X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_n_0));
   NAND2_X1 X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_2 (.A1(
      X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_n_2), .A2(X_Count[3]), 
      .ZN(X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_n_1));
   INV_X1 X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_3 (.A(
      X_Counter_genblk1_3_counterBits_n_2), .ZN(
      X_Counter_genblk1_3_counterBits_Q_reg_enable_mux_n_2));
   NAND2_X1 X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_0 (.A1(
      X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_n_1), .A2(
      X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_n_0), .ZN(n_0_135));
   NAND2_X1 X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_1 (.A1(
      X_Counter_genblk1_4_counterBits_n_2), .A2(
      X_Counter_genblk1_4_counterBits_n_4), .ZN(
      X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_n_0));
   NAND2_X1 X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_2 (.A1(
      X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_n_2), .A2(X_Count[4]), 
      .ZN(X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_n_1));
   INV_X1 X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_3 (.A(
      X_Counter_genblk1_4_counterBits_n_2), .ZN(
      X_Counter_genblk1_4_counterBits_Q_reg_enable_mux_n_2));
   NAND2_X1 X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_0 (.A1(
      X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_n_1), .A2(
      X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_n_0), .ZN(n_0_180));
   NAND2_X1 X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_1 (.A1(
      X_Counter_genblk1_5_counterBits_n_2), .A2(
      X_Counter_genblk1_5_counterBits_n_4), .ZN(
      X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_n_0));
   NAND2_X1 X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_2 (.A1(
      X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_n_2), .A2(X_Count[5]), 
      .ZN(X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_n_1));
   INV_X1 X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_3 (.A(
      X_Counter_genblk1_5_counterBits_n_2), .ZN(
      X_Counter_genblk1_5_counterBits_Q_reg_enable_mux_n_2));
   NAND2_X1 X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_0 (.A1(
      X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_n_1), .A2(
      X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_n_0), .ZN(n_0_181));
   NAND2_X1 X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_1 (.A1(
      X_Counter_genblk1_6_counterBits_n_2), .A2(
      X_Counter_genblk1_6_counterBits_n_4), .ZN(
      X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_n_0));
   NAND2_X1 X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_2 (.A1(
      X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_n_2), .A2(X_Count[6]), 
      .ZN(X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_n_1));
   INV_X1 X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_3 (.A(
      X_Counter_genblk1_6_counterBits_n_2), .ZN(
      X_Counter_genblk1_6_counterBits_Q_reg_enable_mux_n_2));
   NAND2_X1 X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_0 (.A1(
      X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_n_1), .A2(
      X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_n_0), .ZN(n_0_182));
   NAND2_X1 X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_1 (.A1(
      X_Counter_genblk1_7_counterBits_n_2), .A2(
      X_Counter_genblk1_7_counterBits_n_4), .ZN(
      X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_n_0));
   NAND2_X1 X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_2 (.A1(
      X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_n_2), .A2(X_Count[7]), 
      .ZN(X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_n_1));
   INV_X1 X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_3 (.A(
      X_Counter_genblk1_7_counterBits_n_2), .ZN(
      X_Counter_genblk1_7_counterBits_Q_reg_enable_mux_n_2));
   MUX2_X1 T_Counter_firstBit_Q_reg_enable_mux_0 (.A(T_Count[0]), .B(
      T_Counter_firstBit_n_4), .S(T_Counter_firstBit_n_2), .Z(n_0_184));
   MUX2_X1 T_Counter_genblk1_1_counterBits_Q_reg_enable_mux_0 (.A(T_Count[1]), 
      .B(T_Counter_genblk1_1_counterBits_n_4), .S(
      T_Counter_genblk1_1_counterBits_n_2), .Z(n_0_185));
   MUX2_X1 T_Counter_genblk1_2_counterBits_Q_reg_enable_mux_0 (.A(T_Count[2]), 
      .B(T_Counter_genblk1_2_counterBits_n_4), .S(
      T_Counter_genblk1_2_counterBits_n_2), .Z(n_0_186));
   MUX2_X1 T_Counter_genblk1_3_counterBits_Q_reg_enable_mux_0 (.A(T_Count[3]), 
      .B(T_Counter_genblk1_3_counterBits_n_4), .S(
      T_Counter_genblk1_3_counterBits_n_2), .Z(n_0_187));
   MUX2_X1 T_Counter_genblk1_4_counterBits_Q_reg_enable_mux_0 (.A(T_Count[4]), 
      .B(T_Counter_genblk1_4_counterBits_n_4), .S(
      T_Counter_genblk1_4_counterBits_n_2), .Z(n_0_188));
   MUX2_X1 T_Counter_genblk1_5_counterBits_Q_reg_enable_mux_0 (.A(T_Count[5]), 
      .B(T_Counter_genblk1_5_counterBits_n_4), .S(
      T_Counter_genblk1_5_counterBits_n_2), .Z(n_0_189));
   MUX2_X1 T_Counter_genblk1_6_counterBits_Q_reg_enable_mux_0 (.A(T_Count[6]), 
      .B(T_Counter_genblk1_6_counterBits_n_4), .S(
      T_Counter_genblk1_6_counterBits_n_2), .Z(n_0_190));
   MUX2_X1 T_Counter_genblk1_7_counterBits_Q_reg_enable_mux_0 (.A(T_Count[7]), 
      .B(T_Counter_genblk1_7_counterBits_n_4), .S(
      T_Counter_genblk1_7_counterBits_n_2), .Z(n_0_242));
   MUX2_X1 Init_Counter_firstBit_Q_reg_enable_mux_0 (.A(Init_Count[0]), .B(
      Init_Counter_firstBit_n_4), .S(Init_Counter_firstBit_n_2), .Z(n_0_243));
   MUX2_X1 Init_Counter_genblk1_1_counterBits_Q_reg_enable_mux_0 (.A(
      Init_Count[1]), .B(Init_Counter_genblk1_1_counterBits_n_4), .S(
      Init_Counter_genblk1_1_counterBits_n_2), .Z(n_0_308));
   DFF_X2 \num_of_X_reg[3]  (.D(n_0_169), .CK(n_0_0), .Q(num_of_X[3]), .QN());
   BUF_X1 rt_shieldBuf__1 (.A(Done_Sending), .Z(n_0_136));
   INV_X1 i_0_30_0 (.A(Init_Count[0]), .ZN(n_0_30_0));
   NAND2_X1 i_0_30_1 (.A1(n_0_30_2), .A2(n_0_30_1), .ZN(n_0_138));
   NAND2_X1 i_0_30_2 (.A1(Init_Count_Enable), .A2(n_0_30_4), .ZN(n_0_30_1));
   NAND2_X1 i_0_30_3 (.A1(Sending_Enable), .A2(n_0_30_3), .ZN(n_0_30_2));
   AOI21_X1 i_0_30_4 (.A(n_0_30_4), .B1(n_0_30_0), .B2(Init_Count[1]), .ZN(
      n_0_30_3));
   INV_X1 i_0_30_5 (.A(n_0_139), .ZN(n_0_30_4));
   AND2_X1 i_0_3_0 (.A1(Sending_Enable), .A2(n_0_340), .ZN(n_0_344));
   AOI21_X1 i_0_4_0 (.A(n_0_4_0), .B1(Sending_Enable), .B2(n_0_340), .ZN(n_0_157));
   NAND4_X1 i_0_4_1 (.A1(n_0_156), .A2(n_0_141), .A3(n_0_155), .A4(n_0_4_1), 
      .ZN(n_0_4_0));
   INV_X1 i_0_4_2 (.A(RST), .ZN(n_0_4_1));
   INV_X1 i_0_5_0 (.A(n_0_139), .ZN(n_0_5_0));
   NAND2_X1 i_0_5_1 (.A1(T_Count_Enable), .A2(n_0_5_0), .ZN(n_0_5_1));
   INV_X1 i_0_5_2 (.A(n_0_5_1), .ZN(n_0_5_2));
   NOR2_X1 i_0_5_3 (.A1(Partial_Data_Count[0]), .A2(n_0_5_0), .ZN(n_0_5_3));
   NAND2_X1 i_0_5_4 (.A1(n_0_343), .A2(n_0_5_3), .ZN(n_0_5_4));
   NOR2_X1 i_0_5_5 (.A1(n_0_5_4), .A2(n_0_141), .ZN(n_0_5_5));
   AOI21_X1 i_0_5_6 (.A(n_0_5_2), .B1(n_0_155), .B2(n_0_5_5), .ZN(n_0_5_6));
   INV_X1 i_0_5_7 (.A(n_0_5_4), .ZN(n_0_5_7));
   NAND2_X1 i_0_5_8 (.A1(n_0_155), .A2(n_0_5_7), .ZN(n_0_5_8));
   OAI21_X1 i_0_5_9 (.A(n_0_5_6), .B1(n_0_5_8), .B2(n_0_156), .ZN(n_0_5_9));
   INV_X1 i_0_5_10 (.A(n_0_5_9), .ZN(n_0_5_10));
   INV_X1 i_0_5_11 (.A(Sending_Enable), .ZN(n_0_5_11));
   INV_X1 i_0_5_12 (.A(n_0_340), .ZN(n_0_5_12));
   NOR2_X1 i_0_5_13 (.A1(n_0_5_4), .A2(n_0_5_12), .ZN(n_0_5_13));
   NAND2_X1 i_0_5_14 (.A1(n_0_155), .A2(n_0_5_13), .ZN(n_0_5_14));
   OAI21_X1 i_0_5_15 (.A(n_0_5_10), .B1(n_0_5_11), .B2(n_0_5_14), .ZN(n_0_345));
   NAND4_X1 i_0_6_0 (.A1(n_0_156), .A2(n_0_141), .A3(n_0_155), .A4(n_0_139), 
      .ZN(n_0_6_0));
   OAI21_X1 i_0_6_1 (.A(n_0_6_5), .B1(n_0_6_2), .B2(n_0_139), .ZN(n_0_6_1));
   INV_X1 i_0_6_2 (.A(X_Count_Enable), .ZN(n_0_6_2));
   NAND2_X1 i_0_6_3 (.A1(n_0_6_4), .A2(n_0_340), .ZN(n_0_6_3));
   INV_X1 i_0_6_4 (.A(n_0_6_5), .ZN(n_0_6_4));
   NAND4_X1 i_0_6_5 (.A1(n_0_343), .A2(n_0_6_6), .A3(n_0_139), .A4(T_OR_X[0]), 
      .ZN(n_0_6_5));
   INV_X1 i_0_6_6 (.A(Partial_Data_Count[0]), .ZN(n_0_6_6));
   NAND2_X1 i_0_6_7 (.A1(n_0_6_0), .A2(n_0_6_1), .ZN(n_0_6_7));
   INV_X1 i_0_6_8 (.A(Sending_Enable), .ZN(n_0_6_8));
   OAI21_X1 i_0_6_9 (.A(n_0_6_7), .B1(n_0_6_8), .B2(n_0_6_3), .ZN(n_0_346));
   AOI21_X1 i_0_7_0 (.A(n_0_7_0), .B1(Sending_Enable), .B2(n_0_7_6), .ZN(n_0_347));
   AOI21_X1 i_0_7_1 (.A(n_0_7_3), .B1(n_0_154), .B2(n_0_7_1), .ZN(n_0_7_0));
   INV_X1 i_0_7_2 (.A(n_0_7_2), .ZN(n_0_7_1));
   NAND2_X1 i_0_7_3 (.A1(T_OR_X[0]), .A2(n_0_139), .ZN(n_0_7_2));
   INV_X1 i_0_7_4 (.A(n_0_7_4), .ZN(n_0_7_3));
   NAND2_X1 i_0_7_5 (.A1(RAM_Address_A[12]), .A2(n_0_7_5), .ZN(n_0_7_4));
   INV_X1 i_0_7_6 (.A(n_0_139), .ZN(n_0_7_5));
   INV_X1 i_0_7_7 (.A(n_0_7_7), .ZN(n_0_7_6));
   NAND2_X1 i_0_7_8 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_7_7));
   INV_X1 i_0_8_0 (.A(n_0_139), .ZN(n_0_8_0));
   NAND2_X1 i_0_8_1 (.A1(RAM_Address_A[11]), .A2(n_0_8_0), .ZN(n_0_8_1));
   NAND2_X1 i_0_8_2 (.A1(n_0_8_1), .A2(n_0_8_0), .ZN(n_0_8_2));
   INV_X1 i_0_8_3 (.A(n_0_8_2), .ZN(n_0_8_3));
   INV_X1 i_0_8_4 (.A(T_OR_X[0]), .ZN(n_0_8_4));
   AOI21_X1 i_0_8_5 (.A(n_0_8_3), .B1(n_0_8_4), .B2(n_0_8_1), .ZN(n_0_8_5));
   INV_X1 i_0_8_6 (.A(n_0_8_1), .ZN(n_0_8_6));
   OAI21_X1 i_0_8_7 (.A(n_0_8_5), .B1(n_0_153), .B2(n_0_8_6), .ZN(n_0_8_7));
   NAND2_X1 i_0_8_8 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_8_8));
   INV_X1 i_0_8_9 (.A(n_0_8_8), .ZN(n_0_8_9));
   AOI21_X1 i_0_8_10 (.A(n_0_8_7), .B1(Sending_Enable), .B2(n_0_8_9), .ZN(
      n_0_348));
   AOI21_X1 i_0_9_0 (.A(n_0_9_0), .B1(Sending_Enable), .B2(n_0_9_6), .ZN(n_0_349));
   AOI21_X1 i_0_9_1 (.A(n_0_9_3), .B1(n_0_152), .B2(n_0_9_1), .ZN(n_0_9_0));
   INV_X1 i_0_9_2 (.A(n_0_9_2), .ZN(n_0_9_1));
   NAND2_X1 i_0_9_3 (.A1(T_OR_X[0]), .A2(n_0_139), .ZN(n_0_9_2));
   INV_X1 i_0_9_4 (.A(n_0_9_4), .ZN(n_0_9_3));
   NAND2_X1 i_0_9_5 (.A1(RAM_Address_A[10]), .A2(n_0_9_5), .ZN(n_0_9_4));
   INV_X1 i_0_9_6 (.A(n_0_139), .ZN(n_0_9_5));
   INV_X1 i_0_9_7 (.A(n_0_9_7), .ZN(n_0_9_6));
   NAND2_X1 i_0_9_8 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_9_7));
   AOI21_X1 i_0_10_0 (.A(n_0_10_0), .B1(Sending_Enable), .B2(n_0_10_6), .ZN(
      n_0_350));
   AOI21_X1 i_0_10_1 (.A(n_0_10_3), .B1(n_0_151), .B2(n_0_10_1), .ZN(n_0_10_0));
   INV_X1 i_0_10_2 (.A(n_0_10_2), .ZN(n_0_10_1));
   NAND2_X1 i_0_10_3 (.A1(T_OR_X[0]), .A2(n_0_139), .ZN(n_0_10_2));
   INV_X1 i_0_10_4 (.A(n_0_10_4), .ZN(n_0_10_3));
   NAND2_X1 i_0_10_5 (.A1(RAM_Address_A[9]), .A2(n_0_10_5), .ZN(n_0_10_4));
   INV_X1 i_0_10_6 (.A(n_0_139), .ZN(n_0_10_5));
   INV_X1 i_0_10_7 (.A(n_0_10_7), .ZN(n_0_10_6));
   NAND2_X1 i_0_10_8 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_10_7));
   INV_X1 i_0_11_0 (.A(n_0_139), .ZN(n_0_11_0));
   NAND2_X1 i_0_11_1 (.A1(RAM_Address_A[8]), .A2(n_0_11_0), .ZN(n_0_11_1));
   INV_X1 i_0_11_2 (.A(n_0_11_1), .ZN(n_0_11_2));
   NOR2_X1 i_0_11_3 (.A1(T_OR_X[0]), .A2(n_0_11_0), .ZN(n_0_11_3));
   AOI21_X1 i_0_11_4 (.A(n_0_11_2), .B1(n_0_165), .B2(n_0_11_3), .ZN(n_0_11_4));
   INV_X1 i_0_11_5 (.A(n_0_11_4), .ZN(n_0_11_5));
   NAND2_X1 i_0_11_6 (.A1(T_OR_X[0]), .A2(n_0_139), .ZN(n_0_11_6));
   INV_X1 i_0_11_7 (.A(n_0_11_6), .ZN(n_0_11_7));
   AOI21_X1 i_0_11_8 (.A(n_0_11_5), .B1(n_0_150), .B2(n_0_11_7), .ZN(n_0_11_8));
   NAND2_X1 i_0_11_9 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_11_9));
   INV_X1 i_0_11_10 (.A(n_0_11_9), .ZN(n_0_11_10));
   AOI21_X1 i_0_11_11 (.A(n_0_11_8), .B1(Sending_Enable), .B2(n_0_11_10), 
      .ZN(n_0_351));
   INV_X1 i_0_12_0 (.A(n_0_139), .ZN(n_0_12_0));
   NAND2_X1 i_0_12_1 (.A1(RAM_Address_A[7]), .A2(n_0_12_0), .ZN(n_0_12_1));
   INV_X1 i_0_12_2 (.A(n_0_12_1), .ZN(n_0_12_2));
   NOR2_X1 i_0_12_3 (.A1(T_OR_X[0]), .A2(n_0_12_0), .ZN(n_0_12_3));
   AOI21_X1 i_0_12_4 (.A(n_0_12_2), .B1(n_0_164), .B2(n_0_12_3), .ZN(n_0_12_4));
   INV_X1 i_0_12_5 (.A(n_0_12_4), .ZN(n_0_12_5));
   NAND2_X1 i_0_12_6 (.A1(T_OR_X[0]), .A2(n_0_139), .ZN(n_0_12_6));
   INV_X1 i_0_12_7 (.A(n_0_12_6), .ZN(n_0_12_7));
   AOI21_X1 i_0_12_8 (.A(n_0_12_5), .B1(n_0_149), .B2(n_0_12_7), .ZN(n_0_12_8));
   NAND2_X1 i_0_12_9 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_12_9));
   INV_X1 i_0_12_10 (.A(n_0_12_9), .ZN(n_0_12_10));
   AOI21_X1 i_0_12_11 (.A(n_0_12_8), .B1(Sending_Enable), .B2(n_0_12_10), 
      .ZN(n_0_352));
   INV_X1 i_0_13_0 (.A(n_0_139), .ZN(n_0_13_0));
   NAND2_X1 i_0_13_1 (.A1(RAM_Address_A[6]), .A2(n_0_13_0), .ZN(n_0_13_1));
   INV_X1 i_0_13_2 (.A(n_0_13_1), .ZN(n_0_13_2));
   NOR2_X1 i_0_13_3 (.A1(T_OR_X[0]), .A2(n_0_13_0), .ZN(n_0_13_3));
   AOI21_X1 i_0_13_4 (.A(n_0_13_2), .B1(n_0_163), .B2(n_0_13_3), .ZN(n_0_13_4));
   INV_X1 i_0_13_5 (.A(n_0_13_4), .ZN(n_0_13_5));
   NAND2_X1 i_0_13_6 (.A1(T_OR_X[0]), .A2(n_0_139), .ZN(n_0_13_6));
   INV_X1 i_0_13_7 (.A(n_0_13_6), .ZN(n_0_13_7));
   AOI21_X1 i_0_13_8 (.A(n_0_13_5), .B1(n_0_148), .B2(n_0_13_7), .ZN(n_0_13_8));
   NAND2_X1 i_0_13_9 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_13_9));
   INV_X1 i_0_13_10 (.A(n_0_13_9), .ZN(n_0_13_10));
   AOI21_X1 i_0_13_11 (.A(n_0_13_8), .B1(Sending_Enable), .B2(n_0_13_10), 
      .ZN(n_0_353));
   INV_X1 i_0_14_0 (.A(n_0_139), .ZN(n_0_14_0));
   NAND2_X1 i_0_14_1 (.A1(RAM_Address_A[5]), .A2(n_0_14_0), .ZN(n_0_14_1));
   INV_X1 i_0_14_2 (.A(n_0_14_1), .ZN(n_0_14_2));
   NOR2_X1 i_0_14_3 (.A1(T_OR_X[0]), .A2(n_0_14_0), .ZN(n_0_14_3));
   AOI21_X1 i_0_14_4 (.A(n_0_14_2), .B1(n_0_162), .B2(n_0_14_3), .ZN(n_0_14_4));
   INV_X1 i_0_14_5 (.A(n_0_14_4), .ZN(n_0_14_5));
   NAND2_X1 i_0_14_6 (.A1(T_OR_X[0]), .A2(n_0_139), .ZN(n_0_14_6));
   INV_X1 i_0_14_7 (.A(n_0_14_6), .ZN(n_0_14_7));
   AOI21_X1 i_0_14_8 (.A(n_0_14_5), .B1(n_0_147), .B2(n_0_14_7), .ZN(n_0_14_8));
   NAND2_X1 i_0_14_9 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_14_9));
   INV_X1 i_0_14_10 (.A(n_0_14_9), .ZN(n_0_14_10));
   AOI21_X1 i_0_14_11 (.A(n_0_14_8), .B1(Sending_Enable), .B2(n_0_14_10), 
      .ZN(n_0_354));
   INV_X1 i_0_15_0 (.A(n_0_139), .ZN(n_0_15_0));
   NAND2_X1 i_0_15_1 (.A1(RAM_Address_A[4]), .A2(n_0_15_0), .ZN(n_0_15_1));
   INV_X1 i_0_15_2 (.A(n_0_15_1), .ZN(n_0_15_2));
   NOR2_X1 i_0_15_3 (.A1(T_OR_X[0]), .A2(n_0_15_0), .ZN(n_0_15_3));
   AOI21_X1 i_0_15_4 (.A(n_0_15_2), .B1(n_0_161), .B2(n_0_15_3), .ZN(n_0_15_4));
   INV_X1 i_0_15_5 (.A(n_0_15_4), .ZN(n_0_15_5));
   NAND2_X1 i_0_15_6 (.A1(T_OR_X[0]), .A2(n_0_139), .ZN(n_0_15_6));
   INV_X1 i_0_15_7 (.A(n_0_15_6), .ZN(n_0_15_7));
   AOI21_X1 i_0_15_8 (.A(n_0_15_5), .B1(n_0_146), .B2(n_0_15_7), .ZN(n_0_15_8));
   NAND2_X1 i_0_15_9 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_15_9));
   INV_X1 i_0_15_10 (.A(n_0_15_9), .ZN(n_0_15_10));
   AOI21_X1 i_0_15_11 (.A(n_0_15_8), .B1(Sending_Enable), .B2(n_0_15_10), 
      .ZN(n_0_355));
   INV_X1 i_0_16_0 (.A(n_0_139), .ZN(n_0_16_0));
   NAND2_X1 i_0_16_1 (.A1(RAM_Address_A[3]), .A2(n_0_16_0), .ZN(n_0_16_1));
   INV_X1 i_0_16_2 (.A(n_0_16_1), .ZN(n_0_16_2));
   NOR2_X1 i_0_16_3 (.A1(T_OR_X[0]), .A2(n_0_16_0), .ZN(n_0_16_3));
   AOI21_X1 i_0_16_4 (.A(n_0_16_2), .B1(n_0_160), .B2(n_0_16_3), .ZN(n_0_16_4));
   INV_X1 i_0_16_5 (.A(n_0_16_4), .ZN(n_0_16_5));
   NAND2_X1 i_0_16_6 (.A1(T_OR_X[0]), .A2(n_0_139), .ZN(n_0_16_6));
   INV_X1 i_0_16_7 (.A(n_0_16_6), .ZN(n_0_16_7));
   AOI21_X1 i_0_16_8 (.A(n_0_16_5), .B1(n_0_145), .B2(n_0_16_7), .ZN(n_0_16_8));
   NAND2_X1 i_0_16_9 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_16_9));
   INV_X1 i_0_16_10 (.A(n_0_16_9), .ZN(n_0_16_10));
   AOI21_X1 i_0_16_11 (.A(n_0_16_8), .B1(Sending_Enable), .B2(n_0_16_10), 
      .ZN(n_0_356));
   INV_X1 i_0_17_0 (.A(n_0_139), .ZN(n_0_17_0));
   NAND2_X1 i_0_17_1 (.A1(RAM_Address_A[2]), .A2(n_0_17_0), .ZN(n_0_17_1));
   INV_X1 i_0_17_2 (.A(n_0_17_1), .ZN(n_0_17_2));
   NOR2_X1 i_0_17_3 (.A1(T_OR_X[0]), .A2(n_0_17_0), .ZN(n_0_17_3));
   AOI21_X1 i_0_17_4 (.A(n_0_17_2), .B1(n_0_159), .B2(n_0_17_3), .ZN(n_0_17_4));
   INV_X1 i_0_17_5 (.A(n_0_17_4), .ZN(n_0_17_5));
   NAND2_X1 i_0_17_6 (.A1(T_OR_X[0]), .A2(n_0_139), .ZN(n_0_17_6));
   INV_X1 i_0_17_7 (.A(n_0_17_6), .ZN(n_0_17_7));
   AOI21_X1 i_0_17_8 (.A(n_0_17_5), .B1(n_0_144), .B2(n_0_17_7), .ZN(n_0_17_8));
   NAND2_X1 i_0_17_9 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_17_9));
   INV_X1 i_0_17_10 (.A(n_0_17_9), .ZN(n_0_17_10));
   AOI21_X1 i_0_17_11 (.A(n_0_17_8), .B1(Sending_Enable), .B2(n_0_17_10), 
      .ZN(n_0_357));
   INV_X1 i_0_19_0 (.A(n_0_139), .ZN(n_0_19_0));
   NAND2_X1 i_0_19_1 (.A1(RAM_Address_A[1]), .A2(n_0_19_0), .ZN(n_0_19_1));
   INV_X1 i_0_19_2 (.A(n_0_19_1), .ZN(n_0_19_2));
   NOR2_X1 i_0_19_3 (.A1(T_OR_X[0]), .A2(n_0_19_0), .ZN(n_0_19_3));
   AOI21_X1 i_0_19_4 (.A(n_0_19_2), .B1(n_0_158), .B2(n_0_19_3), .ZN(n_0_19_4));
   INV_X1 i_0_19_5 (.A(n_0_19_4), .ZN(n_0_19_5));
   NAND2_X1 i_0_19_6 (.A1(T_OR_X[0]), .A2(n_0_139), .ZN(n_0_19_6));
   INV_X1 i_0_19_7 (.A(n_0_19_6), .ZN(n_0_19_7));
   AOI21_X1 i_0_19_8 (.A(n_0_19_5), .B1(n_0_143), .B2(n_0_19_7), .ZN(n_0_19_8));
   NAND2_X1 i_0_19_9 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_19_9));
   INV_X1 i_0_19_10 (.A(n_0_19_9), .ZN(n_0_19_10));
   AOI21_X1 i_0_19_11 (.A(n_0_19_8), .B1(Sending_Enable), .B2(n_0_19_10), 
      .ZN(n_0_358));
   NAND3_X1 i_0_21_0 (.A1(n_0_343), .A2(n_0_340), .A3(n_0_139), .ZN(n_0_21_0));
   NAND4_X1 i_0_21_1 (.A1(n_0_156), .A2(n_0_155), .A3(n_0_141), .A4(n_0_139), 
      .ZN(n_0_21_1));
   MUX2_X1 i_0_21_2 (.A(_64data_Enable), .B(n_0_343), .S(n_0_139), .Z(n_0_21_2));
   NAND2_X1 i_0_21_3 (.A1(n_0_21_1), .A2(n_0_21_2), .ZN(n_0_21_3));
   INV_X1 i_0_21_4 (.A(Sending_Enable), .ZN(n_0_21_4));
   OAI21_X1 i_0_21_5 (.A(n_0_21_3), .B1(n_0_21_4), .B2(n_0_21_0), .ZN(n_0_359));
   NAND3_X1 i_0_26_3 (.A1(n_0_155), .A2(n_0_340), .A3(n_0_26_3), .ZN(n_0_26_2));
   INV_X1 i_0_26_4 (.A(n_0_26_9), .ZN(n_0_26_3));
   OAI21_X1 i_0_26_6 (.A(n_0_139), .B1(n_0_155), .B2(T_OR_X[0]), .ZN(n_0_26_5));
   AOI21_X1 i_0_26_7 (.A(n_0_26_7), .B1(n_0_156), .B2(n_0_141), .ZN(n_0_26_6));
   INV_X1 i_0_26_8 (.A(n_0_155), .ZN(n_0_26_7));
   OAI21_X1 i_0_26_9 (.A(n_0_26_9), .B1(n_0_26_0), .B2(n_0_139), .ZN(n_0_26_8));
   NAND3_X1 i_0_26_10 (.A1(n_0_343), .A2(n_0_26_10), .A3(n_0_139), .ZN(n_0_26_9));
   INV_X1 i_0_26_11 (.A(Partial_Data_Count[0]), .ZN(n_0_26_10));
   INV_X1 i_0_26_12 (.A(T_OR_X_Enable), .ZN(n_0_26_0));
   OAI21_X1 i_0_26_0 (.A(n_0_26_8), .B1(n_0_26_6), .B2(n_0_26_5), .ZN(n_0_26_1));
   INV_X1 i_0_26_1 (.A(Sending_Enable), .ZN(n_0_26_4));
   OAI21_X1 i_0_26_2 (.A(n_0_26_1), .B1(n_0_26_4), .B2(n_0_26_2), .ZN(n_0_364));
   NAND2_X1 i_0_18_2 (.A1(RAM_Address_A[0]), .A2(n_0_18_2), .ZN(n_0_18_1));
   INV_X1 i_0_18_4 (.A(T_OR_X[0]), .ZN(n_0_18_0));
   AOI22_X1 i_0_18_6 (.A1(n_0_142), .A2(T_OR_X[0]), .B1(n_0_140), .B2(n_0_18_0), 
      .ZN(n_0_18_3));
   INV_X1 i_0_18_0 (.A(n_0_18_1), .ZN(n_0_18_4));
   INV_X1 i_0_18_1 (.A(n_0_18_3), .ZN(n_0_18_5));
   INV_X1 i_0_18_3 (.A(n_0_139), .ZN(n_0_18_2));
   NAND2_X1 i_0_18_5 (.A1(n_0_18_7), .A2(n_0_18_6), .ZN(n_0_365));
   AOI21_X1 i_0_18_7 (.A(n_0_18_4), .B1(n_0_18_5), .B2(n_0_139), .ZN(n_0_18_6));
   NAND2_X1 i_0_18_8 (.A1(Sending_Enable), .A2(n_0_18_8), .ZN(n_0_18_7));
   INV_X1 i_0_18_9 (.A(n_0_18_9), .ZN(n_0_18_8));
   NAND2_X1 i_0_18_10 (.A1(n_0_340), .A2(n_0_139), .ZN(n_0_18_9));
   DFF_X1 T_OR_X_Enable_reg (.D(n_0_364), .CK(n_0_137), .Q(T_OR_X_Enable), .QN());
   DFF_X2 Done_Sending_reg (.D(n_0_157), .CK(n_0_137), .Q(Done_Sending), .QN());
   DFF_X1 _64data_Enable_reg (.D(n_0_359), .CK(n_0_137), .Q(_64data_Enable), 
      .QN());
   DFF_X1 T_Count_Enable_reg (.D(n_0_345), .CK(n_0_137), .Q(T_Count_Enable), 
      .QN());
   DFF_X1 X_Count_Enable_reg (.D(n_0_346), .CK(n_0_137), .Q(X_Count_Enable), 
      .QN());
   DFF_X1 Init_Count_Enable_reg (.D(n_0_138), .CK(n_0_137), .Q(Init_Count_Enable), 
      .QN());
   DFF_X1 \RAM_Address_A_reg[11]  (.D(n_0_348), .CK(n_0_137), .Q(
      RAM_Address_A[11]), .QN());
   DFF_X1 \RAM_Address_A_reg[10]  (.D(n_0_349), .CK(n_0_137), .Q(
      RAM_Address_A[10]), .QN());
   DFF_X1 \RAM_Address_A_reg[12]  (.D(n_0_347), .CK(n_0_137), .Q(
      RAM_Address_A[12]), .QN());
   DFF_X1 \RAM_Address_A_reg[7]  (.D(n_0_352), .CK(n_0_137), .Q(RAM_Address_A[7]), 
      .QN());
   DFF_X1 \RAM_Address_A_reg[6]  (.D(n_0_353), .CK(n_0_137), .Q(RAM_Address_A[6]), 
      .QN());
   DFF_X1 \RAM_Address_A_reg[5]  (.D(n_0_354), .CK(n_0_137), .Q(RAM_Address_A[5]), 
      .QN());
   DFF_X1 \RAM_Address_A_reg[4]  (.D(n_0_355), .CK(n_0_137), .Q(RAM_Address_A[4]), 
      .QN());
   DFF_X1 \RAM_Address_A_reg[3]  (.D(n_0_356), .CK(n_0_137), .Q(RAM_Address_A[3]), 
      .QN());
   DFF_X1 \RAM_Address_A_reg[2]  (.D(n_0_357), .CK(n_0_137), .Q(RAM_Address_A[2]), 
      .QN());
   DFF_X1 \RAM_Address_A_reg[1]  (.D(n_0_358), .CK(n_0_137), .Q(RAM_Address_A[1]), 
      .QN());
   DFF_X1 \RAM_Address_A_reg[9]  (.D(n_0_350), .CK(n_0_137), .Q(RAM_Address_A[9]), 
      .QN());
   DFF_X1 \RAM_Address_A_reg[8]  (.D(n_0_351), .CK(n_0_137), .Q(RAM_Address_A[8]), 
      .QN());
   DFF_X1 \RAM_Address_A_reg[0]  (.D(n_0_365), .CK(n_0_137), .Q(RAM_Address_A[0]), 
      .QN());
endmodule
