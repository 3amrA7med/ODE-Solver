/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Apr 24 21:28:52 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3015471426 */

module add_sub_cs(sub, in1, in2, cin, out, cout, invalid);
   input sub;
   input [15:0]in1;
   input [15:0]in2;
   input cin;
   output [15:0]out;
   output cout;
   output invalid;

   wire n_0_11_0;
   wire n_0_11_1;
   wire n_0_11_2;
   wire n_0_11_3;
   wire n_0_11_4;
   wire n_0_117;
   wire n_0_47_0;
   wire n_0_47_1;
   wire n_0_47_2;
   wire n_0_47_3;
   wire n_0_43;
   wire n_0_32_0;
   wire n_0_32_1;
   wire n_0_0;
   wire n_0_13_0;
   wire n_0_13_1;
   wire n_0_13_2;
   wire n_0_51;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_67_0;
   wire n_0_67_1;
   wire n_0_67_2;
   wire n_0_67_3;
   wire n_0_5;
   wire n_0_6;
   wire n_0_69_0;
   wire n_0_69_1;
   wire n_0_69_2;
   wire n_0_69_3;
   wire n_0_7;
   wire n_0_70_0;
   wire n_0_70_1;
   wire n_0_70_2;
   wire n_0_70_3;
   wire n_0_8;
   wire n_0_43_0;
   wire n_0_43_1;
   wire n_0_10;
   wire n_0_45_0;
   wire n_0_45_1;
   wire n_0_11;
   wire n_0_56_0;
   wire n_0_56_1;
   wire n_0_12;
   wire n_0_17_0;
   wire n_0_17_1;
   wire n_0_14;
   wire n_0_55;
   wire n_0_56;
   wire n_0_29_0;
   wire n_0_29_1;
   wire n_0_29_2;
   wire n_0_57;
   wire n_0_51_0;
   wire n_0_51_1;
   wire n_0_51_2;
   wire n_0_61;
   wire n_0_62;
   wire n_0_64;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_97_0;
   wire n_0_97_1;
   wire n_0_97_2;
   wire n_0_72;
   wire n_0_97_3;
   wire n_0_73;
   wire n_0_74;
   wire n_0_76;
   wire n_0_77;
   wire n_0_79;
   wire n_0_80;
   wire n_0_97_4;
   wire n_0_97_5;
   wire n_0_97_6;
   wire n_0_97_7;
   wire n_0_97_8;
   wire n_0_97_9;
   wire n_0_97_10;
   wire n_0_97_11;
   wire n_0_75;
   wire n_0_78;
   wire n_0_6_0;
   wire n_0_6_1;
   wire n_0_6_2;
   wire n_0_96;
   wire n_0_50_0;
   wire n_0_50_1;
   wire n_0_50_2;
   wire n_0_50_3;
   wire n_0_50_4;
   wire n_0_50_5;
   wire n_0_50_6;
   wire n_0_97;
   wire n_0_84_4;
   wire n_0_101;
   wire n_0_84_0;
   wire n_0_84_1;
   wire n_0_84_2;
   wire n_0_84_3;
   wire n_0_84_5;
   wire n_0_84_6;
   wire n_0_84_7;
   wire n_0_84_8;
   wire n_0_101_0;
   wire n_0_101_1;
   wire n_0_102;
   wire n_0_109;
   wire n_0_5_0;
   wire n_0_5_1;
   wire n_0_5_6;
   wire n_0_5_2;
   wire n_0_5_5;
   wire n_0_5_8;
   wire n_0_5_3;
   wire n_0_5_4;
   wire n_0_5_7;
   wire n_0_7_0;
   wire n_0_7_6;
   wire n_0_7_13;
   wire n_0_7_1;
   wire n_0_7_2;
   wire n_0_7_3;
   wire n_0_7_4;
   wire n_0_7_5;
   wire n_0_7_7;
   wire n_0_7_8;
   wire n_0_7_9;
   wire n_0_7_10;
   wire n_0_7_11;
   wire n_0_7_12;
   wire n_0_7_19;
   wire n_0_7_14;
   wire n_0_7_15;
   wire n_0_7_16;
   wire n_0_7_17;
   wire n_0_7_18;
   wire n_0_7_34;
   wire n_0_7_20;
   wire n_0_7_21;
   wire n_0_7_22;
   wire n_0_7_23;
   wire n_0_7_24;
   wire n_0_7_25;
   wire n_0_7_26;
   wire n_0_7_27;
   wire n_0_7_28;
   wire n_0_7_29;
   wire n_0_7_30;
   wire n_0_7_31;
   wire n_0_7_32;
   wire n_0_7_33;
   wire n_0_7_38;
   wire n_0_7_35;
   wire n_0_7_36;
   wire n_0_7_37;
   wire n_0_7_39;
   wire n_0_7_40;
   wire n_0_7_41;
   wire n_0_7_43;
   wire n_0_7_45;
   wire n_0_7_44;
   wire n_0_7_48;
   wire n_0_7_49;
   wire n_0_7_50;
   wire n_0_7_51;
   wire n_0_7_52;
   wire n_0_7_55;
   wire n_0_7_53;
   wire n_0_7_57;
   wire n_0_7_58;
   wire n_0_7_59;
   wire n_0_7_60;
   wire n_0_7_61;
   wire n_0_7_54;
   wire n_0_7_64;
   wire n_0_7_65;
   wire n_0_7_56;
   wire n_0_7_70;
   wire n_0_7_62;
   wire n_0_7_73;
   wire n_0_7_74;
   wire n_0_7_75;
   wire n_0_7_76;
   wire n_0_7_77;
   wire n_0_7_63;
   wire n_0_7_80;
   wire n_0_7_81;
   wire n_0_7_82;
   wire n_0_7_83;
   wire n_0_7_84;
   wire n_0_7_85;
   wire n_0_7_86;
   wire n_0_7_87;
   wire n_0_7_88;
   wire n_0_7_89;
   wire n_0_7_90;
   wire n_0_7_92;
   wire n_0_7_93;
   wire n_0_7_94;
   wire n_0_7_95;
   wire n_0_7_96;
   wire n_0_7_97;
   wire n_0_7_98;
   wire n_0_7_99;
   wire n_0_7_100;
   wire n_0_7_101;
   wire n_0_7_102;
   wire n_0_7_103;
   wire n_0_7_104;
   wire n_0_7_105;
   wire n_0_7_66;
   wire n_0_7_108;
   wire n_0_7_109;
   wire n_0_7_110;
   wire n_0_7_111;
   wire n_0_7_112;
   wire n_0_7_113;
   wire n_0_7_114;
   wire n_0_7_115;
   wire n_0_7_116;
   wire n_0_7_117;
   wire n_0_7_118;
   wire n_0_7_119;
   wire n_0_7_120;
   wire n_0_7_121;
   wire n_0_7_122;
   wire n_0_7_123;
   wire n_0_7_124;
   wire n_0_7_125;
   wire n_0_7_126;
   wire n_0_7_127;
   wire n_0_7_128;
   wire n_0_7_129;
   wire n_0_7_130;
   wire n_0_7_131;
   wire n_0_7_133;
   wire n_0_7_134;
   wire n_0_7_135;
   wire n_0_7_136;
   wire n_0_7_67;
   wire n_0_7_138;
   wire n_0_7_139;
   wire n_0_7_140;
   wire n_0_7_141;
   wire n_0_7_142;
   wire n_0_7_143;
   wire n_0_7_144;
   wire n_0_7_145;
   wire n_0_7_146;
   wire n_0_7_147;
   wire n_0_7_68;
   wire n_0_7_151;
   wire n_0_7_152;
   wire n_0_7_153;
   wire n_0_7_154;
   wire n_0_7_155;
   wire n_0_7_156;
   wire n_0_7_157;
   wire n_0_7_158;
   wire n_0_7_159;
   wire n_0_7_160;
   wire n_0_7_162;
   wire n_0_7_163;
   wire n_0_7_69;
   wire n_0_7_165;
   wire n_0_7_166;
   wire n_0_7_78;
   wire n_0_7_79;
   wire n_0_7_91;
   wire n_0_7_106;
   wire n_0_7_107;
   wire n_0_7_132;
   wire n_0_7_137;
   wire n_0_7_148;
   wire n_0_7_149;
   wire n_0_7_150;
   wire n_0_7_161;
   wire n_0_7_164;
   wire n_0_7_167;
   wire n_0_7_168;
   wire n_0_7_46;
   wire n_0_7_71;
   wire n_0_7_72;
   wire n_0_7_169;
   wire n_0_7_170;
   wire n_0_7_42;
   wire n_0_7_47;
   wire n_0_7_171;
   wire n_0_18;
   wire n_0_3_0;
   wire n_0_3_1;
   wire n_0_3_2;
   wire n_0_3_3;
   wire n_0_65;
   wire n_0_67;
   wire n_0_20_0;
   wire n_0_95;
   wire n_0_20_1;
   wire n_0_99;
   wire n_0_20_2;
   wire n_0_20_3;
   wire n_0_98;
   wire n_0_20_4;
   wire n_0_20_5;
   wire n_0_20_6;
   wire n_0_20_7;
   wire n_0_20_8;
   wire n_0_20_9;
   wire n_0_20_10;
   wire n_0_20_11;
   wire n_0_20_12;
   wire n_0_100;
   wire n_0_18_0;
   wire n_0_18_1;
   wire n_0_18_2;
   wire n_0_18_3;
   wire n_0_18_4;
   wire n_0_18_5;
   wire n_0_18_6;
   wire n_0_18_7;
   wire n_0_103;
   wire n_0_25_0;
   wire n_0_25_1;
   wire n_0_25_2;
   wire n_0_25_3;
   wire n_0_111;
   wire n_0_25_4;
   wire n_0_116;
   wire n_0_25_5;
   wire n_0_25_6;
   wire n_0_112;
   wire n_0_110;
   wire n_0_108;
   wire n_0_25_7;
   wire n_0_107;
   wire n_0_25_8;
   wire n_0_25_9;
   wire n_0_25_10;
   wire n_0_25_11;
   wire n_0_25_12;
   wire n_0_25_13;
   wire n_0_25_14;
   wire n_0_106;
   wire n_0_25_15;
   wire n_0_23_0;
   wire n_0_23_1;
   wire n_0_13;
   wire n_0_23_2;
   wire n_0_23_3;
   wire n_0_9;
   wire n_0_130;
   wire n_0_128;
   wire n_0_23_4;
   wire n_0_125;
   wire n_0_23_5;
   wire n_0_23_6;
   wire n_0_23_7;
   wire n_0_23_8;
   wire n_0_23_9;
   wire n_0_23_10;
   wire n_0_23_11;
   wire n_0_23_12;
   wire n_0_120;
   wire n_0_23_13;
   wire n_0_23_14;
   wire n_0_1;
   wire n_0_23_15;
   wire n_0_2_0;
   wire n_0_2_1;
   wire n_0_2_2;
   wire n_0_2_3;
   wire n_0_2_4;
   wire n_0_2_5;
   wire n_0_2_6;
   wire n_0_2_7;
   wire n_0_2_8;
   wire n_0_2_9;
   wire n_0_2_10;
   wire n_0_20;
   wire n_0_2_11;
   wire n_0_2_12;
   wire n_0_19;
   wire n_0_15;
   wire n_0_16;
   wire n_0_2_13;
   wire n_0_2_14;
   wire n_0_2_15;
   wire n_0_2_16;
   wire n_0_2_17;
   wire n_0_17;
   wire n_0_8_49;
   wire n_0_8_50;
   wire n_0_8_0;
   wire n_0_8_51;
   wire n_0_8_2;
   wire n_0_8_57;
   wire n_0_8_61;
   wire n_0_8_6;
   wire n_0_8_7;
   wire n_0_8_8;
   wire n_0_8_9;
   wire n_0_8_12;
   wire n_0_8_62;
   wire n_0_8_14;
   wire n_0_8_77;
   wire n_0_8_78;
   wire n_0_91;
   wire n_0_8_18;
   wire n_0_88;
   wire n_0_8_19;
   wire n_0_87;
   wire n_0_8_20;
   wire n_0_8_21;
   wire n_0_86;
   wire n_0_8_22;
   wire n_0_85;
   wire n_0_8_26;
   wire n_0_8_31;
   wire n_0_92;
   wire n_0_8_33;
   wire n_0_8_87;
   wire n_0_8_95;
   wire n_0_127;
   wire n_0_8_99;
   wire n_0_8_100;
   wire n_0_54;
   wire n_0_8_1;
   wire n_0_8_3;
   wire n_0_8_4;
   wire n_0_8_5;
   wire n_0_8_10;
   wire n_0_8_11;
   wire n_0_124;
   wire n_0_8_13;
   wire n_0_8_16;
   wire n_0_8_102;
   wire n_0_8_15;
   wire n_0_8_103;
   wire n_0_122;
   wire n_0_8_17;
   wire n_0_8_23;
   wire n_0_113;
   wire n_0_8_24;
   wire n_0_8_25;
   wire n_0_8_27;
   wire n_0_8_28;
   wire n_0_123;
   wire n_0_8_29;
   wire n_0_8_30;
   wire n_0_8_580;
   wire n_0_8_32;
   wire n_0_8_110;
   wire n_0_8_34;
   wire n_0_8_35;
   wire n_0_8_595;
   wire n_0_8_36;
   wire n_0_119;
   wire n_0_8_37;
   wire n_0_8_38;
   wire n_0_121;
   wire n_0_8_39;
   wire n_0_8_40;
   wire n_0_35;
   wire n_0_8_63;
   wire n_0_8_64;
   wire n_0_8_65;
   wire n_0_8_66;
   wire n_0_38;
   wire n_0_8_67;
   wire n_0_8_68;
   wire n_0_8_69;
   wire n_0_8_70;
   wire n_0_39;
   wire n_0_8_71;
   wire n_0_8_72;
   wire n_0_8_73;
   wire n_0_8_74;
   wire n_0_8_41;
   wire n_0_8_42;
   wire n_0_50;
   wire n_0_8_43;
   wire n_0_37;
   wire n_0_8_44;
   wire n_0_44;
   wire n_0_8_45;
   wire n_0_58;
   wire n_0_8_150;
   wire n_0_8_46;
   wire n_0_8_587;
   wire n_0_8_588;
   wire n_0_8_155;
   wire n_0_8_47;
   wire n_0_8_48;
   wire n_0_8_175;
   wire n_0_8_189;
   wire n_0_46;
   wire n_0_8_52;
   wire n_0_8_53;
   wire n_0_47;
   wire n_0_8_54;
   wire n_0_8_55;
   wire n_0_48;
   wire n_0_8_56;
   wire n_0_8_232;
   wire n_0_8_85;
   wire n_0_8_86;
   wire n_0_32;
   wire n_0_8_88;
   wire n_0_8_89;
   wire n_0_8_90;
   wire n_0_8_91;
   wire n_0_8_58;
   wire n_0_8_92;
   wire n_0_8_59;
   wire n_0_8_60;
   wire n_0_8_93;
   wire n_0_8_233;
   wire n_0_8_234;
   wire n_0_8_94;
   wire n_0_8_75;
   wire n_0_8_76;
   wire n_0_8_235;
   wire n_0_8_96;
   wire n_0_8_79;
   wire n_0_8_97;
   wire n_0_8_98;
   wire n_0_8_101;
   wire n_0_8_107;
   wire n_0_8_80;
   wire n_0_8_109;
   wire n_0_8_81;
   wire n_0_8_82;
   wire n_0_8_83;
   wire n_0_8_84;
   wire n_0_8_243;
   wire n_0_8_245;
   wire n_0_8_249;
   wire n_0_8_104;
   wire n_0_8_111;
   wire n_0_8_112;
   wire n_0_8_114;
   wire n_0_8_115;
   wire n_0_8_116;
   wire n_0_8_117;
   wire n_0_8_118;
   wire n_0_8_119;
   wire n_0_8_121;
   wire n_0_8_122;
   wire n_0_8_123;
   wire n_0_8_124;
   wire n_0_8_125;
   wire n_0_8_126;
   wire n_0_8_127;
   wire n_0_8_128;
   wire n_0_8_129;
   wire n_0_8_130;
   wire n_0_8_131;
   wire n_0_8_132;
   wire n_0_8_133;
   wire n_0_8_134;
   wire n_0_8_135;
   wire n_0_8_136;
   wire n_0_8_137;
   wire n_0_8_138;
   wire n_0_8_139;
   wire n_0_8_140;
   wire n_0_8_143;
   wire n_0_8_144;
   wire n_0_8_105;
   wire n_0_8_250;
   wire n_0_8_589;
   wire n_0_8_106;
   wire n_0_8_169;
   wire n_0_8_108;
   wire n_0_8_113;
   wire n_0_8_120;
   wire n_0_8_590;
   wire n_0_8_591;
   wire n_0_8_172;
   wire n_0_8_148;
   wire n_0_8_157;
   wire n_0_8_158;
   wire n_0_8_141;
   wire n_0_8_170;
   wire n_0_8_171;
   wire n_0_8_146;
   wire n_0_8_600;
   wire n_0_8_601;
   wire n_0_8_177;
   wire n_0_8_142;
   wire n_0_8_182;
   wire n_0_8_183;
   wire n_0_8_145;
   wire n_0_8_185;
   wire n_0_8_147;
   wire n_0_8_188;
   wire n_0_8_251;
   wire n_0_8_190;
   wire n_0_8_191;
   wire n_0_8_149;
   wire n_0_8_151;
   wire n_0_8_152;
   wire n_0_8_592;
   wire n_0_8_593;
   wire n_0_8_153;
   wire n_0_8_154;
   wire n_0_8_258;
   wire n_0_8_156;
   wire n_0_8_159;
   wire n_0_8_160;
   wire n_0_8_163;
   wire n_0_8_164;
   wire n_0_8_161;
   wire n_0_8_162;
   wire n_0_8_165;
   wire n_0_8_166;
   wire n_0_45;
   wire n_0_8_167;
   wire n_0_8_168;
   wire n_0_8_173;
   wire n_0_8_174;
   wire n_0_8_179;
   wire n_0_8_180;
   wire n_0_8_181;
   wire n_0_8_184;
   wire n_0_8_186;
   wire n_0_8_187;
   wire n_0_49;
   wire n_0_8_192;
   wire n_0_8_193;
   wire n_0_8_194;
   wire n_0_8_195;
   wire n_0_8_196;
   wire n_0_8_197;
   wire n_0_8_198;
   wire n_0_8_199;
   wire n_0_8_200;
   wire n_0_8_201;
   wire n_0_60;
   wire n_0_8_202;
   wire n_0_8_203;
   wire n_0_8_204;
   wire n_0_8_205;
   wire n_0_8_206;
   wire n_0_8_207;
   wire n_0_8_208;
   wire n_0_93;
   wire n_0_8_209;
   wire n_0_8_210;
   wire n_0_8_211;
   wire n_0_8_212;
   wire n_0_8_213;
   wire n_0_8_214;
   wire n_0_8_215;
   wire n_0_8_261;
   wire n_0_8_176;
   wire n_0_8_178;
   wire n_0_53;
   wire n_0_8_216;
   wire n_0_8_217;
   wire n_0_8_218;
   wire n_0_8_219;
   wire n_0_8_220;
   wire n_0_8_221;
   wire n_0_8_222;
   wire n_0_8_223;
   wire n_0_8_224;
   wire n_0_8_225;
   wire n_0_8_226;
   wire n_0_8_227;
   wire n_0_8_228;
   wire n_0_8_229;
   wire n_0_8_230;
   wire n_0_8_231;
   wire n_0_8_262;
   wire n_0_8_263;
   wire n_0_8_236;
   wire n_0_8_237;
   wire n_0_8_238;
   wire n_0_8_268;
   wire n_0_8_239;
   wire n_0_26;
   wire n_0_8_240;
   wire n_0_27;
   wire n_0_8_241;
   wire n_0_29;
   wire n_0_8_242;
   wire n_0_24;
   wire n_0_41;
   wire n_0_8_244;
   wire n_0_8_276;
   wire n_0_8_594;
   wire n_0_8_286;
   wire n_0_8_287;
   wire n_0_8_246;
   wire n_0_8_247;
   wire n_0_8_248;
   wire n_0_8_292;
   wire n_0_8_294;
   wire n_0_8_309;
   wire n_0_8_252;
   wire n_0_8_253;
   wire n_0_8_254;
   wire n_0_8_255;
   wire n_0_8_256;
   wire n_0_8_257;
   wire n_0_8_315;
   wire n_0_8_316;
   wire n_0_8_259;
   wire n_0_8_260;
   wire n_0_8_320;
   wire n_0_8_321;
   wire n_0_8_264;
   wire n_0_8_265;
   wire n_0_8_266;
   wire n_0_8_267;
   wire n_0_8_342;
   wire n_0_8_269;
   wire n_0_8_270;
   wire n_0_8_271;
   wire n_0_8_272;
   wire n_0_8_273;
   wire n_0_8_274;
   wire n_0_8_275;
   wire n_0_8_343;
   wire n_0_8_277;
   wire n_0_8_278;
   wire n_0_8_279;
   wire n_0_8_280;
   wire n_0_8_281;
   wire n_0_8_282;
   wire n_0_8_283;
   wire n_0_8_284;
   wire n_0_8_285;
   wire n_0_8_344;
   wire n_0_8_345;
   wire n_0_8_288;
   wire n_0_8_289;
   wire n_0_8_291;
   wire n_0_8_347;
   wire n_0_8_295;
   wire n_0_8_296;
   wire n_0_8_297;
   wire n_0_8_298;
   wire n_0_8_299;
   wire n_0_8_300;
   wire n_0_8_301;
   wire n_0_8_302;
   wire n_0_8_303;
   wire n_0_8_304;
   wire n_0_8_305;
   wire n_0_8_306;
   wire n_0_28;
   wire n_0_8_307;
   wire n_0_8_308;
   wire n_0_8_310;
   wire n_0_8_311;
   wire n_0_8_312;
   wire n_0_8_313;
   wire n_0_8_314;
   wire n_0_8_348;
   wire n_0_8_317;
   wire n_0_8_318;
   wire n_0_8_319;
   wire n_0_8_322;
   wire n_0_8_323;
   wire n_0_8_324;
   wire n_0_8_325;
   wire n_0_8_326;
   wire n_0_8_327;
   wire n_0_8_328;
   wire n_0_8_329;
   wire n_0_8_330;
   wire n_0_8_331;
   wire n_0_8_332;
   wire n_0_8_333;
   wire n_0_8_334;
   wire n_0_8_335;
   wire n_0_8_336;
   wire n_0_8_337;
   wire n_0_8_338;
   wire n_0_8_339;
   wire n_0_8_340;
   wire n_0_8_361;
   wire n_0_8_341;
   wire n_0_8_362;
   wire n_0_8_372;
   wire n_0_8_597;
   wire n_0_8_373;
   wire n_0_8_374;
   wire n_0_8_346;
   wire n_0_8_375;
   wire n_0_8_376;
   wire n_0_8_349;
   wire n_0_8_350;
   wire n_0_8_351;
   wire n_0_8_352;
   wire n_0_8_353;
   wire n_0_8_354;
   wire n_0_8_355;
   wire n_0_8_356;
   wire n_0_8_357;
   wire n_0_8_358;
   wire n_0_8_359;
   wire n_0_8_360;
   wire n_0_8_377;
   wire n_0_8_363;
   wire n_0_8_364;
   wire n_0_8_365;
   wire n_0_8_634;
   wire n_0_8_366;
   wire n_0_8_367;
   wire n_0_8_368;
   wire n_0_8_369;
   wire n_0_8_370;
   wire n_0_8_371;
   wire n_0_8_635;
   wire n_0_8_378;
   wire n_0_8_383;
   wire n_0_8_390;
   wire n_0_8_391;
   wire n_0_8_393;
   wire n_0_8_379;
   wire n_0_8_380;
   wire n_0_8_381;
   wire n_0_8_382;
   wire n_0_8_638;
   wire n_0_8_639;
   wire n_0_8_400;
   wire n_0_8_384;
   wire n_0_8_385;
   wire n_0_8_386;
   wire n_0_8_640;
   wire n_0_8_387;
   wire n_0_8_388;
   wire n_0_8_389;
   wire n_0_8_641;
   wire n_0_8_642;
   wire n_0_8_403;
   wire n_0_8_404;
   wire n_0_8_392;
   wire n_0_8_405;
   wire n_0_8_394;
   wire n_0_8_395;
   wire n_0_8_396;
   wire n_0_8_397;
   wire n_0_8_398;
   wire n_0_8_399;
   wire n_0_8_406;
   wire n_0_8_401;
   wire n_0_8_402;
   wire n_0_8_414;
   wire n_0_8_455;
   wire n_0_8_407;
   wire n_0_8_408;
   wire n_0_8_409;
   wire n_0_8_410;
   wire n_0_8_411;
   wire n_0_8_412;
   wire n_0_8_485;
   wire n_0_8_413;
   wire n_0_8_415;
   wire n_0_8_416;
   wire n_0_8_417;
   wire n_0_8_418;
   wire n_0_8_419;
   wire n_0_8_420;
   wire n_0_8_421;
   wire n_0_36;
   wire n_0_8_422;
   wire n_0_8_423;
   wire n_0_8_424;
   wire n_0_8_425;
   wire n_0_8_426;
   wire n_0_8_427;
   wire n_0_8_428;
   wire n_0_8_429;
   wire n_0_8_430;
   wire n_0_8_431;
   wire n_0_8_432;
   wire n_0_8_433;
   wire n_0_8_434;
   wire n_0_8_435;
   wire n_0_8_436;
   wire n_0_8_437;
   wire n_0_8_438;
   wire n_0_8_439;
   wire n_0_8_440;
   wire n_0_8_441;
   wire n_0_8_442;
   wire n_0_8_443;
   wire n_0_8_444;
   wire n_0_8_445;
   wire n_0_33;
   wire n_0_8_644;
   wire n_0_8_446;
   wire n_0_8_447;
   wire n_0_8_448;
   wire n_0_8_449;
   wire n_0_8_450;
   wire n_0_8_451;
   wire n_0_8_452;
   wire n_0_8_453;
   wire n_0_8_454;
   wire n_0_8_456;
   wire n_0_8_457;
   wire n_0_8_458;
   wire n_0_8_459;
   wire n_0_8_460;
   wire n_0_8_464;
   wire n_0_8_465;
   wire n_0_8_466;
   wire n_0_8_467;
   wire n_0_8_468;
   wire n_0_8_469;
   wire n_0_8_470;
   wire n_0_8_471;
   wire n_0_8_472;
   wire n_0_8_473;
   wire n_0_8_474;
   wire n_0_8_475;
   wire n_0_8_476;
   wire n_0_8_477;
   wire n_0_8_700;
   wire n_0_8_479;
   wire n_0_8_480;
   wire n_0_8_481;
   wire n_0_30;
   wire n_0_8_482;
   wire n_0_8_483;
   wire n_0_8_484;
   wire n_0_8_486;
   wire n_0_8_487;
   wire n_0_8_492;
   wire n_0_8_488;
   wire n_0_8_604;
   wire n_0_8_495;
   wire n_0_8_496;
   wire n_0_8_497;
   wire n_0_8_498;
   wire n_0_8_499;
   wire n_0_8_500;
   wire n_0_8_501;
   wire n_0_8_489;
   wire n_0_8_503;
   wire n_0_8_493;
   wire n_0_8_502;
   wire n_0_8_702;
   wire n_0_8_511;
   wire n_0_8_513;
   wire n_0_8_514;
   wire n_0_8_515;
   wire n_0_8_504;
   wire n_0_8_507;
   wire n_0_8_508;
   wire n_0_8_520;
   wire n_0_8_521;
   wire n_0_8_649;
   wire n_0_8_526;
   wire n_0_8_527;
   wire n_0_8_528;
   wire n_0_8_529;
   wire n_0_8_530;
   wire n_0_8_531;
   wire n_0_8_509;
   wire n_0_8_516;
   wire n_0_8_517;
   wire n_0_8_518;
   wire n_0_8_537;
   wire n_0_8_540;
   wire n_0_8_519;
   wire n_0_8_542;
   wire n_0_8_534;
   wire n_0_8_535;
   wire n_0_8_548;
   wire n_0_8_549;
   wire n_0_8_550;
   wire n_0_8_536;
   wire n_0_8_538;
   wire n_0_8_539;
   wire n_0_8_541;
   wire n_0_8_544;
   wire n_0_8_545;
   wire n_0_8_653;
   wire n_0_8_654;
   wire n_0_8_582;
   wire n_0_8_583;
   wire n_0_8_546;
   wire n_0_8_606;
   wire n_0_8_547;
   wire n_0_8_608;
   wire n_0_8_556;
   wire n_0_8_611;
   wire n_0_8_613;
   wire n_0_8_585;
   wire n_0_8_614;
   wire n_0_8_615;
   wire n_0_8_616;
   wire n_0_8_617;
   wire n_0_8_618;
   wire n_0_8_619;
   wire n_0_8_620;
   wire n_0_8_621;
   wire n_0_8_586;
   wire n_0_8_622;
   wire n_0_8_623;
   wire n_0_8_624;
   wire n_0_8_625;
   wire n_0_8_626;
   wire n_0_8_627;
   wire n_0_8_628;
   wire n_0_8_629;
   wire n_0_8_631;
   wire n_0_8_632;
   wire n_0_8_557;
   wire n_0_8_558;
   wire n_0_8_560;
   wire n_0_8_562;
   wire n_0_8_461;
   wire n_0_8_462;
   wire n_0_8_463;
   wire n_0_8_478;
   wire n_0_8_490;
   wire n_0_8_491;
   wire n_0_8_494;
   wire n_0_8_505;
   wire n_0_8_506;
   wire n_0_8_510;
   wire n_0_8_512;
   wire n_0_8_522;
   wire n_0_8_523;
   wire n_0_8_524;
   wire n_0_8_525;
   wire n_0_8_532;
   wire n_0_8_533;
   wire n_0_8_543;
   wire n_0_8_551;
   wire n_0_8_552;
   wire n_0_8_565;
   wire n_0_8_574;
   wire n_0_8_575;
   wire n_0_8_576;
   wire n_0_8_577;
   wire n_0_8_663;
   wire n_0_8_578;
   wire n_0_8_579;
   wire n_0_8_581;
   wire n_0_8_563;
   wire n_0_8_564;
   wire n_0_8_666;
   wire n_0_8_667;
   wire n_0_8_668;
   wire n_0_8_669;
   wire n_0_8_670;
   wire n_0_8_671;
   wire n_0_8_672;
   wire n_0_8_673;
   wire n_0_8_566;
   wire n_0_8_675;
   wire n_0_8_676;
   wire n_0_8_567;
   wire n_0_8_679;
   wire n_0_8_680;
   wire n_0_8_681;
   wire n_0_8_683;
   wire n_0_8_684;
   wire n_0_8_686;
   wire n_0_8_687;
   wire n_0_8_688;
   wire n_0_8_568;
   wire n_0_8_569;
   wire n_0_8_695;
   wire n_0_34;
   wire n_0_21;
   wire n_0_8_711;
   wire n_0_8_712;
   wire n_0_8_570;
   wire n_0_8_571;
   wire n_0_8_715;
   wire n_0_8_648;
   wire n_0_8_716;
   wire n_0_8_717;
   wire n_0_8_572;
   wire n_0_8_719;
   wire n_0_8_573;
   wire n_0_8_724;
   wire n_0_8_725;
   wire n_0_8_726;
   wire n_0_8_584;
   wire n_0_8_596;
   wire n_0_8_598;
   wire n_0_8_602;
   wire n_0_8_599;
   wire n_0_8_603;
   wire n_0_8_605;
   wire n_0_8_607;
   wire n_0_8_609;
   wire n_0_8_610;
   wire n_0_84;
   wire n_0_42;
   wire n_0_52;
   wire n_0_8_612;
   wire n_0_8_630;
   wire n_0_8_633;
   wire n_0_8_636;
   wire n_0_8_637;
   wire n_0_8_643;
   wire n_0_8_645;
   wire n_0_8_646;
   wire n_0_8_647;
   wire n_0_8_650;
   wire n_0_8_651;
   wire n_0_8_652;
   wire n_0_8_655;
   wire n_0_8_656;
   wire n_0_8_657;
   wire n_0_8_658;
   wire n_0_8_659;
   wire n_0_8_660;
   wire n_0_8_661;
   wire n_0_8_662;
   wire n_0_8_664;
   wire n_0_8_665;
   wire n_0_8_674;
   wire n_0_8_677;
   wire n_0_8_678;
   wire n_0_8_682;
   wire n_0_8_685;
   wire n_0_8_689;
   wire n_0_8_690;
   wire n_0_8_691;
   wire n_0_8_692;
   wire n_0_8_693;
   wire n_0_8_694;
   wire n_0_8_553;
   wire n_0_8_555;
   wire n_0_8_561;
   wire n_0_8_559;
   wire n_0_8_554;
   wire n_0_8_696;
   wire n_0_8_697;
   wire n_0_8_698;
   wire n_0_8_699;
   wire n_0_8_701;
   wire n_0_8_703;
   wire n_0_8_704;
   wire n_0_8_705;
   wire n_0_8_706;
   wire n_0_8_707;
   wire n_0_8_708;
   wire n_0_8_709;
   wire n_0_8_710;
   wire n_0_8_713;
   wire n_0_8_714;
   wire n_0_8_718;
   wire n_0_8_720;
   wire n_0_8_721;
   wire n_0_8_722;
   wire n_0_8_723;
   wire n_0_8_727;
   wire n_0_8_728;
   wire n_0_8_729;
   wire n_0_8_730;
   wire n_0_8_731;
   wire n_0_8_732;
   wire n_0_8_733;
   wire n_0_25;
   wire n_0_8_734;
   wire n_0_8_735;
   wire n_0_8_736;
   wire n_0_8_737;
   wire n_0_8_738;
   wire n_0_8_739;
   wire n_0_59;
   wire n_0_8_740;
   wire n_0_8_741;
   wire n_0_8_742;
   wire n_0_8_743;
   wire n_0_8_744;
   wire n_0_8_745;
   wire n_0_8_746;
   wire n_0_8_747;
   wire n_0_8_748;
   wire n_0_114;
   wire n_0_8_749;
   wire n_0_8_750;
   wire n_0_8_751;
   wire n_0_8_752;
   wire n_0_8_753;
   wire n_0_8_754;
   wire n_0_8_755;
   wire n_0_8_756;
   wire n_0_8_757;
   wire n_0_8_758;
   wire n_0_8_759;
   wire n_0_8_760;
   wire n_0_8_761;
   wire n_0_8_762;
   wire n_0_8_763;
   wire n_0_8_764;
   wire n_0_8_765;
   wire n_0_8_766;
   wire n_0_8_767;
   wire n_0_8_768;
   wire n_0_8_769;
   wire n_0_8_770;
   wire n_0_8_771;
   wire n_0_8_772;
   wire n_0_8_773;
   wire n_0_8_774;
   wire n_0_8_775;
   wire n_0_8_776;
   wire n_0_94;
   wire n_0_8_777;
   wire n_0_8_778;
   wire n_0_8_779;
   wire n_0_8_780;
   wire n_0_8_781;
   wire n_0_8_782;
   wire n_0_8_783;
   wire n_0_8_784;
   wire n_0_40;
   wire n_0_8_785;
   wire n_0_8_786;
   wire n_0_8_787;
   wire n_0_8_788;
   wire n_0_8_789;
   wire n_0_8_790;
   wire n_0_8_791;
   wire n_0_8_792;
   wire n_0_8_793;
   wire n_0_8_794;
   wire n_0_23;
   wire n_0_8_795;
   wire n_0_8_796;
   wire n_0_8_797;
   wire n_0_8_798;
   wire n_0_8_799;
   wire n_0_8_800;
   wire n_0_22;
   wire n_0_8_801;
   wire n_0_8_802;
   wire n_0_63;
   wire n_0_8_803;
   wire n_0_8_804;
   wire n_0_8_805;
   wire n_0_8_806;
   wire n_0_8_807;
   wire n_0_8_808;
   wire n_0_8_809;
   wire n_0_8_810;
   wire n_0_8_811;
   wire n_0_8_812;
   wire n_0_8_290;
   wire n_0_8_293;
   wire n_0_8_813;
   wire n_0_8_814;
   wire n_0_8_815;
   wire n_0_8_816;
   wire n_0_8_817;
   wire n_0_8_818;
   wire n_0_8_819;
   wire n_0_8_820;
   wire n_0_8_821;
   wire n_0_8_822;
   wire n_0_8_823;
   wire n_0_8_824;
   wire n_0_8_825;
   wire n_0_8_826;
   wire n_0_8_827;
   wire n_0_8_828;
   wire n_0_8_829;
   wire n_0_8_830;
   wire n_0_8_831;
   wire n_0_8_832;
   wire n_0_8_833;
   wire n_0_8_834;
   wire n_0_8_835;
   wire n_0_8_836;
   wire n_0_8_837;
   wire n_0_8_838;
   wire n_0_8_839;
   wire n_0_8_840;
   wire n_0_8_841;
   wire n_0_8_842;
   wire n_0_8_843;
   wire n_0_8_844;
   wire n_0_8_845;
   wire n_0_8_846;
   wire n_0_8_847;
   wire n_0_8_848;
   wire n_0_8_849;
   wire n_0_8_850;
   wire n_0_8_851;
   wire n_0_8_852;
   wire n_0_8_853;
   wire n_0_8_854;
   wire n_0_8_855;
   wire n_0_8_856;
   wire n_0_8_857;
   wire n_0_8_858;
   wire n_0_8_859;
   wire n_0_8_860;
   wire n_0_8_861;
   wire n_0_8_862;
   wire n_0_31;
   wire n_0_8_863;
   wire n_0_8_864;
   wire n_0_129;
   wire n_0_83;
   wire n_0_66;
   wire n_0_0_0;
   wire n_0_81;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_89;
   wire n_0_0_6;
   wire n_0_90;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_82;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_1_2;
   wire n_0_1_3;
   wire n_0_1_4;
   wire n_0_1_5;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_1_8;
   wire n_0_1_9;
   wire n_0_1_10;
   wire n_0_126;
   wire n_0_1_11;
   wire n_0_1_12;
   wire n_0_118;
   wire n_0_1_13;
   wire n_0_115;
   wire n_0_104;
   wire n_0_105;
   wire n_0_1_14;
   wire n_0_1_15;
   wire n_0_1_16;
   wire n_0_1_17;
   wire n_0_1_18;
   wire n_0_1_19;

   NAND2_X1 i_0_11_0 (.A1(n_0_11_0), .A2(n_0_11_1), .ZN(out[10]));
   NAND2_X1 i_0_11_1 (.A1(n_0_11_3), .A2(n_0_51), .ZN(n_0_11_0));
   NAND2_X1 i_0_11_2 (.A1(n_0_97), .A2(n_0_71), .ZN(n_0_11_1));
   NAND2_X1 i_0_11_3 (.A1(n_0_11_2), .A2(n_0_11_4), .ZN(out[11]));
   NAND2_X1 i_0_11_4 (.A1(n_0_11_3), .A2(n_0_2), .ZN(n_0_11_2));
   INV_X1 i_0_11_5 (.A(n_0_97), .ZN(n_0_11_3));
   NAND2_X1 i_0_11_6 (.A1(n_0_97), .A2(n_0_3), .ZN(n_0_11_4));
   NAND2_X1 i_0_47_0 (.A1(n_0_47_0), .A2(n_0_47_2), .ZN(n_0_117));
   NAND2_X1 i_0_47_1 (.A1(n_0_47_1), .A2(n_0_44), .ZN(n_0_47_0));
   INV_X1 i_0_47_2 (.A(n_0_105), .ZN(n_0_47_1));
   NAND2_X1 i_0_47_3 (.A1(n_0_105), .A2(n_0_47_3), .ZN(n_0_47_2));
   INV_X1 i_0_47_4 (.A(n_0_44), .ZN(n_0_47_3));
   NAND2_X1 i_0_32_0 (.A1(n_0_32_1), .A2(n_0_32_0), .ZN(n_0_43));
   NAND2_X1 i_0_32_1 (.A1(n_0_105), .A2(n_0_44), .ZN(n_0_32_0));
   NAND2_X1 i_0_32_2 (.A1(n_0_0), .A2(n_0_117), .ZN(n_0_32_1));
   AND2_X1 i_0_63_0 (.A1(n_0_104), .A2(n_0_37), .ZN(n_0_0));
   INV_X1 i_0_13_0 (.A(n_0_96), .ZN(n_0_13_0));
   AOI22_X1 i_0_13_1 (.A1(n_0_13_0), .A2(n_0_74), .B1(n_0_70), .B2(n_0_96), 
      .ZN(n_0_13_1));
   INV_X1 i_0_13_2 (.A(n_0_13_1), .ZN(out[8]));
   AOI22_X1 i_0_13_3 (.A1(n_0_13_0), .A2(n_0_61), .B1(n_0_96), .B2(n_0_62), 
      .ZN(n_0_13_2));
   INV_X1 i_0_13_4 (.A(n_0_13_2), .ZN(out[9]));
   XOR2_X1 i_0_14_0 (.A(n_0_37), .B(n_0_104), .Z(n_0_51));
   XOR2_X1 i_0_15_0 (.A(n_0_117), .B(n_0_0), .Z(n_0_2));
   XOR2_X1 i_0_16_0 (.A(n_0_115), .B(n_0_118), .Z(n_0_3));
   NAND2_X1 i_0_67_0 (.A1(n_0_67_2), .A2(n_0_67_0), .ZN(n_0_4));
   NAND2_X1 i_0_67_1 (.A1(n_0_17), .A2(n_0_67_1), .ZN(n_0_67_0));
   INV_X1 i_0_67_2 (.A(n_0_19), .ZN(n_0_67_1));
   NAND2_X1 i_0_67_3 (.A1(n_0_67_3), .A2(n_0_19), .ZN(n_0_67_2));
   INV_X1 i_0_67_4 (.A(n_0_17), .ZN(n_0_67_3));
   INV_X1 i_0_4_0 (.A(n_0_109), .ZN(n_0_5));
   NAND2_X1 i_0_69_0 (.A1(n_0_69_0), .A2(n_0_69_2), .ZN(n_0_6));
   NAND2_X1 i_0_69_1 (.A1(n_0_69_1), .A2(n_0_58), .ZN(n_0_69_0));
   INV_X1 i_0_69_2 (.A(n_0_16), .ZN(n_0_69_1));
   NAND2_X1 i_0_69_3 (.A1(n_0_16), .A2(n_0_69_3), .ZN(n_0_69_2));
   INV_X1 i_0_69_4 (.A(n_0_58), .ZN(n_0_69_3));
   NAND2_X1 i_0_70_0 (.A1(n_0_70_2), .A2(n_0_70_0), .ZN(n_0_7));
   NAND2_X1 i_0_70_1 (.A1(n_0_6), .A2(n_0_70_1), .ZN(n_0_70_0));
   INV_X1 i_0_70_2 (.A(n_0_64), .ZN(n_0_70_1));
   NAND2_X1 i_0_70_3 (.A1(n_0_70_3), .A2(n_0_64), .ZN(n_0_70_2));
   INV_X1 i_0_70_4 (.A(n_0_6), .ZN(n_0_70_3));
   NAND2_X1 i_0_43_0 (.A1(n_0_43_0), .A2(n_0_43_1), .ZN(n_0_8));
   NAND2_X1 i_0_43_1 (.A1(n_0_119), .A2(n_0_122), .ZN(n_0_43_0));
   NAND2_X1 i_0_43_2 (.A1(n_0_121), .A2(n_0_60), .ZN(n_0_43_1));
   NAND2_X1 i_0_45_0 (.A1(n_0_45_1), .A2(n_0_45_0), .ZN(n_0_10));
   NAND2_X1 i_0_45_1 (.A1(n_0_83), .A2(n_0_49), .ZN(n_0_45_0));
   NAND2_X1 i_0_45_2 (.A1(n_0_66), .A2(n_0_89), .ZN(n_0_45_1));
   NAND2_X1 i_0_56_0 (.A1(n_0_56_1), .A2(n_0_56_0), .ZN(n_0_11));
   NAND2_X1 i_0_56_1 (.A1(n_0_16), .A2(n_0_58), .ZN(n_0_56_0));
   NAND2_X1 i_0_56_2 (.A1(n_0_6), .A2(n_0_64), .ZN(n_0_56_1));
   XOR2_X1 i_0_74_0 (.A(n_0_66), .B(n_0_82), .Z(n_0_12));
   INV_X1 i_0_17_0 (.A(n_0_119), .ZN(n_0_17_0));
   INV_X1 i_0_17_1 (.A(n_0_114), .ZN(n_0_17_1));
   OAI22_X1 i_0_17_2 (.A1(n_0_17_0), .A2(n_0_114), .B1(n_0_17_1), .B2(n_0_119), 
      .ZN(n_0_14));
   OR2_X1 i_0_21_0 (.A1(cin), .A2(sub), .ZN(n_0_55));
   XOR2_X1 i_0_28_0 (.A(n_0_85), .B(n_0_86), .Z(n_0_56));
   INV_X1 i_0_29_0 (.A(n_0_18), .ZN(n_0_29_0));
   AOI22_X1 i_0_29_1 (.A1(n_0_29_0), .A2(n_0_79), .B1(n_0_78), .B2(n_0_18), 
      .ZN(n_0_29_1));
   INV_X1 i_0_29_2 (.A(n_0_29_1), .ZN(out[4]));
   AOI22_X1 i_0_29_3 (.A1(n_0_29_0), .A2(n_0_80), .B1(n_0_18), .B2(n_0_56), 
      .ZN(n_0_29_2));
   INV_X1 i_0_29_4 (.A(n_0_29_2), .ZN(out[5]));
   XOR2_X1 i_0_31_0 (.A(n_0_125), .B(n_0_128), .Z(n_0_57));
   INV_X1 i_0_51_0 (.A(n_0_92), .ZN(n_0_51_0));
   AOI22_X1 i_0_51_1 (.A1(n_0_51_0), .A2(n_0_76), .B1(n_0_75), .B2(n_0_92), 
      .ZN(n_0_51_1));
   INV_X1 i_0_51_2 (.A(n_0_51_1), .ZN(out[6]));
   AOI22_X1 i_0_51_3 (.A1(n_0_51_0), .A2(n_0_77), .B1(n_0_92), .B2(n_0_57), 
      .ZN(n_0_51_2));
   INV_X1 i_0_51_4 (.A(n_0_51_2), .ZN(out[7]));
   XOR2_X1 i_0_52_0 (.A(n_0_107), .B(n_0_112), .Z(n_0_61));
   XOR2_X1 i_0_54_0 (.A(n_0_107), .B(n_0_108), .Z(n_0_62));
   OR2_X1 i_0_72_0 (.A1(n_0_15), .A2(n_0_53), .ZN(n_0_64));
   XOR2_X1 i_0_89_0 (.A(n_0_93), .B(n_0_65), .Z(n_0_68));
   INV_X1 i_0_94_0 (.A(n_0_68), .ZN(n_0_69));
   INV_X1 i_0_95_0 (.A(n_0_110), .ZN(n_0_70));
   INV_X1 i_0_96_0 (.A(n_0_51), .ZN(n_0_71));
   NAND2_X1 i_0_97_0 (.A1(in1[12]), .A2(n_0_67), .ZN(n_0_97_0));
   INV_X1 i_0_97_1 (.A(n_0_97_0), .ZN(n_0_97_1));
   OAI22_X1 i_0_97_2 (.A1(n_0_97_1), .A2(n_0_95), .B1(in1[12]), .B2(n_0_67), 
      .ZN(n_0_97_2));
   INV_X1 i_0_97_3 (.A(n_0_97_2), .ZN(n_0_72));
   NAND2_X1 i_0_97_4 (.A1(n_0_98), .A2(n_0_102), .ZN(n_0_97_3));
   NAND2_X1 i_0_97_5 (.A1(n_0_97_0), .A2(n_0_97_3), .ZN(n_0_73));
   XOR2_X1 i_0_97_6 (.A(n_0_48), .B(n_0_111), .Z(n_0_74));
   XOR2_X1 i_0_97_7 (.A(n_0_46), .B(n_0_1), .Z(n_0_76));
   XOR2_X1 i_0_97_8 (.A(n_0_9), .B(n_0_125), .Z(n_0_77));
   XOR2_X1 i_0_97_9 (.A(n_0_42), .B(n_0_88), .Z(n_0_79));
   XOR2_X1 i_0_97_10 (.A(n_0_91), .B(n_0_85), .Z(n_0_80));
   XOR2_X1 i_0_97_11 (.A(n_0_55), .B(n_0_35), .Z(out[0]));
   XOR2_X1 i_0_97_12 (.A(n_0_38), .B(n_0_39), .Z(out[1]));
   XNOR2_X1 i_0_97_13 (.A(n_0_124), .B(n_0_129), .ZN(n_0_97_4));
   INV_X1 i_0_97_14 (.A(n_0_52), .ZN(n_0_97_5));
   AOI22_X1 i_0_97_15 (.A1(n_0_97_4), .A2(n_0_97_5), .B1(n_0_127), .B2(n_0_52), 
      .ZN(out[2]));
   XNOR2_X1 i_0_97_16 (.A(n_0_54), .B(n_0_22), .ZN(n_0_97_6));
   XNOR2_X1 i_0_97_17 (.A(n_0_23), .B(n_0_84), .ZN(n_0_97_7));
   AOI22_X1 i_0_97_18 (.A1(n_0_97_6), .A2(n_0_52), .B1(n_0_97_7), .B2(n_0_97_5), 
      .ZN(out[3]));
   OR2_X1 i_0_97_19 (.A1(n_0_34), .A2(n_0_21), .ZN(n_0_97_8));
   AOI22_X1 i_0_97_20 (.A1(n_0_97_8), .A2(in2[13]), .B1(in1[13]), .B2(n_0_32), 
      .ZN(n_0_97_9));
   INV_X1 i_0_97_21 (.A(n_0_97_9), .ZN(out[13]));
   AOI22_X1 i_0_97_22 (.A1(n_0_97_8), .A2(in2[14]), .B1(n_0_32), .B2(in1[14]), 
      .ZN(n_0_97_10));
   INV_X1 i_0_97_23 (.A(n_0_97_10), .ZN(out[14]));
   AOI22_X1 i_0_97_24 (.A1(n_0_97_8), .A2(in2[15]), .B1(n_0_32), .B2(in1[15]), 
      .ZN(n_0_97_11));
   INV_X1 i_0_97_25 (.A(n_0_97_11), .ZN(out[15]));
   INV_X1 i_0_97_26 (.A(n_0_130), .ZN(n_0_75));
   INV_X1 i_0_97_27 (.A(n_0_87), .ZN(n_0_78));
   INV_X1 i_0_6_0 (.A(n_0_92), .ZN(n_0_6_0));
   NAND2_X1 i_0_6_1 (.A1(n_0_6_0), .A2(n_0_13), .ZN(n_0_6_1));
   NAND2_X1 i_0_6_2 (.A1(n_0_92), .A2(n_0_120), .ZN(n_0_6_2));
   NAND2_X1 i_0_6_3 (.A1(n_0_6_1), .A2(n_0_6_2), .ZN(n_0_96));
   INV_X1 i_0_50_0 (.A(n_0_92), .ZN(n_0_50_0));
   NAND2_X1 i_0_50_1 (.A1(n_0_50_0), .A2(n_0_13), .ZN(n_0_50_1));
   NAND2_X1 i_0_50_2 (.A1(n_0_92), .A2(n_0_120), .ZN(n_0_50_2));
   NAND2_X1 i_0_50_3 (.A1(n_0_50_1), .A2(n_0_50_2), .ZN(n_0_50_3));
   INV_X1 i_0_50_4 (.A(n_0_50_3), .ZN(n_0_50_4));
   NAND2_X1 i_0_50_5 (.A1(n_0_116), .A2(n_0_50_4), .ZN(n_0_50_5));
   NAND2_X1 i_0_50_6 (.A1(n_0_106), .A2(n_0_50_3), .ZN(n_0_50_6));
   NAND2_X1 i_0_50_7 (.A1(n_0_50_5), .A2(n_0_50_6), .ZN(n_0_97));
   INV_X1 i_0_84_3 (.A(n_0_93), .ZN(n_0_84_4));
   NAND2_X1 i_0_84_0 (.A1(n_0_84_1), .A2(n_0_84_0), .ZN(n_0_101));
   NAND2_X1 i_0_84_1 (.A1(n_0_84_4), .A2(n_0_98), .ZN(n_0_84_0));
   NAND3_X1 i_0_84_2 (.A1(n_0_84_2), .A2(n_0_93), .A3(n_0_84_6), .ZN(n_0_84_1));
   NAND2_X1 i_0_84_4 (.A1(n_0_84_5), .A2(n_0_84_3), .ZN(n_0_84_2));
   INV_X1 i_0_84_5 (.A(n_0_84_7), .ZN(n_0_84_3));
   INV_X1 i_0_84_6 (.A(n_0_41), .ZN(n_0_84_5));
   NAND2_X1 i_0_84_7 (.A1(n_0_41), .A2(n_0_84_7), .ZN(n_0_84_6));
   XNOR2_X1 i_0_84_8 (.A(n_0_98), .B(n_0_84_8), .ZN(n_0_84_7));
   INV_X1 i_0_84_9 (.A(sub), .ZN(n_0_84_8));
   XNOR2_X1 i_0_101_0 (.A(sub), .B(n_0_41), .ZN(n_0_101_0));
   INV_X1 i_0_101_1 (.A(n_0_93), .ZN(n_0_101_1));
   NOR2_X1 i_0_101_2 (.A1(n_0_101_0), .A2(n_0_101_1), .ZN(n_0_102));
   NAND2_X1 i_0_5_0 (.A1(n_0_5_7), .A2(n_0_5_5), .ZN(n_0_109));
   INV_X1 i_0_5_1 (.A(n_0_30), .ZN(n_0_5_0));
   NAND2_X1 i_0_5_2 (.A1(n_0_5_6), .A2(n_0_30), .ZN(n_0_5_1));
   INV_X1 i_0_5_7 (.A(sub), .ZN(n_0_5_6));
   NAND2_X1 i_0_5_3 (.A1(n_0_5_0), .A2(sub), .ZN(n_0_5_2));
   NAND3_X1 i_0_5_4 (.A1(n_0_5_1), .A2(n_0_5_8), .A3(n_0_53), .ZN(n_0_5_5));
   NAND2_X1 i_0_5_5 (.A1(n_0_5_0), .A2(sub), .ZN(n_0_5_8));
   NAND2_X1 i_0_5_6 (.A1(n_0_5_2), .A2(n_0_5_1), .ZN(n_0_5_3));
   INV_X1 i_0_5_8 (.A(n_0_53), .ZN(n_0_5_4));
   NAND2_X1 i_0_5_9 (.A1(n_0_5_3), .A2(n_0_5_4), .ZN(n_0_5_7));
   INV_X1 i_0_7_0 (.A(n_0_4), .ZN(n_0_7_0));
   INV_X1 i_0_7_1 (.A(n_0_20), .ZN(n_0_7_6));
   BUF_X1 rt_shieldBuf__1__1__1 (.A(n_0_5), .Z(n_0_7_13));
   NAND2_X1 i_0_7_6 (.A1(n_0_7_2), .A2(n_0_7_1), .ZN(out[12]));
   NAND2_X1 i_0_7_7 (.A1(n_0_7_117), .A2(n_0_7_13), .ZN(n_0_7_1));
   NAND2_X1 i_0_7_8 (.A1(n_0_7_90), .A2(n_0_7_3), .ZN(n_0_7_2));
   INV_X1 i_0_7_9 (.A(n_0_7_13), .ZN(n_0_7_3));
   OAI21_X1 i_0_7_2 (.A(n_0_7_5), .B1(n_0_7_9), .B2(n_0_20), .ZN(n_0_7_4));
   NAND2_X1 i_0_7_3 (.A1(n_0_7_11), .A2(n_0_20), .ZN(n_0_7_5));
   OAI21_X1 i_0_7_4 (.A(n_0_7_8), .B1(n_0_7_48), .B2(n_0_7_11), .ZN(n_0_7_7));
   NAND2_X1 i_0_7_5 (.A1(n_0_7_9), .A2(n_0_7_48), .ZN(n_0_7_8));
   INV_X1 i_0_7_10 (.A(n_0_7_10), .ZN(n_0_7_9));
   OAI21_X1 i_0_7_16 (.A(n_0_7_25), .B1(n_0_81), .B2(n_0_113), .ZN(n_0_7_10));
   OAI21_X1 i_0_7_11 (.A(n_0_7_12), .B1(n_0_10), .B2(n_0_113), .ZN(n_0_7_11));
   NAND2_X1 i_0_7_19 (.A1(n_0_10), .A2(n_0_7_89), .ZN(n_0_7_12));
   XNOR2_X1 i_0_7_12 (.A(n_0_7_14), .B(n_0_69), .ZN(n_0_7_19));
   OAI21_X1 i_0_7_21 (.A(n_0_7_15), .B1(n_0_7_17), .B2(n_0_8), .ZN(n_0_7_14));
   OAI211_X1 i_0_7_22 (.A(n_0_7_16), .B(n_0_8), .C1(n_0_113), .C2(n_0_100), 
      .ZN(n_0_7_15));
   NAND2_X1 i_0_7_23 (.A1(n_0_113), .A2(n_0_7_87), .ZN(n_0_7_16));
   OAI21_X1 i_0_7_24 (.A(n_0_7_18), .B1(n_0_113), .B2(n_0_7_82), .ZN(n_0_7_17));
   NAND2_X1 i_0_7_25 (.A1(n_0_113), .A2(n_0_100), .ZN(n_0_7_18));
   OAI21_X1 i_0_7_13 (.A(n_0_7_20), .B1(n_0_7_24), .B2(n_0_7_28), .ZN(n_0_7_34));
   NAND4_X1 i_0_7_27 (.A1(n_0_7_23), .A2(n_0_7_22), .A3(n_0_7_65), .A4(n_0_7_21), 
      .ZN(n_0_7_20));
   NAND2_X1 i_0_7_28 (.A1(n_0_81), .A2(n_0_7_27), .ZN(n_0_7_21));
   NAND3_X1 i_0_7_29 (.A1(n_0_7_67), .A2(n_0_7_75), .A3(n_0_7_26), .ZN(n_0_7_22));
   NAND3_X1 i_0_7_30 (.A1(n_0_7_67), .A2(n_0_113), .A3(n_0_7_30), .ZN(n_0_7_23));
   OAI22_X1 i_0_7_31 (.A1(n_0_7_25), .A2(n_0_7_26), .B1(n_0_81), .B2(n_0_7_27), 
      .ZN(n_0_7_24));
   NAND2_X1 i_0_7_32 (.A1(n_0_81), .A2(n_0_7_89), .ZN(n_0_7_25));
   XNOR2_X1 i_0_7_33 (.A(n_0_101), .B(n_0_100), .ZN(n_0_7_26));
   XNOR2_X1 i_0_7_34 (.A(n_0_103), .B(n_0_100), .ZN(n_0_7_27));
   OAI21_X1 i_0_7_35 (.A(n_0_10), .B1(n_0_7_29), .B2(n_0_7_30), .ZN(n_0_7_28));
   NAND2_X1 i_0_7_36 (.A1(n_0_81), .A2(n_0_8), .ZN(n_0_7_29));
   XNOR2_X1 i_0_7_37 (.A(n_0_99), .B(n_0_100), .ZN(n_0_7_30));
   OAI21_X1 i_0_7_38 (.A(n_0_7_32), .B1(n_0_7_48), .B2(n_0_7_33), .ZN(n_0_7_31));
   NAND2_X1 i_0_7_39 (.A1(n_0_7_33), .A2(n_0_20), .ZN(n_0_7_32));
   XNOR2_X1 i_0_7_40 (.A(n_0_5), .B(n_0_103), .ZN(n_0_7_33));
   OAI211_X1 i_0_7_14 (.A(n_0_7_36), .B(n_0_7_35), .C1(n_0_7_67), .C2(n_0_7_37), 
      .ZN(n_0_7_38));
   NOR2_X1 i_0_7_42 (.A1(n_0_11), .A2(n_0_20), .ZN(n_0_7_35));
   NAND2_X1 i_0_7_43 (.A1(n_0_7_40), .A2(n_0_7_67), .ZN(n_0_7_36));
   NAND2_X1 i_0_7_44 (.A1(n_0_7_43), .A2(n_0_7_44), .ZN(n_0_7_37));
   AOI21_X1 i_0_7_15 (.A(n_0_7_6), .B1(n_0_7_40), .B2(n_0_7_65), .ZN(n_0_7_39));
   OAI21_X1 i_0_7_47 (.A(n_0_7_41), .B1(n_0_7_45), .B2(n_0_7_75), .ZN(n_0_7_40));
   NAND2_X1 i_0_7_48 (.A1(n_0_7_171), .A2(n_0_7_75), .ZN(n_0_7_41));
   NAND2_X1 i_0_7_51 (.A1(n_0_7_45), .A2(n_0_8), .ZN(n_0_7_43));
   XNOR2_X1 i_0_7_50 (.A(n_0_99), .B(n_0_103), .ZN(n_0_7_45));
   NAND2_X1 i_0_7_53 (.A1(n_0_7_42), .A2(n_0_7_89), .ZN(n_0_7_44));
   INV_X1 i_0_7_18 (.A(n_0_11), .ZN(n_0_7_48));
   NAND2_X1 i_0_7_20 (.A1(n_0_7_73), .A2(n_0_7_74), .ZN(n_0_7_49));
   NAND3_X1 i_0_7_26 (.A1(n_0_7_51), .A2(n_0_11), .A3(n_0_7_56), .ZN(n_0_7_50));
   XNOR2_X1 i_0_7_41 (.A(n_0_7), .B(n_0_5), .ZN(n_0_7_51));
   OAI211_X1 i_0_7_17 (.A(n_0_7_55), .B(n_0_7_160), .C1(n_0_7_112), .C2(n_0_81), 
      .ZN(n_0_7_52));
   NAND2_X1 i_0_7_46 (.A1(n_0_7_58), .A2(n_0_81), .ZN(n_0_7_55));
   OAI211_X1 i_0_7_45 (.A(n_0_7_57), .B(n_0_20), .C1(n_0_7_112), .C2(n_0_10), 
      .ZN(n_0_7_53));
   NAND2_X1 i_0_7_49 (.A1(n_0_7_58), .A2(n_0_10), .ZN(n_0_7_57));
   OAI21_X1 i_0_7_70 (.A(n_0_7_59), .B1(n_0_7_108), .B2(n_0_7_89), .ZN(n_0_7_58));
   NAND2_X1 i_0_7_71 (.A1(n_0_7_60), .A2(n_0_7_89), .ZN(n_0_7_59));
   XNOR2_X1 i_0_7_72 (.A(n_0_101), .B(n_0_7_61), .ZN(n_0_7_60));
   INV_X1 i_0_7_73 (.A(in1[12]), .ZN(n_0_7_61));
   XNOR2_X1 i_0_7_74 (.A(n_0_67), .B(in1[12]), .ZN(n_0_7_54));
   NAND2_X1 i_0_7_55 (.A1(n_0_7_62), .A2(n_0_7_65), .ZN(n_0_7_64));
   INV_X1 i_0_7_52 (.A(n_0_10), .ZN(n_0_7_65));
   XNOR2_X1 i_0_7_54 (.A(n_0_90), .B(n_0_5), .ZN(n_0_7_56));
   NAND2_X1 i_0_7_75 (.A1(n_0_7_69), .A2(n_0_10), .ZN(n_0_7_70));
   NAND3_X1 i_0_7_76 (.A1(n_0_7_76), .A2(n_0_7_74), .A3(n_0_7_73), .ZN(n_0_7_62));
   NAND2_X1 i_0_7_56 (.A1(n_0_7_84), .A2(n_0_113), .ZN(n_0_7_73));
   NAND3_X1 i_0_7_57 (.A1(n_0_7_83), .A2(n_0_7_75), .A3(n_0_7_81), .ZN(n_0_7_74));
   INV_X1 i_0_7_58 (.A(n_0_113), .ZN(n_0_7_75));
   INV_X1 i_0_7_60 (.A(n_0_7_77), .ZN(n_0_7_76));
   XNOR2_X1 i_0_7_61 (.A(n_0_14), .B(n_0_5), .ZN(n_0_7_77));
   XNOR2_X1 i_0_7_59 (.A(n_0_12), .B(n_0_5), .ZN(n_0_7_63));
   NAND2_X1 i_0_7_102 (.A1(n_0_7_83), .A2(n_0_7_81), .ZN(n_0_7_80));
   NAND2_X1 i_0_7_62 (.A1(n_0_5), .A2(n_0_7_82), .ZN(n_0_7_81));
   INV_X1 i_0_7_104 (.A(n_0_101), .ZN(n_0_7_82));
   NAND2_X1 i_0_7_63 (.A1(n_0_7_88), .A2(n_0_101), .ZN(n_0_7_83));
   NAND2_X1 i_0_7_64 (.A1(n_0_7_86), .A2(n_0_7_85), .ZN(n_0_7_84));
   NAND2_X1 i_0_7_107 (.A1(n_0_99), .A2(n_0_5), .ZN(n_0_7_85));
   NAND2_X1 i_0_7_108 (.A1(n_0_7_87), .A2(n_0_7_88), .ZN(n_0_7_86));
   INV_X1 i_0_7_109 (.A(n_0_99), .ZN(n_0_7_87));
   INV_X1 i_0_7_110 (.A(n_0_5), .ZN(n_0_7_88));
   INV_X1 i_0_7_90 (.A(n_0_8), .ZN(n_0_7_89));
   INV_X1 i_0_7_65 (.A(n_0_7_117), .ZN(n_0_7_90));
   NAND3_X1 i_0_7_66 (.A1(n_0_7_63), .A2(n_0_7_48), .A3(n_0_7_51), .ZN(n_0_7_92));
   INV_X1 i_0_7_117 (.A(n_0_7_89), .ZN(n_0_7_93));
   INV_X1 i_0_7_118 (.A(n_0_7_84), .ZN(n_0_7_94));
   OAI211_X1 i_0_7_67 (.A(n_0_7_57), .B(n_0_11), .C1(n_0_7_112), .C2(n_0_10), 
      .ZN(n_0_7_95));
   OAI211_X1 i_0_7_68 (.A(n_0_7_55), .B(n_0_7_48), .C1(n_0_7_112), .C2(n_0_81), 
      .ZN(n_0_7_96));
   XNOR2_X1 i_0_7_124 (.A(n_0_123), .B(n_0_5), .ZN(n_0_7_97));
   NAND2_X1 i_0_7_125 (.A1(n_0_7_80), .A2(n_0_7_89), .ZN(n_0_7_98));
   NAND2_X1 i_0_7_126 (.A1(n_0_7_89), .A2(n_0_7_80), .ZN(n_0_7_99));
   XNOR2_X1 i_0_7_127 (.A(n_0_123), .B(n_0_5), .ZN(n_0_7_100));
   NAND2_X1 i_0_7_128 (.A1(n_0_7_99), .A2(n_0_7_100), .ZN(n_0_7_101));
   INV_X1 i_0_7_69 (.A(n_0_7_101), .ZN(n_0_7_102));
   NAND2_X1 i_0_7_77 (.A1(n_0_7_94), .A2(n_0_7_93), .ZN(n_0_7_103));
   NAND3_X1 i_0_7_78 (.A1(n_0_7_96), .A2(n_0_7_95), .A3(n_0_7_54), .ZN(n_0_7_104));
   NOR2_X1 i_0_7_79 (.A1(n_0_7_153), .A2(n_0_7_50), .ZN(n_0_7_105));
   INV_X1 i_0_7_80 (.A(n_0_7_31), .ZN(n_0_7_66));
   XNOR2_X1 i_0_7_140 (.A(n_0_99), .B(in1[12]), .ZN(n_0_7_108));
   INV_X1 i_0_7_141 (.A(n_0_7_75), .ZN(n_0_7_109));
   INV_X1 i_0_7_142 (.A(in1[12]), .ZN(n_0_7_110));
   XNOR2_X1 i_0_7_143 (.A(n_0_99), .B(n_0_7_110), .ZN(n_0_7_111));
   OAI22_X1 i_0_7_81 (.A1(n_0_7_109), .A2(n_0_7_60), .B1(n_0_7_75), .B2(
      n_0_7_111), .ZN(n_0_7_112));
   NAND2_X1 i_0_7_82 (.A1(n_0_7_105), .A2(n_0_7_104), .ZN(n_0_7_113));
   INV_X1 i_0_7_151 (.A(n_0_116), .ZN(n_0_7_114));
   INV_X1 i_0_7_152 (.A(n_0_13), .ZN(n_0_7_115));
   INV_X1 i_0_7_153 (.A(n_0_106), .ZN(n_0_7_116));
   NAND2_X1 i_0_7_83 (.A1(n_0_7_128), .A2(n_0_7_126), .ZN(n_0_7_117));
   INV_X1 i_0_7_155 (.A(n_0_92), .ZN(n_0_7_118));
   INV_X1 i_0_7_156 (.A(n_0_7_115), .ZN(n_0_7_119));
   NAND2_X1 i_0_7_157 (.A1(n_0_92), .A2(n_0_120), .ZN(n_0_7_120));
   NAND2_X1 i_0_7_158 (.A1(n_0_43), .A2(n_0_7_114), .ZN(n_0_7_121));
   NAND2_X1 i_0_7_159 (.A1(n_0_116), .A2(n_0_126), .ZN(n_0_7_122));
   NAND2_X1 i_0_7_84 (.A1(n_0_7_121), .A2(n_0_7_122), .ZN(n_0_7_123));
   NAND2_X1 i_0_7_85 (.A1(n_0_7_118), .A2(n_0_7_119), .ZN(n_0_7_124));
   NAND2_X1 i_0_7_86 (.A1(n_0_92), .A2(n_0_120), .ZN(n_0_7_125));
   NAND3_X1 i_0_7_87 (.A1(n_0_7_123), .A2(n_0_7_124), .A3(n_0_7_125), .ZN(
      n_0_7_126));
   OAI21_X1 i_0_7_88 (.A(n_0_7_120), .B1(n_0_92), .B2(n_0_7_115), .ZN(n_0_7_127));
   NAND2_X1 i_0_7_89 (.A1(n_0_7_127), .A2(n_0_7_131), .ZN(n_0_7_128));
   NAND2_X1 i_0_7_166 (.A1(n_0_7_116), .A2(n_0_43), .ZN(n_0_7_129));
   NAND2_X1 i_0_7_167 (.A1(n_0_106), .A2(n_0_126), .ZN(n_0_7_130));
   NAND2_X1 i_0_7_91 (.A1(n_0_7_129), .A2(n_0_7_130), .ZN(n_0_7_131));
   OAI21_X1 i_0_7_92 (.A(n_0_7_144), .B1(n_0_7_117), .B2(n_0_7_4), .ZN(n_0_7_133));
   INV_X1 i_0_7_93 (.A(n_0_7_117), .ZN(n_0_7_134));
   INV_X1 i_0_7_94 (.A(n_0_7_4), .ZN(n_0_7_135));
   NAND2_X1 i_0_7_97 (.A1(n_0_7_49), .A2(n_0_7_77), .ZN(n_0_7_136));
   INV_X1 i_0_7_100 (.A(n_0_81), .ZN(n_0_7_67));
   NAND2_X1 i_0_7_99 (.A1(n_0_7_102), .A2(n_0_7_103), .ZN(n_0_7_138));
   INV_X1 i_0_7_133 (.A(n_0_81), .ZN(n_0_7_139));
   NAND3_X1 i_0_7_101 (.A1(n_0_7_77), .A2(n_0_7_49), .A3(n_0_7_139), .ZN(
      n_0_7_140));
   NAND2_X1 i_0_7_165 (.A1(n_0_7_103), .A2(n_0_81), .ZN(n_0_7_141));
   INV_X1 i_0_7_135 (.A(n_0_7_141), .ZN(n_0_7_142));
   NAND2_X1 i_0_7_103 (.A1(n_0_7_142), .A2(n_0_7_102), .ZN(n_0_7_143));
   NAND2_X1 i_0_7_105 (.A1(n_0_7_117), .A2(n_0_7_7), .ZN(n_0_7_144));
   NAND2_X1 i_0_7_106 (.A1(n_0_7_135), .A2(n_0_7_134), .ZN(n_0_7_145));
   INV_X1 i_0_7_95 (.A(n_0_73), .ZN(n_0_7_146));
   AOI21_X1 i_0_7_111 (.A(n_0_7_146), .B1(n_0_7_117), .B2(n_0_7_7), .ZN(
      n_0_7_147));
   NAND3_X1 i_0_7_96 (.A1(n_0_7_168), .A2(n_0_7_64), .A3(n_0_7_70), .ZN(n_0_7_68));
   NAND2_X1 i_0_7_115 (.A1(n_0_7_136), .A2(n_0_7_65), .ZN(n_0_7_151));
   NAND2_X1 i_0_7_116 (.A1(n_0_7_138), .A2(n_0_10), .ZN(n_0_7_152));
   NAND2_X1 i_0_7_119 (.A1(n_0_7_151), .A2(n_0_7_152), .ZN(n_0_7_153));
   NAND2_X1 i_0_7_120 (.A1(n_0_7_133), .A2(n_0_72), .ZN(n_0_7_154));
   NAND2_X1 i_0_7_122 (.A1(n_0_7_145), .A2(n_0_7_147), .ZN(n_0_7_155));
   NAND2_X1 i_0_7_123 (.A1(n_0_7_154), .A2(n_0_7_155), .ZN(cout));
   NAND3_X1 i_0_7_129 (.A1(n_0_7_96), .A2(n_0_7_95), .A3(n_0_7_54), .ZN(
      n_0_7_156));
   INV_X1 i_0_7_130 (.A(n_0_7_92), .ZN(n_0_7_157));
   NAND2_X1 i_0_7_131 (.A1(n_0_7_143), .A2(n_0_7_140), .ZN(n_0_7_158));
   NAND3_X1 i_0_7_134 (.A1(n_0_7_156), .A2(n_0_7_157), .A3(n_0_7_158), .ZN(
      n_0_7_159));
   INV_X1 i_0_7_112 (.A(n_0_20), .ZN(n_0_7_160));
   INV_X1 i_0_7_121 (.A(n_0_7_97), .ZN(n_0_7_162));
   OAI21_X1 i_0_7_132 (.A(n_0_7_98), .B1(n_0_7_84), .B2(n_0_7_89), .ZN(n_0_7_163));
   NAND2_X1 i_0_7_138 (.A1(n_0_7_162), .A2(n_0_7_163), .ZN(n_0_7_69));
   NAND3_X1 i_0_7_136 (.A1(n_0_7_159), .A2(n_0_7_113), .A3(n_0_7_117), .ZN(
      n_0_7_165));
   NAND2_X1 i_0_7_137 (.A1(n_0_7_106), .A2(n_0_7_90), .ZN(n_0_7_166));
   NAND3_X1 i_0_7_139 (.A1(n_0_7_165), .A2(n_0_7_166), .A3(n_0_7_148), .ZN(
      invalid));
   NAND2_X1 i_0_7_144 (.A1(n_0_7_68), .A2(n_0_7_164), .ZN(n_0_7_78));
   NAND3_X1 i_0_7_145 (.A1(n_0_7_52), .A2(n_0_7_53), .A3(n_0_7_54), .ZN(n_0_7_79));
   XNOR2_X1 i_0_7_147 (.A(n_0_7_13), .B(n_0_7_0), .ZN(n_0_7_91));
   NAND3_X1 i_0_7_148 (.A1(n_0_7_78), .A2(n_0_7_79), .A3(n_0_7_91), .ZN(
      n_0_7_106));
   NAND2_X1 i_0_7_149 (.A1(n_0_7_19), .A2(n_0_7_34), .ZN(n_0_7_107));
   NAND2_X1 i_0_7_150 (.A1(n_0_7_38), .A2(n_0_7_66), .ZN(n_0_7_132));
   NAND2_X1 i_0_7_160 (.A1(n_0_7_170), .A2(n_0_7_39), .ZN(n_0_7_137));
   AOI21_X1 i_0_7_161 (.A(n_0_7_107), .B1(n_0_7_132), .B2(n_0_7_137), .ZN(
      n_0_7_148));
   NAND2_X1 i_0_7_168 (.A1(n_0_7_62), .A2(n_0_7_67), .ZN(n_0_7_149));
   NAND2_X1 i_0_7_169 (.A1(n_0_7_69), .A2(n_0_81), .ZN(n_0_7_150));
   NOR2_X1 i_0_7_170 (.A1(n_0_20), .A2(n_0_7_63), .ZN(n_0_7_161));
   NAND3_X1 i_0_7_171 (.A1(n_0_7_149), .A2(n_0_7_150), .A3(n_0_7_161), .ZN(
      n_0_7_164));
   INV_X1 i_0_7_98 (.A(n_0_20), .ZN(n_0_7_167));
   NOR2_X1 i_0_7_114 (.A1(n_0_7_56), .A2(n_0_7_167), .ZN(n_0_7_168));
   INV_X1 i_0_7_113 (.A(n_0_7_44), .ZN(n_0_7_46));
   NAND2_X1 i_0_7_146 (.A1(n_0_7_46), .A2(n_0_11), .ZN(n_0_7_71));
   NAND2_X1 i_0_7_154 (.A1(n_0_7_43), .A2(n_0_10), .ZN(n_0_7_72));
   NAND2_X1 i_0_7_164 (.A1(n_0_7_72), .A2(n_0_11), .ZN(n_0_7_169));
   NAND2_X1 i_0_7_162 (.A1(n_0_7_71), .A2(n_0_7_169), .ZN(n_0_7_170));
   XNOR2_X1 i_0_7_163 (.A(n_0_101), .B(n_0_103), .ZN(n_0_7_42));
   INV_X1 i_0_7_172 (.A(n_0_101), .ZN(n_0_7_47));
   XNOR2_X1 i_0_7_173 (.A(n_0_103), .B(n_0_7_47), .ZN(n_0_7_171));
   NAND3_X1 i_0_3_0 (.A1(n_0_3_1), .A2(n_0_3_3), .A3(n_0_3_0), .ZN(n_0_18));
   NAND2_X1 i_0_3_1 (.A1(n_0_63), .A2(n_0_40), .ZN(n_0_3_0));
   NAND3_X1 i_0_3_2 (.A1(n_0_3_2), .A2(n_0_84), .A3(n_0_23), .ZN(n_0_3_1));
   INV_X1 i_0_3_3 (.A(n_0_52), .ZN(n_0_3_2));
   NAND3_X1 i_0_3_4 (.A1(n_0_52), .A2(n_0_22), .A3(n_0_54), .ZN(n_0_3_3));
   INV_X1 i_0_20_0 (.A(n_0_20_1), .ZN(n_0_65));
   INV_X1 i_0_20_1 (.A(n_0_20_0), .ZN(n_0_67));
   XNOR2_X1 i_0_20_2 (.A(in2[12]), .B(sub), .ZN(n_0_20_0));
   NAND2_X1 i_0_20_3 (.A1(n_0_20_1), .A2(n_0_20_12), .ZN(n_0_95));
   XNOR2_X1 i_0_20_4 (.A(n_0_41), .B(sub), .ZN(n_0_20_1));
   INV_X1 i_0_20_5 (.A(n_0_20_2), .ZN(n_0_99));
   NAND2_X1 i_0_20_6 (.A1(n_0_20_4), .A2(n_0_20_3), .ZN(n_0_20_2));
   NAND2_X1 i_0_20_7 (.A1(n_0_93), .A2(n_0_98), .ZN(n_0_20_3));
   XNOR2_X1 i_0_20_8 (.A(n_0_20_7), .B(sub), .ZN(n_0_98));
   NAND2_X1 i_0_20_9 (.A1(n_0_20_5), .A2(n_0_20_12), .ZN(n_0_20_4));
   NAND2_X1 i_0_20_10 (.A1(n_0_20_6), .A2(n_0_20_9), .ZN(n_0_20_5));
   NAND2_X1 i_0_20_11 (.A1(n_0_20_8), .A2(n_0_20_7), .ZN(n_0_20_6));
   INV_X1 i_0_20_12 (.A(n_0_20_10), .ZN(n_0_20_7));
   INV_X1 i_0_20_13 (.A(n_0_41), .ZN(n_0_20_8));
   NAND2_X1 i_0_20_14 (.A1(n_0_41), .A2(n_0_20_10), .ZN(n_0_20_9));
   XNOR2_X1 i_0_20_15 (.A(n_0_20_11), .B(in2[12]), .ZN(n_0_20_10));
   INV_X1 i_0_20_16 (.A(in1[12]), .ZN(n_0_20_11));
   INV_X1 i_0_20_17 (.A(n_0_93), .ZN(n_0_20_12));
   XNOR2_X1 i_0_42_0 (.A(n_0_59), .B(n_0_94), .ZN(n_0_100));
   INV_X1 i_0_18_3 (.A(sub), .ZN(n_0_18_0));
   INV_X1 i_0_18_2 (.A(sub), .ZN(n_0_18_1));
   INV_X1 i_0_18_0 (.A(n_0_18_0), .ZN(n_0_18_2));
   XNOR2_X1 i_0_18_1 (.A(n_0_33), .B(n_0_18_2), .ZN(n_0_18_3));
   INV_X1 i_0_18_4 (.A(n_0_45), .ZN(n_0_18_4));
   NAND2_X1 i_0_18_5 (.A1(n_0_18_3), .A2(n_0_18_4), .ZN(n_0_18_5));
   XNOR2_X1 i_0_18_6 (.A(n_0_33), .B(n_0_18_1), .ZN(n_0_18_6));
   NAND2_X1 i_0_18_7 (.A1(n_0_18_6), .A2(n_0_45), .ZN(n_0_18_7));
   NAND2_X1 i_0_18_8 (.A1(n_0_18_5), .A2(n_0_18_7), .ZN(n_0_103));
   INV_X1 i_0_25_0 (.A(sub), .ZN(n_0_25_0));
   XNOR2_X1 i_0_25_1 (.A(n_0_29), .B(n_0_25_0), .ZN(n_0_25_1));
   NAND2_X1 i_0_25_2 (.A1(n_0_25_1), .A2(n_0_50), .ZN(n_0_25_2));
   NOR2_X1 i_0_25_3 (.A1(n_0_25_1), .A2(n_0_50), .ZN(n_0_25_3));
   XNOR2_X1 i_0_25_4 (.A(n_0_28), .B(n_0_25_0), .ZN(n_0_111));
   NAND2_X1 i_0_25_5 (.A1(n_0_111), .A2(n_0_48), .ZN(n_0_25_4));
   OAI21_X1 i_0_25_6 (.A(n_0_25_2), .B1(n_0_25_3), .B2(n_0_25_4), .ZN(n_0_116));
   XNOR2_X1 i_0_25_7 (.A(n_0_28), .B(sub), .ZN(n_0_25_5));
   INV_X1 i_0_25_8 (.A(n_0_48), .ZN(n_0_25_6));
   NOR2_X1 i_0_25_9 (.A1(n_0_25_5), .A2(n_0_25_6), .ZN(n_0_112));
   XNOR2_X1 i_0_25_10 (.A(n_0_25_5), .B(n_0_48), .ZN(n_0_110));
   NAND2_X1 i_0_25_11 (.A1(n_0_25_5), .A2(n_0_25_6), .ZN(n_0_108));
   XNOR2_X1 i_0_25_12 (.A(n_0_29), .B(sub), .ZN(n_0_25_7));
   XNOR2_X1 i_0_25_13 (.A(n_0_25_7), .B(n_0_50), .ZN(n_0_107));
   INV_X1 i_0_25_14 (.A(n_0_29), .ZN(n_0_25_8));
   NOR2_X1 i_0_25_15 (.A1(n_0_28), .A2(n_0_25_0), .ZN(n_0_25_9));
   AOI21_X1 i_0_25_16 (.A(n_0_25_9), .B1(n_0_48), .B2(sub), .ZN(n_0_25_10));
   OAI22_X1 i_0_25_17 (.A1(n_0_25_15), .A2(n_0_25_8), .B1(n_0_25_10), .B2(n_0_29), 
      .ZN(n_0_25_11));
   INV_X1 i_0_25_18 (.A(n_0_25_11), .ZN(n_0_25_12));
   NAND3_X1 i_0_25_19 (.A1(n_0_25_7), .A2(n_0_25_5), .A3(n_0_25_6), .ZN(
      n_0_25_13));
   NAND2_X1 i_0_25_20 (.A1(n_0_25_13), .A2(n_0_50), .ZN(n_0_25_14));
   NAND2_X1 i_0_25_21 (.A1(n_0_25_12), .A2(n_0_25_14), .ZN(n_0_106));
   OAI21_X1 i_0_25_22 (.A(n_0_25_0), .B1(n_0_48), .B2(n_0_28), .ZN(n_0_25_15));
   INV_X1 i_0_23_0 (.A(sub), .ZN(n_0_23_0));
   NAND2_X1 i_0_23_1 (.A1(n_0_23_13), .A2(n_0_47), .ZN(n_0_23_1));
   OAI21_X1 i_0_23_2 (.A(n_0_23_1), .B1(n_0_23_14), .B2(n_0_23_15), .ZN(n_0_13));
   XNOR2_X1 i_0_23_7 (.A(n_0_26), .B(sub), .ZN(n_0_23_2));
   INV_X1 i_0_23_8 (.A(n_0_46), .ZN(n_0_23_3));
   NOR2_X1 i_0_23_9 (.A1(n_0_23_2), .A2(n_0_23_3), .ZN(n_0_9));
   XNOR2_X1 i_0_23_10 (.A(n_0_23_2), .B(n_0_46), .ZN(n_0_130));
   NAND2_X1 i_0_23_11 (.A1(n_0_23_2), .A2(n_0_23_3), .ZN(n_0_128));
   XNOR2_X1 i_0_23_12 (.A(n_0_27), .B(sub), .ZN(n_0_23_4));
   XNOR2_X1 i_0_23_13 (.A(n_0_23_4), .B(n_0_47), .ZN(n_0_125));
   OAI21_X1 i_0_23_14 (.A(n_0_47), .B1(n_0_23_13), .B2(n_0_1), .ZN(n_0_23_5));
   OAI21_X1 i_0_23_15 (.A(n_0_46), .B1(n_0_23_13), .B2(n_0_47), .ZN(n_0_23_6));
   INV_X1 i_0_23_16 (.A(n_0_27), .ZN(n_0_23_7));
   INV_X1 i_0_23_17 (.A(n_0_26), .ZN(n_0_23_8));
   NAND3_X1 i_0_23_18 (.A1(n_0_23_7), .A2(n_0_23_8), .A3(sub), .ZN(n_0_23_9));
   NAND3_X1 i_0_23_19 (.A1(n_0_27), .A2(n_0_26), .A3(n_0_23_0), .ZN(n_0_23_10));
   NAND2_X1 i_0_23_20 (.A1(n_0_23_9), .A2(n_0_23_10), .ZN(n_0_23_11));
   INV_X1 i_0_23_21 (.A(n_0_23_11), .ZN(n_0_23_12));
   NAND3_X1 i_0_23_22 (.A1(n_0_23_5), .A2(n_0_23_6), .A3(n_0_23_12), .ZN(n_0_120));
   XNOR2_X1 i_0_23_3 (.A(n_0_27), .B(n_0_23_0), .ZN(n_0_23_13));
   NOR2_X1 i_0_23_4 (.A1(n_0_23_13), .A2(n_0_47), .ZN(n_0_23_14));
   XNOR2_X1 i_0_23_5 (.A(n_0_26), .B(n_0_23_0), .ZN(n_0_1));
   NAND2_X1 i_0_23_6 (.A1(n_0_1), .A2(n_0_46), .ZN(n_0_23_15));
   NAND2_X1 i_0_2_1 (.A1(n_0_2_14), .A2(n_0_58), .ZN(n_0_2_0));
   INV_X1 i_0_2_2 (.A(n_0_30), .ZN(n_0_2_1));
   NAND2_X1 i_0_2_3 (.A1(n_0_2_1), .A2(n_0_53), .ZN(n_0_2_2));
   NOR2_X1 i_0_2_4 (.A1(n_0_2_14), .A2(n_0_58), .ZN(n_0_2_3));
   OAI21_X1 i_0_2_5 (.A(n_0_2_0), .B1(n_0_2_2), .B2(n_0_2_3), .ZN(n_0_2_4));
   NAND2_X1 i_0_2_6 (.A1(n_0_2_4), .A2(sub), .ZN(n_0_2_5));
   NAND2_X1 i_0_2_7 (.A1(n_0_58), .A2(n_0_31), .ZN(n_0_2_6));
   NOR2_X1 i_0_2_8 (.A1(n_0_58), .A2(n_0_31), .ZN(n_0_2_7));
   NAND2_X1 i_0_2_9 (.A1(n_0_53), .A2(n_0_30), .ZN(n_0_2_8));
   OAI21_X1 i_0_2_10 (.A(n_0_2_6), .B1(n_0_2_7), .B2(n_0_2_8), .ZN(n_0_2_9));
   NAND2_X1 i_0_2_11 (.A1(n_0_2_9), .A2(n_0_2_16), .ZN(n_0_2_10));
   NAND2_X1 i_0_2_12 (.A1(n_0_2_5), .A2(n_0_2_10), .ZN(n_0_20));
   XNOR2_X1 i_0_2_13 (.A(sub), .B(n_0_30), .ZN(n_0_2_11));
   INV_X1 i_0_2_14 (.A(n_0_53), .ZN(n_0_2_12));
   NOR2_X1 i_0_2_15 (.A1(n_0_2_11), .A2(n_0_2_12), .ZN(n_0_19));
   XNOR2_X1 i_0_2_18 (.A(n_0_2_16), .B(n_0_30), .ZN(n_0_15));
   NAND2_X1 i_0_2_0 (.A1(n_0_2_13), .A2(n_0_2_15), .ZN(n_0_16));
   NAND2_X1 i_0_2_16 (.A1(n_0_2_14), .A2(sub), .ZN(n_0_2_13));
   INV_X1 i_0_2_17 (.A(n_0_31), .ZN(n_0_2_14));
   NAND2_X1 i_0_2_19 (.A1(n_0_31), .A2(n_0_2_16), .ZN(n_0_2_15));
   INV_X1 i_0_2_23 (.A(sub), .ZN(n_0_2_16));
   XNOR2_X1 i_0_2_20 (.A(n_0_31), .B(sub), .ZN(n_0_2_17));
   XNOR2_X1 i_0_2_21 (.A(n_0_2_17), .B(n_0_58), .ZN(n_0_17));
   NAND2_X1 i_0_8_1 (.A1(n_0_8_803), .A2(n_0_40), .ZN(n_0_8_49));
   INV_X1 i_0_8_4 (.A(n_0_40), .ZN(n_0_8_50));
   INV_X1 i_0_8_6 (.A(n_0_8_812), .ZN(n_0_8_0));
   NAND2_X1 i_0_8_7 (.A1(n_0_8_0), .A2(n_0_8_788), .ZN(n_0_8_51));
   INV_X1 i_0_8_8 (.A(n_0_8_268), .ZN(n_0_8_2));
   NAND2_X1 i_0_8_9 (.A1(n_0_8_2), .A2(n_0_8_232), .ZN(n_0_8_57));
   NOR2_X1 i_0_8_10 (.A1(n_0_8_0), .A2(n_0_8_788), .ZN(n_0_8_61));
   NAND2_X1 i_0_8_11 (.A1(n_0_8_788), .A2(n_0_8_812), .ZN(n_0_8_6));
   NOR2_X1 i_0_8_12 (.A1(n_0_8_788), .A2(n_0_8_812), .ZN(n_0_8_7));
   NAND2_X1 i_0_8_13 (.A1(n_0_8_268), .A2(n_0_8_232), .ZN(n_0_8_8));
   OAI21_X1 i_0_8_14 (.A(n_0_8_6), .B1(n_0_8_7), .B2(n_0_8_8), .ZN(n_0_8_9));
   NAND2_X1 i_0_8_16 (.A1(n_0_8_2), .A2(n_0_8_21), .ZN(n_0_8_12));
   NAND2_X1 i_0_8_2 (.A1(n_0_8_12), .A2(n_0_8_18), .ZN(n_0_8_62));
   NAND2_X1 i_0_8_18 (.A1(n_0_8_21), .A2(n_0_8_268), .ZN(n_0_8_14));
   NAND2_X1 i_0_8_15 (.A1(n_0_8_14), .A2(sub), .ZN(n_0_8_77));
   NAND2_X1 i_0_8_17 (.A1(n_0_63), .A2(n_0_40), .ZN(n_0_8_78));
   NOR2_X1 i_0_8_22 (.A1(n_0_8_20), .A2(n_0_8_810), .ZN(n_0_91));
   INV_X1 i_0_8_23 (.A(sub), .ZN(n_0_8_18));
   XNOR2_X1 i_0_8_24 (.A(n_0_8_18), .B(n_0_8_268), .ZN(n_0_88));
   XNOR2_X1 i_0_8_25 (.A(n_0_8_268), .B(n_0_42), .ZN(n_0_8_19));
   XNOR2_X1 i_0_8_26 (.A(n_0_8_19), .B(sub), .ZN(n_0_87));
   XNOR2_X1 i_0_8_27 (.A(sub), .B(n_0_8_268), .ZN(n_0_8_20));
   INV_X1 i_0_8_28 (.A(n_0_8_232), .ZN(n_0_8_21));
   NAND2_X1 i_0_8_29 (.A1(n_0_8_20), .A2(n_0_8_810), .ZN(n_0_86));
   XNOR2_X1 i_0_8_30 (.A(n_0_8_812), .B(n_0_8_788), .ZN(n_0_8_22));
   XNOR2_X1 i_0_8_31 (.A(n_0_8_22), .B(sub), .ZN(n_0_85));
   NAND2_X1 i_0_8_20 (.A1(n_0_8_800), .A2(n_0_8_596), .ZN(n_0_8_26));
   NAND2_X1 i_0_8_21 (.A1(n_0_8_9), .A2(n_0_8_18), .ZN(n_0_8_31));
   NAND4_X1 i_0_8_35 (.A1(n_0_8_33), .A2(n_0_8_735), .A3(n_0_8_31), .A4(
      n_0_8_857), .ZN(n_0_92));
   NAND4_X1 i_0_8_36 (.A1(n_0_8_26), .A2(n_0_8_824), .A3(n_0_8_852), .A4(
      n_0_8_853), .ZN(n_0_8_33));
   NAND2_X1 i_0_8_41 (.A1(n_0_8_806), .A2(n_0_40), .ZN(n_0_8_87));
   INV_X1 i_0_8_43 (.A(n_0_40), .ZN(n_0_8_95));
   XNOR2_X1 i_0_8_44 (.A(n_0_124), .B(n_0_8_11), .ZN(n_0_127));
   NAND2_X1 i_0_8_45 (.A1(n_0_8_3), .A2(n_0_8_1), .ZN(n_0_8_99));
   NAND3_X1 i_0_8_19 (.A1(n_0_8_13), .A2(sub), .A3(n_0_8_864), .ZN(n_0_8_100));
   NAND3_X1 i_0_8_47 (.A1(n_0_8_3), .A2(n_0_8_11), .A3(n_0_8_1), .ZN(n_0_54));
   NAND3_X1 i_0_8_48 (.A1(n_0_8_721), .A2(sub), .A3(n_0_8_5), .ZN(n_0_8_1));
   NAND2_X1 i_0_8_49 (.A1(n_0_8_4), .A2(n_0_8_10), .ZN(n_0_8_3));
   NAND2_X1 i_0_8_50 (.A1(n_0_8_721), .A2(n_0_8_5), .ZN(n_0_8_4));
   NAND2_X1 i_0_8_51 (.A1(n_0_8_863), .A2(in2[2]), .ZN(n_0_8_5));
   INV_X1 i_0_8_52 (.A(sub), .ZN(n_0_8_10));
   INV_X1 i_0_8_53 (.A(n_0_8_155), .ZN(n_0_8_11));
   BUF_X1 rt_shieldBuf__1__1__12 (.A(n_0_8_99), .Z(n_0_124));
   NAND2_X1 i_0_8_34 (.A1(n_0_8_485), .A2(n_0_8_714), .ZN(n_0_8_13));
   NAND2_X1 i_0_8_56 (.A1(n_0_8_714), .A2(n_0_8_10), .ZN(n_0_8_16));
   INV_X1 i_0_8_57 (.A(n_0_8_16), .ZN(n_0_8_102));
   NAND2_X1 i_0_8_61 (.A1(n_0_8_10), .A2(in2[3]), .ZN(n_0_8_15));
   INV_X1 i_0_8_62 (.A(n_0_8_15), .ZN(n_0_8_103));
   NAND2_X1 i_0_8_64 (.A1(n_0_8_29), .A2(n_0_8_30), .ZN(n_0_122));
   NAND2_X1 i_0_8_65 (.A1(n_0_121), .A2(n_0_60), .ZN(n_0_8_17));
   NOR2_X1 i_0_8_66 (.A1(n_0_121), .A2(n_0_60), .ZN(n_0_8_23));
   OAI21_X1 i_0_8_67 (.A(n_0_8_17), .B1(n_0_8_23), .B2(n_0_8_35), .ZN(n_0_113));
   XNOR2_X1 i_0_8_68 (.A(n_0_8_837), .B(n_0_8_768), .ZN(n_0_8_24));
   XNOR2_X1 i_0_8_69 (.A(n_0_8_24), .B(n_0_60), .ZN(n_0_8_25));
   NAND2_X1 i_0_8_70 (.A1(n_0_8_25), .A2(n_0_8_30), .ZN(n_0_8_27));
   NAND2_X1 i_0_8_71 (.A1(n_0_8_40), .A2(n_0_59), .ZN(n_0_8_28));
   NAND2_X1 i_0_8_72 (.A1(n_0_8_27), .A2(n_0_8_28), .ZN(n_0_123));
   XNOR2_X1 i_0_8_73 (.A(n_0_8_768), .B(sub), .ZN(n_0_8_29));
   INV_X1 i_0_8_74 (.A(n_0_59), .ZN(n_0_8_30));
   INV_X1 i_0_8_75 (.A(sub), .ZN(n_0_8_580));
   BUF_X1 i_0_8_76 (.A(n_0_8_580), .Z(n_0_8_32));
   INV_X1 i_0_8_77 (.A(sub), .ZN(n_0_8_110));
   XNOR2_X1 i_0_8_78 (.A(n_0_8_768), .B(n_0_8_110), .ZN(n_0_8_34));
   NAND2_X1 i_0_8_79 (.A1(n_0_8_34), .A2(n_0_59), .ZN(n_0_8_35));
   INV_X1 i_0_8_80 (.A(n_0_8_580), .ZN(n_0_8_595));
   NAND2_X1 i_0_8_5 (.A1(n_0_8_683), .A2(n_0_60), .ZN(n_0_8_36));
   NAND2_X1 i_0_8_82 (.A1(n_0_8_38), .A2(n_0_8_36), .ZN(n_0_119));
   INV_X1 i_0_8_83 (.A(n_0_60), .ZN(n_0_8_37));
   NAND2_X1 i_0_8_84 (.A1(n_0_8_684), .A2(n_0_8_37), .ZN(n_0_8_38));
   XNOR2_X1 i_0_8_85 (.A(n_0_8_837), .B(n_0_8_32), .ZN(n_0_121));
   XNOR2_X1 i_0_8_86 (.A(n_0_8_837), .B(n_0_8_32), .ZN(n_0_8_39));
   XNOR2_X1 i_0_8_87 (.A(n_0_8_39), .B(n_0_60), .ZN(n_0_8_40));
   NAND2_X1 i_0_8_88 (.A1(n_0_8_64), .A2(n_0_8_63), .ZN(n_0_35));
   NAND2_X1 i_0_8_89 (.A1(n_0_8_66), .A2(sub), .ZN(n_0_8_63));
   NAND2_X1 i_0_8_90 (.A1(n_0_8_65), .A2(n_0_8_41), .ZN(n_0_8_64));
   INV_X1 i_0_8_91 (.A(n_0_8_66), .ZN(n_0_8_65));
   XNOR2_X1 i_0_8_92 (.A(n_0_8_169), .B(n_0_8_151), .ZN(n_0_8_66));
   INV_X1 i_0_8_93 (.A(n_0_8_67), .ZN(n_0_38));
   OAI21_X1 i_0_8_94 (.A(n_0_8_68), .B1(n_0_8_151), .B2(n_0_8_695), .ZN(n_0_8_67));
   OAI21_X1 i_0_8_95 (.A(n_0_8_69), .B1(sub), .B2(n_0_8_149), .ZN(n_0_8_68));
   INV_X1 i_0_8_96 (.A(n_0_8_70), .ZN(n_0_8_69));
   OAI21_X1 i_0_8_97 (.A(n_0_8_191), .B1(n_0_8_169), .B2(n_0_8_41), .ZN(n_0_8_70));
   NAND2_X1 i_0_8_98 (.A1(n_0_8_71), .A2(n_0_8_73), .ZN(n_0_39));
   NAND2_X1 i_0_8_99 (.A1(n_0_8_72), .A2(sub), .ZN(n_0_8_71));
   NAND2_X1 i_0_8_100 (.A1(n_0_8_74), .A2(n_0_8_190), .ZN(n_0_8_72));
   NAND3_X1 i_0_8_101 (.A1(n_0_8_74), .A2(n_0_8_41), .A3(n_0_8_190), .ZN(
      n_0_8_73));
   NAND2_X1 i_0_8_102 (.A1(n_0_8_141), .A2(n_0_8_631), .ZN(n_0_8_74));
   INV_X1 i_0_8_103 (.A(sub), .ZN(n_0_8_41));
   AOI22_X1 i_0_8_104 (.A1(n_0_8_46), .A2(in1[9]), .B1(n_0_8_619), .B2(n_0_8_96), 
      .ZN(n_0_8_42));
   INV_X1 i_0_8_105 (.A(n_0_8_42), .ZN(n_0_50));
   AOI22_X1 i_0_8_106 (.A1(n_0_8_46), .A2(in1[10]), .B1(n_0_8_619), .B2(n_0_8_97), 
      .ZN(n_0_8_43));
   INV_X1 i_0_8_107 (.A(n_0_8_43), .ZN(n_0_37));
   AOI22_X1 i_0_8_108 (.A1(n_0_8_46), .A2(in1[11]), .B1(n_0_8_619), .B2(n_0_8_98), 
      .ZN(n_0_8_44));
   INV_X1 i_0_8_109 (.A(n_0_8_44), .ZN(n_0_44));
   NAND2_X1 i_0_8_110 (.A1(n_0_8_619), .A2(n_0_8_101), .ZN(n_0_8_45));
   NAND2_X1 i_0_8_111 (.A1(n_0_8_263), .A2(n_0_8_45), .ZN(n_0_58));
   NAND2_X1 i_0_8_112 (.A1(n_0_34), .A2(n_0_8_107), .ZN(n_0_8_150));
   BUF_X1 rt_shieldBuf__1__1__0 (.A(n_0_8_177), .Z(n_0_8_46));
   INV_X1 i_0_8_113 (.A(n_0_21), .ZN(n_0_8_587));
   INV_X1 i_0_8_114 (.A(n_0_8_714), .ZN(n_0_8_588));
   NAND2_X1 i_0_8_115 (.A1(n_0_8_47), .A2(n_0_8_48), .ZN(n_0_8_155));
   OAI21_X1 i_0_8_116 (.A(in1[2]), .B1(n_0_8_714), .B2(n_0_21), .ZN(n_0_8_47));
   NAND2_X1 i_0_8_117 (.A1(n_0_8_134), .A2(n_0_34), .ZN(n_0_8_48));
   OAI21_X1 i_0_8_118 (.A(in1[5]), .B1(n_0_8_714), .B2(n_0_8_620), .ZN(n_0_8_175));
   NAND2_X1 i_0_8_119 (.A1(n_0_8_92), .A2(n_0_34), .ZN(n_0_8_189));
   NAND2_X1 i_0_8_120 (.A1(n_0_8_52), .A2(n_0_8_53), .ZN(n_0_46));
   OAI21_X1 i_0_8_121 (.A(in1[6]), .B1(n_0_32), .B2(n_0_8_620), .ZN(n_0_8_52));
   NAND2_X1 i_0_8_122 (.A1(n_0_8_93), .A2(n_0_8_619), .ZN(n_0_8_53));
   NAND2_X1 i_0_8_123 (.A1(n_0_8_54), .A2(n_0_8_55), .ZN(n_0_47));
   OAI21_X1 i_0_8_124 (.A(in1[7]), .B1(n_0_32), .B2(n_0_8_620), .ZN(n_0_8_54));
   NAND2_X1 i_0_8_125 (.A1(n_0_8_94), .A2(n_0_8_619), .ZN(n_0_8_55));
   NAND2_X1 i_0_8_126 (.A1(n_0_8_851), .A2(n_0_8_56), .ZN(n_0_48));
   NAND2_X1 i_0_8_127 (.A1(in1[8]), .A2(n_0_8_177), .ZN(n_0_8_56));
   NAND2_X1 i_0_8_129 (.A1(n_0_8_85), .A2(n_0_8_86), .ZN(n_0_8_232));
   NAND2_X1 i_0_8_130 (.A1(n_0_8_109), .A2(n_0_34), .ZN(n_0_8_85));
   OAI21_X1 i_0_8_131 (.A(in1[4]), .B1(n_0_8_714), .B2(n_0_21), .ZN(n_0_8_86));
   BUF_X1 rt_shieldBuf__1__1__7 (.A(n_0_8_714), .Z(n_0_32));
   INV_X1 i_0_8_132 (.A(in1[4]), .ZN(n_0_8_88));
   INV_X1 i_0_8_133 (.A(in1[0]), .ZN(n_0_8_89));
   INV_X1 i_0_8_134 (.A(in1[5]), .ZN(n_0_8_90));
   INV_X1 i_0_8_135 (.A(in1[1]), .ZN(n_0_8_91));
   OAI22_X1 i_0_8_136 (.A1(n_0_8_131), .A2(n_0_8_562), .B1(n_0_8_80), .B2(
      n_0_8_262), .ZN(n_0_8_58));
   AOI22_X1 i_0_8_137 (.A1(n_0_8_129), .A2(n_0_8_564), .B1(n_0_8_58), .B2(
      n_0_8_756), .ZN(n_0_8_92));
   AOI22_X1 i_0_8_138 (.A1(n_0_8_178), .A2(n_0_8_755), .B1(n_0_8_112), .B2(
      n_0_8_563), .ZN(n_0_8_59));
   OAI22_X1 i_0_8_139 (.A1(n_0_8_126), .A2(n_0_8_262), .B1(n_0_8_59), .B2(
      n_0_8_562), .ZN(n_0_8_60));
   AOI22_X1 i_0_8_140 (.A1(n_0_8_60), .A2(n_0_8_756), .B1(n_0_8_58), .B2(
      n_0_8_564), .ZN(n_0_8_93));
   AOI22_X1 i_0_8_141 (.A1(n_0_8_176), .A2(n_0_8_755), .B1(n_0_8_245), .B2(
      n_0_8_563), .ZN(n_0_8_233));
   OAI22_X1 i_0_8_142 (.A1(n_0_8_131), .A2(n_0_8_262), .B1(n_0_8_233), .B2(
      n_0_8_562), .ZN(n_0_8_234));
   AOI22_X1 i_0_8_143 (.A1(n_0_8_60), .A2(n_0_8_250), .B1(n_0_8_234), .B2(
      n_0_8_756), .ZN(n_0_8_94));
   INV_X1 i_0_8_144 (.A(in1[8]), .ZN(n_0_8_75));
   AOI22_X1 i_0_8_145 (.A1(n_0_8_75), .A2(n_0_8_755), .B1(n_0_8_88), .B2(
      n_0_8_563), .ZN(n_0_8_76));
   OAI22_X1 i_0_8_146 (.A1(n_0_8_59), .A2(n_0_8_262), .B1(n_0_8_76), .B2(
      n_0_8_562), .ZN(n_0_8_235));
   AOI22_X1 i_0_8_149 (.A1(n_0_8_235), .A2(n_0_8_564), .B1(n_0_8_811), .B2(
      n_0_8_756), .ZN(n_0_8_96));
   OAI22_X1 i_0_8_150 (.A1(n_0_8_76), .A2(n_0_8_262), .B1(n_0_8_228), .B2(
      n_0_8_562), .ZN(n_0_8_79));
   AOI22_X1 i_0_8_3 (.A1(n_0_8_811), .A2(n_0_8_250), .B1(n_0_8_79), .B2(
      n_0_8_120), .ZN(n_0_8_97));
   AOI22_X1 i_0_8_152 (.A1(n_0_8_79), .A2(n_0_8_564), .B1(n_0_8_218), .B2(
      n_0_8_120), .ZN(n_0_8_98));
   AOI22_X1 i_0_8_153 (.A1(n_0_8_227), .A2(n_0_8_250), .B1(n_0_8_165), .B2(
      n_0_8_756), .ZN(n_0_8_101));
   AOI22_X1 i_0_8_154 (.A1(n_0_8_161), .A2(n_0_8_564), .B1(n_0_8_162), .B2(
      n_0_8_756), .ZN(n_0_8_107));
   NOR2_X1 i_0_8_155 (.A1(n_0_8_563), .A2(n_0_8_245), .ZN(n_0_8_80));
   AOI21_X1 i_0_8_156 (.A(n_0_8_81), .B1(n_0_8_756), .B2(n_0_8_129), .ZN(
      n_0_8_109));
   AOI21_X1 i_0_8_157 (.A(n_0_8_756), .B1(n_0_8_83), .B2(n_0_8_82), .ZN(n_0_8_81));
   OAI21_X1 i_0_8_158 (.A(n_0_8_262), .B1(n_0_8_563), .B2(n_0_8_245), .ZN(
      n_0_8_82));
   OAI21_X1 i_0_8_159 (.A(n_0_8_562), .B1(n_0_8_563), .B2(n_0_8_84), .ZN(
      n_0_8_83));
   INV_X1 i_0_8_160 (.A(in1[1]), .ZN(n_0_8_84));
   NAND2_X1 i_0_8_161 (.A1(n_0_8_104), .A2(n_0_8_762), .ZN(n_0_8_243));
   INV_X1 i_0_8_162 (.A(in1[3]), .ZN(n_0_8_245));
   NAND2_X1 i_0_8_163 (.A1(n_0_8_562), .A2(in1[1]), .ZN(n_0_8_249));
   NAND3_X1 i_0_8_164 (.A1(n_0_8_119), .A2(n_0_8_755), .A3(n_0_8_564), .ZN(
      n_0_8_104));
   NAND2_X1 i_0_8_165 (.A1(n_0_8_562), .A2(in1[0]), .ZN(n_0_8_111));
   INV_X1 i_0_8_166 (.A(in1[2]), .ZN(n_0_8_112));
   NAND2_X1 i_0_8_167 (.A1(n_0_8_563), .A2(n_0_8_89), .ZN(n_0_8_114));
   INV_X1 i_0_8_168 (.A(n_0_8_563), .ZN(n_0_8_115));
   INV_X1 i_0_8_169 (.A(n_0_8_88), .ZN(n_0_8_116));
   INV_X1 i_0_8_170 (.A(n_0_8_89), .ZN(n_0_8_117));
   NAND2_X1 i_0_8_171 (.A1(n_0_8_116), .A2(n_0_8_117), .ZN(n_0_8_118));
   OAI21_X1 i_0_8_172 (.A(n_0_8_111), .B1(n_0_8_562), .B2(n_0_8_112), .ZN(
      n_0_8_119));
   INV_X1 i_0_8_173 (.A(n_0_8_562), .ZN(n_0_8_121));
   INV_X1 i_0_8_174 (.A(n_0_8_112), .ZN(n_0_8_122));
   NAND2_X1 i_0_8_175 (.A1(n_0_8_121), .A2(n_0_8_122), .ZN(n_0_8_123));
   NAND2_X1 i_0_8_176 (.A1(n_0_8_111), .A2(n_0_8_123), .ZN(n_0_8_124));
   NOR2_X1 i_0_8_177 (.A1(n_0_8_563), .A2(n_0_8_564), .ZN(n_0_8_125));
   NAND3_X1 i_0_8_178 (.A1(n_0_8_135), .A2(n_0_8_136), .A3(n_0_8_118), .ZN(
      n_0_8_126));
   INV_X1 i_0_8_179 (.A(n_0_8_118), .ZN(n_0_8_127));
   OAI21_X1 i_0_8_180 (.A(n_0_8_562), .B1(n_0_8_563), .B2(n_0_8_112), .ZN(
      n_0_8_128));
   NAND2_X1 i_0_8_181 (.A1(n_0_8_140), .A2(n_0_8_128), .ZN(n_0_8_129));
   INV_X1 i_0_8_182 (.A(n_0_8_563), .ZN(n_0_8_130));
   AOI22_X1 i_0_8_183 (.A1(n_0_8_90), .A2(n_0_8_755), .B1(n_0_8_91), .B2(
      n_0_8_563), .ZN(n_0_8_131));
   NAND2_X1 i_0_8_184 (.A1(n_0_8_124), .A2(n_0_8_125), .ZN(n_0_8_132));
   NAND4_X1 i_0_8_185 (.A1(n_0_8_130), .A2(n_0_8_262), .A3(n_0_8_564), .A4(
      in1[1]), .ZN(n_0_8_133));
   NAND2_X1 i_0_8_186 (.A1(n_0_8_132), .A2(n_0_8_133), .ZN(n_0_8_134));
   NAND2_X1 i_0_8_187 (.A1(n_0_8_563), .A2(n_0_8_114), .ZN(n_0_8_135));
   NAND2_X1 i_0_8_188 (.A1(n_0_8_115), .A2(n_0_8_116), .ZN(n_0_8_136));
   NAND2_X1 i_0_8_189 (.A1(n_0_8_114), .A2(n_0_8_563), .ZN(n_0_8_137));
   NAND2_X1 i_0_8_190 (.A1(n_0_8_115), .A2(n_0_8_116), .ZN(n_0_8_138));
   NOR2_X1 i_0_8_191 (.A1(n_0_8_562), .A2(n_0_8_127), .ZN(n_0_8_139));
   NAND3_X1 i_0_8_192 (.A1(n_0_8_137), .A2(n_0_8_138), .A3(n_0_8_139), .ZN(
      n_0_8_140));
   INV_X1 i_0_8_193 (.A(n_0_8_563), .ZN(n_0_8_143));
   INV_X1 i_0_8_194 (.A(n_0_8_562), .ZN(n_0_8_144));
   NAND2_X1 i_0_8_195 (.A1(n_0_8_143), .A2(n_0_8_144), .ZN(n_0_8_105));
   BUF_X1 rt_shieldBuf__1__1__9 (.A(n_0_8_564), .Z(n_0_8_250));
   INV_X1 i_0_8_196 (.A(sub), .ZN(n_0_8_589));
   NAND2_X1 i_0_8_197 (.A1(n_0_8_606), .A2(n_0_8_589), .ZN(n_0_8_106));
   BUF_X1 rt_shieldBuf__1__1__10 (.A(n_0_8_673), .Z(n_0_8_169));
   INV_X1 i_0_8_198 (.A(n_0_34), .ZN(n_0_8_108));
   NAND2_X1 i_0_8_199 (.A1(n_0_8_151), .A2(n_0_55), .ZN(n_0_8_113));
   BUF_X1 rt_shieldBuf__1__1__13 (.A(n_0_8_756), .Z(n_0_8_120));
   NAND2_X1 i_0_8_200 (.A1(n_0_8_671), .A2(n_0_8_172), .ZN(n_0_8_590));
   OAI21_X1 i_0_8_201 (.A(in1[1]), .B1(n_0_8_714), .B2(n_0_21), .ZN(n_0_8_591));
   NOR2_X1 i_0_8_202 (.A1(n_0_8_108), .A2(n_0_8_105), .ZN(n_0_8_172));
   OAI21_X1 i_0_8_203 (.A(in1[1]), .B1(n_0_8_714), .B2(n_0_21), .ZN(n_0_8_148));
   OAI21_X1 i_0_8_204 (.A(n_0_8_148), .B1(n_0_8_108), .B2(n_0_8_105), .ZN(
      n_0_8_157));
   NAND3_X1 i_0_8_205 (.A1(n_0_8_148), .A2(n_0_8_171), .A3(n_0_8_170), .ZN(
      n_0_8_158));
   NAND2_X1 i_0_8_206 (.A1(n_0_8_157), .A2(n_0_8_158), .ZN(n_0_8_141));
   NAND2_X1 i_0_8_207 (.A1(n_0_8_146), .A2(in1[1]), .ZN(n_0_8_170));
   NAND2_X1 i_0_8_208 (.A1(n_0_8_564), .A2(in1[0]), .ZN(n_0_8_171));
   INV_X1 i_0_8_209 (.A(n_0_8_564), .ZN(n_0_8_146));
   INV_X1 i_0_8_210 (.A(in1[0]), .ZN(n_0_8_600));
   INV_X1 i_0_8_211 (.A(in1[1]), .ZN(n_0_8_601));
   NAND2_X1 i_0_8_212 (.A1(n_0_8_588), .A2(n_0_8_587), .ZN(n_0_8_177));
   INV_X1 i_0_8_213 (.A(in1[0]), .ZN(n_0_8_142));
   INV_X1 i_0_8_214 (.A(n_0_55), .ZN(n_0_8_182));
   NAND2_X1 i_0_8_215 (.A1(n_0_8_621), .A2(n_0_8_182), .ZN(n_0_8_183));
   INV_X1 i_0_8_216 (.A(n_0_8_183), .ZN(n_0_8_145));
   INV_X1 i_0_8_217 (.A(n_0_8_142), .ZN(n_0_8_185));
   NOR2_X1 i_0_8_218 (.A1(n_0_55), .A2(n_0_8_185), .ZN(n_0_8_147));
   NAND2_X1 i_0_8_219 (.A1(n_0_8_616), .A2(n_0_8_106), .ZN(n_0_8_188));
   NAND2_X1 i_0_8_220 (.A1(n_0_8_159), .A2(n_0_8_188), .ZN(n_0_8_251));
   NAND2_X1 i_0_8_221 (.A1(n_0_8_585), .A2(n_0_8_606), .ZN(n_0_8_190));
   NAND2_X1 i_0_8_222 (.A1(n_0_8_151), .A2(n_0_8_695), .ZN(n_0_8_191));
   INV_X1 i_0_8_223 (.A(n_0_8_673), .ZN(n_0_8_149));
   OAI21_X1 i_0_8_224 (.A(n_0_8_621), .B1(n_0_8_588), .B2(n_0_8_142), .ZN(
      n_0_8_151));
   INV_X1 i_0_8_225 (.A(n_0_8_142), .ZN(n_0_8_152));
   NOR2_X1 i_0_8_226 (.A1(n_0_55), .A2(n_0_8_152), .ZN(n_0_8_592));
   INV_X1 i_0_8_227 (.A(n_0_55), .ZN(n_0_8_593));
   NAND3_X1 i_0_8_228 (.A1(n_0_8_614), .A2(n_0_8_237), .A3(n_0_8_113), .ZN(
      n_0_8_153));
   AOI21_X1 i_0_8_229 (.A(n_0_8_41), .B1(n_0_8_141), .B2(n_0_8_606), .ZN(
      n_0_8_154));
   NAND2_X1 i_0_8_230 (.A1(n_0_8_153), .A2(n_0_8_154), .ZN(n_0_8_258));
   NAND2_X1 i_0_8_231 (.A1(n_0_8_151), .A2(n_0_55), .ZN(n_0_8_156));
   NAND3_X1 i_0_8_232 (.A1(n_0_8_615), .A2(n_0_8_164), .A3(n_0_8_156), .ZN(
      n_0_8_159));
   NAND2_X1 i_0_8_233 (.A1(n_0_8_145), .A2(n_0_8_588), .ZN(n_0_8_160));
   NAND2_X1 i_0_8_234 (.A1(n_0_8_621), .A2(n_0_8_147), .ZN(n_0_8_163));
   NAND3_X1 i_0_8_235 (.A1(n_0_8_673), .A2(n_0_8_160), .A3(n_0_8_163), .ZN(
      n_0_8_164));
   NAND2_X1 i_0_8_236 (.A1(n_0_8_193), .A2(n_0_8_195), .ZN(n_0_8_161));
   AOI21_X1 i_0_8_237 (.A(n_0_8_203), .B1(n_0_8_207), .B2(n_0_8_562), .ZN(
      n_0_8_162));
   OAI22_X1 i_0_8_238 (.A1(n_0_8_562), .A2(n_0_8_181), .B1(n_0_8_219), .B2(
      n_0_8_262), .ZN(n_0_8_165));
   INV_X1 i_0_8_239 (.A(in1[9]), .ZN(n_0_8_166));
   NAND2_X1 i_0_8_240 (.A1(n_0_8_167), .A2(n_0_8_263), .ZN(n_0_45));
   NAND4_X1 i_0_8_241 (.A1(n_0_8_179), .A2(n_0_8_168), .A3(n_0_34), .A4(
      n_0_8_187), .ZN(n_0_8_167));
   NAND2_X1 i_0_8_242 (.A1(n_0_8_174), .A2(n_0_8_173), .ZN(n_0_8_168));
   INV_X1 i_0_8_243 (.A(n_0_8_214), .ZN(n_0_8_173));
   INV_X1 i_0_8_244 (.A(n_0_8_219), .ZN(n_0_8_174));
   NAND3_X1 i_0_8_245 (.A1(n_0_8_186), .A2(n_0_8_564), .A3(n_0_8_180), .ZN(
      n_0_8_179));
   INV_X1 i_0_8_246 (.A(n_0_8_181), .ZN(n_0_8_180));
   NAND2_X1 i_0_8_247 (.A1(n_0_8_208), .A2(n_0_8_184), .ZN(n_0_8_181));
   NAND2_X1 i_0_8_248 (.A1(n_0_8_563), .A2(in1[9]), .ZN(n_0_8_184));
   INV_X1 i_0_8_249 (.A(n_0_8_562), .ZN(n_0_8_186));
   OAI21_X1 i_0_8_250 (.A(n_0_8_756), .B1(n_0_8_197), .B2(n_0_8_200), .ZN(
      n_0_8_187));
   OAI211_X1 i_0_8_251 (.A(n_0_8_263), .B(n_0_8_192), .C1(n_0_8_196), .C2(
      n_0_8_201), .ZN(n_0_49));
   NAND4_X1 i_0_8_252 (.A1(n_0_8_193), .A2(n_0_34), .A3(n_0_8_756), .A4(
      n_0_8_195), .ZN(n_0_8_192));
   OAI211_X1 i_0_8_253 (.A(n_0_8_194), .B(n_0_8_563), .C1(n_0_8_221), .C2(
      n_0_8_562), .ZN(n_0_8_193));
   NAND2_X1 i_0_8_254 (.A1(n_0_8_562), .A2(in1[9]), .ZN(n_0_8_194));
   INV_X1 i_0_8_255 (.A(n_0_8_200), .ZN(n_0_8_195));
   OR2_X1 i_0_8_256 (.A1(n_0_8_197), .A2(n_0_8_200), .ZN(n_0_8_196));
   AOI21_X1 i_0_8_257 (.A(n_0_8_755), .B1(n_0_8_198), .B2(n_0_8_199), .ZN(
      n_0_8_197));
   NAND2_X1 i_0_8_258 (.A1(n_0_8_262), .A2(n_0_8_230), .ZN(n_0_8_198));
   NAND2_X1 i_0_8_259 (.A1(n_0_8_562), .A2(n_0_8_75), .ZN(n_0_8_199));
   NOR2_X1 i_0_8_260 (.A1(n_0_8_563), .A2(in1[12]), .ZN(n_0_8_200));
   NAND2_X1 i_0_8_261 (.A1(n_0_34), .A2(n_0_8_564), .ZN(n_0_8_201));
   NAND4_X1 i_0_8_81 (.A1(n_0_8_206), .A2(n_0_8_263), .A3(n_0_8_204), .A4(
      n_0_8_202), .ZN(n_0_60));
   NAND2_X1 i_0_8_263 (.A1(n_0_34), .A2(n_0_8_203), .ZN(n_0_8_202));
   NOR2_X1 i_0_8_264 (.A1(n_0_8_562), .A2(n_0_8_215), .ZN(n_0_8_203));
   NAND4_X1 i_0_8_265 (.A1(n_0_8_205), .A2(n_0_34), .A3(n_0_8_562), .A4(
      n_0_8_756), .ZN(n_0_8_204));
   NAND2_X1 i_0_8_266 (.A1(n_0_8_208), .A2(n_0_8_211), .ZN(n_0_8_205));
   NAND4_X1 i_0_8_267 (.A1(n_0_8_207), .A2(n_0_34), .A3(n_0_8_562), .A4(
      n_0_8_564), .ZN(n_0_8_206));
   OAI21_X1 i_0_8_268 (.A(n_0_8_208), .B1(n_0_8_230), .B2(n_0_8_755), .ZN(
      n_0_8_207));
   NAND2_X1 i_0_8_269 (.A1(n_0_8_755), .A2(in1[12]), .ZN(n_0_8_208));
   NAND2_X1 i_0_8_270 (.A1(n_0_8_209), .A2(n_0_8_263), .ZN(n_0_93));
   NAND2_X1 i_0_8_271 (.A1(n_0_8_210), .A2(n_0_34), .ZN(n_0_8_209));
   OAI22_X1 i_0_8_272 (.A1(n_0_8_212), .A2(n_0_8_215), .B1(n_0_8_214), .B2(
      n_0_8_211), .ZN(n_0_8_210));
   NAND2_X1 i_0_8_273 (.A1(n_0_8_563), .A2(in1[11]), .ZN(n_0_8_211));
   INV_X1 i_0_8_274 (.A(n_0_8_213), .ZN(n_0_8_212));
   NAND3_X1 i_0_8_275 (.A1(n_0_8_564), .A2(n_0_8_563), .A3(n_0_8_562), .ZN(
      n_0_8_213));
   NAND2_X1 i_0_8_276 (.A1(n_0_8_564), .A2(n_0_8_562), .ZN(n_0_8_214));
   INV_X1 i_0_8_277 (.A(in1[12]), .ZN(n_0_8_215));
   INV_X1 i_0_8_278 (.A(n_0_8_223), .ZN(n_0_8_261));
   INV_X1 i_0_8_279 (.A(in1[7]), .ZN(n_0_8_176));
   INV_X1 i_0_8_280 (.A(in1[6]), .ZN(n_0_8_178));
   NAND2_X1 i_0_8_281 (.A1(n_0_8_216), .A2(n_0_8_263), .ZN(n_0_53));
   NAND3_X1 i_0_8_282 (.A1(n_0_8_217), .A2(n_0_34), .A3(n_0_8_226), .ZN(
      n_0_8_216));
   NAND2_X1 i_0_8_283 (.A1(n_0_8_564), .A2(n_0_8_218), .ZN(n_0_8_217));
   OAI21_X1 i_0_8_284 (.A(n_0_8_222), .B1(n_0_8_562), .B2(n_0_8_219), .ZN(
      n_0_8_218));
   OAI21_X1 i_0_8_285 (.A(n_0_8_220), .B1(n_0_8_221), .B2(n_0_8_563), .ZN(
      n_0_8_219));
   NAND2_X1 i_0_8_286 (.A1(n_0_8_563), .A2(in1[7]), .ZN(n_0_8_220));
   INV_X1 i_0_8_287 (.A(in1[11]), .ZN(n_0_8_221));
   NAND2_X1 i_0_8_288 (.A1(n_0_8_223), .A2(n_0_8_562), .ZN(n_0_8_222));
   OAI21_X1 i_0_8_289 (.A(n_0_8_224), .B1(n_0_8_563), .B2(n_0_8_225), .ZN(
      n_0_8_223));
   NAND2_X1 i_0_8_290 (.A1(n_0_8_563), .A2(n_0_8_90), .ZN(n_0_8_224));
   INV_X1 i_0_8_291 (.A(n_0_8_166), .ZN(n_0_8_225));
   NAND2_X1 i_0_8_292 (.A1(n_0_8_227), .A2(n_0_8_756), .ZN(n_0_8_226));
   OAI21_X1 i_0_8_293 (.A(n_0_8_231), .B1(n_0_8_262), .B2(n_0_8_228), .ZN(
      n_0_8_227));
   OAI21_X1 i_0_8_294 (.A(n_0_8_229), .B1(n_0_8_230), .B2(n_0_8_563), .ZN(
      n_0_8_228));
   NAND2_X1 i_0_8_295 (.A1(n_0_8_563), .A2(in1[6]), .ZN(n_0_8_229));
   INV_X1 i_0_8_296 (.A(in1[10]), .ZN(n_0_8_230));
   OAI211_X1 i_0_8_297 (.A(n_0_8_208), .B(n_0_8_262), .C1(n_0_8_755), .C2(
      n_0_8_75), .ZN(n_0_8_231));
   INV_X1 i_0_8_298 (.A(n_0_8_562), .ZN(n_0_8_262));
   NAND2_X1 i_0_8_299 (.A1(n_0_8_177), .A2(in1[12]), .ZN(n_0_8_263));
   INV_X1 i_0_8_300 (.A(n_0_8_673), .ZN(n_0_8_236));
   NAND2_X1 i_0_8_301 (.A1(n_0_8_629), .A2(n_0_8_236), .ZN(n_0_8_237));
   OAI21_X1 i_0_8_302 (.A(in2[4]), .B1(n_0_34), .B2(n_0_8_400), .ZN(n_0_8_238));
   NAND2_X1 i_0_8_303 (.A1(n_0_8_238), .A2(n_0_8_282), .ZN(n_0_8_268));
   OAI21_X1 i_0_8_304 (.A(in2[6]), .B1(n_0_34), .B2(n_0_8_620), .ZN(n_0_8_239));
   NAND2_X1 i_0_8_305 (.A1(n_0_8_239), .A2(n_0_8_439), .ZN(n_0_26));
   OAI21_X1 i_0_8_306 (.A(in2[7]), .B1(n_0_34), .B2(n_0_8_620), .ZN(n_0_8_240));
   NAND2_X1 i_0_8_307 (.A1(n_0_8_240), .A2(n_0_8_285), .ZN(n_0_27));
   OAI21_X1 i_0_8_308 (.A(in2[9]), .B1(n_0_8_276), .B2(n_0_8_400), .ZN(n_0_8_241));
   NAND2_X1 i_0_8_309 (.A1(n_0_8_241), .A2(n_0_8_325), .ZN(n_0_29));
   OAI21_X1 i_0_8_310 (.A(in2[10]), .B1(n_0_8_276), .B2(n_0_8_400), .ZN(
      n_0_8_242));
   NAND2_X1 i_0_8_311 (.A1(n_0_8_242), .A2(n_0_8_681), .ZN(n_0_24));
   NAND2_X1 i_0_8_313 (.A1(n_0_8_858), .A2(n_0_8_307), .ZN(n_0_41));
   INV_X1 i_0_8_314 (.A(in2[0]), .ZN(n_0_8_244));
   BUF_X1 rt_shieldBuf__1 (.A(n_0_34), .Z(n_0_8_276));
   INV_X1 i_0_8_315 (.A(in2[10]), .ZN(n_0_8_594));
   INV_X1 i_0_8_316 (.A(in2[11]), .ZN(n_0_8_286));
   INV_X1 i_0_8_317 (.A(in2[12]), .ZN(n_0_8_287));
   INV_X1 i_0_8_318 (.A(in2[7]), .ZN(n_0_8_246));
   INV_X1 i_0_8_319 (.A(in2[9]), .ZN(n_0_8_247));
   INV_X1 i_0_8_320 (.A(in2[5]), .ZN(n_0_8_248));
   INV_X1 i_0_8_59 (.A(in2[3]), .ZN(n_0_8_292));
   INV_X1 i_0_8_322 (.A(in2[8]), .ZN(n_0_8_294));
   INV_X1 i_0_8_323 (.A(in2[4]), .ZN(n_0_8_309));
   INV_X1 i_0_8_324 (.A(in2[0]), .ZN(n_0_8_252));
   INV_X1 i_0_8_325 (.A(in2[2]), .ZN(n_0_8_253));
   INV_X1 i_0_8_326 (.A(in2[1]), .ZN(n_0_8_254));
   INV_X1 i_0_8_327 (.A(in2[6]), .ZN(n_0_8_255));
   BUF_X1 i_0_8_328 (.A(n_0_8_246), .Z(n_0_8_256));
   BUF_X1 i_0_8_329 (.A(n_0_8_247), .Z(n_0_8_257));
   BUF_X1 i_0_8_330 (.A(n_0_8_294), .Z(n_0_8_315));
   BUF_X1 i_0_8_38 (.A(n_0_8_829), .Z(n_0_8_316));
   BUF_X1 i_0_8_333 (.A(n_0_8_255), .Z(n_0_8_259));
   OAI21_X1 i_0_8_334 (.A(n_0_8_394), .B1(n_0_8_413), .B2(n_0_8_633), .ZN(
      n_0_8_260));
   INV_X1 i_0_8_40 (.A(in1[15]), .ZN(n_0_8_320));
   INV_X1 i_0_8_42 (.A(in2[15]), .ZN(n_0_8_321));
   INV_X1 i_0_8_32 (.A(in1[14]), .ZN(n_0_8_264));
   NAND2_X1 i_0_8_338 (.A1(n_0_8_364), .A2(n_0_8_357), .ZN(n_0_8_265));
   INV_X1 i_0_8_339 (.A(in2[13]), .ZN(n_0_8_266));
   NOR2_X1 i_0_8_340 (.A1(n_0_8_266), .A2(in1[13]), .ZN(n_0_8_267));
   NAND2_X1 i_0_8_63 (.A1(n_0_8_265), .A2(n_0_8_267), .ZN(n_0_8_342));
   NAND2_X1 i_0_8_33 (.A1(n_0_8_264), .A2(in2[14]), .ZN(n_0_8_269));
   NAND2_X1 i_0_8_60 (.A1(n_0_8_275), .A2(n_0_8_269), .ZN(n_0_8_270));
   NAND2_X1 i_0_8_331 (.A1(n_0_8_321), .A2(in1[15]), .ZN(n_0_8_271));
   NAND2_X1 i_0_8_335 (.A1(n_0_8_320), .A2(in2[15]), .ZN(n_0_8_272));
   INV_X1 i_0_8_346 (.A(in1[13]), .ZN(n_0_8_273));
   INV_X1 i_0_8_336 (.A(in1[13]), .ZN(n_0_8_274));
   NAND2_X1 i_0_8_128 (.A1(n_0_8_274), .A2(in2[13]), .ZN(n_0_8_275));
   NAND3_X1 i_0_8_349 (.A1(n_0_8_571), .A2(in2[1]), .A3(n_0_8_636), .ZN(
      n_0_8_343));
   INV_X1 i_0_8_350 (.A(in2[1]), .ZN(n_0_8_277));
   INV_X1 i_0_8_351 (.A(in2[0]), .ZN(n_0_8_278));
   NAND2_X1 i_0_8_352 (.A1(n_0_8_436), .A2(n_0_8_404), .ZN(n_0_8_279));
   INV_X1 i_0_8_353 (.A(n_0_8_714), .ZN(n_0_8_280));
   AOI21_X1 i_0_8_354 (.A(n_0_8_280), .B1(n_0_8_260), .B2(n_0_8_844), .ZN(
      n_0_8_281));
   NAND2_X1 i_0_8_355 (.A1(n_0_8_279), .A2(n_0_8_281), .ZN(n_0_8_282));
   NAND2_X1 i_0_8_356 (.A1(n_0_8_477), .A2(n_0_8_844), .ZN(n_0_8_283));
   NAND2_X1 i_0_8_357 (.A1(n_0_8_422), .A2(n_0_8_404), .ZN(n_0_8_284));
   NAND3_X1 i_0_8_358 (.A1(n_0_8_283), .A2(n_0_8_284), .A3(n_0_8_714), .ZN(
      n_0_8_285));
   NAND2_X1 i_0_8_151 (.A1(n_0_8_418), .A2(n_0_8_404), .ZN(n_0_8_344));
   NAND2_X1 i_0_8_337 (.A1(n_0_8_436), .A2(n_0_8_844), .ZN(n_0_8_345));
   NAND2_X1 i_0_8_361 (.A1(n_0_21), .A2(in2[1]), .ZN(n_0_8_288));
   INV_X1 i_0_8_362 (.A(n_0_8_288), .ZN(n_0_8_289));
   NAND2_X1 i_0_8_364 (.A1(n_0_21), .A2(in2[5]), .ZN(n_0_8_291));
   INV_X1 i_0_8_365 (.A(n_0_8_291), .ZN(n_0_8_347));
   NAND2_X1 i_0_8_369 (.A1(n_0_8_571), .A2(n_0_8_294), .ZN(n_0_8_295));
   NAND2_X1 i_0_8_370 (.A1(n_0_8_832), .A2(n_0_8_309), .ZN(n_0_8_296));
   NAND2_X1 i_0_8_371 (.A1(n_0_8_295), .A2(n_0_8_296), .ZN(n_0_8_297));
   INV_X1 i_0_8_372 (.A(n_0_8_633), .ZN(n_0_8_298));
   NAND2_X1 i_0_8_373 (.A1(n_0_8_571), .A2(n_0_8_255), .ZN(n_0_8_299));
   NAND2_X1 i_0_8_374 (.A1(n_0_8_832), .A2(n_0_8_253), .ZN(n_0_8_300));
   NAND2_X1 i_0_8_375 (.A1(n_0_8_299), .A2(n_0_8_300), .ZN(n_0_8_301));
   INV_X1 i_0_8_377 (.A(in2[12]), .ZN(n_0_8_302));
   NAND3_X1 i_0_8_378 (.A1(n_0_8_430), .A2(n_0_8_356), .A3(n_0_8_535), .ZN(
      n_0_8_303));
   NAND2_X1 i_0_8_379 (.A1(n_0_21), .A2(in2[8]), .ZN(n_0_8_304));
   INV_X1 i_0_8_380 (.A(n_0_8_304), .ZN(n_0_8_305));
   AOI21_X1 i_0_8_381 (.A(n_0_8_305), .B1(n_0_34), .B2(in2[8]), .ZN(n_0_8_306));
   NAND2_X1 i_0_8_382 (.A1(n_0_8_303), .A2(n_0_8_306), .ZN(n_0_28));
   NAND2_X1 i_0_8_359 (.A1(n_0_8_809), .A2(n_0_8_714), .ZN(n_0_8_307));
   NAND2_X1 i_0_8_384 (.A1(n_0_8_571), .A2(n_0_8_246), .ZN(n_0_8_308));
   NAND2_X1 i_0_8_386 (.A1(n_0_8_308), .A2(n_0_8_830), .ZN(n_0_8_310));
   INV_X1 i_0_8_387 (.A(n_0_8_633), .ZN(n_0_8_311));
   NAND2_X1 i_0_8_342 (.A1(n_0_8_571), .A2(n_0_8_248), .ZN(n_0_8_312));
   NAND2_X1 i_0_8_389 (.A1(n_0_8_312), .A2(n_0_8_453), .ZN(n_0_8_313));
   INV_X1 i_0_8_345 (.A(in2[13]), .ZN(n_0_8_314));
   INV_X1 i_0_8_391 (.A(in2[12]), .ZN(n_0_8_348));
   INV_X1 i_0_8_392 (.A(in1[14]), .ZN(n_0_8_317));
   INV_X1 i_0_8_343 (.A(n_0_8_571), .ZN(n_0_8_318));
   INV_X1 i_0_8_394 (.A(n_0_8_278), .ZN(n_0_8_319));
   INV_X1 i_0_8_395 (.A(n_0_8_714), .ZN(n_0_8_322));
   AOI21_X1 i_0_8_396 (.A(n_0_8_322), .B1(n_0_8_349), .B2(n_0_8_844), .ZN(
      n_0_8_323));
   INV_X1 i_0_8_397 (.A(n_0_8_404), .ZN(n_0_8_324));
   OAI21_X1 i_0_8_398 (.A(n_0_8_323), .B1(n_0_8_451), .B2(n_0_8_324), .ZN(
      n_0_8_325));
   INV_X1 i_0_8_344 (.A(n_0_8_368), .ZN(n_0_8_326));
   INV_X1 i_0_8_400 (.A(n_0_8_257), .ZN(n_0_8_327));
   NAND2_X1 i_0_8_388 (.A1(n_0_8_326), .A2(n_0_8_327), .ZN(n_0_8_328));
   INV_X1 i_0_8_393 (.A(n_0_8_636), .ZN(n_0_8_329));
   NAND3_X1 i_0_8_399 (.A1(n_0_8_328), .A2(n_0_8_367), .A3(n_0_8_329), .ZN(
      n_0_8_330));
   INV_X1 i_0_8_401 (.A(n_0_8_785), .ZN(n_0_8_331));
   INV_X1 i_0_8_405 (.A(n_0_8_348), .ZN(n_0_8_332));
   NAND2_X1 i_0_8_402 (.A1(n_0_8_331), .A2(n_0_8_332), .ZN(n_0_8_333));
   NAND2_X1 i_0_8_403 (.A1(n_0_8_340), .A2(n_0_8_286), .ZN(n_0_8_334));
   INV_X1 i_0_8_404 (.A(n_0_8_571), .ZN(n_0_8_335));
   INV_X1 i_0_8_406 (.A(n_0_8_340), .ZN(n_0_8_336));
   OAI21_X1 i_0_8_407 (.A(n_0_8_334), .B1(n_0_8_335), .B2(n_0_8_336), .ZN(
      n_0_8_337));
   NAND2_X1 i_0_8_408 (.A1(n_0_8_333), .A2(n_0_8_337), .ZN(n_0_8_338));
   NAND2_X1 i_0_8_409 (.A1(n_0_8_330), .A2(n_0_8_338), .ZN(n_0_8_339));
   NAND2_X1 i_0_8_413 (.A1(n_0_8_342), .A2(n_0_8_377), .ZN(n_0_8_340));
   NOR2_X1 i_0_8_414 (.A1(n_0_8_287), .A2(n_0_8_633), .ZN(n_0_8_361));
   INV_X1 i_0_8_415 (.A(n_0_8_633), .ZN(n_0_8_341));
   NAND2_X1 i_0_8_416 (.A1(n_0_8_341), .A2(n_0_8_287), .ZN(n_0_8_362));
   INV_X1 i_0_8_417 (.A(n_0_8_318), .ZN(n_0_8_372));
   INV_X1 i_0_8_418 (.A(n_0_8_302), .ZN(n_0_8_597));
   INV_X1 i_0_8_419 (.A(n_0_8_611), .ZN(n_0_8_373));
   NAND2_X1 i_0_8_410 (.A1(n_0_8_339), .A2(n_0_8_844), .ZN(n_0_8_374));
   INV_X1 i_0_8_421 (.A(n_0_8_714), .ZN(n_0_8_346));
   AOI21_X1 i_0_8_422 (.A(n_0_8_346), .B1(n_0_8_843), .B2(n_0_8_821), .ZN(
      n_0_8_375));
   INV_X1 i_0_8_423 (.A(in2[12]), .ZN(n_0_8_376));
   NAND2_X1 i_0_8_425 (.A1(n_0_8_350), .A2(n_0_8_351), .ZN(n_0_8_349));
   NAND2_X1 i_0_8_426 (.A1(n_0_8_297), .A2(n_0_8_298), .ZN(n_0_8_350));
   NAND2_X1 i_0_8_427 (.A1(n_0_8_301), .A2(n_0_8_633), .ZN(n_0_8_351));
   NAND2_X1 i_0_8_428 (.A1(n_0_8_298), .A2(n_0_8_404), .ZN(n_0_8_352));
   INV_X1 i_0_8_429 (.A(n_0_8_352), .ZN(n_0_8_353));
   NAND2_X1 i_0_8_430 (.A1(n_0_8_633), .A2(n_0_8_404), .ZN(n_0_8_354));
   INV_X1 i_0_8_431 (.A(n_0_8_354), .ZN(n_0_8_355));
   AOI22_X1 i_0_8_432 (.A1(n_0_8_297), .A2(n_0_8_353), .B1(n_0_8_301), .B2(
      n_0_8_355), .ZN(n_0_8_356));
   NAND2_X1 i_0_8_433 (.A1(n_0_8_317), .A2(in2[14]), .ZN(n_0_8_357));
   NAND2_X1 i_0_8_434 (.A1(n_0_8_796), .A2(in1[14]), .ZN(n_0_8_358));
   NAND2_X1 i_0_8_435 (.A1(n_0_8_317), .A2(in2[14]), .ZN(n_0_8_359));
   NAND2_X1 i_0_8_436 (.A1(n_0_8_273), .A2(in2[13]), .ZN(n_0_8_360));
   NAND3_X1 i_0_8_385 (.A1(n_0_8_358), .A2(n_0_8_359), .A3(n_0_8_360), .ZN(
      n_0_8_377));
   INV_X1 i_0_8_438 (.A(in2[14]), .ZN(n_0_8_363));
   NAND2_X1 i_0_8_439 (.A1(n_0_8_363), .A2(in1[14]), .ZN(n_0_8_364));
   INV_X1 i_0_8_440 (.A(n_0_8_256), .ZN(n_0_8_365));
   AOI21_X1 i_0_8_148 (.A(n_0_8_365), .B1(n_0_8_519), .B2(n_0_8_517), .ZN(
      n_0_8_634));
   OAI22_X1 i_0_8_312 (.A1(n_0_8_371), .A2(n_0_8_633), .B1(n_0_8_567), .B2(
      n_0_8_383), .ZN(n_0_8_366));
   NAND2_X1 i_0_8_411 (.A1(n_0_8_368), .A2(in2[12]), .ZN(n_0_8_367));
   BUF_X1 i_0_8_412 (.A(n_0_8_571), .Z(n_0_8_368));
   INV_X1 i_0_8_420 (.A(n_0_8_571), .ZN(n_0_8_369));
   INV_X1 i_0_8_446 (.A(in2[12]), .ZN(n_0_8_370));
   OAI22_X1 i_0_8_321 (.A1(n_0_8_369), .A2(n_0_8_370), .B1(n_0_8_571), .B2(
      n_0_8_257), .ZN(n_0_8_371));
   AOI21_X1 i_0_8_448 (.A(n_0_8_289), .B1(n_0_34), .B2(in2[1]), .ZN(n_0_8_635));
   AOI22_X1 i_0_8_437 (.A1(n_0_8_594), .A2(n_0_8_368), .B1(n_0_8_259), .B2(
      n_0_8_832), .ZN(n_0_8_378));
   BUF_X1 i_0_8_0 (.A(n_0_8_636), .Z(n_0_8_383));
   INV_X1 i_0_8_451 (.A(n_0_8_633), .ZN(n_0_8_390));
   INV_X1 i_0_8_452 (.A(n_0_8_376), .ZN(n_0_8_391));
   NOR2_X1 i_0_8_453 (.A1(n_0_8_259), .A2(n_0_8_376), .ZN(n_0_8_393));
   INV_X1 i_0_8_454 (.A(n_0_8_594), .ZN(n_0_8_379));
   NOR2_X1 i_0_8_455 (.A1(n_0_8_636), .A2(n_0_8_379), .ZN(n_0_8_380));
   NAND2_X1 i_0_8_37 (.A1(n_0_8_368), .A2(n_0_8_380), .ZN(n_0_8_381));
   NAND2_X1 i_0_8_54 (.A1(n_0_8_655), .A2(n_0_8_381), .ZN(n_0_8_382));
   INV_X1 i_0_8_458 (.A(n_0_8_244), .ZN(n_0_8_638));
   NAND2_X1 i_0_8_459 (.A1(n_0_21), .A2(n_0_8_638), .ZN(n_0_8_639));
   BUF_X1 rt_shieldBuf__1__1__4 (.A(n_0_21), .Z(n_0_8_400));
   INV_X1 i_0_8_460 (.A(n_0_8_277), .ZN(n_0_8_384));
   XNOR2_X1 i_0_8_461 (.A(n_0_8_278), .B(n_0_8_384), .ZN(n_0_8_385));
   NOR2_X1 i_0_8_462 (.A1(n_0_8_385), .A2(n_0_8_319), .ZN(n_0_8_386));
   NOR2_X1 i_0_8_463 (.A1(n_0_8_458), .A2(n_0_8_386), .ZN(n_0_8_640));
   INV_X1 i_0_8_464 (.A(in2[13]), .ZN(n_0_8_387));
   XNOR2_X1 i_0_8_465 (.A(n_0_8_277), .B(n_0_8_387), .ZN(n_0_8_388));
   XNOR2_X1 i_0_8_466 (.A(n_0_8_388), .B(n_0_8_405), .ZN(n_0_8_389));
   NAND2_X1 i_0_8_467 (.A1(n_0_8_389), .A2(n_0_8_385), .ZN(n_0_8_641));
   INV_X1 i_0_8_468 (.A(n_0_8_633), .ZN(n_0_8_642));
   OAI21_X1 i_0_8_469 (.A(n_0_8_392), .B1(n_0_8_431), .B2(n_0_8_633), .ZN(
      n_0_8_403));
   XNOR2_X1 i_0_8_55 (.A(n_0_8_405), .B(n_0_8_314), .ZN(n_0_8_404));
   OAI21_X1 i_0_8_471 (.A(n_0_8_633), .B1(n_0_8_537), .B2(n_0_8_252), .ZN(
      n_0_8_392));
   INV_X1 i_0_8_445 (.A(in1[13]), .ZN(n_0_8_405));
   OAI21_X1 i_0_8_473 (.A(n_0_8_633), .B1(n_0_8_537), .B2(n_0_8_254), .ZN(
      n_0_8_394));
   NOR2_X1 i_0_8_347 (.A1(in2[13]), .A2(in1[13]), .ZN(n_0_8_395));
   NAND2_X1 i_0_8_348 (.A1(in2[13]), .A2(in1[13]), .ZN(n_0_8_396));
   INV_X1 i_0_8_390 (.A(n_0_8_396), .ZN(n_0_8_397));
   MUX2_X1 i_0_8_474 (.A(n_0_8_395), .B(n_0_8_397), .S(n_0_8_314), .Z(n_0_8_398));
   XNOR2_X1 i_0_8_475 (.A(in1[13]), .B(in2[13]), .ZN(n_0_8_399));
   INV_X1 i_0_8_476 (.A(n_0_8_292), .ZN(n_0_8_406));
   NAND2_X1 i_0_8_477 (.A1(n_0_8_399), .A2(n_0_8_406), .ZN(n_0_8_401));
   AOI21_X1 i_0_8_478 (.A(n_0_8_398), .B1(n_0_8_608), .B2(n_0_8_456), .ZN(
      n_0_8_402));
   XNOR2_X1 i_0_8_482 (.A(n_0_8_314), .B(in1[13]), .ZN(n_0_8_414));
   INV_X1 i_0_8_483 (.A(n_0_8_253), .ZN(n_0_8_455));
   INV_X1 i_0_8_484 (.A(n_0_8_252), .ZN(n_0_8_407));
   INV_X1 i_0_8_485 (.A(n_0_8_254), .ZN(n_0_8_408));
   OAI21_X1 i_0_8_479 (.A(n_0_8_407), .B1(n_0_8_414), .B2(n_0_8_408), .ZN(
      n_0_8_409));
   NAND2_X1 i_0_8_480 (.A1(n_0_8_399), .A2(n_0_8_408), .ZN(n_0_8_410));
   NAND2_X1 i_0_8_481 (.A1(n_0_8_409), .A2(n_0_8_410), .ZN(n_0_8_411));
   AOI22_X1 i_0_8_486 (.A1(n_0_8_754), .A2(n_0_8_608), .B1(n_0_8_633), .B2(
      n_0_8_411), .ZN(n_0_8_412));
   OAI21_X1 i_0_8_487 (.A(n_0_8_402), .B1(n_0_8_412), .B2(n_0_8_537), .ZN(
      n_0_8_485));
   NOR2_X1 i_0_8_491 (.A1(n_0_8_832), .A2(n_0_8_292), .ZN(n_0_8_413));
   INV_X1 i_0_8_493 (.A(n_0_8_292), .ZN(n_0_8_415));
   NAND2_X1 i_0_8_367 (.A1(n_0_8_831), .A2(n_0_8_415), .ZN(n_0_8_416));
   NAND2_X1 i_0_8_450 (.A1(n_0_8_416), .A2(n_0_8_633), .ZN(n_0_8_417));
   OAI21_X1 i_0_8_492 (.A(n_0_8_417), .B1(n_0_8_454), .B2(n_0_8_633), .ZN(
      n_0_8_418));
   NAND2_X1 i_0_8_497 (.A1(n_0_21), .A2(in2[12]), .ZN(n_0_8_419));
   INV_X1 i_0_8_498 (.A(n_0_8_419), .ZN(n_0_8_420));
   AOI21_X1 i_0_8_499 (.A(n_0_8_420), .B1(n_0_34), .B2(in2[12]), .ZN(n_0_8_421));
   NAND2_X1 i_0_8_447 (.A1(n_0_8_550), .A2(n_0_8_421), .ZN(n_0_36));
   NAND2_X1 i_0_8_501 (.A1(n_0_8_423), .A2(n_0_8_424), .ZN(n_0_8_422));
   NAND2_X1 i_0_8_502 (.A1(n_0_8_310), .A2(n_0_8_311), .ZN(n_0_8_423));
   NAND2_X1 i_0_8_503 (.A1(n_0_8_313), .A2(n_0_8_633), .ZN(n_0_8_424));
   XNOR2_X1 i_0_8_504 (.A(n_0_8_405), .B(n_0_8_526), .ZN(n_0_8_425));
   NAND2_X1 i_0_8_505 (.A1(n_0_8_311), .A2(n_0_8_425), .ZN(n_0_8_426));
   INV_X1 i_0_8_506 (.A(n_0_8_426), .ZN(n_0_8_427));
   NAND2_X1 i_0_8_507 (.A1(n_0_8_633), .A2(n_0_8_425), .ZN(n_0_8_428));
   INV_X1 i_0_8_508 (.A(n_0_8_428), .ZN(n_0_8_429));
   AOI22_X1 i_0_8_509 (.A1(n_0_8_310), .A2(n_0_8_427), .B1(n_0_8_313), .B2(
      n_0_8_429), .ZN(n_0_8_430));
   NOR2_X1 i_0_8_510 (.A1(n_0_8_537), .A2(n_0_8_253), .ZN(n_0_8_431));
   INV_X1 i_0_8_511 (.A(n_0_8_537), .ZN(n_0_8_432));
   INV_X1 i_0_8_512 (.A(n_0_8_253), .ZN(n_0_8_433));
   NAND2_X1 i_0_8_513 (.A1(n_0_8_432), .A2(n_0_8_433), .ZN(n_0_8_434));
   NAND2_X1 i_0_8_514 (.A1(n_0_8_434), .A2(n_0_8_633), .ZN(n_0_8_435));
   OAI21_X1 i_0_8_515 (.A(n_0_8_435), .B1(n_0_8_457), .B2(n_0_8_633), .ZN(
      n_0_8_436));
   NAND2_X1 i_0_8_516 (.A1(n_0_8_477), .A2(n_0_8_404), .ZN(n_0_8_437));
   NAND2_X1 i_0_8_517 (.A1(n_0_8_418), .A2(n_0_8_844), .ZN(n_0_8_438));
   NAND3_X1 i_0_8_518 (.A1(n_0_8_437), .A2(n_0_8_438), .A3(n_0_8_714), .ZN(
      n_0_8_439));
   NAND2_X1 i_0_8_519 (.A1(n_0_8_482), .A2(n_0_8_821), .ZN(n_0_8_440));
   INV_X1 i_0_8_520 (.A(n_0_8_440), .ZN(n_0_8_441));
   NAND2_X1 i_0_8_521 (.A1(n_0_8_495), .A2(n_0_8_441), .ZN(n_0_8_442));
   INV_X1 i_0_8_522 (.A(n_0_8_714), .ZN(n_0_8_443));
   NAND3_X1 i_0_8_523 (.A1(n_0_8_482), .A2(n_0_8_483), .A3(n_0_8_443), .ZN(
      n_0_8_444));
   NAND3_X1 i_0_8_524 (.A1(n_0_8_442), .A2(n_0_8_481), .A3(n_0_8_444), .ZN(
      n_0_8_445));
   INV_X1 i_0_8_525 (.A(n_0_8_445), .ZN(n_0_33));
   OAI22_X1 i_0_8_526 (.A1(n_0_8_542), .A2(n_0_8_633), .B1(n_0_8_452), .B2(
      n_0_8_636), .ZN(n_0_8_644));
   INV_X1 i_0_8_527 (.A(n_0_8_452), .ZN(n_0_8_446));
   INV_X1 i_0_8_528 (.A(n_0_8_636), .ZN(n_0_8_447));
   NAND2_X1 i_0_8_529 (.A1(n_0_8_446), .A2(n_0_8_447), .ZN(n_0_8_448));
   NAND2_X1 i_0_8_530 (.A1(n_0_8_448), .A2(n_0_8_542), .ZN(n_0_8_449));
   AOI22_X1 i_0_8_531 (.A1(n_0_8_452), .A2(n_0_8_633), .B1(n_0_8_636), .B2(
      n_0_8_633), .ZN(n_0_8_450));
   NAND2_X1 i_0_8_532 (.A1(n_0_8_449), .A2(n_0_8_450), .ZN(n_0_8_451));
   AOI22_X1 i_0_8_449 (.A1(n_0_8_571), .A2(n_0_8_246), .B1(n_0_8_749), .B2(
      n_0_8_292), .ZN(n_0_8_452));
   NAND2_X1 i_0_8_534 (.A1(n_0_8_749), .A2(n_0_8_254), .ZN(n_0_8_453));
   AOI22_X1 i_0_8_494 (.A1(n_0_8_571), .A2(n_0_8_248), .B1(n_0_8_749), .B2(
      n_0_8_254), .ZN(n_0_8_454));
   NOR2_X1 i_0_8_489 (.A1(n_0_8_749), .A2(n_0_8_401), .ZN(n_0_8_456));
   AOI22_X1 i_0_8_488 (.A1(n_0_8_571), .A2(n_0_8_309), .B1(n_0_8_749), .B2(
      n_0_8_252), .ZN(n_0_8_457));
   NAND2_X1 i_0_8_538 (.A1(n_0_8_459), .A2(n_0_8_460), .ZN(n_0_8_458));
   NAND4_X1 i_0_8_535 (.A1(n_0_8_664), .A2(n_0_8_677), .A3(n_0_8_674), .A4(
      n_0_8_665), .ZN(n_0_8_459));
   NAND2_X1 i_0_8_540 (.A1(n_0_8_511), .A2(n_0_8_700), .ZN(n_0_8_460));
   NAND2_X1 i_0_8_495 (.A1(n_0_8_498), .A2(n_0_8_497), .ZN(n_0_8_464));
   NAND2_X1 i_0_8_496 (.A1(n_0_8_796), .A2(in1[14]), .ZN(n_0_8_465));
   NAND2_X1 i_0_8_536 (.A1(n_0_8_320), .A2(in2[15]), .ZN(n_0_8_466));
   NAND2_X1 i_0_8_537 (.A1(n_0_8_321), .A2(in1[15]), .ZN(n_0_8_467));
   NAND2_X1 i_0_8_545 (.A1(n_0_8_571), .A2(n_0_8_255), .ZN(n_0_8_468));
   NAND2_X1 i_0_8_546 (.A1(n_0_8_749), .A2(n_0_8_253), .ZN(n_0_8_469));
   NAND2_X1 i_0_8_547 (.A1(n_0_8_468), .A2(n_0_8_469), .ZN(n_0_8_470));
   INV_X1 i_0_8_548 (.A(n_0_8_633), .ZN(n_0_8_471));
   NAND2_X1 i_0_8_549 (.A1(n_0_8_470), .A2(n_0_8_471), .ZN(n_0_8_472));
   NAND2_X1 i_0_8_550 (.A1(n_0_8_571), .A2(n_0_8_309), .ZN(n_0_8_473));
   NAND2_X1 i_0_8_551 (.A1(n_0_8_749), .A2(n_0_8_252), .ZN(n_0_8_474));
   NAND2_X1 i_0_8_552 (.A1(n_0_8_473), .A2(n_0_8_474), .ZN(n_0_8_475));
   NAND2_X1 i_0_8_553 (.A1(n_0_8_475), .A2(n_0_8_633), .ZN(n_0_8_476));
   NAND2_X1 i_0_8_554 (.A1(n_0_8_472), .A2(n_0_8_476), .ZN(n_0_8_477));
   NAND2_X1 i_0_8_424 (.A1(n_0_8_271), .A2(n_0_8_272), .ZN(n_0_8_700));
   NAND2_X1 i_0_8_539 (.A1(n_0_8_272), .A2(n_0_8_271), .ZN(n_0_8_479));
   OAI22_X1 i_0_8_557 (.A1(n_0_8_371), .A2(n_0_8_633), .B1(n_0_8_567), .B2(
      n_0_8_383), .ZN(n_0_8_480));
   NAND2_X1 i_0_8_558 (.A1(n_0_8_662), .A2(n_0_8_480), .ZN(n_0_8_481));
   NAND2_X1 i_0_8_341 (.A1(n_0_8_530), .A2(n_0_8_858), .ZN(n_0_30));
   AOI21_X1 i_0_8_560 (.A(n_0_8_521), .B1(n_0_34), .B2(in2[12]), .ZN(n_0_8_482));
   NAND2_X1 i_0_8_561 (.A1(n_0_8_484), .A2(n_0_8_714), .ZN(n_0_8_483));
   INV_X1 i_0_8_562 (.A(n_0_8_844), .ZN(n_0_8_484));
   NAND2_X1 i_0_8_563 (.A1(n_0_34), .A2(in2[12]), .ZN(n_0_8_486));
   NAND2_X1 i_0_8_564 (.A1(n_0_8_778), .A2(n_0_8_714), .ZN(n_0_8_487));
   NAND2_X1 i_0_8_565 (.A1(n_0_21), .A2(in2[12]), .ZN(n_0_8_492));
   INV_X1 i_0_8_566 (.A(n_0_8_492), .ZN(n_0_8_488));
   OAI22_X1 i_0_8_500 (.A1(n_0_8_318), .A2(n_0_8_302), .B1(n_0_8_571), .B2(
      n_0_8_594), .ZN(n_0_8_604));
   OAI22_X1 i_0_8_568 (.A1(n_0_8_618), .A2(n_0_8_383), .B1(n_0_8_496), .B2(
      n_0_8_633), .ZN(n_0_8_495));
   OAI22_X1 i_0_8_569 (.A1(n_0_8_318), .A2(n_0_8_302), .B1(n_0_8_571), .B2(
      n_0_8_594), .ZN(n_0_8_496));
   NAND2_X1 i_0_8_541 (.A1(n_0_8_499), .A2(in2[14]), .ZN(n_0_8_497));
   NAND2_X1 i_0_8_542 (.A1(n_0_8_500), .A2(in2[13]), .ZN(n_0_8_498));
   INV_X1 i_0_8_572 (.A(in1[14]), .ZN(n_0_8_499));
   INV_X1 i_0_8_573 (.A(in1[13]), .ZN(n_0_8_500));
   INV_X1 i_0_8_574 (.A(in1[14]), .ZN(n_0_8_501));
   NAND2_X1 i_0_8_533 (.A1(n_0_8_501), .A2(in2[14]), .ZN(n_0_8_489));
   INV_X1 i_0_8_576 (.A(in1[13]), .ZN(n_0_8_503));
   NAND2_X1 i_0_8_555 (.A1(n_0_8_503), .A2(in2[13]), .ZN(n_0_8_493));
   NAND2_X1 i_0_8_543 (.A1(n_0_8_779), .A2(n_0_8_821), .ZN(n_0_8_502));
   NAND2_X1 i_0_8_441 (.A1(n_0_8_270), .A2(n_0_8_798), .ZN(n_0_8_702));
   NAND2_X1 i_0_8_544 (.A1(n_0_8_270), .A2(n_0_8_798), .ZN(n_0_8_511));
   INV_X1 i_0_8_582 (.A(n_0_8_247), .ZN(n_0_8_513));
   NOR2_X1 i_0_8_570 (.A1(n_0_8_715), .A2(n_0_8_513), .ZN(n_0_8_514));
   INV_X1 i_0_8_584 (.A(n_0_8_248), .ZN(n_0_8_515));
   NAND2_X1 i_0_8_442 (.A1(n_0_8_382), .A2(n_0_8_566), .ZN(n_0_8_504));
   NAND2_X1 i_0_8_443 (.A1(n_0_8_366), .A2(n_0_8_821), .ZN(n_0_8_507));
   NAND2_X1 i_0_8_588 (.A1(n_0_21), .A2(in2[12]), .ZN(n_0_8_508));
   NAND2_X1 i_0_8_589 (.A1(n_0_21), .A2(in2[12]), .ZN(n_0_8_520));
   INV_X1 i_0_8_590 (.A(n_0_8_520), .ZN(n_0_8_521));
   INV_X1 i_0_8_591 (.A(n_0_8_714), .ZN(n_0_8_649));
   BUF_X1 rt_shieldBuf__1__1__3 (.A(in2[13]), .Z(n_0_8_526));
   NAND2_X1 i_0_8_366 (.A1(n_0_8_382), .A2(n_0_8_821), .ZN(n_0_8_527));
   INV_X1 i_0_8_456 (.A(n_0_8_714), .ZN(n_0_8_528));
   AOI21_X1 i_0_8_457 (.A(n_0_8_528), .B1(n_0_8_676), .B2(n_0_8_844), .ZN(
      n_0_8_529));
   NAND2_X1 i_0_8_470 (.A1(n_0_8_527), .A2(n_0_8_529), .ZN(n_0_8_530));
   INV_X1 i_0_8_596 (.A(n_0_8_259), .ZN(n_0_8_531));
   AOI21_X1 i_0_8_597 (.A(n_0_8_531), .B1(n_0_8_519), .B2(n_0_8_517), .ZN(
      n_0_8_509));
   NAND4_X1 i_0_8_571 (.A1(n_0_8_464), .A2(n_0_8_465), .A3(n_0_8_466), .A4(
      n_0_8_467), .ZN(n_0_8_516));
   NAND4_X1 i_0_8_577 (.A1(n_0_8_464), .A2(n_0_8_465), .A3(n_0_8_466), .A4(
      n_0_8_467), .ZN(n_0_8_517));
   NAND2_X1 i_0_8_575 (.A1(n_0_8_511), .A2(n_0_8_479), .ZN(n_0_8_518));
   NAND2_X1 i_0_8_581 (.A1(n_0_8_519), .A2(n_0_8_459), .ZN(n_0_8_537));
   OAI22_X1 i_0_8_603 (.A1(n_0_8_518), .A2(n_0_8_515), .B1(n_0_8_516), .B2(
      n_0_8_515), .ZN(n_0_8_540));
   NAND2_X1 i_0_8_578 (.A1(n_0_8_511), .A2(n_0_8_479), .ZN(n_0_8_519));
   NOR2_X1 i_0_8_605 (.A1(n_0_8_514), .A2(n_0_8_540), .ZN(n_0_8_542));
   NOR2_X1 i_0_8_559 (.A1(n_0_8_514), .A2(n_0_8_540), .ZN(n_0_8_534));
   BUF_X1 rt_shieldBuf__1__1__5 (.A(n_0_8_714), .Z(n_0_8_535));
   NAND2_X1 i_0_8_580 (.A1(n_0_8_339), .A2(n_0_8_821), .ZN(n_0_8_548));
   NAND2_X1 i_0_8_583 (.A1(n_0_8_632), .A2(n_0_8_844), .ZN(n_0_8_549));
   NAND3_X1 i_0_8_600 (.A1(n_0_8_548), .A2(n_0_8_549), .A3(n_0_8_714), .ZN(
      n_0_8_550));
   INV_X1 i_0_8_601 (.A(in1[14]), .ZN(n_0_8_536));
   INV_X1 i_0_8_611 (.A(in1[15]), .ZN(n_0_8_538));
   INV_X1 i_0_8_612 (.A(in1[14]), .ZN(n_0_8_539));
   INV_X1 i_0_8_613 (.A(in1[15]), .ZN(n_0_8_541));
   INV_X1 i_0_8_614 (.A(in1[13]), .ZN(n_0_8_544));
   INV_X1 i_0_8_615 (.A(in2[13]), .ZN(n_0_8_545));
   INV_X1 i_0_8_616 (.A(in1[15]), .ZN(n_0_8_653));
   INV_X1 i_0_8_617 (.A(in2[15]), .ZN(n_0_8_654));
   NAND3_X1 i_0_8_618 (.A1(n_0_8_658), .A2(n_0_8_657), .A3(n_0_8_656), .ZN(
      n_0_8_582));
   NAND3_X1 i_0_8_619 (.A1(n_0_8_693), .A2(n_0_8_692), .A3(n_0_8_694), .ZN(
      n_0_8_583));
   NAND2_X1 i_0_8_620 (.A1(n_0_8_583), .A2(n_0_8_582), .ZN(n_0_8_546));
   NAND2_X1 i_0_8_621 (.A1(n_0_8_688), .A2(n_0_8_635), .ZN(n_0_8_606));
   INV_X1 i_0_8_592 (.A(n_0_8_612), .ZN(n_0_8_547));
   INV_X1 i_0_8_602 (.A(n_0_8_547), .ZN(n_0_8_608));
   OAI21_X1 i_0_8_608 (.A(n_0_8_547), .B1(n_0_8_571), .B2(n_0_8_594), .ZN(
      n_0_8_556));
   NAND2_X1 i_0_8_625 (.A1(n_0_8_547), .A2(n_0_8_597), .ZN(n_0_8_611));
   NAND2_X1 i_0_8_626 (.A1(n_0_8_590), .A2(n_0_8_591), .ZN(n_0_8_613));
   NAND2_X1 i_0_8_627 (.A1(n_0_8_590), .A2(n_0_8_591), .ZN(n_0_8_585));
   NAND2_X1 i_0_8_628 (.A1(n_0_8_631), .A2(n_0_8_613), .ZN(n_0_8_614));
   NAND2_X1 i_0_8_629 (.A1(n_0_8_613), .A2(n_0_8_606), .ZN(n_0_8_615));
   NAND2_X1 i_0_8_630 (.A1(n_0_8_585), .A2(n_0_8_589), .ZN(n_0_8_616));
   OAI22_X1 i_0_8_609 (.A1(n_0_8_572), .A2(n_0_8_376), .B1(n_0_8_571), .B2(
      n_0_8_315), .ZN(n_0_8_617));
   OAI22_X1 i_0_8_632 (.A1(n_0_8_572), .A2(n_0_8_376), .B1(n_0_8_571), .B2(
      n_0_8_315), .ZN(n_0_8_618));
   BUF_X1 rt_shieldBuf__1__1__6 (.A(n_0_34), .Z(n_0_8_619));
   BUF_X1 rt_shieldBuf__1__1__8 (.A(n_0_21), .Z(n_0_8_620));
   NAND2_X1 i_0_8_633 (.A1(n_0_8_586), .A2(in1[0]), .ZN(n_0_8_621));
   INV_X1 i_0_8_634 (.A(n_0_8_587), .ZN(n_0_8_586));
   INV_X1 i_0_8_635 (.A(n_0_8_587), .ZN(n_0_8_622));
   NAND2_X1 i_0_8_636 (.A1(n_0_8_622), .A2(in1[0]), .ZN(n_0_8_623));
   INV_X1 i_0_8_637 (.A(n_0_8_593), .ZN(n_0_8_624));
   NOR2_X1 i_0_8_638 (.A1(n_0_8_592), .A2(n_0_8_624), .ZN(n_0_8_625));
   NAND3_X1 i_0_8_639 (.A1(n_0_8_588), .A2(n_0_8_623), .A3(n_0_8_625), .ZN(
      n_0_8_626));
   NAND2_X1 i_0_8_640 (.A1(n_0_8_623), .A2(n_0_8_592), .ZN(n_0_8_627));
   NAND2_X1 i_0_8_641 (.A1(n_0_8_626), .A2(n_0_8_627), .ZN(n_0_8_628));
   INV_X1 i_0_8_642 (.A(n_0_8_628), .ZN(n_0_8_629));
   INV_X1 i_0_8_643 (.A(n_0_8_687), .ZN(n_0_8_631));
   OAI22_X1 i_0_8_610 (.A1(n_0_8_604), .A2(n_0_8_633), .B1(n_0_8_617), .B2(
      n_0_8_383), .ZN(n_0_8_632));
   NAND2_X1 i_0_8_645 (.A1(n_0_8_769), .A2(n_0_8_770), .ZN(n_0_8_557));
   INV_X1 i_0_8_646 (.A(n_0_8_844), .ZN(n_0_8_558));
   NAND2_X1 i_0_8_647 (.A1(n_0_8_821), .A2(n_0_8_287), .ZN(n_0_8_560));
   INV_X1 i_0_8_648 (.A(n_0_8_461), .ZN(n_0_8_562));
   NAND2_X1 i_0_8_649 (.A1(n_0_8_463), .A2(n_0_8_462), .ZN(n_0_8_461));
   NAND3_X1 i_0_8_650 (.A1(n_0_8_505), .A2(n_0_8_506), .A3(n_0_8_532), .ZN(
      n_0_8_462));
   NAND3_X1 i_0_8_651 (.A1(n_0_8_478), .A2(n_0_8_663), .A3(in1[13]), .ZN(
      n_0_8_463));
   NAND2_X1 i_0_8_652 (.A1(n_0_8_505), .A2(n_0_8_532), .ZN(n_0_8_478));
   INV_X1 i_0_8_653 (.A(in2[15]), .ZN(n_0_8_490));
   INV_X1 i_0_8_654 (.A(in1[15]), .ZN(n_0_8_491));
   INV_X1 i_0_8_655 (.A(in2[14]), .ZN(n_0_8_494));
   NAND2_X1 i_0_8_656 (.A1(n_0_8_494), .A2(in1[14]), .ZN(n_0_8_505));
   NAND2_X1 i_0_8_657 (.A1(n_0_8_663), .A2(in1[13]), .ZN(n_0_8_506));
   NAND2_X1 i_0_8_658 (.A1(n_0_8_494), .A2(in1[14]), .ZN(n_0_8_510));
   INV_X1 i_0_8_659 (.A(in1[14]), .ZN(n_0_8_512));
   NAND2_X1 i_0_8_660 (.A1(n_0_8_491), .A2(in2[15]), .ZN(n_0_8_522));
   NAND2_X1 i_0_8_661 (.A1(n_0_8_490), .A2(in1[15]), .ZN(n_0_8_523));
   INV_X1 i_0_8_662 (.A(in1[14]), .ZN(n_0_8_524));
   NAND2_X1 i_0_8_663 (.A1(n_0_8_524), .A2(in2[14]), .ZN(n_0_8_525));
   NAND2_X1 i_0_8_664 (.A1(n_0_8_512), .A2(in2[14]), .ZN(n_0_8_532));
   NAND2_X1 i_0_8_665 (.A1(n_0_8_576), .A2(n_0_8_510), .ZN(n_0_8_533));
   NAND2_X1 i_0_8_666 (.A1(n_0_8_523), .A2(n_0_8_522), .ZN(n_0_8_543));
   NAND2_X1 i_0_8_667 (.A1(n_0_8_512), .A2(in2[14]), .ZN(n_0_8_551));
   NAND2_X1 i_0_8_668 (.A1(n_0_8_494), .A2(in1[14]), .ZN(n_0_8_552));
   NAND2_X1 i_0_8_669 (.A1(n_0_8_491), .A2(in2[15]), .ZN(n_0_8_565));
   NAND2_X1 i_0_8_670 (.A1(n_0_8_490), .A2(in1[15]), .ZN(n_0_8_574));
   INV_X1 i_0_8_671 (.A(in2[13]), .ZN(n_0_8_575));
   NAND2_X1 i_0_8_672 (.A1(n_0_8_575), .A2(in1[13]), .ZN(n_0_8_576));
   NAND3_X1 i_0_8_673 (.A1(n_0_8_525), .A2(n_0_8_575), .A3(in1[13]), .ZN(
      n_0_8_577));
   INV_X1 i_0_8_674 (.A(in2[13]), .ZN(n_0_8_663));
   NAND4_X1 i_0_8_675 (.A1(n_0_8_577), .A2(n_0_8_552), .A3(n_0_8_565), .A4(
      n_0_8_574), .ZN(n_0_8_578));
   NAND3_X1 i_0_8_676 (.A1(n_0_8_533), .A2(n_0_8_543), .A3(n_0_8_551), .ZN(
      n_0_8_579));
   NAND2_X1 i_0_8_677 (.A1(n_0_8_578), .A2(n_0_8_579), .ZN(n_0_8_581));
   INV_X1 i_0_8_678 (.A(n_0_8_581), .ZN(n_0_8_563));
   XNOR2_X1 i_0_8_679 (.A(n_0_8_663), .B(in1[13]), .ZN(n_0_8_564));
   XNOR2_X1 i_0_8_680 (.A(n_0_8_601), .B(n_0_8_600), .ZN(n_0_8_666));
   INV_X1 i_0_8_681 (.A(n_0_8_600), .ZN(n_0_8_667));
   NAND2_X1 i_0_8_682 (.A1(n_0_8_666), .A2(n_0_8_667), .ZN(n_0_8_668));
   XNOR2_X1 i_0_8_683 (.A(n_0_8_600), .B(in1[13]), .ZN(n_0_8_669));
   XNOR2_X1 i_0_8_684 (.A(n_0_8_669), .B(n_0_8_663), .ZN(n_0_8_670));
   OAI21_X1 i_0_8_685 (.A(n_0_8_668), .B1(n_0_8_670), .B2(n_0_8_666), .ZN(
      n_0_8_671));
   INV_X1 i_0_8_686 (.A(n_0_8_638), .ZN(n_0_8_672));
   OAI21_X1 i_0_8_687 (.A(n_0_8_639), .B1(n_0_8_711), .B2(n_0_8_672), .ZN(
      n_0_8_673));
   BUF_X1 rt_shieldBuf__1__1__2 (.A(n_0_8_844), .Z(n_0_8_566));
   AOI21_X1 i_0_8_567 (.A(n_0_8_634), .B1(n_0_8_571), .B2(n_0_8_286), .ZN(
      n_0_8_675));
   OAI22_X1 i_0_8_587 (.A1(n_0_8_675), .A2(n_0_8_633), .B1(n_0_8_383), .B2(
      n_0_8_534), .ZN(n_0_8_676));
   AOI21_X1 i_0_8_490 (.A(n_0_8_634), .B1(n_0_8_571), .B2(n_0_8_286), .ZN(
      n_0_8_567));
   NAND2_X1 i_0_8_691 (.A1(n_0_8_644), .A2(n_0_8_844), .ZN(n_0_8_679));
   INV_X1 i_0_8_692 (.A(n_0_8_649), .ZN(n_0_8_680));
   NAND3_X1 i_0_8_693 (.A1(n_0_8_603), .A2(n_0_8_679), .A3(n_0_8_680), .ZN(
      n_0_8_681));
   XNOR2_X1 i_0_8_368 (.A(n_0_8_729), .B(n_0_8_595), .ZN(n_0_8_683));
   XNOR2_X1 i_0_8_695 (.A(n_0_8_729), .B(n_0_8_580), .ZN(n_0_8_684));
   NAND4_X1 i_0_8_697 (.A1(n_0_8_714), .A2(n_0_8_642), .A3(n_0_8_641), .A4(
      n_0_8_640), .ZN(n_0_8_686));
   NAND2_X1 i_0_8_698 (.A1(n_0_8_686), .A2(n_0_8_635), .ZN(n_0_8_687));
   NAND4_X1 i_0_8_699 (.A1(n_0_8_714), .A2(n_0_8_642), .A3(n_0_8_641), .A4(
      n_0_8_640), .ZN(n_0_8_688));
   NAND2_X1 i_0_8_700 (.A1(n_0_8_653), .A2(n_0_8_654), .ZN(n_0_8_568));
   NAND2_X1 i_0_8_701 (.A1(in2[15]), .A2(in1[15]), .ZN(n_0_8_569));
   BUF_X1 rt_shieldBuf__1__1__11 (.A(n_0_55), .Z(n_0_8_695));
   INV_X1 i_0_8_593 (.A(n_0_8_711), .ZN(n_0_34));
   INV_X1 i_0_8_598 (.A(n_0_8_660), .ZN(n_0_21));
   NAND2_X1 i_0_8_595 (.A1(n_0_8_713), .A2(n_0_8_660), .ZN(n_0_8_711));
   NAND3_X1 i_0_8_705 (.A1(n_0_8_658), .A2(n_0_8_657), .A3(n_0_8_656), .ZN(
      n_0_8_712));
   NAND2_X1 i_0_8_604 (.A1(n_0_8_691), .A2(n_0_8_712), .ZN(n_0_8_570));
   INV_X1 i_0_8_556 (.A(n_0_8_715), .ZN(n_0_8_571));
   NAND2_X1 i_0_8_585 (.A1(n_0_8_648), .A2(n_0_8_690), .ZN(n_0_8_715));
   NAND2_X1 i_0_8_586 (.A1(n_0_8_702), .A2(n_0_8_700), .ZN(n_0_8_648));
   NAND2_X1 i_0_8_690 (.A1(n_0_8_702), .A2(n_0_8_700), .ZN(n_0_8_716));
   NAND4_X1 i_0_8_711 (.A1(n_0_8_664), .A2(n_0_8_677), .A3(n_0_8_674), .A4(
      n_0_8_665), .ZN(n_0_8_717));
   NAND2_X1 i_0_8_712 (.A1(n_0_8_716), .A2(n_0_8_717), .ZN(n_0_8_572));
   NAND2_X1 i_0_8_360 (.A1(n_0_8_822), .A2(n_0_8_633), .ZN(n_0_8_719));
   INV_X1 i_0_8_363 (.A(n_0_8_719), .ZN(n_0_8_573));
   NAND2_X1 i_0_8_717 (.A1(n_0_8_787), .A2(n_0_8_633), .ZN(n_0_8_724));
   INV_X1 i_0_8_718 (.A(n_0_8_821), .ZN(n_0_8_725));
   NOR2_X1 i_0_8_719 (.A1(n_0_8_361), .A2(n_0_8_725), .ZN(n_0_8_726));
   NAND2_X1 i_0_8_376 (.A1(n_0_8_724), .A2(n_0_8_726), .ZN(n_0_8_584));
   NAND2_X1 i_0_8_721 (.A1(n_0_8_258), .A2(n_0_8_251), .ZN(n_0_8_596));
   NAND2_X1 i_0_8_722 (.A1(n_0_8_258), .A2(n_0_8_251), .ZN(n_0_8_598));
   OAI22_X1 i_0_8_631 (.A1(n_0_8_316), .A2(n_0_8_383), .B1(n_0_8_378), .B2(
      n_0_8_633), .ZN(n_0_8_602));
   NAND2_X1 i_0_8_702 (.A1(n_0_8_602), .A2(n_0_8_566), .ZN(n_0_8_599));
   NAND2_X1 i_0_8_703 (.A1(n_0_8_605), .A2(n_0_8_821), .ZN(n_0_8_603));
   OAI22_X1 i_0_8_708 (.A1(n_0_8_316), .A2(n_0_8_383), .B1(n_0_8_378), .B2(
      n_0_8_633), .ZN(n_0_8_605));
   NAND2_X1 i_0_8_623 (.A1(n_0_8_570), .A2(n_0_8_103), .ZN(n_0_8_607));
   INV_X1 i_0_8_706 (.A(n_0_8_607), .ZN(n_0_8_609));
   OAI22_X1 i_0_8_332 (.A1(n_0_8_485), .A2(n_0_8_609), .B1(n_0_8_102), .B2(
      n_0_8_609), .ZN(n_0_8_610));
   NAND2_X1 i_0_8_731 (.A1(n_0_8_87), .A2(n_0_8_805), .ZN(n_0_84));
   BUF_X1 rt_shieldBuf__1__1__14 (.A(n_0_8_232), .Z(n_0_42));
   BUF_X1 rt_shieldBuf__1__1__15 (.A(n_0_8_596), .Z(n_0_52));
   NAND2_X1 i_0_8_728 (.A1(n_0_8_342), .A2(n_0_8_377), .ZN(n_0_8_612));
   NAND2_X1 i_0_8_724 (.A1(n_0_8_342), .A2(n_0_8_377), .ZN(n_0_8_630));
   INV_X1 i_0_8_606 (.A(n_0_8_630), .ZN(n_0_8_633));
   INV_X1 i_0_8_726 (.A(n_0_8_547), .ZN(n_0_8_636));
   INV_X1 i_0_8_594 (.A(n_0_8_572), .ZN(n_0_8_637));
   INV_X1 i_0_8_740 (.A(n_0_8_393), .ZN(n_0_8_643));
   INV_X1 i_0_8_741 (.A(n_0_8_391), .ZN(n_0_8_645));
   OAI21_X1 i_0_8_709 (.A(n_0_8_643), .B1(n_0_8_547), .B2(n_0_8_645), .ZN(
      n_0_8_646));
   OAI21_X1 i_0_8_733 (.A(n_0_8_637), .B1(n_0_8_827), .B2(n_0_8_646), .ZN(
      n_0_8_647));
   OAI21_X1 i_0_8_710 (.A(n_0_8_390), .B1(n_0_8_571), .B2(n_0_8_315), .ZN(
      n_0_8_650));
   NAND2_X1 i_0_8_745 (.A1(n_0_8_633), .A2(n_0_8_509), .ZN(n_0_8_651));
   NAND2_X1 i_0_8_738 (.A1(n_0_8_650), .A2(n_0_8_651), .ZN(n_0_8_652));
   NAND2_X1 i_0_8_622 (.A1(n_0_8_647), .A2(n_0_8_652), .ZN(n_0_8_655));
   NAND2_X1 i_0_8_748 (.A1(n_0_8_763), .A2(n_0_8_764), .ZN(n_0_8_656));
   NAND2_X1 i_0_8_749 (.A1(n_0_8_736), .A2(n_0_8_737), .ZN(n_0_8_657));
   NAND2_X1 i_0_8_750 (.A1(n_0_8_568), .A2(n_0_8_569), .ZN(n_0_8_658));
   NAND2_X1 i_0_8_751 (.A1(n_0_8_569), .A2(n_0_8_568), .ZN(n_0_8_659));
   NAND3_X1 i_0_8_752 (.A1(n_0_8_659), .A2(n_0_8_767), .A3(n_0_8_739), .ZN(
      n_0_8_660));
   NAND3_X1 i_0_8_753 (.A1(n_0_8_487), .A2(n_0_8_486), .A3(n_0_8_508), .ZN(
      n_0_8_661));
   INV_X1 i_0_8_754 (.A(n_0_8_661), .ZN(n_0_8_662));
   NAND2_X1 i_0_8_734 (.A1(n_0_8_489), .A2(n_0_8_493), .ZN(n_0_8_664));
   NAND2_X1 i_0_8_735 (.A1(n_0_8_320), .A2(in2[15]), .ZN(n_0_8_665));
   NAND2_X1 i_0_8_736 (.A1(n_0_8_321), .A2(in1[15]), .ZN(n_0_8_674));
   NAND2_X1 i_0_8_755 (.A1(n_0_8_796), .A2(in1[14]), .ZN(n_0_8_677));
   NAND2_X1 i_0_8_730 (.A1(n_0_8_493), .A2(n_0_8_489), .ZN(n_0_8_678));
   NAND2_X1 i_0_8_737 (.A1(n_0_8_796), .A2(in1[14]), .ZN(n_0_8_682));
   NAND2_X1 i_0_8_744 (.A1(n_0_8_320), .A2(in2[15]), .ZN(n_0_8_685));
   NAND2_X1 i_0_8_759 (.A1(n_0_8_321), .A2(in1[15]), .ZN(n_0_8_689));
   NAND4_X1 i_0_8_607 (.A1(n_0_8_678), .A2(n_0_8_682), .A3(n_0_8_685), .A4(
      n_0_8_689), .ZN(n_0_8_690));
   NAND3_X1 i_0_8_764 (.A1(n_0_8_692), .A2(n_0_8_693), .A3(n_0_8_694), .ZN(
      n_0_8_691));
   NAND2_X1 i_0_8_765 (.A1(n_0_8_553), .A2(n_0_8_555), .ZN(n_0_8_692));
   NAND3_X1 i_0_8_766 (.A1(n_0_8_561), .A2(n_0_8_559), .A3(in1[13]), .ZN(
      n_0_8_693));
   NAND2_X1 i_0_8_767 (.A1(n_0_8_554), .A2(in1[15]), .ZN(n_0_8_694));
   NOR2_X1 i_0_8_768 (.A1(n_0_8_536), .A2(in2[14]), .ZN(n_0_8_553));
   NAND2_X1 i_0_8_769 (.A1(n_0_8_538), .A2(in2[15]), .ZN(n_0_8_555));
   NAND2_X1 i_0_8_770 (.A1(n_0_8_541), .A2(in2[15]), .ZN(n_0_8_561));
   NAND2_X1 i_0_8_771 (.A1(n_0_8_539), .A2(in2[14]), .ZN(n_0_8_559));
   INV_X1 i_0_8_772 (.A(in2[15]), .ZN(n_0_8_554));
   INV_X1 i_0_8_773 (.A(in1[15]), .ZN(n_0_8_696));
   NAND3_X1 i_0_8_774 (.A1(n_0_8_539), .A2(n_0_8_696), .A3(in2[14]), .ZN(
      n_0_8_697));
   INV_X1 i_0_8_775 (.A(in1[13]), .ZN(n_0_8_698));
   NAND2_X1 i_0_8_776 (.A1(n_0_8_696), .A2(n_0_8_698), .ZN(n_0_8_699));
   INV_X1 i_0_8_777 (.A(in2[15]), .ZN(n_0_8_701));
   NAND3_X1 i_0_8_778 (.A1(n_0_8_697), .A2(n_0_8_699), .A3(n_0_8_701), .ZN(
      n_0_8_703));
   NAND2_X1 i_0_8_779 (.A1(n_0_8_538), .A2(in2[15]), .ZN(n_0_8_704));
   NOR2_X1 i_0_8_780 (.A1(n_0_8_536), .A2(in2[14]), .ZN(n_0_8_705));
   NAND2_X1 i_0_8_781 (.A1(n_0_8_704), .A2(n_0_8_705), .ZN(n_0_8_706));
   NAND2_X1 i_0_8_782 (.A1(n_0_8_539), .A2(in2[14]), .ZN(n_0_8_707));
   NOR2_X1 i_0_8_783 (.A1(n_0_8_541), .A2(n_0_8_698), .ZN(n_0_8_708));
   NAND2_X1 i_0_8_784 (.A1(n_0_8_707), .A2(n_0_8_708), .ZN(n_0_8_709));
   NAND3_X1 i_0_8_58 (.A1(n_0_8_703), .A2(n_0_8_706), .A3(n_0_8_709), .ZN(
      n_0_8_710));
   INV_X1 i_0_8_444 (.A(n_0_8_710), .ZN(n_0_8_713));
   INV_X1 i_0_8_644 (.A(n_0_8_546), .ZN(n_0_8_714));
   NAND2_X1 i_0_8_788 (.A1(n_0_8_403), .A2(n_0_8_404), .ZN(n_0_8_718));
   AOI21_X1 i_0_8_789 (.A(n_0_8_546), .B1(n_0_8_343), .B2(n_0_8_844), .ZN(
      n_0_8_720));
   NAND2_X1 i_0_8_790 (.A1(n_0_8_718), .A2(n_0_8_720), .ZN(n_0_8_721));
   NAND3_X1 i_0_8_579 (.A1(n_0_8_848), .A2(n_0_8_584), .A3(n_0_8_714), .ZN(
      n_0_8_722));
   NAND2_X1 i_0_8_794 (.A1(n_0_21), .A2(in2[12]), .ZN(n_0_8_723));
   INV_X1 i_0_8_795 (.A(n_0_8_723), .ZN(n_0_8_727));
   AOI21_X1 i_0_8_694 (.A(n_0_8_727), .B1(n_0_34), .B2(in2[12]), .ZN(n_0_8_728));
   NAND2_X1 i_0_8_720 (.A1(n_0_8_722), .A2(n_0_8_728), .ZN(n_0_8_729));
   NAND2_X1 i_0_8_727 (.A1(n_0_8_502), .A2(n_0_8_535), .ZN(n_0_8_730));
   INV_X1 i_0_8_729 (.A(n_0_8_730), .ZN(n_0_8_731));
   NAND2_X1 i_0_8_761 (.A1(n_0_8_599), .A2(n_0_8_731), .ZN(n_0_8_732));
   AOI22_X1 i_0_8_798 (.A1(n_0_8_276), .A2(in2[11]), .B1(n_0_8_400), .B2(in2[11]), 
      .ZN(n_0_8_733));
   NAND2_X1 i_0_8_799 (.A1(n_0_8_732), .A2(n_0_8_733), .ZN(n_0_25));
   OAI21_X1 i_0_8_803 (.A(n_0_8_51), .B1(n_0_8_61), .B2(n_0_8_57), .ZN(n_0_8_734));
   NAND2_X1 i_0_8_707 (.A1(n_0_8_734), .A2(sub), .ZN(n_0_8_735));
   NAND2_X1 i_0_8_805 (.A1(in2[14]), .A2(in1[14]), .ZN(n_0_8_736));
   NAND2_X1 i_0_8_806 (.A1(n_0_8_791), .A2(n_0_8_790), .ZN(n_0_8_737));
   NAND2_X1 i_0_8_807 (.A1(in2[14]), .A2(in1[14]), .ZN(n_0_8_738));
   NAND2_X1 i_0_8_808 (.A1(n_0_8_794), .A2(n_0_8_738), .ZN(n_0_8_739));
   NAND2_X1 i_0_8_809 (.A1(n_0_8_263), .A2(n_0_8_150), .ZN(n_0_59));
   INV_X1 i_0_8_810 (.A(n_0_8_263), .ZN(n_0_8_740));
   NAND2_X1 i_0_8_811 (.A1(n_0_8_740), .A2(sub), .ZN(n_0_8_741));
   INV_X1 i_0_8_812 (.A(sub), .ZN(n_0_8_742));
   OAI21_X1 i_0_8_813 (.A(n_0_8_741), .B1(n_0_8_150), .B2(n_0_8_742), .ZN(
      n_0_8_743));
   INV_X1 i_0_8_814 (.A(n_0_8_557), .ZN(n_0_8_744));
   NAND2_X1 i_0_8_815 (.A1(n_0_8_743), .A2(n_0_8_744), .ZN(n_0_8_745));
   NAND2_X1 i_0_8_816 (.A1(n_0_8_740), .A2(n_0_8_742), .ZN(n_0_8_746));
   OAI21_X1 i_0_8_817 (.A(n_0_8_746), .B1(n_0_8_150), .B2(sub), .ZN(n_0_8_747));
   NAND2_X1 i_0_8_818 (.A1(n_0_8_747), .A2(n_0_8_557), .ZN(n_0_8_748));
   NAND2_X1 i_0_8_819 (.A1(n_0_8_745), .A2(n_0_8_748), .ZN(n_0_114));
   NAND2_X1 i_0_8_757 (.A1(n_0_8_516), .A2(n_0_8_518), .ZN(n_0_8_749));
   NAND2_X1 i_0_8_821 (.A1(n_0_8_406), .A2(n_0_8_455), .ZN(n_0_8_750));
   INV_X1 i_0_8_822 (.A(n_0_8_750), .ZN(n_0_8_751));
   NAND3_X1 i_0_8_758 (.A1(n_0_8_518), .A2(n_0_8_516), .A3(n_0_8_751), .ZN(
      n_0_8_752));
   NAND2_X1 i_0_8_787 (.A1(n_0_8_414), .A2(n_0_8_455), .ZN(n_0_8_753));
   NAND2_X1 i_0_8_820 (.A1(n_0_8_752), .A2(n_0_8_753), .ZN(n_0_8_754));
   INV_X1 i_0_8_826 (.A(n_0_8_563), .ZN(n_0_8_755));
   INV_X1 i_0_8_827 (.A(n_0_8_564), .ZN(n_0_8_756));
   INV_X1 i_0_8_828 (.A(n_0_8_562), .ZN(n_0_8_757));
   INV_X1 i_0_8_829 (.A(n_0_8_245), .ZN(n_0_8_758));
   NAND2_X1 i_0_8_830 (.A1(n_0_8_757), .A2(n_0_8_758), .ZN(n_0_8_759));
   NAND2_X1 i_0_8_831 (.A1(n_0_8_249), .A2(n_0_8_759), .ZN(n_0_8_760));
   NOR2_X1 i_0_8_832 (.A1(n_0_8_564), .A2(n_0_8_563), .ZN(n_0_8_761));
   NAND2_X1 i_0_8_833 (.A1(n_0_8_760), .A2(n_0_8_761), .ZN(n_0_8_762));
   NAND2_X1 i_0_8_834 (.A1(in2[13]), .A2(in1[13]), .ZN(n_0_8_763));
   NAND2_X1 i_0_8_835 (.A1(n_0_8_545), .A2(n_0_8_544), .ZN(n_0_8_764));
   NAND2_X1 i_0_8_836 (.A1(n_0_8_544), .A2(n_0_8_545), .ZN(n_0_8_765));
   NAND2_X1 i_0_8_837 (.A1(in2[13]), .A2(in1[13]), .ZN(n_0_8_766));
   NAND2_X1 i_0_8_838 (.A1(n_0_8_765), .A2(n_0_8_766), .ZN(n_0_8_767));
   NAND2_X1 i_0_8_839 (.A1(n_0_8_769), .A2(n_0_8_770), .ZN(n_0_8_768));
   NAND2_X1 i_0_8_840 (.A1(n_0_8_374), .A2(n_0_8_375), .ZN(n_0_8_769));
   AOI21_X1 i_0_8_841 (.A(n_0_8_488), .B1(n_0_34), .B2(in2[12]), .ZN(n_0_8_770));
   NAND2_X1 i_0_8_842 (.A1(n_0_8_374), .A2(n_0_8_375), .ZN(n_0_8_771));
   INV_X1 i_0_8_843 (.A(n_0_8_771), .ZN(n_0_8_772));
   NAND2_X1 i_0_8_844 (.A1(n_0_34), .A2(in2[12]), .ZN(n_0_8_773));
   INV_X1 i_0_8_845 (.A(n_0_8_110), .ZN(n_0_8_774));
   XNOR2_X1 i_0_8_846 (.A(n_0_8_488), .B(n_0_8_774), .ZN(n_0_8_775));
   MUX2_X1 i_0_8_847 (.A(n_0_8_774), .B(n_0_8_775), .S(n_0_8_773), .Z(n_0_8_776));
   OAI22_X1 i_0_8_848 (.A1(n_0_8_772), .A2(n_0_8_776), .B1(n_0_8_771), .B2(
      n_0_8_774), .ZN(n_0_94));
   INV_X1 i_0_8_850 (.A(n_0_8_526), .ZN(n_0_8_777));
   XNOR2_X1 i_0_8_851 (.A(n_0_8_795), .B(n_0_8_777), .ZN(n_0_8_778));
   OAI22_X1 i_0_8_853 (.A1(n_0_8_567), .A2(n_0_8_633), .B1(n_0_8_534), .B2(
      n_0_8_383), .ZN(n_0_8_779));
   NAND2_X1 i_0_8_854 (.A1(n_0_21), .A2(in1[3]), .ZN(n_0_8_780));
   INV_X1 i_0_8_855 (.A(n_0_8_714), .ZN(n_0_8_781));
   INV_X1 i_0_8_856 (.A(in1[3]), .ZN(n_0_8_782));
   OAI21_X1 i_0_8_857 (.A(n_0_8_780), .B1(n_0_8_781), .B2(n_0_8_782), .ZN(
      n_0_8_783));
   AOI21_X1 i_0_8_858 (.A(n_0_8_783), .B1(n_0_8_243), .B2(n_0_34), .ZN(n_0_8_784));
   INV_X1 i_0_8_859 (.A(n_0_8_784), .ZN(n_0_40));
   INV_X1 i_0_8_860 (.A(n_0_8_571), .ZN(n_0_8_785));
   INV_X1 i_0_8_762 (.A(n_0_8_571), .ZN(n_0_8_786));
   OAI22_X1 i_0_8_599 (.A1(n_0_8_786), .A2(n_0_8_348), .B1(n_0_8_571), .B2(
      n_0_8_286), .ZN(n_0_8_787));
   NAND2_X1 i_0_8_863 (.A1(n_0_8_175), .A2(n_0_8_189), .ZN(n_0_8_788));
   NAND2_X1 i_0_8_804 (.A1(n_0_8_189), .A2(n_0_8_175), .ZN(n_0_8_789));
   INV_X1 i_0_8_866 (.A(in1[14]), .ZN(n_0_8_790));
   INV_X1 i_0_8_867 (.A(in2[14]), .ZN(n_0_8_791));
   INV_X1 i_0_8_868 (.A(in1[14]), .ZN(n_0_8_792));
   INV_X1 i_0_8_869 (.A(in2[14]), .ZN(n_0_8_793));
   NAND2_X1 i_0_8_870 (.A1(n_0_8_792), .A2(n_0_8_793), .ZN(n_0_8_794));
   BUF_X1 rt_shieldBuf__1__1__16 (.A(n_0_8_838), .Z(n_0_23));
   BUF_X1 rt_shieldBuf__1__1__17 (.A(n_0_8_405), .Z(n_0_8_795));
   INV_X1 i_0_8_801 (.A(in2[14]), .ZN(n_0_8_796));
   INV_X1 i_0_8_802 (.A(in2[14]), .ZN(n_0_8_797));
   NAND2_X1 i_0_8_624 (.A1(n_0_8_797), .A2(in1[14]), .ZN(n_0_8_798));
   NAND2_X1 i_0_8_39 (.A1(n_0_8_49), .A2(n_0_8_804), .ZN(n_0_8_799));
   NAND2_X1 i_0_8_865 (.A1(n_0_8_799), .A2(n_0_54), .ZN(n_0_8_800));
   NAND2_X1 i_0_8_874 (.A1(n_0_8_49), .A2(n_0_8_804), .ZN(n_0_22));
   INV_X1 i_0_8_871 (.A(n_0_8_789), .ZN(n_0_8_801));
   NAND2_X1 i_0_8_46 (.A1(n_0_8_610), .A2(n_0_8_100), .ZN(n_0_8_802));
   NAND2_X1 i_0_8_383 (.A1(n_0_8_610), .A2(n_0_8_100), .ZN(n_0_63));
   INV_X1 i_0_8_715 (.A(n_0_63), .ZN(n_0_8_803));
   NAND2_X1 i_0_8_716 (.A1(n_0_63), .A2(n_0_8_50), .ZN(n_0_8_804));
   NAND2_X1 i_0_8_756 (.A1(n_0_8_802), .A2(n_0_8_95), .ZN(n_0_8_805));
   INV_X1 i_0_8_852 (.A(n_0_8_802), .ZN(n_0_8_806));
   NAND2_X1 i_0_8_713 (.A1(n_0_8_573), .A2(n_0_8_787), .ZN(n_0_8_807));
   AOI22_X1 i_0_8_714 (.A1(n_0_8_558), .A2(n_0_8_560), .B1(n_0_8_822), .B2(
      n_0_8_361), .ZN(n_0_8_808));
   NAND2_X1 i_0_8_763 (.A1(n_0_8_807), .A2(n_0_8_808), .ZN(n_0_8_809));
   BUF_X1 rt_shieldBuf__1__1__18 (.A(n_0_8_21), .Z(n_0_8_810));
   OAI22_X1 i_0_8_873 (.A1(n_0_8_261), .A2(n_0_8_562), .B1(n_0_8_233), .B2(
      n_0_8_262), .ZN(n_0_8_811));
   NAND2_X1 i_0_8_849 (.A1(n_0_8_290), .A2(n_0_8_293), .ZN(n_0_8_812));
   NAND3_X1 i_0_8_861 (.A1(n_0_8_344), .A2(n_0_8_345), .A3(n_0_8_714), .ZN(
      n_0_8_290));
   AOI21_X1 i_0_8_862 (.A(n_0_8_347), .B1(n_0_34), .B2(in2[5]), .ZN(n_0_8_293));
   NAND3_X1 i_0_8_864 (.A1(n_0_8_344), .A2(n_0_8_345), .A3(n_0_8_714), .ZN(
      n_0_8_813));
   INV_X1 i_0_8_875 (.A(n_0_8_813), .ZN(n_0_8_814));
   NAND2_X1 i_0_8_876 (.A1(n_0_8_814), .A2(sub), .ZN(n_0_8_815));
   NAND2_X1 i_0_8_877 (.A1(n_0_34), .A2(in2[5]), .ZN(n_0_8_816));
   INV_X1 i_0_8_878 (.A(sub), .ZN(n_0_8_817));
   XNOR2_X1 i_0_8_879 (.A(n_0_8_347), .B(n_0_8_817), .ZN(n_0_8_818));
   MUX2_X1 i_0_8_880 (.A(n_0_8_817), .B(n_0_8_818), .S(n_0_8_816), .Z(n_0_8_819));
   OAI21_X1 i_0_8_881 (.A(n_0_8_815), .B1(n_0_8_819), .B2(n_0_8_814), .ZN(
      n_0_8_820));
   BUF_X1 i_0_8_688 (.A(n_0_8_404), .Z(n_0_8_821));
   NAND2_X1 i_0_8_872 (.A1(n_0_8_404), .A2(n_0_8_287), .ZN(n_0_8_822));
   INV_X1 i_0_8_723 (.A(n_0_8_598), .ZN(n_0_8_823));
   NAND2_X1 i_0_8_732 (.A1(n_0_8_842), .A2(n_0_8_823), .ZN(n_0_8_824));
   INV_X1 i_0_8_825 (.A(n_0_8_376), .ZN(n_0_8_825));
   NAND3_X1 i_0_8_882 (.A1(n_0_8_519), .A2(n_0_8_517), .A3(n_0_8_825), .ZN(
      n_0_8_826));
   INV_X1 i_0_8_883 (.A(n_0_8_826), .ZN(n_0_8_827));
   NAND2_X1 i_0_8_696 (.A1(n_0_8_517), .A2(n_0_8_519), .ZN(n_0_8_828));
   AOI22_X1 i_0_8_791 (.A1(n_0_8_571), .A2(n_0_8_294), .B1(n_0_8_828), .B2(
      n_0_8_309), .ZN(n_0_8_829));
   NAND2_X1 i_0_8_792 (.A1(n_0_8_828), .A2(n_0_8_292), .ZN(n_0_8_830));
   INV_X1 i_0_8_824 (.A(n_0_8_832), .ZN(n_0_8_831));
   NAND2_X1 i_0_8_884 (.A1(n_0_8_517), .A2(n_0_8_519), .ZN(n_0_8_832));
   NAND3_X1 i_0_8_746 (.A1(n_0_8_848), .A2(n_0_8_584), .A3(n_0_8_714), .ZN(
      n_0_8_833));
   NAND2_X1 i_0_8_747 (.A1(n_0_21), .A2(in2[12]), .ZN(n_0_8_834));
   INV_X1 i_0_8_885 (.A(n_0_8_834), .ZN(n_0_8_835));
   AOI21_X1 i_0_8_886 (.A(n_0_8_835), .B1(n_0_34), .B2(in2[12]), .ZN(n_0_8_836));
   NAND2_X1 i_0_8_887 (.A1(n_0_8_833), .A2(n_0_8_836), .ZN(n_0_8_837));
   AND2_X1 i_0_8_796 (.A1(n_0_8_99), .A2(n_0_129), .ZN(n_0_8_838));
   NAND2_X1 i_0_8_797 (.A1(n_0_8_87), .A2(n_0_8_805), .ZN(n_0_8_839));
   NAND2_X1 i_0_8_800 (.A1(n_0_8_99), .A2(n_0_8_155), .ZN(n_0_8_840));
   INV_X1 i_0_8_888 (.A(n_0_8_840), .ZN(n_0_8_841));
   NAND2_X1 i_0_8_889 (.A1(n_0_8_839), .A2(n_0_8_841), .ZN(n_0_8_842));
   AOI22_X1 i_0_8_262 (.A1(n_0_8_373), .A2(n_0_8_372), .B1(n_0_8_556), .B2(
      n_0_8_362), .ZN(n_0_8_843));
   XNOR2_X1 i_0_8_689 (.A(n_0_8_405), .B(in2[13]), .ZN(n_0_8_844));
   NAND2_X1 i_0_8_793 (.A1(n_0_8_372), .A2(n_0_8_373), .ZN(n_0_8_845));
   NAND2_X1 i_0_8_890 (.A1(n_0_8_556), .A2(n_0_8_362), .ZN(n_0_8_846));
   XNOR2_X1 i_0_8_891 (.A(n_0_8_795), .B(n_0_8_526), .ZN(n_0_8_847));
   NAND3_X1 i_0_8_892 (.A1(n_0_8_845), .A2(n_0_8_846), .A3(n_0_8_847), .ZN(
      n_0_8_848));
   NAND2_X1 i_0_8_147 (.A1(n_0_8_250), .A2(n_0_8_234), .ZN(n_0_8_849));
   NAND2_X1 i_0_8_472 (.A1(n_0_8_235), .A2(n_0_8_756), .ZN(n_0_8_850));
   NAND3_X1 i_0_8_893 (.A1(n_0_8_849), .A2(n_0_8_850), .A3(n_0_34), .ZN(
      n_0_8_851));
   NAND2_X1 i_0_8_742 (.A1(n_0_8_820), .A2(n_0_8_801), .ZN(n_0_8_852));
   NAND2_X1 i_0_8_743 (.A1(n_0_8_62), .A2(n_0_8_77), .ZN(n_0_8_853));
   NAND2_X1 i_0_8_760 (.A1(n_0_8_62), .A2(n_0_8_77), .ZN(n_0_8_854));
   NAND2_X1 i_0_8_823 (.A1(n_0_8_820), .A2(n_0_8_801), .ZN(n_0_8_855));
   INV_X1 i_0_8_894 (.A(n_0_8_78), .ZN(n_0_8_856));
   NAND3_X1 i_0_8_895 (.A1(n_0_8_854), .A2(n_0_8_855), .A3(n_0_8_856), .ZN(
      n_0_8_857));
   OAI21_X1 i_0_8_704 (.A(in2[12]), .B1(n_0_34), .B2(n_0_21), .ZN(n_0_8_858));
   NAND3_X1 i_0_8_785 (.A1(n_0_8_507), .A2(n_0_8_504), .A3(n_0_8_714), .ZN(
      n_0_8_859));
   NAND2_X1 i_0_8_786 (.A1(n_0_21), .A2(in2[12]), .ZN(n_0_8_860));
   INV_X1 i_0_8_896 (.A(n_0_8_860), .ZN(n_0_8_861));
   AOI21_X1 i_0_8_897 (.A(n_0_8_861), .B1(n_0_34), .B2(in2[12]), .ZN(n_0_8_862));
   NAND2_X1 i_0_8_898 (.A1(n_0_8_859), .A2(n_0_8_862), .ZN(n_0_31));
   OR2_X1 i_0_8_725 (.A1(n_0_34), .A2(n_0_21), .ZN(n_0_8_863));
   OAI21_X1 i_0_8_739 (.A(in2[3]), .B1(n_0_34), .B2(n_0_21), .ZN(n_0_8_864));
   BUF_X1 rt_shieldBuf__1__1__19 (.A(n_0_8_155), .Z(n_0_129));
   XNOR2_X1 i_0_0_0 (.A(n_0_0_20), .B(n_0_36), .ZN(n_0_83));
   NAND2_X1 i_0_0_1 (.A1(n_0_0_0), .A2(n_0_0_31), .ZN(n_0_66));
   NAND2_X1 i_0_0_2 (.A1(n_0_0_23), .A2(n_0_0_15), .ZN(n_0_0_0));
   NAND2_X1 i_0_0_4 (.A1(n_0_0_4), .A2(n_0_0_1), .ZN(n_0_81));
   NAND2_X1 i_0_0_5 (.A1(n_0_0_2), .A2(n_0_0_23), .ZN(n_0_0_1));
   NAND2_X1 i_0_0_7 (.A1(n_0_0_3), .A2(n_0_0_15), .ZN(n_0_0_2));
   NAND2_X1 i_0_0_8 (.A1(n_0_45), .A2(n_0_33), .ZN(n_0_0_3));
   NAND2_X1 i_0_0_9 (.A1(n_0_0_5), .A2(n_0_0_17), .ZN(n_0_0_4));
   OAI21_X1 i_0_0_11 (.A(n_0_0_29), .B1(n_0_0_13), .B2(n_0_33), .ZN(n_0_0_5));
   NAND2_X1 i_0_0_15 (.A1(n_0_0_6), .A2(n_0_0_13), .ZN(n_0_89));
   NAND2_X1 i_0_0_16 (.A1(n_0_0_24), .A2(n_0_0_25), .ZN(n_0_0_6));
   NAND2_X1 i_0_0_19 (.A1(n_0_0_7), .A2(n_0_0_11), .ZN(n_0_90));
   NAND3_X1 i_0_0_20 (.A1(n_0_0_10), .A2(n_0_0_9), .A3(n_0_0_8), .ZN(n_0_0_7));
   NAND2_X1 i_0_0_21 (.A1(n_0_0_13), .A2(n_0_0_26), .ZN(n_0_0_8));
   NAND2_X1 i_0_0_23 (.A1(n_0_45), .A2(sub), .ZN(n_0_0_9));
   NAND2_X1 i_0_0_24 (.A1(n_0_0_16), .A2(n_0_0_15), .ZN(n_0_0_10));
   NAND4_X1 i_0_0_25 (.A1(n_0_0_12), .A2(n_0_0_14), .A3(n_0_0_16), .A4(n_0_0_15), 
      .ZN(n_0_0_11));
   NAND2_X1 i_0_0_26 (.A1(n_0_0_13), .A2(n_0_33), .ZN(n_0_0_12));
   INV_X1 i_0_0_27 (.A(n_0_45), .ZN(n_0_0_13));
   NAND2_X1 i_0_0_28 (.A1(n_0_45), .A2(n_0_0_20), .ZN(n_0_0_14));
   NAND2_X1 i_0_0_6 (.A1(n_0_36), .A2(n_0_49), .ZN(n_0_0_15));
   NAND2_X1 i_0_0_31 (.A1(n_0_0_18), .A2(n_0_0_19), .ZN(n_0_0_16));
   AOI21_X1 i_0_0_34 (.A(n_0_0_20), .B1(n_0_36), .B2(n_0_0_19), .ZN(n_0_0_17));
   INV_X1 i_0_0_18 (.A(n_0_36), .ZN(n_0_0_18));
   INV_X1 i_0_0_22 (.A(n_0_49), .ZN(n_0_0_19));
   INV_X1 i_0_0_30 (.A(sub), .ZN(n_0_0_20));
   NAND2_X1 i_0_0_35 (.A1(n_0_36), .A2(n_0_0_20), .ZN(n_0_0_21));
   NAND2_X1 i_0_0_36 (.A1(n_0_49), .A2(n_0_0_20), .ZN(n_0_0_22));
   NAND2_X1 i_0_0_37 (.A1(n_0_0_21), .A2(n_0_0_22), .ZN(n_0_0_23));
   NAND2_X1 i_0_0_13 (.A1(n_0_0_26), .A2(n_0_0_20), .ZN(n_0_0_24));
   NAND2_X1 i_0_0_14 (.A1(n_0_33), .A2(sub), .ZN(n_0_0_25));
   INV_X1 i_0_0_33 (.A(n_0_33), .ZN(n_0_0_26));
   NAND2_X1 i_0_0_39 (.A1(n_0_0_26), .A2(sub), .ZN(n_0_0_27));
   NAND2_X1 i_0_0_41 (.A1(n_0_33), .A2(n_0_0_20), .ZN(n_0_0_28));
   AOI21_X1 i_0_0_42 (.A(n_0_0_13), .B1(n_0_0_27), .B2(n_0_0_28), .ZN(n_0_82));
   NAND2_X1 i_0_0_3 (.A1(n_0_0_18), .A2(n_0_49), .ZN(n_0_0_29));
   NAND2_X1 i_0_0_10 (.A1(n_0_0_19), .A2(n_0_36), .ZN(n_0_0_30));
   NAND3_X1 i_0_0_12 (.A1(n_0_0_29), .A2(n_0_0_30), .A3(sub), .ZN(n_0_0_31));
   INV_X1 i_0_1_0 (.A(n_0_24), .ZN(n_0_1_0));
   OAI21_X1 i_0_1_1 (.A(n_0_1_0), .B1(n_0_1_17), .B2(n_0_44), .ZN(n_0_1_1));
   OAI21_X1 i_0_1_2 (.A(n_0_44), .B1(n_0_1_17), .B2(n_0_37), .ZN(n_0_1_2));
   NAND2_X1 i_0_1_3 (.A1(n_0_1_17), .A2(n_0_37), .ZN(n_0_1_3));
   NAND3_X1 i_0_1_4 (.A1(n_0_1_1), .A2(n_0_1_2), .A3(n_0_1_3), .ZN(n_0_1_4));
   NAND2_X1 i_0_1_5 (.A1(n_0_1_4), .A2(sub), .ZN(n_0_1_5));
   OAI21_X1 i_0_1_6 (.A(n_0_44), .B1(n_0_25), .B2(n_0_37), .ZN(n_0_1_6));
   OAI21_X1 i_0_1_7 (.A(n_0_24), .B1(n_0_44), .B2(n_0_25), .ZN(n_0_1_7));
   NAND2_X1 i_0_1_8 (.A1(n_0_25), .A2(n_0_37), .ZN(n_0_1_8));
   NAND3_X1 i_0_1_9 (.A1(n_0_1_6), .A2(n_0_1_7), .A3(n_0_1_8), .ZN(n_0_1_9));
   NAND2_X1 i_0_1_10 (.A1(n_0_1_9), .A2(n_0_1_15), .ZN(n_0_1_10));
   NAND2_X1 i_0_1_11 (.A1(n_0_1_5), .A2(n_0_1_10), .ZN(n_0_126));
   XNOR2_X1 i_0_1_12 (.A(sub), .B(n_0_1_19), .ZN(n_0_1_11));
   INV_X1 i_0_1_13 (.A(n_0_37), .ZN(n_0_1_12));
   NAND2_X1 i_0_1_14 (.A1(n_0_1_11), .A2(n_0_1_12), .ZN(n_0_118));
   XNOR2_X1 i_0_1_15 (.A(n_0_1_18), .B(n_0_44), .ZN(n_0_1_13));
   XNOR2_X1 i_0_1_16 (.A(n_0_1_13), .B(sub), .ZN(n_0_115));
   XNOR2_X1 i_0_1_17 (.A(n_0_1_15), .B(n_0_24), .ZN(n_0_104));
   NAND2_X1 i_0_1_18 (.A1(n_0_1_16), .A2(n_0_1_14), .ZN(n_0_105));
   NAND2_X1 i_0_1_19 (.A1(n_0_25), .A2(n_0_1_15), .ZN(n_0_1_14));
   INV_X1 i_0_1_20 (.A(sub), .ZN(n_0_1_15));
   NAND2_X1 i_0_1_21 (.A1(n_0_1_17), .A2(sub), .ZN(n_0_1_16));
   INV_X1 i_0_1_22 (.A(n_0_25), .ZN(n_0_1_17));
   BUF_X1 rt_shieldBuf__1__1__20 (.A(n_0_25), .Z(n_0_1_18));
   BUF_X1 rt_shieldBuf__1__1__21 (.A(n_0_24), .Z(n_0_1_19));
endmodule
